module tuple (
  output [2:0] out1,
  output [3:0] out2,
  output [3:0] out3,
  output [3:0] out4,
  output [2:0] out5,
  output [2:0] out6
);

assign out1 = 3'd7;
assign out2 = 4'd8;
assign out3 = 4'd9;
assign out4 = 4'd10;
assign out5 = 3'd7;
assign out6 = 3'd6;

endmodule
