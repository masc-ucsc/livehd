module package_Anon_46(
  input  [19:0] io_x_ppn,
  input         io_x_u,
  input         io_x_ae,
  input         io_x_sw,
  input         io_x_sx,
  input         io_x_sr,
  input         io_x_pw,
  input         io_x_px,
  input         io_x_pr,
  input         io_x_pal,
  input         io_x_paa,
  input         io_x_eff,
  input         io_x_c,
  output [19:0] io_y_ppn,
  output        io_y_u,
  output        io_y_ae,
  output        io_y_sw,
  output        io_y_sx,
  output        io_y_sr,
  output        io_y_pw,
  output        io_y_px,
  output        io_y_pr,
  output        io_y_pal,
  output        io_y_paa,
  output        io_y_eff,
  output        io_y_c
);
  assign io_y_ppn = io_x_ppn; // @[package.scala 218:12]
  assign io_y_u = io_x_u; // @[package.scala 218:12]
  assign io_y_ae = io_x_ae; // @[package.scala 218:12]
  assign io_y_sw = io_x_sw; // @[package.scala 218:12]
  assign io_y_sx = io_x_sx; // @[package.scala 218:12]
  assign io_y_sr = io_x_sr; // @[package.scala 218:12]
  assign io_y_pw = io_x_pw; // @[package.scala 218:12]
  assign io_y_px = io_x_px; // @[package.scala 218:12]
  assign io_y_pr = io_x_pr; // @[package.scala 218:12]
  assign io_y_pal = io_x_pal; // @[package.scala 218:12]
  assign io_y_paa = io_x_paa; // @[package.scala 218:12]
  assign io_y_eff = io_x_eff; // @[package.scala 218:12]
  assign io_y_c = io_x_c; // @[package.scala 218:12]
endmodule
module PMPChecker_1(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  input  [1:0]  io_size,
  output        io_r,
  output        io_w,
  output        io_x
);
  wire  default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  wire [5:0] _T_3 = 6'h7 << io_size; // @[package.scala 189:77]
  wire [2:0] _T_5 = ~_T_3[2:0]; // @[package.scala 189:46]
  wire [31:0] _GEN_0 = {{29'd0}, _T_5}; // @[PMP.scala 70:26]
  wire [31:0] _T_6 = io_pmp_7_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [31:0] _T_8 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_9 = ~_T_8; // @[PMP.scala 62:29]
  wire [31:0] _T_10 = _T_9 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_11 = ~_T_10; // @[PMP.scala 62:27]
  wire [28:0] _T_14 = io_addr[31:3] ^ _T_11[31:3]; // @[PMP.scala 65:47]
  wire [28:0] _T_15 = ~io_pmp_7_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_16 = _T_14 & _T_15; // @[PMP.scala 65:52]
  wire  _T_17 = _T_16 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_25 = io_addr[2:0] ^ _T_11[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_26 = ~_T_6[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_27 = _T_25 & _T_26; // @[PMP.scala 65:52]
  wire  _T_28 = _T_27 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_29 = _T_17 & _T_28; // @[PMP.scala 73:16]
  wire [31:0] _T_36 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_37 = ~_T_36; // @[PMP.scala 62:29]
  wire [31:0] _T_38 = _T_37 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_39 = ~_T_38; // @[PMP.scala 62:27]
  wire  _T_41 = io_addr[31:3] < _T_39[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_48 = io_addr[31:3] ^ _T_39[31:3]; // @[PMP.scala 83:41]
  wire  _T_49 = _T_48 == 29'h0; // @[PMP.scala 83:69]
  wire [2:0] _T_51 = io_addr[2:0] | _T_5; // @[PMP.scala 84:42]
  wire  _T_57 = _T_51 < _T_39[2:0]; // @[PMP.scala 84:53]
  wire  _T_59 = _T_41 | _T_49 & _T_57; // @[PMP.scala 85:16]
  wire  _T_60 = ~_T_59; // @[PMP.scala 90:5]
  wire  _T_67 = io_addr[31:3] < _T_11[31:3]; // @[PMP.scala 82:39]
  wire  _T_75 = _T_14 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_83 = io_addr[2:0] < _T_11[2:0]; // @[PMP.scala 84:53]
  wire  _T_85 = _T_67 | _T_75 & _T_83; // @[PMP.scala 85:16]
  wire  _T_86 = _T_60 & _T_85; // @[PMP.scala 96:48]
  wire  _T_88 = io_pmp_7_cfg_a[1] ? _T_29 : io_pmp_7_cfg_a[0] & _T_86; // @[PMP.scala 134:8]
  wire  _T_90 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_109 = ~io_addr[2:0]; // @[PMP.scala 125:125]
  wire [2:0] _T_110 = _T_39[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_112 = _T_49 & _T_110 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_128 = _T_11[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_130 = _T_75 & _T_128 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_132 = ~(_T_112 | _T_130); // @[PMP.scala 127:24]
  wire [2:0] _T_134 = ~io_pmp_7_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_135 = _T_5 & _T_134; // @[PMP.scala 128:32]
  wire  _T_136 = _T_135 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_138 = io_pmp_7_cfg_a[1] ? _T_136 : _T_132; // @[PMP.scala 129:8]
  wire  _T_191 = _T_138 & (io_pmp_7_cfg_r | _T_90); // @[PMP.scala 183:26]
  wire  _T_193 = _T_138 & (io_pmp_7_cfg_w | _T_90); // @[PMP.scala 184:26]
  wire  _T_195 = _T_138 & (io_pmp_7_cfg_x | _T_90); // @[PMP.scala 185:26]
  wire  _T_196_cfg_x = _T_88 ? _T_195 : default_; // @[PMP.scala 186:8]
  wire  _T_196_cfg_w = _T_88 ? _T_193 : default_; // @[PMP.scala 186:8]
  wire  _T_196_cfg_r = _T_88 ? _T_191 : default_; // @[PMP.scala 186:8]
  wire [31:0] _T_202 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_211 = ~io_pmp_6_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_212 = _T_48 & _T_211; // @[PMP.scala 65:52]
  wire  _T_213 = _T_212 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_221 = io_addr[2:0] ^ _T_39[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_222 = ~_T_202[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_223 = _T_221 & _T_222; // @[PMP.scala 65:52]
  wire  _T_224 = _T_223 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_225 = _T_213 & _T_224; // @[PMP.scala 73:16]
  wire [31:0] _T_232 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_233 = ~_T_232; // @[PMP.scala 62:29]
  wire [31:0] _T_234 = _T_233 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_235 = ~_T_234; // @[PMP.scala 62:27]
  wire  _T_237 = io_addr[31:3] < _T_235[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_244 = io_addr[31:3] ^ _T_235[31:3]; // @[PMP.scala 83:41]
  wire  _T_245 = _T_244 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_253 = _T_51 < _T_235[2:0]; // @[PMP.scala 84:53]
  wire  _T_255 = _T_237 | _T_245 & _T_253; // @[PMP.scala 85:16]
  wire  _T_256 = ~_T_255; // @[PMP.scala 90:5]
  wire  _T_279 = io_addr[2:0] < _T_39[2:0]; // @[PMP.scala 84:53]
  wire  _T_281 = _T_41 | _T_49 & _T_279; // @[PMP.scala 85:16]
  wire  _T_282 = _T_256 & _T_281; // @[PMP.scala 96:48]
  wire  _T_284 = io_pmp_6_cfg_a[1] ? _T_225 : io_pmp_6_cfg_a[0] & _T_282; // @[PMP.scala 134:8]
  wire  _T_286 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_306 = _T_235[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_308 = _T_245 & _T_306 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_324 = _T_39[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_326 = _T_49 & _T_324 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_328 = ~(_T_308 | _T_326); // @[PMP.scala 127:24]
  wire [2:0] _T_330 = ~io_pmp_6_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_331 = _T_5 & _T_330; // @[PMP.scala 128:32]
  wire  _T_332 = _T_331 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_334 = io_pmp_6_cfg_a[1] ? _T_332 : _T_328; // @[PMP.scala 129:8]
  wire  _T_387 = _T_334 & (io_pmp_6_cfg_r | _T_286); // @[PMP.scala 183:26]
  wire  _T_389 = _T_334 & (io_pmp_6_cfg_w | _T_286); // @[PMP.scala 184:26]
  wire  _T_391 = _T_334 & (io_pmp_6_cfg_x | _T_286); // @[PMP.scala 185:26]
  wire  _T_392_cfg_x = _T_284 ? _T_391 : _T_196_cfg_x; // @[PMP.scala 186:8]
  wire  _T_392_cfg_w = _T_284 ? _T_389 : _T_196_cfg_w; // @[PMP.scala 186:8]
  wire  _T_392_cfg_r = _T_284 ? _T_387 : _T_196_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_398 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_407 = ~io_pmp_5_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_408 = _T_244 & _T_407; // @[PMP.scala 65:52]
  wire  _T_409 = _T_408 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_417 = io_addr[2:0] ^ _T_235[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_418 = ~_T_398[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_419 = _T_417 & _T_418; // @[PMP.scala 65:52]
  wire  _T_420 = _T_419 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_421 = _T_409 & _T_420; // @[PMP.scala 73:16]
  wire [31:0] _T_428 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_429 = ~_T_428; // @[PMP.scala 62:29]
  wire [31:0] _T_430 = _T_429 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_431 = ~_T_430; // @[PMP.scala 62:27]
  wire  _T_433 = io_addr[31:3] < _T_431[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_440 = io_addr[31:3] ^ _T_431[31:3]; // @[PMP.scala 83:41]
  wire  _T_441 = _T_440 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_449 = _T_51 < _T_431[2:0]; // @[PMP.scala 84:53]
  wire  _T_451 = _T_433 | _T_441 & _T_449; // @[PMP.scala 85:16]
  wire  _T_452 = ~_T_451; // @[PMP.scala 90:5]
  wire  _T_475 = io_addr[2:0] < _T_235[2:0]; // @[PMP.scala 84:53]
  wire  _T_477 = _T_237 | _T_245 & _T_475; // @[PMP.scala 85:16]
  wire  _T_478 = _T_452 & _T_477; // @[PMP.scala 96:48]
  wire  _T_480 = io_pmp_5_cfg_a[1] ? _T_421 : io_pmp_5_cfg_a[0] & _T_478; // @[PMP.scala 134:8]
  wire  _T_482 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_502 = _T_431[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_504 = _T_441 & _T_502 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_520 = _T_235[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_522 = _T_245 & _T_520 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_524 = ~(_T_504 | _T_522); // @[PMP.scala 127:24]
  wire [2:0] _T_526 = ~io_pmp_5_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_527 = _T_5 & _T_526; // @[PMP.scala 128:32]
  wire  _T_528 = _T_527 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_530 = io_pmp_5_cfg_a[1] ? _T_528 : _T_524; // @[PMP.scala 129:8]
  wire  _T_583 = _T_530 & (io_pmp_5_cfg_r | _T_482); // @[PMP.scala 183:26]
  wire  _T_585 = _T_530 & (io_pmp_5_cfg_w | _T_482); // @[PMP.scala 184:26]
  wire  _T_587 = _T_530 & (io_pmp_5_cfg_x | _T_482); // @[PMP.scala 185:26]
  wire  _T_588_cfg_x = _T_480 ? _T_587 : _T_392_cfg_x; // @[PMP.scala 186:8]
  wire  _T_588_cfg_w = _T_480 ? _T_585 : _T_392_cfg_w; // @[PMP.scala 186:8]
  wire  _T_588_cfg_r = _T_480 ? _T_583 : _T_392_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_594 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_603 = ~io_pmp_4_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_604 = _T_440 & _T_603; // @[PMP.scala 65:52]
  wire  _T_605 = _T_604 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_613 = io_addr[2:0] ^ _T_431[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_614 = ~_T_594[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_615 = _T_613 & _T_614; // @[PMP.scala 65:52]
  wire  _T_616 = _T_615 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_617 = _T_605 & _T_616; // @[PMP.scala 73:16]
  wire [31:0] _T_624 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_625 = ~_T_624; // @[PMP.scala 62:29]
  wire [31:0] _T_626 = _T_625 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_627 = ~_T_626; // @[PMP.scala 62:27]
  wire  _T_629 = io_addr[31:3] < _T_627[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_636 = io_addr[31:3] ^ _T_627[31:3]; // @[PMP.scala 83:41]
  wire  _T_637 = _T_636 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_645 = _T_51 < _T_627[2:0]; // @[PMP.scala 84:53]
  wire  _T_647 = _T_629 | _T_637 & _T_645; // @[PMP.scala 85:16]
  wire  _T_648 = ~_T_647; // @[PMP.scala 90:5]
  wire  _T_671 = io_addr[2:0] < _T_431[2:0]; // @[PMP.scala 84:53]
  wire  _T_673 = _T_433 | _T_441 & _T_671; // @[PMP.scala 85:16]
  wire  _T_674 = _T_648 & _T_673; // @[PMP.scala 96:48]
  wire  _T_676 = io_pmp_4_cfg_a[1] ? _T_617 : io_pmp_4_cfg_a[0] & _T_674; // @[PMP.scala 134:8]
  wire  _T_678 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_698 = _T_627[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_700 = _T_637 & _T_698 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_716 = _T_431[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_718 = _T_441 & _T_716 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_720 = ~(_T_700 | _T_718); // @[PMP.scala 127:24]
  wire [2:0] _T_722 = ~io_pmp_4_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_723 = _T_5 & _T_722; // @[PMP.scala 128:32]
  wire  _T_724 = _T_723 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_726 = io_pmp_4_cfg_a[1] ? _T_724 : _T_720; // @[PMP.scala 129:8]
  wire  _T_779 = _T_726 & (io_pmp_4_cfg_r | _T_678); // @[PMP.scala 183:26]
  wire  _T_781 = _T_726 & (io_pmp_4_cfg_w | _T_678); // @[PMP.scala 184:26]
  wire  _T_783 = _T_726 & (io_pmp_4_cfg_x | _T_678); // @[PMP.scala 185:26]
  wire  _T_784_cfg_x = _T_676 ? _T_783 : _T_588_cfg_x; // @[PMP.scala 186:8]
  wire  _T_784_cfg_w = _T_676 ? _T_781 : _T_588_cfg_w; // @[PMP.scala 186:8]
  wire  _T_784_cfg_r = _T_676 ? _T_779 : _T_588_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_790 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_799 = ~io_pmp_3_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_800 = _T_636 & _T_799; // @[PMP.scala 65:52]
  wire  _T_801 = _T_800 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_809 = io_addr[2:0] ^ _T_627[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_810 = ~_T_790[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_811 = _T_809 & _T_810; // @[PMP.scala 65:52]
  wire  _T_812 = _T_811 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_813 = _T_801 & _T_812; // @[PMP.scala 73:16]
  wire [31:0] _T_820 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_821 = ~_T_820; // @[PMP.scala 62:29]
  wire [31:0] _T_822 = _T_821 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_823 = ~_T_822; // @[PMP.scala 62:27]
  wire  _T_825 = io_addr[31:3] < _T_823[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_832 = io_addr[31:3] ^ _T_823[31:3]; // @[PMP.scala 83:41]
  wire  _T_833 = _T_832 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_841 = _T_51 < _T_823[2:0]; // @[PMP.scala 84:53]
  wire  _T_843 = _T_825 | _T_833 & _T_841; // @[PMP.scala 85:16]
  wire  _T_844 = ~_T_843; // @[PMP.scala 90:5]
  wire  _T_867 = io_addr[2:0] < _T_627[2:0]; // @[PMP.scala 84:53]
  wire  _T_869 = _T_629 | _T_637 & _T_867; // @[PMP.scala 85:16]
  wire  _T_870 = _T_844 & _T_869; // @[PMP.scala 96:48]
  wire  _T_872 = io_pmp_3_cfg_a[1] ? _T_813 : io_pmp_3_cfg_a[0] & _T_870; // @[PMP.scala 134:8]
  wire  _T_874 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_894 = _T_823[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_896 = _T_833 & _T_894 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_912 = _T_627[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_914 = _T_637 & _T_912 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_916 = ~(_T_896 | _T_914); // @[PMP.scala 127:24]
  wire [2:0] _T_918 = ~io_pmp_3_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_919 = _T_5 & _T_918; // @[PMP.scala 128:32]
  wire  _T_920 = _T_919 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_922 = io_pmp_3_cfg_a[1] ? _T_920 : _T_916; // @[PMP.scala 129:8]
  wire  _T_975 = _T_922 & (io_pmp_3_cfg_r | _T_874); // @[PMP.scala 183:26]
  wire  _T_977 = _T_922 & (io_pmp_3_cfg_w | _T_874); // @[PMP.scala 184:26]
  wire  _T_979 = _T_922 & (io_pmp_3_cfg_x | _T_874); // @[PMP.scala 185:26]
  wire  _T_980_cfg_x = _T_872 ? _T_979 : _T_784_cfg_x; // @[PMP.scala 186:8]
  wire  _T_980_cfg_w = _T_872 ? _T_977 : _T_784_cfg_w; // @[PMP.scala 186:8]
  wire  _T_980_cfg_r = _T_872 ? _T_975 : _T_784_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_986 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_995 = ~io_pmp_2_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_996 = _T_832 & _T_995; // @[PMP.scala 65:52]
  wire  _T_997 = _T_996 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1005 = io_addr[2:0] ^ _T_823[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1006 = ~_T_986[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1007 = _T_1005 & _T_1006; // @[PMP.scala 65:52]
  wire  _T_1008 = _T_1007 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1009 = _T_997 & _T_1008; // @[PMP.scala 73:16]
  wire [31:0] _T_1016 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_1017 = ~_T_1016; // @[PMP.scala 62:29]
  wire [31:0] _T_1018 = _T_1017 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_1019 = ~_T_1018; // @[PMP.scala 62:27]
  wire  _T_1021 = io_addr[31:3] < _T_1019[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_1028 = io_addr[31:3] ^ _T_1019[31:3]; // @[PMP.scala 83:41]
  wire  _T_1029 = _T_1028 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_1037 = _T_51 < _T_1019[2:0]; // @[PMP.scala 84:53]
  wire  _T_1039 = _T_1021 | _T_1029 & _T_1037; // @[PMP.scala 85:16]
  wire  _T_1040 = ~_T_1039; // @[PMP.scala 90:5]
  wire  _T_1063 = io_addr[2:0] < _T_823[2:0]; // @[PMP.scala 84:53]
  wire  _T_1065 = _T_825 | _T_833 & _T_1063; // @[PMP.scala 85:16]
  wire  _T_1066 = _T_1040 & _T_1065; // @[PMP.scala 96:48]
  wire  _T_1068 = io_pmp_2_cfg_a[1] ? _T_1009 : io_pmp_2_cfg_a[0] & _T_1066; // @[PMP.scala 134:8]
  wire  _T_1070 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1090 = _T_1019[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_1092 = _T_1029 & _T_1090 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_1108 = _T_823[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1110 = _T_833 & _T_1108 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1112 = ~(_T_1092 | _T_1110); // @[PMP.scala 127:24]
  wire [2:0] _T_1114 = ~io_pmp_2_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1115 = _T_5 & _T_1114; // @[PMP.scala 128:32]
  wire  _T_1116 = _T_1115 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1118 = io_pmp_2_cfg_a[1] ? _T_1116 : _T_1112; // @[PMP.scala 129:8]
  wire  _T_1171 = _T_1118 & (io_pmp_2_cfg_r | _T_1070); // @[PMP.scala 183:26]
  wire  _T_1173 = _T_1118 & (io_pmp_2_cfg_w | _T_1070); // @[PMP.scala 184:26]
  wire  _T_1175 = _T_1118 & (io_pmp_2_cfg_x | _T_1070); // @[PMP.scala 185:26]
  wire  _T_1176_cfg_x = _T_1068 ? _T_1175 : _T_980_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_w = _T_1068 ? _T_1173 : _T_980_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_r = _T_1068 ? _T_1171 : _T_980_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1182 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_1191 = ~io_pmp_1_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_1192 = _T_1028 & _T_1191; // @[PMP.scala 65:52]
  wire  _T_1193 = _T_1192 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1201 = io_addr[2:0] ^ _T_1019[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1202 = ~_T_1182[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1203 = _T_1201 & _T_1202; // @[PMP.scala 65:52]
  wire  _T_1204 = _T_1203 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1205 = _T_1193 & _T_1204; // @[PMP.scala 73:16]
  wire [31:0] _T_1212 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_1213 = ~_T_1212; // @[PMP.scala 62:29]
  wire [31:0] _T_1214 = _T_1213 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_1215 = ~_T_1214; // @[PMP.scala 62:27]
  wire  _T_1217 = io_addr[31:3] < _T_1215[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_1224 = io_addr[31:3] ^ _T_1215[31:3]; // @[PMP.scala 83:41]
  wire  _T_1225 = _T_1224 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_1233 = _T_51 < _T_1215[2:0]; // @[PMP.scala 84:53]
  wire  _T_1235 = _T_1217 | _T_1225 & _T_1233; // @[PMP.scala 85:16]
  wire  _T_1236 = ~_T_1235; // @[PMP.scala 90:5]
  wire  _T_1259 = io_addr[2:0] < _T_1019[2:0]; // @[PMP.scala 84:53]
  wire  _T_1261 = _T_1021 | _T_1029 & _T_1259; // @[PMP.scala 85:16]
  wire  _T_1262 = _T_1236 & _T_1261; // @[PMP.scala 96:48]
  wire  _T_1264 = io_pmp_1_cfg_a[1] ? _T_1205 : io_pmp_1_cfg_a[0] & _T_1262; // @[PMP.scala 134:8]
  wire  _T_1266 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1286 = _T_1215[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_1288 = _T_1225 & _T_1286 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_1304 = _T_1019[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1306 = _T_1029 & _T_1304 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1308 = ~(_T_1288 | _T_1306); // @[PMP.scala 127:24]
  wire [2:0] _T_1310 = ~io_pmp_1_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1311 = _T_5 & _T_1310; // @[PMP.scala 128:32]
  wire  _T_1312 = _T_1311 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1314 = io_pmp_1_cfg_a[1] ? _T_1312 : _T_1308; // @[PMP.scala 129:8]
  wire  _T_1367 = _T_1314 & (io_pmp_1_cfg_r | _T_1266); // @[PMP.scala 183:26]
  wire  _T_1369 = _T_1314 & (io_pmp_1_cfg_w | _T_1266); // @[PMP.scala 184:26]
  wire  _T_1371 = _T_1314 & (io_pmp_1_cfg_x | _T_1266); // @[PMP.scala 185:26]
  wire  _T_1372_cfg_x = _T_1264 ? _T_1371 : _T_1176_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_w = _T_1264 ? _T_1369 : _T_1176_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_r = _T_1264 ? _T_1367 : _T_1176_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1378 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_1387 = ~io_pmp_0_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_1388 = _T_1224 & _T_1387; // @[PMP.scala 65:52]
  wire  _T_1389 = _T_1388 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1397 = io_addr[2:0] ^ _T_1215[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1398 = ~_T_1378[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1399 = _T_1397 & _T_1398; // @[PMP.scala 65:52]
  wire  _T_1400 = _T_1399 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1401 = _T_1389 & _T_1400; // @[PMP.scala 73:16]
  wire  _T_1455 = io_addr[2:0] < _T_1215[2:0]; // @[PMP.scala 84:53]
  wire  _T_1457 = _T_1217 | _T_1225 & _T_1455; // @[PMP.scala 85:16]
  wire  _T_1460 = io_pmp_0_cfg_a[1] ? _T_1401 : io_pmp_0_cfg_a[0] & _T_1457; // @[PMP.scala 134:8]
  wire  _T_1462 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1500 = _T_1215[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1502 = _T_1225 & _T_1500 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1504 = ~_T_1502; // @[PMP.scala 127:24]
  wire [2:0] _T_1506 = ~io_pmp_0_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1507 = _T_5 & _T_1506; // @[PMP.scala 128:32]
  wire  _T_1508 = _T_1507 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1510 = io_pmp_0_cfg_a[1] ? _T_1508 : _T_1504; // @[PMP.scala 129:8]
  wire  _T_1563 = _T_1510 & (io_pmp_0_cfg_r | _T_1462); // @[PMP.scala 183:26]
  wire  _T_1565 = _T_1510 & (io_pmp_0_cfg_w | _T_1462); // @[PMP.scala 184:26]
  wire  _T_1567 = _T_1510 & (io_pmp_0_cfg_x | _T_1462); // @[PMP.scala 185:26]
  assign io_r = _T_1460 ? _T_1563 : _T_1372_cfg_r; // @[PMP.scala 186:8]
  assign io_w = _T_1460 ? _T_1565 : _T_1372_cfg_w; // @[PMP.scala 186:8]
  assign io_x = _T_1460 ? _T_1567 : _T_1372_cfg_x; // @[PMP.scala 186:8]
endmodule
module NBDTLB(
  input         clock,
  input         reset,
  output        io_req_0_ready,
  input         io_req_0_valid,
  input  [39:0] io_req_0_bits_vaddr,
  input         io_req_0_bits_passthrough,
  input  [1:0]  io_req_0_bits_size,
  input  [4:0]  io_req_0_bits_cmd,
  output        io_miss_rdy,
  output        io_resp_0_miss,
  output [31:0] io_resp_0_paddr,
  output        io_resp_0_pf_ld,
  output        io_resp_0_pf_st,
  output        io_resp_0_pf_inst,
  output        io_resp_0_ae_ld,
  output        io_resp_0_ae_st,
  output        io_resp_0_ae_inst,
  output        io_resp_0_ma_ld,
  output        io_resp_0_ma_st,
  output        io_resp_0_ma_inst,
  output        io_resp_0_cacheable,
  output        io_resp_0_must_alloc,
  output        io_resp_0_prefetchable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_sfence_bits_asid,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0]  io_ptw_resp_bits_pte_reserved_for_software,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_fragmented_superpage,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [15:0] io_ptw_ptbr_asid,
  input  [43:0] io_ptw_ptbr_ppn,
  input         io_ptw_status_debug,
  input         io_ptw_status_cease,
  input         io_ptw_status_wfi,
  input  [31:0] io_ptw_status_isa,
  input  [1:0]  io_ptw_status_dprv,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_status_sd,
  input  [26:0] io_ptw_status_zero2,
  input  [1:0]  io_ptw_status_sxl,
  input  [1:0]  io_ptw_status_uxl,
  input         io_ptw_status_sd_rv32,
  input  [7:0]  io_ptw_status_zero1,
  input         io_ptw_status_tsr,
  input         io_ptw_status_tw,
  input         io_ptw_status_tvm,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_status_mprv,
  input  [1:0]  io_ptw_status_xs,
  input  [1:0]  io_ptw_status_fs,
  input  [1:0]  io_ptw_status_mpp,
  input  [1:0]  io_ptw_status_vs,
  input         io_ptw_status_spp,
  input         io_ptw_status_mpie,
  input         io_ptw_status_hpie,
  input         io_ptw_status_spie,
  input         io_ptw_status_upie,
  input         io_ptw_status_mie,
  input         io_ptw_status_hie,
  input         io_ptw_status_sie,
  input         io_ptw_status_uie,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_res,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_res,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_res,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_res,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_res,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_res,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_res,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_res,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_ptw_customCSRs_csrs_0_wen,
  input  [63:0] io_ptw_customCSRs_csrs_0_wdata,
  input  [63:0] io_ptw_customCSRs_csrs_0_value,
  input         io_kill
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  wire [19:0] package_Anon_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_io_y_c; // @[package.scala 213:21]
  wire [1:0] pmp_0_io_prv; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_0_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_0_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_0_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_0_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_0_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_0_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_0_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_1_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_1_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_1_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_1_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_1_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_1_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_1_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_2_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_2_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_2_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_2_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_2_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_2_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_2_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_3_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_3_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_3_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_3_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_3_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_3_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_3_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_4_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_4_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_4_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_4_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_4_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_4_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_4_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_5_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_5_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_5_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_5_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_5_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_5_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_5_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_6_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_6_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_6_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_6_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_6_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_6_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_6_mask; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_7_cfg_l; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_pmp_7_cfg_a; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_7_cfg_x; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_7_cfg_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_pmp_7_cfg_r; // @[tlb.scala 150:40]
  wire [29:0] pmp_0_io_pmp_7_addr; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_pmp_7_mask; // @[tlb.scala 150:40]
  wire [31:0] pmp_0_io_addr; // @[tlb.scala 150:40]
  wire [1:0] pmp_0_io_size; // @[tlb.scala 150:40]
  wire  pmp_0_io_r; // @[tlb.scala 150:40]
  wire  pmp_0_io_w; // @[tlb.scala 150:40]
  wire  pmp_0_io_x; // @[tlb.scala 150:40]
  wire [19:0] package_Anon_1_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_1_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_1_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_1_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_2_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_2_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_2_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_2_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_3_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_3_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_3_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_3_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_4_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_4_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_4_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_4_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_5_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_5_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_5_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_5_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_6_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_6_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_6_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_6_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_7_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_7_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_7_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_7_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_8_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_8_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_8_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_8_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_9_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_9_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_9_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_9_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_10_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_10_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_10_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_10_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_11_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_11_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_11_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_11_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_12_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_12_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_12_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_12_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_13_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_13_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_13_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_13_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_14_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_14_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_14_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_14_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_15_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_15_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_15_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_15_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_16_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_16_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_16_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_16_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_17_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_17_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_17_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_17_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_18_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_18_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_18_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_18_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_19_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_19_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_19_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_19_io_y_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_20_io_x_ppn; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_u; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_ae; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_sw; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_sx; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_sr; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_pw; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_px; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_pr; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_pal; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_paa; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_eff; // @[package.scala 213:21]
  wire  package_Anon_20_io_x_c; // @[package.scala 213:21]
  wire [19:0] package_Anon_20_io_y_ppn; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_u; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_ae; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_sw; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_sx; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_sr; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_pw; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_px; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_pr; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_pal; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_paa; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_eff; // @[package.scala 213:21]
  wire  package_Anon_20_io_y_c; // @[package.scala 213:21]
  reg [26:0] sectored_entries_0_tag; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_0_data_0; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_0_data_1; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_0_data_2; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_0_data_3; // @[tlb.scala 122:29]
  reg  sectored_entries_0_valid_0; // @[tlb.scala 122:29]
  reg  sectored_entries_0_valid_1; // @[tlb.scala 122:29]
  reg  sectored_entries_0_valid_2; // @[tlb.scala 122:29]
  reg  sectored_entries_0_valid_3; // @[tlb.scala 122:29]
  reg [26:0] sectored_entries_1_tag; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_1_data_0; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_1_data_1; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_1_data_2; // @[tlb.scala 122:29]
  reg [33:0] sectored_entries_1_data_3; // @[tlb.scala 122:29]
  reg  sectored_entries_1_valid_0; // @[tlb.scala 122:29]
  reg  sectored_entries_1_valid_1; // @[tlb.scala 122:29]
  reg  sectored_entries_1_valid_2; // @[tlb.scala 122:29]
  reg  sectored_entries_1_valid_3; // @[tlb.scala 122:29]
  reg [1:0] superpage_entries_0_level; // @[tlb.scala 123:30]
  reg [26:0] superpage_entries_0_tag; // @[tlb.scala 123:30]
  reg [33:0] superpage_entries_0_data_0; // @[tlb.scala 123:30]
  reg  superpage_entries_0_valid_0; // @[tlb.scala 123:30]
  reg [1:0] superpage_entries_1_level; // @[tlb.scala 123:30]
  reg [26:0] superpage_entries_1_tag; // @[tlb.scala 123:30]
  reg [33:0] superpage_entries_1_data_0; // @[tlb.scala 123:30]
  reg  superpage_entries_1_valid_0; // @[tlb.scala 123:30]
  reg [1:0] superpage_entries_2_level; // @[tlb.scala 123:30]
  reg [26:0] superpage_entries_2_tag; // @[tlb.scala 123:30]
  reg [33:0] superpage_entries_2_data_0; // @[tlb.scala 123:30]
  reg  superpage_entries_2_valid_0; // @[tlb.scala 123:30]
  reg [1:0] superpage_entries_3_level; // @[tlb.scala 123:30]
  reg [26:0] superpage_entries_3_tag; // @[tlb.scala 123:30]
  reg [33:0] superpage_entries_3_data_0; // @[tlb.scala 123:30]
  reg  superpage_entries_3_valid_0; // @[tlb.scala 123:30]
  reg [1:0] special_entry_level; // @[tlb.scala 124:56]
  reg [26:0] special_entry_tag; // @[tlb.scala 124:56]
  reg [33:0] special_entry_data_0; // @[tlb.scala 124:56]
  reg  special_entry_valid_0; // @[tlb.scala 124:56]
  reg [1:0] state; // @[tlb.scala 129:22]
  reg [26:0] r_refill_tag; // @[tlb.scala 130:25]
  reg [1:0] r_superpage_repl_addr; // @[tlb.scala 131:34]
  reg  r_sectored_repl_addr; // @[tlb.scala 132:33]
  reg  r_sectored_hit_addr; // @[tlb.scala 133:32]
  reg  r_sectored_hit; // @[tlb.scala 134:27]
  wire  priv_s = io_ptw_status_dprv[0]; // @[tlb.scala 137:20]
  wire  priv_uses_vm = io_ptw_status_dprv <= 2'h1; // @[tlb.scala 138:27]
  wire  vm_enabled_0 = io_ptw_ptbr_mode[3] & priv_uses_vm & ~io_req_0_bits_passthrough; // @[tlb.scala 139:109]
  wire [26:0] vpn_0 = io_req_0_bits_vaddr[38:12]; // @[tlb.scala 142:47]
  wire [19:0] refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[tlb.scala 143:44]
  wire  _T_6 = state == 2'h1; // @[package.scala 15:47]
  wire  _T_7 = state == 2'h3; // @[package.scala 15:47]
  wire  invalidate_refill = _T_6 | _T_7; // @[package.scala 64:59]
  wire  _T_27 = special_entry_level < 2'h1; // @[tlb.scala 80:31]
  wire [26:0] _T_29 = _T_27 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _GEN_326 = {{7'd0}, package_Anon_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_30 = _T_29 | _GEN_326; // @[tlb.scala 81:49]
  wire  _T_33 = special_entry_level < 2'h2; // @[tlb.scala 80:31]
  wire [26:0] _T_35 = _T_33 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _T_36 = _T_35 | _GEN_326; // @[tlb.scala 81:49]
  wire [19:0] _T_38 = {package_Anon_io_y_ppn[19:18],_T_30[17:9],_T_36[8:0]}; // @[Cat.scala 29:58]
  wire [27:0] _T_40 = vm_enabled_0 ? {{8'd0}, _T_38} : io_req_0_bits_vaddr[39:12]; // @[tlb.scala 148:20]
  wire [27:0] mpu_ppn_0 = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_40; // @[tlb.scala 147:20]
  wire [39:0] mpu_physaddr_0 = {mpu_ppn_0,io_req_0_bits_vaddr[11:0]}; // @[Cat.scala 29:58]
  wire [39:0] _T_47 = mpu_physaddr_0 ^ 40'h3000; // @[Parameters.scala 137:31]
  wire [40:0] _T_48 = {1'b0,$signed(_T_47)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_50 = $signed(_T_48) & -41'sh1000; // @[Parameters.scala 137:52]
  wire  _T_51 = $signed(_T_50) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_52 = mpu_physaddr_0 ^ 40'h2010000; // @[Parameters.scala 137:31]
  wire [40:0] _T_53 = {1'b0,$signed(_T_52)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_55 = $signed(_T_53) & -41'sh1000; // @[Parameters.scala 137:52]
  wire  _T_56 = $signed(_T_55) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_57 = mpu_physaddr_0 ^ 40'h54000000; // @[Parameters.scala 137:31]
  wire [40:0] _T_58 = {1'b0,$signed(_T_57)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_60 = $signed(_T_58) & -41'sh1000; // @[Parameters.scala 137:52]
  wire  _T_61 = $signed(_T_60) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_62 = mpu_physaddr_0 ^ 40'hc000000; // @[Parameters.scala 137:31]
  wire [40:0] _T_63 = {1'b0,$signed(_T_62)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_65 = $signed(_T_63) & -41'sh4000000; // @[Parameters.scala 137:52]
  wire  _T_66 = $signed(_T_65) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_67 = mpu_physaddr_0 ^ 40'h2000000; // @[Parameters.scala 137:31]
  wire [40:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_70 = $signed(_T_68) & -41'sh10000; // @[Parameters.scala 137:52]
  wire  _T_71 = $signed(_T_70) == 41'sh0; // @[Parameters.scala 137:67]
  wire [40:0] _T_73 = {1'b0,$signed(mpu_physaddr_0)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_75 = $signed(_T_73) & -41'sh1000; // @[Parameters.scala 137:52]
  wire  _T_76 = $signed(_T_75) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_77 = mpu_physaddr_0 ^ 40'h10000; // @[Parameters.scala 137:31]
  wire [40:0] _T_78 = {1'b0,$signed(_T_77)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_80 = $signed(_T_78) & -41'sh10000; // @[Parameters.scala 137:52]
  wire  _T_81 = $signed(_T_80) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_82 = mpu_physaddr_0 ^ 40'h80000000; // @[Parameters.scala 137:31]
  wire [40:0] _T_83 = {1'b0,$signed(_T_82)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_85 = $signed(_T_83) & -41'sh10000000; // @[Parameters.scala 137:52]
  wire  _T_86 = $signed(_T_85) == 41'sh0; // @[Parameters.scala 137:67]
  wire  _T_91 = _T_51 | _T_56 | _T_61 | _T_66 | _T_71; // @[tlb.scala 157:84]
  wire  legal_address_0 = _T_51 | _T_56 | _T_61 | _T_66 | _T_71 | _T_76 | _T_81 | _T_86; // @[tlb.scala 157:84]
  wire [40:0] _T_103 = $signed(_T_83) & 41'sh80000000; // @[Parameters.scala 137:52]
  wire  _T_104 = $signed(_T_103) == 41'sh0; // @[Parameters.scala 137:67]
  wire  cacheable_0 = legal_address_0 & _T_104; // @[tlb.scala 159:22]
  wire  homogeneous_0 = _T_91 | _T_86 | _T_81 | _T_76; // @[TLBPermissions.scala 98:65]
  wire [40:0] _T_170 = $signed(_T_73) & 41'sh86000000; // @[Parameters.scala 137:52]
  wire  _T_171 = $signed(_T_170) == 41'sh0; // @[Parameters.scala 137:67]
  wire  _T_178 = _T_171 | _T_104; // @[TLBPermissions.scala 82:66]
  wire  prot_r_0 = legal_address_0 & pmp_0_io_r; // @[tlb.scala 162:60]
  wire [40:0] _T_209 = $signed(_T_73) & 41'sh82010000; // @[Parameters.scala 137:52]
  wire  _T_210 = $signed(_T_209) == 41'sh0; // @[Parameters.scala 137:67]
  wire [40:0] _T_214 = $signed(_T_68) & 41'sh86000000; // @[Parameters.scala 137:52]
  wire  _T_215 = $signed(_T_214) == 41'sh0; // @[Parameters.scala 137:67]
  wire [39:0] _T_216 = mpu_physaddr_0 ^ 40'h4000000; // @[Parameters.scala 137:31]
  wire [40:0] _T_217 = {1'b0,$signed(_T_216)}; // @[Parameters.scala 137:49]
  wire [40:0] _T_219 = $signed(_T_217) & 41'sh84000000; // @[Parameters.scala 137:52]
  wire  _T_220 = $signed(_T_219) == 41'sh0; // @[Parameters.scala 137:67]
  wire  _T_228 = _T_210 | _T_215 | _T_220 | _T_104; // @[Parameters.scala 528:89]
  wire  _T_238 = legal_address_0 & _T_228; // @[tlb.scala 159:22]
  wire  prot_w_0 = _T_238 & pmp_0_io_w; // @[tlb.scala 163:64]
  wire  _T_338 = legal_address_0 & _T_178; // @[tlb.scala 159:22]
  wire  prot_x_0 = _T_338 & pmp_0_io_x; // @[tlb.scala 166:59]
  wire [40:0] _T_360 = $signed(_T_53) & 41'sh86012000; // @[Parameters.scala 137:52]
  wire  _T_361 = $signed(_T_360) == 41'sh0; // @[Parameters.scala 137:67]
  wire [40:0] _T_365 = $signed(_T_73) & 41'sh82012000; // @[Parameters.scala 137:52]
  wire  _T_366 = $signed(_T_365) == 41'sh0; // @[Parameters.scala 137:67]
  wire [40:0] _T_375 = $signed(_T_68) & 41'sh86010000; // @[Parameters.scala 137:52]
  wire  _T_376 = $signed(_T_375) == 41'sh0; // @[Parameters.scala 137:67]
  wire  _T_379 = _T_361 | _T_366 | _T_220 | _T_376; // @[Parameters.scala 528:89]
  wire  prot_eff_0 = legal_address_0 & _T_379; // @[tlb.scala 159:22]
  wire  _T_387 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1 | sectored_entries_0_valid_2 |
    sectored_entries_0_valid_3; // @[package.scala 64:59]
  wire [26:0] _T_388 = sectored_entries_0_tag ^ vpn_0; // @[tlb.scala 60:43]
  wire  _T_390 = _T_388[26:2] == 25'h0; // @[tlb.scala 60:73]
  wire  sector_hits_0_0 = _T_387 & _T_390; // @[tlb.scala 59:42]
  wire  _T_394 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1 | sectored_entries_1_valid_2 |
    sectored_entries_1_valid_3; // @[package.scala 64:59]
  wire [26:0] _T_395 = sectored_entries_1_tag ^ vpn_0; // @[tlb.scala 60:43]
  wire  _T_397 = _T_395[26:2] == 25'h0; // @[tlb.scala 60:73]
  wire  sector_hits_0_1 = _T_394 & _T_397; // @[tlb.scala 59:42]
  wire  _T_407 = superpage_entries_0_level < 2'h1; // @[tlb.scala 66:30]
  wire  superpage_hits_0_0 = superpage_entries_0_valid_0 & superpage_entries_0_tag[26:18] == vpn_0[26:18] & (_T_407 |
    superpage_entries_0_tag[17:9] == vpn_0[17:9]); // @[tlb.scala 67:31]
  wire  _T_428 = superpage_entries_1_level < 2'h1; // @[tlb.scala 66:30]
  wire  superpage_hits_0_1 = superpage_entries_1_valid_0 & superpage_entries_1_tag[26:18] == vpn_0[26:18] & (_T_428 |
    superpage_entries_1_tag[17:9] == vpn_0[17:9]); // @[tlb.scala 67:31]
  wire  _T_449 = superpage_entries_2_level < 2'h1; // @[tlb.scala 66:30]
  wire  superpage_hits_0_2 = superpage_entries_2_valid_0 & superpage_entries_2_tag[26:18] == vpn_0[26:18] & (_T_449 |
    superpage_entries_2_tag[17:9] == vpn_0[17:9]); // @[tlb.scala 67:31]
  wire  _T_470 = superpage_entries_3_level < 2'h1; // @[tlb.scala 66:30]
  wire  superpage_hits_0_3 = superpage_entries_3_valid_0 & superpage_entries_3_tag[26:18] == vpn_0[26:18] & (_T_470 |
    superpage_entries_3_tag[17:9] == vpn_0[17:9]); // @[tlb.scala 67:31]
  wire  _GEN_1 = 2'h1 == vpn_0[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[tlb.scala 72:{20,20}]
  wire  _GEN_2 = 2'h2 == vpn_0[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[tlb.scala 72:{20,20}]
  wire  _GEN_3 = 2'h3 == vpn_0[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[tlb.scala 72:{20,20}]
  wire  _T_489 = _GEN_3 & _T_390; // @[tlb.scala 72:20]
  wire  hitsVec_0_0 = vm_enabled_0 & _T_489; // @[tlb.scala 171:69]
  wire  _GEN_5 = 2'h1 == vpn_0[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[tlb.scala 72:{20,20}]
  wire  _GEN_6 = 2'h2 == vpn_0[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[tlb.scala 72:{20,20}]
  wire  _GEN_7 = 2'h3 == vpn_0[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[tlb.scala 72:{20,20}]
  wire  _T_495 = _GEN_7 & _T_397; // @[tlb.scala 72:20]
  wire  hitsVec_0_1 = vm_enabled_0 & _T_495; // @[tlb.scala 171:69]
  wire  hitsVec_0_2 = vm_enabled_0 & superpage_hits_0_0; // @[tlb.scala 171:69]
  wire  hitsVec_0_3 = vm_enabled_0 & superpage_hits_0_1; // @[tlb.scala 171:69]
  wire  hitsVec_0_4 = vm_enabled_0 & superpage_hits_0_2; // @[tlb.scala 171:69]
  wire  hitsVec_0_5 = vm_enabled_0 & superpage_hits_0_3; // @[tlb.scala 171:69]
  wire  _T_605 = special_entry_valid_0 & special_entry_tag[26:18] == vpn_0[26:18] & (_T_27 | special_entry_tag[17:9] ==
    vpn_0[17:9]) & (_T_33 | special_entry_tag[8:0] == vpn_0[8:0]); // @[tlb.scala 67:31]
  wire  hitsVec_0_6 = vm_enabled_0 & _T_605; // @[tlb.scala 171:69]
  wire [6:0] real_hits_0 = {hitsVec_0_6,hitsVec_0_5,hitsVec_0_4,hitsVec_0_3,hitsVec_0_2,hitsVec_0_1,hitsVec_0_0}; // @[tlb.scala 172:44]
  wire  _T_614 = ~vm_enabled_0; // @[tlb.scala 173:32]
  wire [7:0] hits_0 = {_T_614,hitsVec_0_6,hitsVec_0_5,hitsVec_0_4,hitsVec_0_3,hitsVec_0_2,hitsVec_0_1,hitsVec_0_0}; // @[Cat.scala 29:58]
  wire [33:0] _GEN_9 = 2'h1 == vpn_0[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[]
  wire [33:0] _GEN_10 = 2'h2 == vpn_0[1:0] ? sectored_entries_0_data_2 : _GEN_9; // @[]
  wire [33:0] _GEN_11 = 2'h3 == vpn_0[1:0] ? sectored_entries_0_data_3 : _GEN_10; // @[]
  wire [33:0] _GEN_13 = 2'h1 == vpn_0[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[]
  wire [33:0] _GEN_14 = 2'h2 == vpn_0[1:0] ? sectored_entries_1_data_2 : _GEN_13; // @[]
  wire [33:0] _GEN_15 = 2'h3 == vpn_0[1:0] ? sectored_entries_1_data_3 : _GEN_14; // @[]
  wire [26:0] _T_673 = _T_407 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _GEN_328 = {{7'd0}, package_Anon_3_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_674 = _T_673 | _GEN_328; // @[tlb.scala 81:49]
  wire [26:0] _T_680 = vpn_0 | _GEN_328; // @[tlb.scala 81:49]
  wire [19:0] _T_682 = {package_Anon_3_io_y_ppn[19:18],_T_674[17:9],_T_680[8:0]}; // @[Cat.scala 29:58]
  wire [26:0] _T_703 = _T_428 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _GEN_330 = {{7'd0}, package_Anon_4_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_704 = _T_703 | _GEN_330; // @[tlb.scala 81:49]
  wire [26:0] _T_710 = vpn_0 | _GEN_330; // @[tlb.scala 81:49]
  wire [19:0] _T_712 = {package_Anon_4_io_y_ppn[19:18],_T_704[17:9],_T_710[8:0]}; // @[Cat.scala 29:58]
  wire [26:0] _T_733 = _T_449 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _GEN_332 = {{7'd0}, package_Anon_5_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_734 = _T_733 | _GEN_332; // @[tlb.scala 81:49]
  wire [26:0] _T_740 = vpn_0 | _GEN_332; // @[tlb.scala 81:49]
  wire [19:0] _T_742 = {package_Anon_5_io_y_ppn[19:18],_T_734[17:9],_T_740[8:0]}; // @[Cat.scala 29:58]
  wire [26:0] _T_763 = _T_470 ? vpn_0 : 27'h0; // @[tlb.scala 81:30]
  wire [26:0] _GEN_334 = {{7'd0}, package_Anon_6_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_764 = _T_763 | _GEN_334; // @[tlb.scala 81:49]
  wire [26:0] _T_770 = vpn_0 | _GEN_334; // @[tlb.scala 81:49]
  wire [19:0] _T_772 = {package_Anon_6_io_y_ppn[19:18],_T_764[17:9],_T_770[8:0]}; // @[Cat.scala 29:58]
  wire [26:0] _GEN_336 = {{7'd0}, package_Anon_7_io_y_ppn}; // @[tlb.scala 81:49]
  wire [26:0] _T_794 = _T_29 | _GEN_336; // @[tlb.scala 81:49]
  wire [26:0] _T_800 = _T_35 | _GEN_336; // @[tlb.scala 81:49]
  wire [19:0] _T_802 = {package_Anon_7_io_y_ppn[19:18],_T_794[17:9],_T_800[8:0]}; // @[Cat.scala 29:58]
  wire [19:0] _T_804 = hitsVec_0_0 ? package_Anon_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_805 = hitsVec_0_1 ? package_Anon_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_806 = hitsVec_0_2 ? _T_682 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_807 = hitsVec_0_3 ? _T_712 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_808 = hitsVec_0_4 ? _T_742 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_809 = hitsVec_0_5 ? _T_772 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_810 = hitsVec_0_6 ? _T_802 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_811 = _T_614 ? vpn_0[19:0] : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _T_812 = _T_804 | _T_805; // @[Mux.scala 27:72]
  wire [19:0] _T_813 = _T_812 | _T_806; // @[Mux.scala 27:72]
  wire [19:0] _T_814 = _T_813 | _T_807; // @[Mux.scala 27:72]
  wire [19:0] _T_815 = _T_814 | _T_808; // @[Mux.scala 27:72]
  wire [19:0] _T_816 = _T_815 | _T_809; // @[Mux.scala 27:72]
  wire [19:0] _T_817 = _T_816 | _T_810; // @[Mux.scala 27:72]
  wire [19:0] ppn_0 = _T_817 | _T_811; // @[Mux.scala 27:72]
  wire  _T_827 = io_ptw_resp_bits_pte_v & (io_ptw_resp_bits_pte_r | io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w) &
    io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52]
  wire  _T_828 = _T_827 & io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35]
  wire  _T_835 = _T_827 & io_ptw_resp_bits_pte_w & io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40]
  wire  _T_841 = _T_827 & io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35]
  wire [6:0] _T_850 = {prot_x_0,prot_r_0,_T_238,_T_238,prot_eff_0,cacheable_0,io_ptw_resp_bits_fragmented_superpage}; // @[tlb.scala 95:26]
  wire [33:0] _T_858 = {refill_ppn,io_ptw_resp_bits_pte_u,io_ptw_resp_bits_pte_g,io_ptw_resp_bits_ae,_T_835,_T_841,
    _T_828,prot_w_0,_T_850}; // @[tlb.scala 95:26]
  wire  _GEN_18 = r_superpage_repl_addr == 2'h0 | superpage_entries_0_valid_0; // @[tlb.scala 199:91 94:18 123:30]
  wire  _GEN_22 = r_superpage_repl_addr == 2'h1 | superpage_entries_1_valid_0; // @[tlb.scala 199:91 94:18 123:30]
  wire  _GEN_26 = r_superpage_repl_addr == 2'h2 | superpage_entries_2_valid_0; // @[tlb.scala 199:91 94:18 123:30]
  wire  _GEN_30 = r_superpage_repl_addr == 2'h3 | superpage_entries_3_valid_0; // @[tlb.scala 199:91 94:18 123:30]
  wire  _T_924 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[tlb.scala 203:22]
  wire  _GEN_32 = ~r_sectored_hit ? 1'h0 : sectored_entries_0_valid_0; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_33 = ~r_sectored_hit ? 1'h0 : sectored_entries_0_valid_1; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_34 = ~r_sectored_hit ? 1'h0 : sectored_entries_0_valid_2; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_35 = ~r_sectored_hit ? 1'h0 : sectored_entries_0_valid_3; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_36 = 2'h0 == r_refill_tag[1:0] | _GEN_32; // @[tlb.scala 94:{18,18}]
  wire  _GEN_37 = 2'h1 == r_refill_tag[1:0] | _GEN_33; // @[tlb.scala 94:{18,18}]
  wire  _GEN_38 = 2'h2 == r_refill_tag[1:0] | _GEN_34; // @[tlb.scala 94:{18,18}]
  wire  _GEN_39 = 2'h3 == r_refill_tag[1:0] | _GEN_35; // @[tlb.scala 94:{18,18}]
  wire [33:0] _GEN_40 = 2'h0 == r_refill_tag[1:0] ? _T_858 : sectored_entries_0_data_0; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_41 = 2'h1 == r_refill_tag[1:0] ? _T_858 : sectored_entries_0_data_1; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_42 = 2'h2 == r_refill_tag[1:0] ? _T_858 : sectored_entries_0_data_2; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_43 = 2'h3 == r_refill_tag[1:0] ? _T_858 : sectored_entries_0_data_3; // @[tlb.scala 95:{17,17} 122:29]
  wire  _GEN_44 = ~_T_924 ? _GEN_36 : sectored_entries_0_valid_0; // @[tlb.scala 122:29 204:74]
  wire  _GEN_45 = ~_T_924 ? _GEN_37 : sectored_entries_0_valid_1; // @[tlb.scala 122:29 204:74]
  wire  _GEN_46 = ~_T_924 ? _GEN_38 : sectored_entries_0_valid_2; // @[tlb.scala 122:29 204:74]
  wire  _GEN_47 = ~_T_924 ? _GEN_39 : sectored_entries_0_valid_3; // @[tlb.scala 122:29 204:74]
  wire  _GEN_54 = ~r_sectored_hit ? 1'h0 : sectored_entries_1_valid_0; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_55 = ~r_sectored_hit ? 1'h0 : sectored_entries_1_valid_1; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_56 = ~r_sectored_hit ? 1'h0 : sectored_entries_1_valid_2; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_57 = ~r_sectored_hit ? 1'h0 : sectored_entries_1_valid_3; // @[tlb.scala 122:29 205:32 98:40]
  wire  _GEN_58 = 2'h0 == r_refill_tag[1:0] | _GEN_54; // @[tlb.scala 94:{18,18}]
  wire  _GEN_59 = 2'h1 == r_refill_tag[1:0] | _GEN_55; // @[tlb.scala 94:{18,18}]
  wire  _GEN_60 = 2'h2 == r_refill_tag[1:0] | _GEN_56; // @[tlb.scala 94:{18,18}]
  wire  _GEN_61 = 2'h3 == r_refill_tag[1:0] | _GEN_57; // @[tlb.scala 94:{18,18}]
  wire [33:0] _GEN_62 = 2'h0 == r_refill_tag[1:0] ? _T_858 : sectored_entries_1_data_0; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_63 = 2'h1 == r_refill_tag[1:0] ? _T_858 : sectored_entries_1_data_1; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_64 = 2'h2 == r_refill_tag[1:0] ? _T_858 : sectored_entries_1_data_2; // @[tlb.scala 95:{17,17} 122:29]
  wire [33:0] _GEN_65 = 2'h3 == r_refill_tag[1:0] ? _T_858 : sectored_entries_1_data_3; // @[tlb.scala 95:{17,17} 122:29]
  wire  _GEN_66 = _T_924 ? _GEN_58 : sectored_entries_1_valid_0; // @[tlb.scala 122:29 204:74]
  wire  _GEN_67 = _T_924 ? _GEN_59 : sectored_entries_1_valid_1; // @[tlb.scala 122:29 204:74]
  wire  _GEN_68 = _T_924 ? _GEN_60 : sectored_entries_1_valid_2; // @[tlb.scala 122:29 204:74]
  wire  _GEN_69 = _T_924 ? _GEN_61 : sectored_entries_1_valid_3; // @[tlb.scala 122:29 204:74]
  wire  _GEN_78 = io_ptw_resp_bits_level < 2'h2 ? _GEN_18 : superpage_entries_0_valid_0; // @[tlb.scala 123:30 198:58]
  wire  _GEN_82 = io_ptw_resp_bits_level < 2'h2 ? _GEN_22 : superpage_entries_1_valid_0; // @[tlb.scala 123:30 198:58]
  wire  _GEN_86 = io_ptw_resp_bits_level < 2'h2 ? _GEN_26 : superpage_entries_2_valid_0; // @[tlb.scala 123:30 198:58]
  wire  _GEN_90 = io_ptw_resp_bits_level < 2'h2 ? _GEN_30 : superpage_entries_3_valid_0; // @[tlb.scala 123:30 198:58]
  wire  _GEN_92 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_valid_0 : _GEN_44; // @[tlb.scala 122:29 198:58]
  wire  _GEN_93 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_valid_1 : _GEN_45; // @[tlb.scala 122:29 198:58]
  wire  _GEN_94 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_valid_2 : _GEN_46; // @[tlb.scala 122:29 198:58]
  wire  _GEN_95 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_valid_3 : _GEN_47; // @[tlb.scala 122:29 198:58]
  wire  _GEN_102 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_1_valid_0 : _GEN_66; // @[tlb.scala 122:29 198:58]
  wire  _GEN_103 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_1_valid_1 : _GEN_67; // @[tlb.scala 122:29 198:58]
  wire  _GEN_104 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_1_valid_2 : _GEN_68; // @[tlb.scala 122:29 198:58]
  wire  _GEN_105 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_1_valid_3 : _GEN_69; // @[tlb.scala 122:29 198:58]
  wire  _GEN_114 = ~io_ptw_resp_bits_homogeneous | special_entry_valid_0; // @[tlb.scala 196:70 94:18 124:56]
  wire  _GEN_118 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_0_valid_0 : _GEN_78; // @[tlb.scala 123:30 196:70]
  wire  _GEN_122 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_1_valid_0 : _GEN_82; // @[tlb.scala 123:30 196:70]
  wire  _GEN_126 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_2_valid_0 : _GEN_86; // @[tlb.scala 123:30 196:70]
  wire  _GEN_130 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_3_valid_0 : _GEN_90; // @[tlb.scala 123:30 196:70]
  wire  _GEN_132 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_valid_0 : _GEN_92; // @[tlb.scala 122:29 196:70]
  wire  _GEN_133 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_valid_1 : _GEN_93; // @[tlb.scala 122:29 196:70]
  wire  _GEN_134 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_valid_2 : _GEN_94; // @[tlb.scala 122:29 196:70]
  wire  _GEN_135 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_valid_3 : _GEN_95; // @[tlb.scala 122:29 196:70]
  wire  _GEN_142 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_1_valid_0 : _GEN_102; // @[tlb.scala 122:29 196:70]
  wire  _GEN_143 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_1_valid_1 : _GEN_103; // @[tlb.scala 122:29 196:70]
  wire  _GEN_144 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_1_valid_2 : _GEN_104; // @[tlb.scala 122:29 196:70]
  wire  _GEN_145 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_1_valid_3 : _GEN_105; // @[tlb.scala 122:29 196:70]
  wire  _GEN_154 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_114 : special_entry_valid_0; // @[tlb.scala 177:42 124:56]
  wire  _GEN_158 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_118 : superpage_entries_0_valid_0; // @[tlb.scala 123:30 177:42]
  wire  _GEN_162 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_122 : superpage_entries_1_valid_0; // @[tlb.scala 123:30 177:42]
  wire  _GEN_166 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_126 : superpage_entries_2_valid_0; // @[tlb.scala 123:30 177:42]
  wire  _GEN_170 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_130 : superpage_entries_3_valid_0; // @[tlb.scala 123:30 177:42]
  wire  _GEN_172 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_132 : sectored_entries_0_valid_0; // @[tlb.scala 122:29 177:42]
  wire  _GEN_173 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_133 : sectored_entries_0_valid_1; // @[tlb.scala 122:29 177:42]
  wire  _GEN_174 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_134 : sectored_entries_0_valid_2; // @[tlb.scala 122:29 177:42]
  wire  _GEN_175 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_135 : sectored_entries_0_valid_3; // @[tlb.scala 122:29 177:42]
  wire  _GEN_182 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_142 : sectored_entries_1_valid_0; // @[tlb.scala 122:29 177:42]
  wire  _GEN_183 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_143 : sectored_entries_1_valid_1; // @[tlb.scala 122:29 177:42]
  wire  _GEN_184 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_144 : sectored_entries_1_valid_2; // @[tlb.scala 122:29 177:42]
  wire  _GEN_185 = io_ptw_resp_valid & ~invalidate_refill ? _GEN_145 : sectored_entries_1_valid_3; // @[tlb.scala 122:29 177:42]
  wire  entries_0_2_ae = package_Anon_10_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_1_ae = package_Anon_9_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_0_ae = package_Anon_8_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_4_ae = package_Anon_12_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_3_ae = package_Anon_11_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_6_ae = package_Anon_14_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire  entries_0_5_ae = package_Anon_13_io_y_ae; // @[tlb.scala 211:{38,38}]
  wire [7:0] ptw_ae_array_0 = {1'h0,entries_0_6_ae,entries_0_5_ae,entries_0_4_ae,entries_0_3_ae,entries_0_2_ae,
    entries_0_1_ae,entries_0_0_ae}; // @[Cat.scala 29:58]
  wire  entries_0_2_u = package_Anon_10_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_1_u = package_Anon_9_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_0_u = package_Anon_8_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_4_u = package_Anon_12_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_3_u = package_Anon_11_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_6_u = package_Anon_14_io_y_u; // @[tlb.scala 211:{38,38}]
  wire  entries_0_5_u = package_Anon_13_io_y_u; // @[tlb.scala 211:{38,38}]
  wire [6:0] _T_1200 = {entries_0_6_u,entries_0_5_u,entries_0_4_u,entries_0_3_u,entries_0_2_u,entries_0_1_u,
    entries_0_0_u}; // @[Cat.scala 29:58]
  wire [6:0] _T_1201 = ~priv_s | io_ptw_status_sum ? _T_1200 : 7'h0; // @[tlb.scala 215:39]
  wire [6:0] _T_1208 = ~_T_1200; // @[tlb.scala 215:117]
  wire [6:0] _T_1209 = priv_s ? _T_1208 : 7'h0; // @[tlb.scala 215:108]
  wire [6:0] priv_rw_ok_0 = _T_1201 | _T_1209; // @[tlb.scala 215:103]
  wire [6:0] priv_x_ok_0 = priv_s ? _T_1208 : _T_1200; // @[tlb.scala 216:39]
  wire  entries_0_2_sr = package_Anon_10_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_1_sr = package_Anon_9_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_0_sr = package_Anon_8_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_4_sr = package_Anon_12_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_3_sr = package_Anon_11_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_6_sr = package_Anon_14_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire  entries_0_5_sr = package_Anon_13_io_y_sr; // @[tlb.scala 211:{38,38}]
  wire [6:0] _T_1230 = {entries_0_6_sr,entries_0_5_sr,entries_0_4_sr,entries_0_3_sr,entries_0_2_sr,entries_0_1_sr,
    entries_0_0_sr}; // @[Cat.scala 29:58]
  wire  entries_0_2_sx = package_Anon_10_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_1_sx = package_Anon_9_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_0_sx = package_Anon_8_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_4_sx = package_Anon_12_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_3_sx = package_Anon_11_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_6_sx = package_Anon_14_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire  entries_0_5_sx = package_Anon_13_io_y_sx; // @[tlb.scala 211:{38,38}]
  wire [6:0] _T_1236 = {entries_0_6_sx,entries_0_5_sx,entries_0_4_sx,entries_0_3_sx,entries_0_2_sx,entries_0_1_sx,
    entries_0_0_sx}; // @[Cat.scala 29:58]
  wire [6:0] _T_1237 = io_ptw_status_mxr ? _T_1236 : 7'h0; // @[tlb.scala 217:98]
  wire [6:0] _T_1238 = _T_1230 | _T_1237; // @[tlb.scala 217:93]
  wire [6:0] _T_1239 = priv_rw_ok_0 & _T_1238; // @[tlb.scala 217:62]
  wire [7:0] r_array_0 = {1'h1,_T_1239}; // @[Cat.scala 29:58]
  wire  entries_0_2_sw = package_Anon_10_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_1_sw = package_Anon_9_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_0_sw = package_Anon_8_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_4_sw = package_Anon_12_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_3_sw = package_Anon_11_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_6_sw = package_Anon_14_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire  entries_0_5_sw = package_Anon_13_io_y_sw; // @[tlb.scala 211:{38,38}]
  wire [6:0] _T_1246 = {entries_0_6_sw,entries_0_5_sw,entries_0_4_sw,entries_0_3_sw,entries_0_2_sw,entries_0_1_sw,
    entries_0_0_sw}; // @[Cat.scala 29:58]
  wire [6:0] _T_1247 = priv_rw_ok_0 & _T_1246; // @[tlb.scala 218:62]
  wire [7:0] w_array_0 = {1'h1,_T_1247}; // @[Cat.scala 29:58]
  wire [6:0] _T_1255 = priv_x_ok_0 & _T_1236; // @[tlb.scala 219:62]
  wire [7:0] x_array_0 = {1'h1,_T_1255}; // @[Cat.scala 29:58]
  wire [1:0] _T_1258 = prot_r_0 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_pr = package_Anon_17_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_pr = package_Anon_16_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_pr = package_Anon_15_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_pr = package_Anon_20_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_pr = package_Anon_19_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_pr = package_Anon_18_io_y_pr; // @[tlb.scala 212:{45,45}]
  wire [7:0] _T_1264 = {_T_1258,normal_entries_0_5_pr,normal_entries_0_4_pr,normal_entries_0_3_pr,normal_entries_0_2_pr,
    normal_entries_0_1_pr,normal_entries_0_0_pr}; // @[Cat.scala 29:58]
  wire [7:0] _T_1265 = ~ptw_ae_array_0; // @[tlb.scala 220:116]
  wire [7:0] pr_array_0 = _T_1264 & _T_1265; // @[tlb.scala 220:114]
  wire [1:0] _T_1268 = prot_w_0 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_pw = package_Anon_17_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_pw = package_Anon_16_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_pw = package_Anon_15_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_pw = package_Anon_20_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_pw = package_Anon_19_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_pw = package_Anon_18_io_y_pw; // @[tlb.scala 212:{45,45}]
  wire [7:0] _T_1274 = {_T_1268,normal_entries_0_5_pw,normal_entries_0_4_pw,normal_entries_0_3_pw,normal_entries_0_2_pw,
    normal_entries_0_1_pw,normal_entries_0_0_pw}; // @[Cat.scala 29:58]
  wire [7:0] pw_array_0 = _T_1274 & _T_1265; // @[tlb.scala 221:114]
  wire [1:0] _T_1278 = prot_x_0 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_px = package_Anon_17_io_y_px; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_px = package_Anon_16_io_y_px; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_px = package_Anon_15_io_y_px; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_px = package_Anon_20_io_y_px; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_px = package_Anon_19_io_y_px; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_px = package_Anon_18_io_y_px; // @[tlb.scala 212:{45,45}]
  wire [7:0] _T_1284 = {_T_1278,normal_entries_0_5_px,normal_entries_0_4_px,normal_entries_0_3_px,normal_entries_0_2_px,
    normal_entries_0_1_px,normal_entries_0_0_px}; // @[Cat.scala 29:58]
  wire [7:0] px_array_0 = _T_1284 & _T_1265; // @[tlb.scala 222:114]
  wire [1:0] _T_1288 = prot_eff_0 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_eff = package_Anon_17_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_eff = package_Anon_16_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_eff = package_Anon_15_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_eff = package_Anon_20_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_eff = package_Anon_19_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_eff = package_Anon_18_io_y_eff; // @[tlb.scala 212:{45,45}]
  wire [7:0] eff_array_0 = {_T_1288,normal_entries_0_5_eff,normal_entries_0_4_eff,normal_entries_0_3_eff,
    normal_entries_0_2_eff,normal_entries_0_1_eff,normal_entries_0_0_eff}; // @[Cat.scala 29:58]
  wire [1:0] _T_1296 = cacheable_0 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_c = package_Anon_17_io_y_c; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_c = package_Anon_16_io_y_c; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_c = package_Anon_15_io_y_c; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_c = package_Anon_20_io_y_c; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_c = package_Anon_19_io_y_c; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_c = package_Anon_18_io_y_c; // @[tlb.scala 212:{45,45}]
  wire [7:0] c_array_0 = {_T_1296,normal_entries_0_5_c,normal_entries_0_4_c,normal_entries_0_3_c,normal_entries_0_2_c,
    normal_entries_0_1_c,normal_entries_0_0_c}; // @[Cat.scala 29:58]
  wire [1:0] _T_1304 = _T_238 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  normal_entries_0_2_paa = package_Anon_17_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_paa = package_Anon_16_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_paa = package_Anon_15_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_paa = package_Anon_20_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_paa = package_Anon_19_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_paa = package_Anon_18_io_y_paa; // @[tlb.scala 212:{45,45}]
  wire [7:0] paa_array_0 = {_T_1304,normal_entries_0_5_paa,normal_entries_0_4_paa,normal_entries_0_3_paa,
    normal_entries_0_2_paa,normal_entries_0_1_paa,normal_entries_0_0_paa}; // @[Cat.scala 29:58]
  wire  normal_entries_0_2_pal = package_Anon_17_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_1_pal = package_Anon_16_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_0_pal = package_Anon_15_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_5_pal = package_Anon_20_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_4_pal = package_Anon_19_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire  normal_entries_0_3_pal = package_Anon_18_io_y_pal; // @[tlb.scala 212:{45,45}]
  wire [7:0] pal_array_0 = {_T_1304,normal_entries_0_5_pal,normal_entries_0_4_pal,normal_entries_0_3_pal,
    normal_entries_0_2_pal,normal_entries_0_1_pal,normal_entries_0_0_pal}; // @[Cat.scala 29:58]
  wire [7:0] paa_array_if_cached_0 = paa_array_0 | c_array_0; // @[tlb.scala 227:56]
  wire [7:0] pal_array_if_cached_0 = pal_array_0 | c_array_0; // @[tlb.scala 228:56]
  wire  _T_1323 = cacheable_0 & homogeneous_0; // @[tlb.scala 229:61]
  wire [1:0] _T_1324 = {_T_1323, 1'h0}; // @[tlb.scala 229:80]
  wire [7:0] prefetchable_array_0 = {_T_1324,normal_entries_0_5_c,normal_entries_0_4_c,normal_entries_0_3_c,
    normal_entries_0_2_c,normal_entries_0_1_c,normal_entries_0_0_c}; // @[Cat.scala 29:58]
  wire [3:0] _T_1331 = 4'h1 << io_req_0_bits_size; // @[OneHot.scala 58:35]
  wire [3:0] _T_1333 = _T_1331 - 4'h1; // @[tlb.scala 231:89]
  wire [39:0] _GEN_346 = {{36'd0}, _T_1333}; // @[tlb.scala 231:56]
  wire [39:0] _T_1334 = io_req_0_bits_vaddr & _GEN_346; // @[tlb.scala 231:56]
  wire  misaligned_0 = |_T_1334; // @[tlb.scala 231:97]
  wire [39:0] _T_1336 = io_req_0_bits_vaddr & 40'hc000000000; // @[tlb.scala 237:46]
  wire  _T_1341 = ~(_T_1336 == 40'h0 | _T_1336 == 40'hc000000000); // @[tlb.scala 238:49]
  wire  bad_va_0 = vm_enabled_0 & _T_1341; // @[tlb.scala 232:134]
  wire  _T_1344 = io_req_0_bits_cmd == 5'h6; // @[package.scala 15:47]
  wire  _T_1345 = io_req_0_bits_cmd == 5'h7; // @[package.scala 15:47]
  wire  cmd_lrsc_0 = _T_1344 | _T_1345; // @[package.scala 64:59]
  wire  _T_1348 = io_req_0_bits_cmd == 5'h4; // @[package.scala 15:47]
  wire  _T_1349 = io_req_0_bits_cmd == 5'h9; // @[package.scala 15:47]
  wire  _T_1350 = io_req_0_bits_cmd == 5'ha; // @[package.scala 15:47]
  wire  _T_1351 = io_req_0_bits_cmd == 5'hb; // @[package.scala 15:47]
  wire  cmd_amo_logical_0 = _T_1348 | _T_1349 | _T_1350 | _T_1351; // @[package.scala 64:59]
  wire  _T_1356 = io_req_0_bits_cmd == 5'h8; // @[package.scala 15:47]
  wire  _T_1357 = io_req_0_bits_cmd == 5'hc; // @[package.scala 15:47]
  wire  _T_1358 = io_req_0_bits_cmd == 5'hd; // @[package.scala 15:47]
  wire  _T_1359 = io_req_0_bits_cmd == 5'he; // @[package.scala 15:47]
  wire  _T_1360 = io_req_0_bits_cmd == 5'hf; // @[package.scala 15:47]
  wire  cmd_amo_arithmetic_0 = _T_1356 | _T_1357 | _T_1358 | _T_1359 | _T_1360; // @[package.scala 64:59]
  wire  _T_1387 = cmd_amo_logical_0 | cmd_amo_arithmetic_0; // @[Consts.scala 80:44]
  wire  cmd_read_0 = io_req_0_bits_cmd == 5'h0 | _T_1344 | _T_1345 | _T_1387; // @[Consts.scala 82:75]
  wire  cmd_write_0 = io_req_0_bits_cmd == 5'h1 | io_req_0_bits_cmd == 5'h11 | _T_1345 | _T_1387; // @[Consts.scala 83:76]
  wire [7:0] _T_1416 = misaligned_0 ? eff_array_0 : 8'h0; // @[tlb.scala 252:8]
  wire [7:0] _T_1417 = ~c_array_0; // @[tlb.scala 253:24]
  wire [7:0] _T_1418 = cmd_lrsc_0 ? _T_1417 : 8'h0; // @[tlb.scala 253:8]
  wire [7:0] ae_array_0 = _T_1416 | _T_1418; // @[tlb.scala 252:43]
  wire [7:0] _T_1420 = ~pr_array_0; // @[tlb.scala 254:66]
  wire [7:0] _T_1421 = ae_array_0 | _T_1420; // @[tlb.scala 254:64]
  wire [7:0] ae_ld_array_0 = cmd_read_0 ? _T_1421 : 8'h0; // @[tlb.scala 254:38]
  wire [7:0] _T_1423 = ~pw_array_0; // @[tlb.scala 256:46]
  wire [7:0] _T_1424 = ae_array_0 | _T_1423; // @[tlb.scala 256:44]
  wire [7:0] _T_1425 = cmd_write_0 ? _T_1424 : 8'h0; // @[tlb.scala 256:8]
  wire [7:0] _T_1426 = ~pal_array_if_cached_0; // @[tlb.scala 257:32]
  wire [7:0] _T_1427 = cmd_amo_logical_0 ? _T_1426 : 8'h0; // @[tlb.scala 257:8]
  wire [7:0] _T_1428 = _T_1425 | _T_1427; // @[tlb.scala 256:65]
  wire [7:0] _T_1429 = ~paa_array_if_cached_0; // @[tlb.scala 258:32]
  wire [7:0] _T_1430 = cmd_amo_arithmetic_0 ? _T_1429 : 8'h0; // @[tlb.scala 258:8]
  wire [7:0] ae_st_array_0 = _T_1428 | _T_1430; // @[tlb.scala 257:62]
  wire [7:0] _T_1432 = ~paa_array_0; // @[tlb.scala 260:32]
  wire [7:0] _T_1433 = cmd_amo_logical_0 ? _T_1432 : 8'h0; // @[tlb.scala 260:8]
  wire [7:0] _T_1434 = ~pal_array_0; // @[tlb.scala 261:32]
  wire [7:0] _T_1435 = cmd_amo_arithmetic_0 ? _T_1434 : 8'h0; // @[tlb.scala 261:8]
  wire [7:0] _T_1436 = _T_1433 | _T_1435; // @[tlb.scala 260:52]
  wire [7:0] _T_1438 = cmd_lrsc_0 ? 8'hff : 8'h0; // @[tlb.scala 262:8]
  wire [7:0] must_alloc_array_0 = _T_1436 | _T_1438; // @[tlb.scala 261:52]
  wire [7:0] _T_1441 = ~eff_array_0; // @[tlb.scala 263:70]
  wire [7:0] ma_ld_array_0 = misaligned_0 & cmd_read_0 ? _T_1441 : 8'h0; // @[tlb.scala 263:38]
  wire [7:0] ma_st_array_0 = misaligned_0 & cmd_write_0 ? _T_1441 : 8'h0; // @[tlb.scala 264:38]
  wire [7:0] _T_1446 = r_array_0 | ptw_ae_array_0; // @[tlb.scala 265:72]
  wire [7:0] _T_1447 = ~_T_1446; // @[tlb.scala 265:59]
  wire [7:0] pf_ld_array_0 = cmd_read_0 ? _T_1447 : 8'h0; // @[tlb.scala 265:38]
  wire [7:0] _T_1449 = w_array_0 | ptw_ae_array_0; // @[tlb.scala 266:72]
  wire [7:0] _T_1450 = ~_T_1449; // @[tlb.scala 266:59]
  wire [7:0] pf_st_array_0 = cmd_write_0 ? _T_1450 : 8'h0; // @[tlb.scala 266:38]
  wire [7:0] _T_1452 = x_array_0 | ptw_ae_array_0; // @[tlb.scala 267:50]
  wire [7:0] pf_inst_array_0 = ~_T_1452; // @[tlb.scala 267:37]
  wire  tlb_hit_0 = |real_hits_0; // @[tlb.scala 269:44]
  wire  tlb_miss_0 = vm_enabled_0 & ~bad_va_0 & ~tlb_hit_0; // @[tlb.scala 270:60]
  reg  _T_1459; // @[Replacement.scala 42:30]
  reg [2:0] _T_1460; // @[Replacement.scala 42:30]
  wire  _T_1462 = sector_hits_0_0 | sector_hits_0_1; // @[package.scala 64:59]
  wire [1:0] _T_1463 = {sector_hits_0_1,sector_hits_0_0}; // @[OneHot.scala 22:45]
  wire [1:0] _T_1465 = {_T_1459, 1'h0}; // @[Replacement.scala 50:28]
  wire [1:0] _T_1469 = _T_1465 | 2'h2; // @[Replacement.scala 54:37]
  wire [1:0] _T_1470 = ~_T_1465; // @[Replacement.scala 54:37]
  wire [1:0] _T_1471 = _T_1470 | 2'h2; // @[Replacement.scala 54:37]
  wire [1:0] _T_1472 = ~_T_1471; // @[Replacement.scala 54:37]
  wire [1:0] _T_1473 = ~_T_1463[1] ? _T_1469 : _T_1472; // @[Replacement.scala 54:37]
  wire  _T_1478 = superpage_hits_0_0 | superpage_hits_0_1 | superpage_hits_0_2 | superpage_hits_0_3; // @[package.scala 64:59]
  wire [3:0] _T_1481 = {superpage_hits_0_3,superpage_hits_0_2,superpage_hits_0_1,superpage_hits_0_0}; // @[OneHot.scala 22:45]
  wire  _T_1484 = |_T_1481[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_1485 = _T_1481[3:2] | _T_1481[1:0]; // @[OneHot.scala 32:28]
  wire [1:0] _T_1487 = {_T_1484,_T_1485[1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1488 = {_T_1460, 1'h0}; // @[Replacement.scala 50:28]
  wire [3:0] _T_1492 = _T_1488 | 4'h2; // @[Replacement.scala 54:37]
  wire [3:0] _T_1493 = ~_T_1488; // @[Replacement.scala 54:37]
  wire [3:0] _T_1494 = _T_1493 | 4'h2; // @[Replacement.scala 54:37]
  wire [3:0] _T_1495 = ~_T_1494; // @[Replacement.scala 54:37]
  wire [3:0] _T_1496 = ~_T_1487[1] ? _T_1492 : _T_1495; // @[Replacement.scala 54:37]
  wire [1:0] _T_1497 = {1'h1,_T_1487[1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1500 = 4'h1 << _T_1497; // @[Replacement.scala 54:37]
  wire [3:0] _T_1501 = _T_1496 | _T_1500; // @[Replacement.scala 54:37]
  wire [3:0] _T_1502 = ~_T_1496; // @[Replacement.scala 54:37]
  wire [3:0] _T_1503 = _T_1502 | _T_1500; // @[Replacement.scala 54:37]
  wire [3:0] _T_1504 = ~_T_1503; // @[Replacement.scala 54:37]
  wire [3:0] _T_1505 = ~_T_1487[0] ? _T_1501 : _T_1504; // @[Replacement.scala 54:37]
  wire  multipleHits_0 = real_hits_0[1] & real_hits_0[2] | real_hits_0[0] & (real_hits_0[1] | real_hits_0[2]) | (
    real_hits_0[3] & real_hits_0[4] | real_hits_0[5] & real_hits_0[6] | (real_hits_0[3] | real_hits_0[4]) & (real_hits_0
    [5] | real_hits_0[6])) | (real_hits_0[0] | (real_hits_0[1] | real_hits_0[2])) & (real_hits_0[3] | real_hits_0[4] | (
    real_hits_0[5] | real_hits_0[6])); // @[Misc.scala 182:49]
  wire  _T_1551 = state == 2'h0; // @[tlb.scala 288:24]
  wire [7:0] _T_1553 = pf_ld_array_0 & hits_0; // @[tlb.scala 291:73]
  wire [7:0] _T_1557 = pf_st_array_0 & hits_0; // @[tlb.scala 292:80]
  wire [7:0] _T_1560 = pf_inst_array_0 & hits_0; // @[tlb.scala 293:58]
  wire [7:0] _T_1563 = ae_ld_array_0 & hits_0; // @[tlb.scala 294:43]
  wire [7:0] _T_1565 = ae_st_array_0 & hits_0; // @[tlb.scala 295:43]
  wire [7:0] _T_1567 = ~px_array_0; // @[tlb.scala 296:28]
  wire [7:0] _T_1568 = _T_1567 & hits_0; // @[tlb.scala 296:43]
  wire [7:0] _T_1570 = ma_ld_array_0 & hits_0; // @[tlb.scala 297:43]
  wire [7:0] _T_1572 = ma_st_array_0 & hits_0; // @[tlb.scala 298:43]
  wire [7:0] _T_1574 = c_array_0 & hits_0; // @[tlb.scala 300:44]
  wire [7:0] _T_1576 = must_alloc_array_0 & hits_0; // @[tlb.scala 301:53]
  wire [7:0] _T_1578 = prefetchable_array_0 & hits_0; // @[tlb.scala 302:55]
  wire  _T_1587 = io_req_0_ready & io_req_0_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_1595 = {{1'd0}, _T_1488[3:1]}; // @[Replacement.scala 65:48]
  wire [1:0] _T_1598 = {1'h1,_T_1595[0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1602 = _T_1488 >> _T_1598; // @[Replacement.scala 65:48]
  wire [2:0] _T_1605 = {1'h1,_T_1595[0],_T_1602[0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1609 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,
    superpage_entries_0_valid_0}; // @[Cat.scala 29:58]
  wire [3:0] _T_1611 = ~_T_1609; // @[tlb.scala 353:43]
  wire [1:0] _T_1616 = _T_1611[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:69]
  wire [1:0] _T_1624 = {{1'd0}, _T_1465[1]}; // @[Replacement.scala 65:48]
  wire [1:0] _T_1627 = {1'h1,_T_1624[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_1635 = {_T_394,_T_387}; // @[Cat.scala 29:58]
  wire [1:0] _T_1637 = ~_T_1635; // @[tlb.scala 353:43]
  wire [1:0] _GEN_212 = _T_1587 & tlb_miss_0 & _T_1551 ? 2'h1 : state; // @[tlb.scala 314:67 315:15 129:22]
  wire [1:0] _GEN_218 = io_sfence_valid ? 2'h0 : _GEN_212; // @[tlb.scala 325:{21,29}]
  wire [1:0] _T_1646 = io_sfence_valid ? 2'h3 : 2'h2; // @[tlb.scala 326:45]
  wire [1:0] _GEN_219 = io_ptw_req_ready ? _T_1646 : _GEN_218; // @[tlb.scala 326:{31,39}]
  wire [1:0] _GEN_220 = io_kill ? 2'h0 : _GEN_219; // @[tlb.scala 327:{22,30}]
  wire  _GEN_224 = 2'h0 == vpn_0[1:0] ? 1'h0 : _GEN_172; // @[tlb.scala 103:{60,60}]
  wire  _GEN_225 = 2'h1 == vpn_0[1:0] ? 1'h0 : _GEN_173; // @[tlb.scala 103:{60,60}]
  wire  _GEN_226 = 2'h2 == vpn_0[1:0] ? 1'h0 : _GEN_174; // @[tlb.scala 103:{60,60}]
  wire  _GEN_227 = 2'h3 == vpn_0[1:0] ? 1'h0 : _GEN_175; // @[tlb.scala 103:{60,60}]
  wire  _GEN_228 = _T_390 ? _GEN_224 : _GEN_172; // @[tlb.scala 103:36]
  wire  _GEN_229 = _T_390 ? _GEN_225 : _GEN_173; // @[tlb.scala 103:36]
  wire  _GEN_230 = _T_390 ? _GEN_226 : _GEN_174; // @[tlb.scala 103:36]
  wire  _GEN_231 = _T_390 ? _GEN_227 : _GEN_175; // @[tlb.scala 103:36]
  wire  _GEN_232 = sectored_entries_0_data_0[0] ? 1'h0 : _GEN_228; // @[tlb.scala 109:{44,48}]
  wire  _GEN_233 = sectored_entries_0_data_1[0] ? 1'h0 : _GEN_229; // @[tlb.scala 109:{44,48}]
  wire  _GEN_234 = sectored_entries_0_data_2[0] ? 1'h0 : _GEN_230; // @[tlb.scala 109:{44,48}]
  wire  _GEN_235 = sectored_entries_0_data_3[0] ? 1'h0 : _GEN_231; // @[tlb.scala 109:{44,48}]
  wire  _GEN_240 = ~sectored_entries_0_data_0[12] ? 1'h0 : _GEN_172; // @[tlb.scala 115:{22,26}]
  wire  _GEN_241 = ~sectored_entries_0_data_1[12] ? 1'h0 : _GEN_173; // @[tlb.scala 115:{22,26}]
  wire  _GEN_242 = ~sectored_entries_0_data_2[12] ? 1'h0 : _GEN_174; // @[tlb.scala 115:{22,26}]
  wire  _GEN_243 = ~sectored_entries_0_data_3[12] ? 1'h0 : _GEN_175; // @[tlb.scala 115:{22,26}]
  wire  _GEN_244 = io_sfence_bits_rs2 & _GEN_240; // @[tlb.scala 341:42 98:40]
  wire  _GEN_245 = io_sfence_bits_rs2 & _GEN_241; // @[tlb.scala 341:42 98:40]
  wire  _GEN_246 = io_sfence_bits_rs2 & _GEN_242; // @[tlb.scala 341:42 98:40]
  wire  _GEN_247 = io_sfence_bits_rs2 & _GEN_243; // @[tlb.scala 341:42 98:40]
  wire  _GEN_252 = 2'h0 == vpn_0[1:0] ? 1'h0 : _GEN_182; // @[tlb.scala 103:{60,60}]
  wire  _GEN_253 = 2'h1 == vpn_0[1:0] ? 1'h0 : _GEN_183; // @[tlb.scala 103:{60,60}]
  wire  _GEN_254 = 2'h2 == vpn_0[1:0] ? 1'h0 : _GEN_184; // @[tlb.scala 103:{60,60}]
  wire  _GEN_255 = 2'h3 == vpn_0[1:0] ? 1'h0 : _GEN_185; // @[tlb.scala 103:{60,60}]
  wire  _GEN_256 = _T_397 ? _GEN_252 : _GEN_182; // @[tlb.scala 103:36]
  wire  _GEN_257 = _T_397 ? _GEN_253 : _GEN_183; // @[tlb.scala 103:36]
  wire  _GEN_258 = _T_397 ? _GEN_254 : _GEN_184; // @[tlb.scala 103:36]
  wire  _GEN_259 = _T_397 ? _GEN_255 : _GEN_185; // @[tlb.scala 103:36]
  wire  _GEN_260 = sectored_entries_1_data_0[0] ? 1'h0 : _GEN_256; // @[tlb.scala 109:{44,48}]
  wire  _GEN_261 = sectored_entries_1_data_1[0] ? 1'h0 : _GEN_257; // @[tlb.scala 109:{44,48}]
  wire  _GEN_262 = sectored_entries_1_data_2[0] ? 1'h0 : _GEN_258; // @[tlb.scala 109:{44,48}]
  wire  _GEN_263 = sectored_entries_1_data_3[0] ? 1'h0 : _GEN_259; // @[tlb.scala 109:{44,48}]
  wire  _GEN_268 = ~sectored_entries_1_data_0[12] ? 1'h0 : _GEN_182; // @[tlb.scala 115:{22,26}]
  wire  _GEN_269 = ~sectored_entries_1_data_1[12] ? 1'h0 : _GEN_183; // @[tlb.scala 115:{22,26}]
  wire  _GEN_270 = ~sectored_entries_1_data_2[12] ? 1'h0 : _GEN_184; // @[tlb.scala 115:{22,26}]
  wire  _GEN_271 = ~sectored_entries_1_data_3[12] ? 1'h0 : _GEN_185; // @[tlb.scala 115:{22,26}]
  wire  _GEN_272 = io_sfence_bits_rs2 & _GEN_268; // @[tlb.scala 341:42 98:40]
  wire  _GEN_273 = io_sfence_bits_rs2 & _GEN_269; // @[tlb.scala 341:42 98:40]
  wire  _GEN_274 = io_sfence_bits_rs2 & _GEN_270; // @[tlb.scala 341:42 98:40]
  wire  _GEN_275 = io_sfence_bits_rs2 & _GEN_271; // @[tlb.scala 341:42 98:40]
  wire  _GEN_281 = ~superpage_entries_0_data_0[12] ? 1'h0 : _GEN_158; // @[tlb.scala 115:{22,26}]
  wire  _GEN_282 = io_sfence_bits_rs2 & _GEN_281; // @[tlb.scala 341:42 98:40]
  wire  _GEN_285 = ~superpage_entries_1_data_0[12] ? 1'h0 : _GEN_162; // @[tlb.scala 115:{22,26}]
  wire  _GEN_286 = io_sfence_bits_rs2 & _GEN_285; // @[tlb.scala 341:42 98:40]
  wire  _GEN_289 = ~superpage_entries_2_data_0[12] ? 1'h0 : _GEN_166; // @[tlb.scala 115:{22,26}]
  wire  _GEN_290 = io_sfence_bits_rs2 & _GEN_289; // @[tlb.scala 341:42 98:40]
  wire  _GEN_293 = ~superpage_entries_3_data_0[12] ? 1'h0 : _GEN_170; // @[tlb.scala 115:{22,26}]
  wire  _GEN_294 = io_sfence_bits_rs2 & _GEN_293; // @[tlb.scala 341:42 98:40]
  wire  _GEN_297 = ~special_entry_data_0[12] ? 1'h0 : _GEN_154; // @[tlb.scala 115:{22,26}]
  wire  _GEN_298 = io_sfence_bits_rs2 & _GEN_297; // @[tlb.scala 341:42 98:40]
  package_Anon_46 package_Anon ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_io_x_ppn),
    .io_x_u(package_Anon_io_x_u),
    .io_x_ae(package_Anon_io_x_ae),
    .io_x_sw(package_Anon_io_x_sw),
    .io_x_sx(package_Anon_io_x_sx),
    .io_x_sr(package_Anon_io_x_sr),
    .io_x_pw(package_Anon_io_x_pw),
    .io_x_px(package_Anon_io_x_px),
    .io_x_pr(package_Anon_io_x_pr),
    .io_x_pal(package_Anon_io_x_pal),
    .io_x_paa(package_Anon_io_x_paa),
    .io_x_eff(package_Anon_io_x_eff),
    .io_x_c(package_Anon_io_x_c),
    .io_y_ppn(package_Anon_io_y_ppn),
    .io_y_u(package_Anon_io_y_u),
    .io_y_ae(package_Anon_io_y_ae),
    .io_y_sw(package_Anon_io_y_sw),
    .io_y_sx(package_Anon_io_y_sx),
    .io_y_sr(package_Anon_io_y_sr),
    .io_y_pw(package_Anon_io_y_pw),
    .io_y_px(package_Anon_io_y_px),
    .io_y_pr(package_Anon_io_y_pr),
    .io_y_pal(package_Anon_io_y_pal),
    .io_y_paa(package_Anon_io_y_paa),
    .io_y_eff(package_Anon_io_y_eff),
    .io_y_c(package_Anon_io_y_c)
  );
  PMPChecker_1 pmp_0 ( // @[tlb.scala 150:40]
    .io_prv(pmp_0_io_prv),
    .io_pmp_0_cfg_l(pmp_0_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_0_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_0_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_0_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_0_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_0_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_0_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_0_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_0_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_0_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_0_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_0_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_0_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_0_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_0_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_0_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_0_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_0_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_0_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_0_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_0_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_0_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_0_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_0_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_0_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_0_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_0_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_0_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_0_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_0_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_0_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_0_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_0_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_0_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_0_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_0_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_0_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_0_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_0_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_0_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_0_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_0_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_0_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_0_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_0_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_0_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_0_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_0_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_0_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_0_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_0_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_0_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_0_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_0_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_0_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_0_io_pmp_7_mask),
    .io_addr(pmp_0_io_addr),
    .io_size(pmp_0_io_size),
    .io_r(pmp_0_io_r),
    .io_w(pmp_0_io_w),
    .io_x(pmp_0_io_x)
  );
  package_Anon_46 package_Anon_1 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_1_io_x_ppn),
    .io_x_u(package_Anon_1_io_x_u),
    .io_x_ae(package_Anon_1_io_x_ae),
    .io_x_sw(package_Anon_1_io_x_sw),
    .io_x_sx(package_Anon_1_io_x_sx),
    .io_x_sr(package_Anon_1_io_x_sr),
    .io_x_pw(package_Anon_1_io_x_pw),
    .io_x_px(package_Anon_1_io_x_px),
    .io_x_pr(package_Anon_1_io_x_pr),
    .io_x_pal(package_Anon_1_io_x_pal),
    .io_x_paa(package_Anon_1_io_x_paa),
    .io_x_eff(package_Anon_1_io_x_eff),
    .io_x_c(package_Anon_1_io_x_c),
    .io_y_ppn(package_Anon_1_io_y_ppn),
    .io_y_u(package_Anon_1_io_y_u),
    .io_y_ae(package_Anon_1_io_y_ae),
    .io_y_sw(package_Anon_1_io_y_sw),
    .io_y_sx(package_Anon_1_io_y_sx),
    .io_y_sr(package_Anon_1_io_y_sr),
    .io_y_pw(package_Anon_1_io_y_pw),
    .io_y_px(package_Anon_1_io_y_px),
    .io_y_pr(package_Anon_1_io_y_pr),
    .io_y_pal(package_Anon_1_io_y_pal),
    .io_y_paa(package_Anon_1_io_y_paa),
    .io_y_eff(package_Anon_1_io_y_eff),
    .io_y_c(package_Anon_1_io_y_c)
  );
  package_Anon_46 package_Anon_2 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_2_io_x_ppn),
    .io_x_u(package_Anon_2_io_x_u),
    .io_x_ae(package_Anon_2_io_x_ae),
    .io_x_sw(package_Anon_2_io_x_sw),
    .io_x_sx(package_Anon_2_io_x_sx),
    .io_x_sr(package_Anon_2_io_x_sr),
    .io_x_pw(package_Anon_2_io_x_pw),
    .io_x_px(package_Anon_2_io_x_px),
    .io_x_pr(package_Anon_2_io_x_pr),
    .io_x_pal(package_Anon_2_io_x_pal),
    .io_x_paa(package_Anon_2_io_x_paa),
    .io_x_eff(package_Anon_2_io_x_eff),
    .io_x_c(package_Anon_2_io_x_c),
    .io_y_ppn(package_Anon_2_io_y_ppn),
    .io_y_u(package_Anon_2_io_y_u),
    .io_y_ae(package_Anon_2_io_y_ae),
    .io_y_sw(package_Anon_2_io_y_sw),
    .io_y_sx(package_Anon_2_io_y_sx),
    .io_y_sr(package_Anon_2_io_y_sr),
    .io_y_pw(package_Anon_2_io_y_pw),
    .io_y_px(package_Anon_2_io_y_px),
    .io_y_pr(package_Anon_2_io_y_pr),
    .io_y_pal(package_Anon_2_io_y_pal),
    .io_y_paa(package_Anon_2_io_y_paa),
    .io_y_eff(package_Anon_2_io_y_eff),
    .io_y_c(package_Anon_2_io_y_c)
  );
  package_Anon_46 package_Anon_3 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_3_io_x_ppn),
    .io_x_u(package_Anon_3_io_x_u),
    .io_x_ae(package_Anon_3_io_x_ae),
    .io_x_sw(package_Anon_3_io_x_sw),
    .io_x_sx(package_Anon_3_io_x_sx),
    .io_x_sr(package_Anon_3_io_x_sr),
    .io_x_pw(package_Anon_3_io_x_pw),
    .io_x_px(package_Anon_3_io_x_px),
    .io_x_pr(package_Anon_3_io_x_pr),
    .io_x_pal(package_Anon_3_io_x_pal),
    .io_x_paa(package_Anon_3_io_x_paa),
    .io_x_eff(package_Anon_3_io_x_eff),
    .io_x_c(package_Anon_3_io_x_c),
    .io_y_ppn(package_Anon_3_io_y_ppn),
    .io_y_u(package_Anon_3_io_y_u),
    .io_y_ae(package_Anon_3_io_y_ae),
    .io_y_sw(package_Anon_3_io_y_sw),
    .io_y_sx(package_Anon_3_io_y_sx),
    .io_y_sr(package_Anon_3_io_y_sr),
    .io_y_pw(package_Anon_3_io_y_pw),
    .io_y_px(package_Anon_3_io_y_px),
    .io_y_pr(package_Anon_3_io_y_pr),
    .io_y_pal(package_Anon_3_io_y_pal),
    .io_y_paa(package_Anon_3_io_y_paa),
    .io_y_eff(package_Anon_3_io_y_eff),
    .io_y_c(package_Anon_3_io_y_c)
  );
  package_Anon_46 package_Anon_4 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_4_io_x_ppn),
    .io_x_u(package_Anon_4_io_x_u),
    .io_x_ae(package_Anon_4_io_x_ae),
    .io_x_sw(package_Anon_4_io_x_sw),
    .io_x_sx(package_Anon_4_io_x_sx),
    .io_x_sr(package_Anon_4_io_x_sr),
    .io_x_pw(package_Anon_4_io_x_pw),
    .io_x_px(package_Anon_4_io_x_px),
    .io_x_pr(package_Anon_4_io_x_pr),
    .io_x_pal(package_Anon_4_io_x_pal),
    .io_x_paa(package_Anon_4_io_x_paa),
    .io_x_eff(package_Anon_4_io_x_eff),
    .io_x_c(package_Anon_4_io_x_c),
    .io_y_ppn(package_Anon_4_io_y_ppn),
    .io_y_u(package_Anon_4_io_y_u),
    .io_y_ae(package_Anon_4_io_y_ae),
    .io_y_sw(package_Anon_4_io_y_sw),
    .io_y_sx(package_Anon_4_io_y_sx),
    .io_y_sr(package_Anon_4_io_y_sr),
    .io_y_pw(package_Anon_4_io_y_pw),
    .io_y_px(package_Anon_4_io_y_px),
    .io_y_pr(package_Anon_4_io_y_pr),
    .io_y_pal(package_Anon_4_io_y_pal),
    .io_y_paa(package_Anon_4_io_y_paa),
    .io_y_eff(package_Anon_4_io_y_eff),
    .io_y_c(package_Anon_4_io_y_c)
  );
  package_Anon_46 package_Anon_5 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_5_io_x_ppn),
    .io_x_u(package_Anon_5_io_x_u),
    .io_x_ae(package_Anon_5_io_x_ae),
    .io_x_sw(package_Anon_5_io_x_sw),
    .io_x_sx(package_Anon_5_io_x_sx),
    .io_x_sr(package_Anon_5_io_x_sr),
    .io_x_pw(package_Anon_5_io_x_pw),
    .io_x_px(package_Anon_5_io_x_px),
    .io_x_pr(package_Anon_5_io_x_pr),
    .io_x_pal(package_Anon_5_io_x_pal),
    .io_x_paa(package_Anon_5_io_x_paa),
    .io_x_eff(package_Anon_5_io_x_eff),
    .io_x_c(package_Anon_5_io_x_c),
    .io_y_ppn(package_Anon_5_io_y_ppn),
    .io_y_u(package_Anon_5_io_y_u),
    .io_y_ae(package_Anon_5_io_y_ae),
    .io_y_sw(package_Anon_5_io_y_sw),
    .io_y_sx(package_Anon_5_io_y_sx),
    .io_y_sr(package_Anon_5_io_y_sr),
    .io_y_pw(package_Anon_5_io_y_pw),
    .io_y_px(package_Anon_5_io_y_px),
    .io_y_pr(package_Anon_5_io_y_pr),
    .io_y_pal(package_Anon_5_io_y_pal),
    .io_y_paa(package_Anon_5_io_y_paa),
    .io_y_eff(package_Anon_5_io_y_eff),
    .io_y_c(package_Anon_5_io_y_c)
  );
  package_Anon_46 package_Anon_6 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_6_io_x_ppn),
    .io_x_u(package_Anon_6_io_x_u),
    .io_x_ae(package_Anon_6_io_x_ae),
    .io_x_sw(package_Anon_6_io_x_sw),
    .io_x_sx(package_Anon_6_io_x_sx),
    .io_x_sr(package_Anon_6_io_x_sr),
    .io_x_pw(package_Anon_6_io_x_pw),
    .io_x_px(package_Anon_6_io_x_px),
    .io_x_pr(package_Anon_6_io_x_pr),
    .io_x_pal(package_Anon_6_io_x_pal),
    .io_x_paa(package_Anon_6_io_x_paa),
    .io_x_eff(package_Anon_6_io_x_eff),
    .io_x_c(package_Anon_6_io_x_c),
    .io_y_ppn(package_Anon_6_io_y_ppn),
    .io_y_u(package_Anon_6_io_y_u),
    .io_y_ae(package_Anon_6_io_y_ae),
    .io_y_sw(package_Anon_6_io_y_sw),
    .io_y_sx(package_Anon_6_io_y_sx),
    .io_y_sr(package_Anon_6_io_y_sr),
    .io_y_pw(package_Anon_6_io_y_pw),
    .io_y_px(package_Anon_6_io_y_px),
    .io_y_pr(package_Anon_6_io_y_pr),
    .io_y_pal(package_Anon_6_io_y_pal),
    .io_y_paa(package_Anon_6_io_y_paa),
    .io_y_eff(package_Anon_6_io_y_eff),
    .io_y_c(package_Anon_6_io_y_c)
  );
  package_Anon_46 package_Anon_7 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_7_io_x_ppn),
    .io_x_u(package_Anon_7_io_x_u),
    .io_x_ae(package_Anon_7_io_x_ae),
    .io_x_sw(package_Anon_7_io_x_sw),
    .io_x_sx(package_Anon_7_io_x_sx),
    .io_x_sr(package_Anon_7_io_x_sr),
    .io_x_pw(package_Anon_7_io_x_pw),
    .io_x_px(package_Anon_7_io_x_px),
    .io_x_pr(package_Anon_7_io_x_pr),
    .io_x_pal(package_Anon_7_io_x_pal),
    .io_x_paa(package_Anon_7_io_x_paa),
    .io_x_eff(package_Anon_7_io_x_eff),
    .io_x_c(package_Anon_7_io_x_c),
    .io_y_ppn(package_Anon_7_io_y_ppn),
    .io_y_u(package_Anon_7_io_y_u),
    .io_y_ae(package_Anon_7_io_y_ae),
    .io_y_sw(package_Anon_7_io_y_sw),
    .io_y_sx(package_Anon_7_io_y_sx),
    .io_y_sr(package_Anon_7_io_y_sr),
    .io_y_pw(package_Anon_7_io_y_pw),
    .io_y_px(package_Anon_7_io_y_px),
    .io_y_pr(package_Anon_7_io_y_pr),
    .io_y_pal(package_Anon_7_io_y_pal),
    .io_y_paa(package_Anon_7_io_y_paa),
    .io_y_eff(package_Anon_7_io_y_eff),
    .io_y_c(package_Anon_7_io_y_c)
  );
  package_Anon_46 package_Anon_8 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_8_io_x_ppn),
    .io_x_u(package_Anon_8_io_x_u),
    .io_x_ae(package_Anon_8_io_x_ae),
    .io_x_sw(package_Anon_8_io_x_sw),
    .io_x_sx(package_Anon_8_io_x_sx),
    .io_x_sr(package_Anon_8_io_x_sr),
    .io_x_pw(package_Anon_8_io_x_pw),
    .io_x_px(package_Anon_8_io_x_px),
    .io_x_pr(package_Anon_8_io_x_pr),
    .io_x_pal(package_Anon_8_io_x_pal),
    .io_x_paa(package_Anon_8_io_x_paa),
    .io_x_eff(package_Anon_8_io_x_eff),
    .io_x_c(package_Anon_8_io_x_c),
    .io_y_ppn(package_Anon_8_io_y_ppn),
    .io_y_u(package_Anon_8_io_y_u),
    .io_y_ae(package_Anon_8_io_y_ae),
    .io_y_sw(package_Anon_8_io_y_sw),
    .io_y_sx(package_Anon_8_io_y_sx),
    .io_y_sr(package_Anon_8_io_y_sr),
    .io_y_pw(package_Anon_8_io_y_pw),
    .io_y_px(package_Anon_8_io_y_px),
    .io_y_pr(package_Anon_8_io_y_pr),
    .io_y_pal(package_Anon_8_io_y_pal),
    .io_y_paa(package_Anon_8_io_y_paa),
    .io_y_eff(package_Anon_8_io_y_eff),
    .io_y_c(package_Anon_8_io_y_c)
  );
  package_Anon_46 package_Anon_9 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_9_io_x_ppn),
    .io_x_u(package_Anon_9_io_x_u),
    .io_x_ae(package_Anon_9_io_x_ae),
    .io_x_sw(package_Anon_9_io_x_sw),
    .io_x_sx(package_Anon_9_io_x_sx),
    .io_x_sr(package_Anon_9_io_x_sr),
    .io_x_pw(package_Anon_9_io_x_pw),
    .io_x_px(package_Anon_9_io_x_px),
    .io_x_pr(package_Anon_9_io_x_pr),
    .io_x_pal(package_Anon_9_io_x_pal),
    .io_x_paa(package_Anon_9_io_x_paa),
    .io_x_eff(package_Anon_9_io_x_eff),
    .io_x_c(package_Anon_9_io_x_c),
    .io_y_ppn(package_Anon_9_io_y_ppn),
    .io_y_u(package_Anon_9_io_y_u),
    .io_y_ae(package_Anon_9_io_y_ae),
    .io_y_sw(package_Anon_9_io_y_sw),
    .io_y_sx(package_Anon_9_io_y_sx),
    .io_y_sr(package_Anon_9_io_y_sr),
    .io_y_pw(package_Anon_9_io_y_pw),
    .io_y_px(package_Anon_9_io_y_px),
    .io_y_pr(package_Anon_9_io_y_pr),
    .io_y_pal(package_Anon_9_io_y_pal),
    .io_y_paa(package_Anon_9_io_y_paa),
    .io_y_eff(package_Anon_9_io_y_eff),
    .io_y_c(package_Anon_9_io_y_c)
  );
  package_Anon_46 package_Anon_10 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_10_io_x_ppn),
    .io_x_u(package_Anon_10_io_x_u),
    .io_x_ae(package_Anon_10_io_x_ae),
    .io_x_sw(package_Anon_10_io_x_sw),
    .io_x_sx(package_Anon_10_io_x_sx),
    .io_x_sr(package_Anon_10_io_x_sr),
    .io_x_pw(package_Anon_10_io_x_pw),
    .io_x_px(package_Anon_10_io_x_px),
    .io_x_pr(package_Anon_10_io_x_pr),
    .io_x_pal(package_Anon_10_io_x_pal),
    .io_x_paa(package_Anon_10_io_x_paa),
    .io_x_eff(package_Anon_10_io_x_eff),
    .io_x_c(package_Anon_10_io_x_c),
    .io_y_ppn(package_Anon_10_io_y_ppn),
    .io_y_u(package_Anon_10_io_y_u),
    .io_y_ae(package_Anon_10_io_y_ae),
    .io_y_sw(package_Anon_10_io_y_sw),
    .io_y_sx(package_Anon_10_io_y_sx),
    .io_y_sr(package_Anon_10_io_y_sr),
    .io_y_pw(package_Anon_10_io_y_pw),
    .io_y_px(package_Anon_10_io_y_px),
    .io_y_pr(package_Anon_10_io_y_pr),
    .io_y_pal(package_Anon_10_io_y_pal),
    .io_y_paa(package_Anon_10_io_y_paa),
    .io_y_eff(package_Anon_10_io_y_eff),
    .io_y_c(package_Anon_10_io_y_c)
  );
  package_Anon_46 package_Anon_11 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_11_io_x_ppn),
    .io_x_u(package_Anon_11_io_x_u),
    .io_x_ae(package_Anon_11_io_x_ae),
    .io_x_sw(package_Anon_11_io_x_sw),
    .io_x_sx(package_Anon_11_io_x_sx),
    .io_x_sr(package_Anon_11_io_x_sr),
    .io_x_pw(package_Anon_11_io_x_pw),
    .io_x_px(package_Anon_11_io_x_px),
    .io_x_pr(package_Anon_11_io_x_pr),
    .io_x_pal(package_Anon_11_io_x_pal),
    .io_x_paa(package_Anon_11_io_x_paa),
    .io_x_eff(package_Anon_11_io_x_eff),
    .io_x_c(package_Anon_11_io_x_c),
    .io_y_ppn(package_Anon_11_io_y_ppn),
    .io_y_u(package_Anon_11_io_y_u),
    .io_y_ae(package_Anon_11_io_y_ae),
    .io_y_sw(package_Anon_11_io_y_sw),
    .io_y_sx(package_Anon_11_io_y_sx),
    .io_y_sr(package_Anon_11_io_y_sr),
    .io_y_pw(package_Anon_11_io_y_pw),
    .io_y_px(package_Anon_11_io_y_px),
    .io_y_pr(package_Anon_11_io_y_pr),
    .io_y_pal(package_Anon_11_io_y_pal),
    .io_y_paa(package_Anon_11_io_y_paa),
    .io_y_eff(package_Anon_11_io_y_eff),
    .io_y_c(package_Anon_11_io_y_c)
  );
  package_Anon_46 package_Anon_12 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_12_io_x_ppn),
    .io_x_u(package_Anon_12_io_x_u),
    .io_x_ae(package_Anon_12_io_x_ae),
    .io_x_sw(package_Anon_12_io_x_sw),
    .io_x_sx(package_Anon_12_io_x_sx),
    .io_x_sr(package_Anon_12_io_x_sr),
    .io_x_pw(package_Anon_12_io_x_pw),
    .io_x_px(package_Anon_12_io_x_px),
    .io_x_pr(package_Anon_12_io_x_pr),
    .io_x_pal(package_Anon_12_io_x_pal),
    .io_x_paa(package_Anon_12_io_x_paa),
    .io_x_eff(package_Anon_12_io_x_eff),
    .io_x_c(package_Anon_12_io_x_c),
    .io_y_ppn(package_Anon_12_io_y_ppn),
    .io_y_u(package_Anon_12_io_y_u),
    .io_y_ae(package_Anon_12_io_y_ae),
    .io_y_sw(package_Anon_12_io_y_sw),
    .io_y_sx(package_Anon_12_io_y_sx),
    .io_y_sr(package_Anon_12_io_y_sr),
    .io_y_pw(package_Anon_12_io_y_pw),
    .io_y_px(package_Anon_12_io_y_px),
    .io_y_pr(package_Anon_12_io_y_pr),
    .io_y_pal(package_Anon_12_io_y_pal),
    .io_y_paa(package_Anon_12_io_y_paa),
    .io_y_eff(package_Anon_12_io_y_eff),
    .io_y_c(package_Anon_12_io_y_c)
  );
  package_Anon_46 package_Anon_13 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_13_io_x_ppn),
    .io_x_u(package_Anon_13_io_x_u),
    .io_x_ae(package_Anon_13_io_x_ae),
    .io_x_sw(package_Anon_13_io_x_sw),
    .io_x_sx(package_Anon_13_io_x_sx),
    .io_x_sr(package_Anon_13_io_x_sr),
    .io_x_pw(package_Anon_13_io_x_pw),
    .io_x_px(package_Anon_13_io_x_px),
    .io_x_pr(package_Anon_13_io_x_pr),
    .io_x_pal(package_Anon_13_io_x_pal),
    .io_x_paa(package_Anon_13_io_x_paa),
    .io_x_eff(package_Anon_13_io_x_eff),
    .io_x_c(package_Anon_13_io_x_c),
    .io_y_ppn(package_Anon_13_io_y_ppn),
    .io_y_u(package_Anon_13_io_y_u),
    .io_y_ae(package_Anon_13_io_y_ae),
    .io_y_sw(package_Anon_13_io_y_sw),
    .io_y_sx(package_Anon_13_io_y_sx),
    .io_y_sr(package_Anon_13_io_y_sr),
    .io_y_pw(package_Anon_13_io_y_pw),
    .io_y_px(package_Anon_13_io_y_px),
    .io_y_pr(package_Anon_13_io_y_pr),
    .io_y_pal(package_Anon_13_io_y_pal),
    .io_y_paa(package_Anon_13_io_y_paa),
    .io_y_eff(package_Anon_13_io_y_eff),
    .io_y_c(package_Anon_13_io_y_c)
  );
  package_Anon_46 package_Anon_14 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_14_io_x_ppn),
    .io_x_u(package_Anon_14_io_x_u),
    .io_x_ae(package_Anon_14_io_x_ae),
    .io_x_sw(package_Anon_14_io_x_sw),
    .io_x_sx(package_Anon_14_io_x_sx),
    .io_x_sr(package_Anon_14_io_x_sr),
    .io_x_pw(package_Anon_14_io_x_pw),
    .io_x_px(package_Anon_14_io_x_px),
    .io_x_pr(package_Anon_14_io_x_pr),
    .io_x_pal(package_Anon_14_io_x_pal),
    .io_x_paa(package_Anon_14_io_x_paa),
    .io_x_eff(package_Anon_14_io_x_eff),
    .io_x_c(package_Anon_14_io_x_c),
    .io_y_ppn(package_Anon_14_io_y_ppn),
    .io_y_u(package_Anon_14_io_y_u),
    .io_y_ae(package_Anon_14_io_y_ae),
    .io_y_sw(package_Anon_14_io_y_sw),
    .io_y_sx(package_Anon_14_io_y_sx),
    .io_y_sr(package_Anon_14_io_y_sr),
    .io_y_pw(package_Anon_14_io_y_pw),
    .io_y_px(package_Anon_14_io_y_px),
    .io_y_pr(package_Anon_14_io_y_pr),
    .io_y_pal(package_Anon_14_io_y_pal),
    .io_y_paa(package_Anon_14_io_y_paa),
    .io_y_eff(package_Anon_14_io_y_eff),
    .io_y_c(package_Anon_14_io_y_c)
  );
  package_Anon_46 package_Anon_15 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_15_io_x_ppn),
    .io_x_u(package_Anon_15_io_x_u),
    .io_x_ae(package_Anon_15_io_x_ae),
    .io_x_sw(package_Anon_15_io_x_sw),
    .io_x_sx(package_Anon_15_io_x_sx),
    .io_x_sr(package_Anon_15_io_x_sr),
    .io_x_pw(package_Anon_15_io_x_pw),
    .io_x_px(package_Anon_15_io_x_px),
    .io_x_pr(package_Anon_15_io_x_pr),
    .io_x_pal(package_Anon_15_io_x_pal),
    .io_x_paa(package_Anon_15_io_x_paa),
    .io_x_eff(package_Anon_15_io_x_eff),
    .io_x_c(package_Anon_15_io_x_c),
    .io_y_ppn(package_Anon_15_io_y_ppn),
    .io_y_u(package_Anon_15_io_y_u),
    .io_y_ae(package_Anon_15_io_y_ae),
    .io_y_sw(package_Anon_15_io_y_sw),
    .io_y_sx(package_Anon_15_io_y_sx),
    .io_y_sr(package_Anon_15_io_y_sr),
    .io_y_pw(package_Anon_15_io_y_pw),
    .io_y_px(package_Anon_15_io_y_px),
    .io_y_pr(package_Anon_15_io_y_pr),
    .io_y_pal(package_Anon_15_io_y_pal),
    .io_y_paa(package_Anon_15_io_y_paa),
    .io_y_eff(package_Anon_15_io_y_eff),
    .io_y_c(package_Anon_15_io_y_c)
  );
  package_Anon_46 package_Anon_16 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_16_io_x_ppn),
    .io_x_u(package_Anon_16_io_x_u),
    .io_x_ae(package_Anon_16_io_x_ae),
    .io_x_sw(package_Anon_16_io_x_sw),
    .io_x_sx(package_Anon_16_io_x_sx),
    .io_x_sr(package_Anon_16_io_x_sr),
    .io_x_pw(package_Anon_16_io_x_pw),
    .io_x_px(package_Anon_16_io_x_px),
    .io_x_pr(package_Anon_16_io_x_pr),
    .io_x_pal(package_Anon_16_io_x_pal),
    .io_x_paa(package_Anon_16_io_x_paa),
    .io_x_eff(package_Anon_16_io_x_eff),
    .io_x_c(package_Anon_16_io_x_c),
    .io_y_ppn(package_Anon_16_io_y_ppn),
    .io_y_u(package_Anon_16_io_y_u),
    .io_y_ae(package_Anon_16_io_y_ae),
    .io_y_sw(package_Anon_16_io_y_sw),
    .io_y_sx(package_Anon_16_io_y_sx),
    .io_y_sr(package_Anon_16_io_y_sr),
    .io_y_pw(package_Anon_16_io_y_pw),
    .io_y_px(package_Anon_16_io_y_px),
    .io_y_pr(package_Anon_16_io_y_pr),
    .io_y_pal(package_Anon_16_io_y_pal),
    .io_y_paa(package_Anon_16_io_y_paa),
    .io_y_eff(package_Anon_16_io_y_eff),
    .io_y_c(package_Anon_16_io_y_c)
  );
  package_Anon_46 package_Anon_17 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_17_io_x_ppn),
    .io_x_u(package_Anon_17_io_x_u),
    .io_x_ae(package_Anon_17_io_x_ae),
    .io_x_sw(package_Anon_17_io_x_sw),
    .io_x_sx(package_Anon_17_io_x_sx),
    .io_x_sr(package_Anon_17_io_x_sr),
    .io_x_pw(package_Anon_17_io_x_pw),
    .io_x_px(package_Anon_17_io_x_px),
    .io_x_pr(package_Anon_17_io_x_pr),
    .io_x_pal(package_Anon_17_io_x_pal),
    .io_x_paa(package_Anon_17_io_x_paa),
    .io_x_eff(package_Anon_17_io_x_eff),
    .io_x_c(package_Anon_17_io_x_c),
    .io_y_ppn(package_Anon_17_io_y_ppn),
    .io_y_u(package_Anon_17_io_y_u),
    .io_y_ae(package_Anon_17_io_y_ae),
    .io_y_sw(package_Anon_17_io_y_sw),
    .io_y_sx(package_Anon_17_io_y_sx),
    .io_y_sr(package_Anon_17_io_y_sr),
    .io_y_pw(package_Anon_17_io_y_pw),
    .io_y_px(package_Anon_17_io_y_px),
    .io_y_pr(package_Anon_17_io_y_pr),
    .io_y_pal(package_Anon_17_io_y_pal),
    .io_y_paa(package_Anon_17_io_y_paa),
    .io_y_eff(package_Anon_17_io_y_eff),
    .io_y_c(package_Anon_17_io_y_c)
  );
  package_Anon_46 package_Anon_18 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_18_io_x_ppn),
    .io_x_u(package_Anon_18_io_x_u),
    .io_x_ae(package_Anon_18_io_x_ae),
    .io_x_sw(package_Anon_18_io_x_sw),
    .io_x_sx(package_Anon_18_io_x_sx),
    .io_x_sr(package_Anon_18_io_x_sr),
    .io_x_pw(package_Anon_18_io_x_pw),
    .io_x_px(package_Anon_18_io_x_px),
    .io_x_pr(package_Anon_18_io_x_pr),
    .io_x_pal(package_Anon_18_io_x_pal),
    .io_x_paa(package_Anon_18_io_x_paa),
    .io_x_eff(package_Anon_18_io_x_eff),
    .io_x_c(package_Anon_18_io_x_c),
    .io_y_ppn(package_Anon_18_io_y_ppn),
    .io_y_u(package_Anon_18_io_y_u),
    .io_y_ae(package_Anon_18_io_y_ae),
    .io_y_sw(package_Anon_18_io_y_sw),
    .io_y_sx(package_Anon_18_io_y_sx),
    .io_y_sr(package_Anon_18_io_y_sr),
    .io_y_pw(package_Anon_18_io_y_pw),
    .io_y_px(package_Anon_18_io_y_px),
    .io_y_pr(package_Anon_18_io_y_pr),
    .io_y_pal(package_Anon_18_io_y_pal),
    .io_y_paa(package_Anon_18_io_y_paa),
    .io_y_eff(package_Anon_18_io_y_eff),
    .io_y_c(package_Anon_18_io_y_c)
  );
  package_Anon_46 package_Anon_19 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_19_io_x_ppn),
    .io_x_u(package_Anon_19_io_x_u),
    .io_x_ae(package_Anon_19_io_x_ae),
    .io_x_sw(package_Anon_19_io_x_sw),
    .io_x_sx(package_Anon_19_io_x_sx),
    .io_x_sr(package_Anon_19_io_x_sr),
    .io_x_pw(package_Anon_19_io_x_pw),
    .io_x_px(package_Anon_19_io_x_px),
    .io_x_pr(package_Anon_19_io_x_pr),
    .io_x_pal(package_Anon_19_io_x_pal),
    .io_x_paa(package_Anon_19_io_x_paa),
    .io_x_eff(package_Anon_19_io_x_eff),
    .io_x_c(package_Anon_19_io_x_c),
    .io_y_ppn(package_Anon_19_io_y_ppn),
    .io_y_u(package_Anon_19_io_y_u),
    .io_y_ae(package_Anon_19_io_y_ae),
    .io_y_sw(package_Anon_19_io_y_sw),
    .io_y_sx(package_Anon_19_io_y_sx),
    .io_y_sr(package_Anon_19_io_y_sr),
    .io_y_pw(package_Anon_19_io_y_pw),
    .io_y_px(package_Anon_19_io_y_px),
    .io_y_pr(package_Anon_19_io_y_pr),
    .io_y_pal(package_Anon_19_io_y_pal),
    .io_y_paa(package_Anon_19_io_y_paa),
    .io_y_eff(package_Anon_19_io_y_eff),
    .io_y_c(package_Anon_19_io_y_c)
  );
  package_Anon_46 package_Anon_20 ( // @[package.scala 213:21]
    .io_x_ppn(package_Anon_20_io_x_ppn),
    .io_x_u(package_Anon_20_io_x_u),
    .io_x_ae(package_Anon_20_io_x_ae),
    .io_x_sw(package_Anon_20_io_x_sw),
    .io_x_sx(package_Anon_20_io_x_sx),
    .io_x_sr(package_Anon_20_io_x_sr),
    .io_x_pw(package_Anon_20_io_x_pw),
    .io_x_px(package_Anon_20_io_x_px),
    .io_x_pr(package_Anon_20_io_x_pr),
    .io_x_pal(package_Anon_20_io_x_pal),
    .io_x_paa(package_Anon_20_io_x_paa),
    .io_x_eff(package_Anon_20_io_x_eff),
    .io_x_c(package_Anon_20_io_x_c),
    .io_y_ppn(package_Anon_20_io_y_ppn),
    .io_y_u(package_Anon_20_io_y_u),
    .io_y_ae(package_Anon_20_io_y_ae),
    .io_y_sw(package_Anon_20_io_y_sw),
    .io_y_sx(package_Anon_20_io_y_sx),
    .io_y_sr(package_Anon_20_io_y_sr),
    .io_y_pw(package_Anon_20_io_y_pw),
    .io_y_px(package_Anon_20_io_y_px),
    .io_y_pr(package_Anon_20_io_y_pr),
    .io_y_pal(package_Anon_20_io_y_pal),
    .io_y_paa(package_Anon_20_io_y_paa),
    .io_y_eff(package_Anon_20_io_y_eff),
    .io_y_c(package_Anon_20_io_y_c)
  );
  assign io_req_0_ready = 1'h1; // @[tlb.scala 290:24]
  assign io_miss_rdy = state == 2'h0; // @[tlb.scala 288:24]
  assign io_resp_0_miss = io_ptw_resp_valid | tlb_miss_0 | multipleHits_0; // @[tlb.scala 303:50]
  assign io_resp_0_paddr = {ppn_0,io_req_0_bits_vaddr[11:0]}; // @[Cat.scala 29:58]
  assign io_resp_0_pf_ld = bad_va_0 & cmd_read_0 | |_T_1553; // @[tlb.scala 291:54]
  assign io_resp_0_pf_st = bad_va_0 & cmd_write_0 | |_T_1557; // @[tlb.scala 292:61]
  assign io_resp_0_pf_inst = bad_va_0 | |_T_1560; // @[tlb.scala 293:37]
  assign io_resp_0_ae_ld = |_T_1563; // @[tlb.scala 294:54]
  assign io_resp_0_ae_st = |_T_1565; // @[tlb.scala 295:54]
  assign io_resp_0_ae_inst = |_T_1568; // @[tlb.scala 296:54]
  assign io_resp_0_ma_ld = |_T_1570; // @[tlb.scala 297:54]
  assign io_resp_0_ma_st = |_T_1572; // @[tlb.scala 298:54]
  assign io_resp_0_ma_inst = 1'h0; // @[tlb.scala 299:24]
  assign io_resp_0_cacheable = |_T_1574; // @[tlb.scala 300:55]
  assign io_resp_0_must_alloc = |_T_1576; // @[tlb.scala 301:64]
  assign io_resp_0_prefetchable = |_T_1578; // @[tlb.scala 302:66]
  assign io_ptw_req_valid = state == 2'h1; // @[tlb.scala 307:29]
  assign io_ptw_req_bits_valid = ~io_kill; // @[tlb.scala 308:28]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[tlb.scala 309:29]
  assign package_Anon_io_x_ppn = special_entry_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_u = special_entry_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_ae = special_entry_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_sw = special_entry_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_sx = special_entry_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_sr = special_entry_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_pw = special_entry_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_px = special_entry_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_pr = special_entry_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_pal = special_entry_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_paa = special_entry_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_eff = special_entry_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_io_x_c = special_entry_data_0[1]; // @[tlb.scala 58:79]
  assign pmp_0_io_prv = io_ptw_resp_valid | io_req_0_bits_passthrough ? 2'h1 : io_ptw_status_dprv; // @[tlb.scala 155:25]
  assign pmp_0_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[tlb.scala 154:19]
  assign pmp_0_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[tlb.scala 154:19]
  assign pmp_0_io_addr = mpu_physaddr_0[31:0]; // @[tlb.scala 152:20]
  assign pmp_0_io_size = io_req_0_bits_size; // @[tlb.scala 153:20]
  assign package_Anon_1_io_x_ppn = _GEN_11[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_u = _GEN_11[13]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_ae = _GEN_11[11]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_sw = _GEN_11[10]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_sx = _GEN_11[9]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_sr = _GEN_11[8]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_pw = _GEN_11[7]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_px = _GEN_11[6]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_pr = _GEN_11[5]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_pal = _GEN_11[4]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_paa = _GEN_11[3]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_eff = _GEN_11[2]; // @[tlb.scala 58:79]
  assign package_Anon_1_io_x_c = _GEN_11[1]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_ppn = _GEN_15[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_u = _GEN_15[13]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_ae = _GEN_15[11]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_sw = _GEN_15[10]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_sx = _GEN_15[9]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_sr = _GEN_15[8]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_pw = _GEN_15[7]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_px = _GEN_15[6]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_pr = _GEN_15[5]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_pal = _GEN_15[4]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_paa = _GEN_15[3]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_eff = _GEN_15[2]; // @[tlb.scala 58:79]
  assign package_Anon_2_io_x_c = _GEN_15[1]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_u = superpage_entries_0_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_ae = superpage_entries_0_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_sw = superpage_entries_0_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_sx = superpage_entries_0_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_sr = superpage_entries_0_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_pw = superpage_entries_0_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_px = superpage_entries_0_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_pr = superpage_entries_0_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_pal = superpage_entries_0_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_paa = superpage_entries_0_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_eff = superpage_entries_0_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_3_io_x_c = superpage_entries_0_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_u = superpage_entries_1_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_ae = superpage_entries_1_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_sw = superpage_entries_1_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_sx = superpage_entries_1_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_sr = superpage_entries_1_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_pw = superpage_entries_1_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_px = superpage_entries_1_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_pr = superpage_entries_1_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_pal = superpage_entries_1_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_paa = superpage_entries_1_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_eff = superpage_entries_1_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_4_io_x_c = superpage_entries_1_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_u = superpage_entries_2_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_ae = superpage_entries_2_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_sw = superpage_entries_2_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_sx = superpage_entries_2_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_sr = superpage_entries_2_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_pw = superpage_entries_2_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_px = superpage_entries_2_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_pr = superpage_entries_2_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_pal = superpage_entries_2_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_paa = superpage_entries_2_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_eff = superpage_entries_2_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_5_io_x_c = superpage_entries_2_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_u = superpage_entries_3_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_ae = superpage_entries_3_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_sw = superpage_entries_3_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_sx = superpage_entries_3_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_sr = superpage_entries_3_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_pw = superpage_entries_3_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_px = superpage_entries_3_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_pr = superpage_entries_3_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_pal = superpage_entries_3_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_paa = superpage_entries_3_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_eff = superpage_entries_3_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_6_io_x_c = superpage_entries_3_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_ppn = special_entry_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_u = special_entry_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_ae = special_entry_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_sw = special_entry_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_sx = special_entry_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_sr = special_entry_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_pw = special_entry_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_px = special_entry_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_pr = special_entry_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_pal = special_entry_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_paa = special_entry_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_eff = special_entry_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_7_io_x_c = special_entry_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_ppn = _GEN_11[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_u = _GEN_11[13]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_ae = _GEN_11[11]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_sw = _GEN_11[10]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_sx = _GEN_11[9]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_sr = _GEN_11[8]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_pw = _GEN_11[7]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_px = _GEN_11[6]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_pr = _GEN_11[5]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_pal = _GEN_11[4]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_paa = _GEN_11[3]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_eff = _GEN_11[2]; // @[tlb.scala 58:79]
  assign package_Anon_8_io_x_c = _GEN_11[1]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_ppn = _GEN_15[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_u = _GEN_15[13]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_ae = _GEN_15[11]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_sw = _GEN_15[10]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_sx = _GEN_15[9]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_sr = _GEN_15[8]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_pw = _GEN_15[7]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_px = _GEN_15[6]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_pr = _GEN_15[5]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_pal = _GEN_15[4]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_paa = _GEN_15[3]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_eff = _GEN_15[2]; // @[tlb.scala 58:79]
  assign package_Anon_9_io_x_c = _GEN_15[1]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_u = superpage_entries_0_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_ae = superpage_entries_0_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_sw = superpage_entries_0_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_sx = superpage_entries_0_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_sr = superpage_entries_0_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_pw = superpage_entries_0_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_px = superpage_entries_0_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_pr = superpage_entries_0_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_pal = superpage_entries_0_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_paa = superpage_entries_0_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_eff = superpage_entries_0_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_10_io_x_c = superpage_entries_0_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_u = superpage_entries_1_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_ae = superpage_entries_1_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_sw = superpage_entries_1_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_sx = superpage_entries_1_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_sr = superpage_entries_1_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_pw = superpage_entries_1_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_px = superpage_entries_1_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_pr = superpage_entries_1_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_pal = superpage_entries_1_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_paa = superpage_entries_1_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_eff = superpage_entries_1_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_11_io_x_c = superpage_entries_1_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_u = superpage_entries_2_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_ae = superpage_entries_2_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_sw = superpage_entries_2_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_sx = superpage_entries_2_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_sr = superpage_entries_2_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_pw = superpage_entries_2_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_px = superpage_entries_2_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_pr = superpage_entries_2_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_pal = superpage_entries_2_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_paa = superpage_entries_2_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_eff = superpage_entries_2_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_12_io_x_c = superpage_entries_2_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_u = superpage_entries_3_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_ae = superpage_entries_3_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_sw = superpage_entries_3_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_sx = superpage_entries_3_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_sr = superpage_entries_3_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_pw = superpage_entries_3_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_px = superpage_entries_3_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_pr = superpage_entries_3_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_pal = superpage_entries_3_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_paa = superpage_entries_3_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_eff = superpage_entries_3_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_13_io_x_c = superpage_entries_3_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_ppn = special_entry_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_u = special_entry_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_ae = special_entry_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_sw = special_entry_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_sx = special_entry_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_sr = special_entry_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_pw = special_entry_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_px = special_entry_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_pr = special_entry_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_pal = special_entry_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_paa = special_entry_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_eff = special_entry_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_14_io_x_c = special_entry_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_ppn = _GEN_11[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_u = _GEN_11[13]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_ae = _GEN_11[11]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_sw = _GEN_11[10]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_sx = _GEN_11[9]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_sr = _GEN_11[8]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_pw = _GEN_11[7]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_px = _GEN_11[6]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_pr = _GEN_11[5]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_pal = _GEN_11[4]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_paa = _GEN_11[3]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_eff = _GEN_11[2]; // @[tlb.scala 58:79]
  assign package_Anon_15_io_x_c = _GEN_11[1]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_ppn = _GEN_15[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_u = _GEN_15[13]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_ae = _GEN_15[11]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_sw = _GEN_15[10]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_sx = _GEN_15[9]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_sr = _GEN_15[8]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_pw = _GEN_15[7]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_px = _GEN_15[6]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_pr = _GEN_15[5]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_pal = _GEN_15[4]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_paa = _GEN_15[3]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_eff = _GEN_15[2]; // @[tlb.scala 58:79]
  assign package_Anon_16_io_x_c = _GEN_15[1]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_u = superpage_entries_0_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_ae = superpage_entries_0_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_sw = superpage_entries_0_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_sx = superpage_entries_0_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_sr = superpage_entries_0_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_pw = superpage_entries_0_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_px = superpage_entries_0_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_pr = superpage_entries_0_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_pal = superpage_entries_0_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_paa = superpage_entries_0_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_eff = superpage_entries_0_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_17_io_x_c = superpage_entries_0_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_u = superpage_entries_1_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_ae = superpage_entries_1_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_sw = superpage_entries_1_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_sx = superpage_entries_1_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_sr = superpage_entries_1_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_pw = superpage_entries_1_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_px = superpage_entries_1_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_pr = superpage_entries_1_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_pal = superpage_entries_1_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_paa = superpage_entries_1_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_eff = superpage_entries_1_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_18_io_x_c = superpage_entries_1_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_u = superpage_entries_2_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_ae = superpage_entries_2_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_sw = superpage_entries_2_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_sx = superpage_entries_2_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_sr = superpage_entries_2_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_pw = superpage_entries_2_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_px = superpage_entries_2_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_pr = superpage_entries_2_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_pal = superpage_entries_2_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_paa = superpage_entries_2_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_eff = superpage_entries_2_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_19_io_x_c = superpage_entries_2_data_0[1]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_u = superpage_entries_3_data_0[13]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_ae = superpage_entries_3_data_0[11]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_sw = superpage_entries_3_data_0[10]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_sx = superpage_entries_3_data_0[9]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_sr = superpage_entries_3_data_0[8]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_pw = superpage_entries_3_data_0[7]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_px = superpage_entries_3_data_0[6]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_pr = superpage_entries_3_data_0[5]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_pal = superpage_entries_3_data_0[4]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_paa = superpage_entries_3_data_0[3]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_eff = superpage_entries_3_data_0[2]; // @[tlb.scala 58:79]
  assign package_Anon_20_io_x_c = superpage_entries_3_data_0[1]; // @[tlb.scala 58:79]
  always @(posedge clock) begin
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (~_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_0_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (~_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_0_data_0 <= _GEN_40;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (~_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_0_data_1 <= _GEN_41;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (~_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_0_data_2 <= _GEN_42;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (~_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_0_data_3 <= _GEN_43;
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_0_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_388[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_0_valid_0 <= _GEN_232;
        end else begin
          sectored_entries_0_valid_0 <= _GEN_228;
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_244;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_0_valid_0 <= _GEN_92;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_0_valid_1 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_388[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_0_valid_1 <= _GEN_233;
        end else begin
          sectored_entries_0_valid_1 <= _GEN_229;
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_245;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_0_valid_1 <= _GEN_93;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_0_valid_2 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_388[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_0_valid_2 <= _GEN_234;
        end else begin
          sectored_entries_0_valid_2 <= _GEN_230;
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_246;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_0_valid_2 <= _GEN_94;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_0_valid_3 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_388[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_0_valid_3 <= _GEN_235;
        end else begin
          sectored_entries_0_valid_3 <= _GEN_231;
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_247;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_0_valid_3 <= _GEN_95;
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_1_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_1_data_0 <= _GEN_62;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_1_data_1 <= _GEN_63;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_1_data_2 <= _GEN_64;
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[tlb.scala 198:58]
          if (_T_924) begin // @[tlb.scala 204:74]
            sectored_entries_1_data_3 <= _GEN_65;
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_1_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_395[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_1_valid_0 <= _GEN_260;
        end else begin
          sectored_entries_1_valid_0 <= _GEN_256;
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_272;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_1_valid_0 <= _GEN_102;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_1_valid_1 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_395[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_1_valid_1 <= _GEN_261;
        end else begin
          sectored_entries_1_valid_1 <= _GEN_257;
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_273;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_1_valid_1 <= _GEN_103;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_1_valid_2 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_395[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_1_valid_2 <= _GEN_262;
        end else begin
          sectored_entries_1_valid_2 <= _GEN_258;
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_274;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_1_valid_2 <= _GEN_104;
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      sectored_entries_1_valid_3 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_395[26:18] == 9'h0) begin // @[tlb.scala 107:73]
          sectored_entries_1_valid_3 <= _GEN_263;
        end else begin
          sectored_entries_1_valid_3 <= _GEN_259;
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_275;
      end
    end else if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        sectored_entries_1_valid_3 <= _GEN_105;
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h0) begin // @[tlb.scala 199:91]
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[tlb.scala 91:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h0) begin // @[tlb.scala 199:91]
            superpage_entries_0_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h0) begin // @[tlb.scala 199:91]
            superpage_entries_0_data_0 <= _T_858; // @[tlb.scala 95:17]
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      superpage_entries_0_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (superpage_hits_0_0) begin // @[tlb.scala 101:26]
          superpage_entries_0_valid_0 <= 1'h0; // @[tlb.scala 98:40]
        end else begin
          superpage_entries_0_valid_0 <= _GEN_158;
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_282;
      end
    end else begin
      superpage_entries_0_valid_0 <= _GEN_158;
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h1) begin // @[tlb.scala 199:91]
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[tlb.scala 91:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h1) begin // @[tlb.scala 199:91]
            superpage_entries_1_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h1) begin // @[tlb.scala 199:91]
            superpage_entries_1_data_0 <= _T_858; // @[tlb.scala 95:17]
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      superpage_entries_1_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (superpage_hits_0_1) begin // @[tlb.scala 101:26]
          superpage_entries_1_valid_0 <= 1'h0; // @[tlb.scala 98:40]
        end else begin
          superpage_entries_1_valid_0 <= _GEN_162;
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_286;
      end
    end else begin
      superpage_entries_1_valid_0 <= _GEN_162;
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h2) begin // @[tlb.scala 199:91]
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[tlb.scala 91:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h2) begin // @[tlb.scala 199:91]
            superpage_entries_2_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h2) begin // @[tlb.scala 199:91]
            superpage_entries_2_data_0 <= _T_858; // @[tlb.scala 95:17]
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      superpage_entries_2_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (superpage_hits_0_2) begin // @[tlb.scala 101:26]
          superpage_entries_2_valid_0 <= 1'h0; // @[tlb.scala 98:40]
        end else begin
          superpage_entries_2_valid_0 <= _GEN_166;
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_290;
      end
    end else begin
      superpage_entries_2_valid_0 <= _GEN_166;
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h3) begin // @[tlb.scala 199:91]
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[tlb.scala 91:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h3) begin // @[tlb.scala 199:91]
            superpage_entries_3_tag <= r_refill_tag; // @[tlb.scala 90:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[tlb.scala 196:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[tlb.scala 198:58]
          if (r_superpage_repl_addr == 2'h3) begin // @[tlb.scala 199:91]
            superpage_entries_3_data_0 <= _T_858; // @[tlb.scala 95:17]
          end
        end
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      superpage_entries_3_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (superpage_hits_0_3) begin // @[tlb.scala 101:26]
          superpage_entries_3_valid_0 <= 1'h0; // @[tlb.scala 98:40]
        end else begin
          superpage_entries_3_valid_0 <= _GEN_170;
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_294;
      end
    end else begin
      superpage_entries_3_valid_0 <= _GEN_170;
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (~io_ptw_resp_bits_homogeneous) begin // @[tlb.scala 196:70]
        special_entry_level <= io_ptw_resp_bits_level; // @[tlb.scala 91:18]
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (~io_ptw_resp_bits_homogeneous) begin // @[tlb.scala 196:70]
        special_entry_tag <= r_refill_tag; // @[tlb.scala 90:16]
      end
    end
    if (io_ptw_resp_valid & ~invalidate_refill) begin // @[tlb.scala 177:42]
      if (~io_ptw_resp_bits_homogeneous) begin // @[tlb.scala 196:70]
        special_entry_data_0 <= _T_858; // @[tlb.scala 95:17]
      end
    end
    if (multipleHits_0 | reset) begin // @[tlb.scala 346:45]
      special_entry_valid_0 <= 1'h0; // @[tlb.scala 98:40]
    end else if (io_sfence_valid) begin // @[tlb.scala 336:19]
      if (io_sfence_bits_rs1) begin // @[tlb.scala 340:37]
        if (_T_605) begin // @[tlb.scala 101:26]
          special_entry_valid_0 <= 1'h0; // @[tlb.scala 98:40]
        end else begin
          special_entry_valid_0 <= _GEN_154;
        end
      end else begin
        special_entry_valid_0 <= _GEN_298;
      end
    end else begin
      special_entry_valid_0 <= _GEN_154;
    end
    if (reset) begin // @[tlb.scala 129:22]
      state <= 2'h0; // @[tlb.scala 129:22]
    end else if (io_ptw_resp_valid) begin // @[tlb.scala 332:30]
      state <= 2'h0; // @[tlb.scala 333:13]
    end else if (state == 2'h2 & io_sfence_valid) begin // @[tlb.scala 329:39]
      state <= 2'h3; // @[tlb.scala 330:13]
    end else if (_T_6) begin // @[tlb.scala 324:32]
      state <= _GEN_220;
    end else begin
      state <= _GEN_212;
    end
    if (_T_1587 & tlb_miss_0 & _T_1551) begin // @[tlb.scala 314:67]
      r_refill_tag <= vpn_0; // @[tlb.scala 316:22]
    end
    if (_T_1587 & tlb_miss_0 & _T_1551) begin // @[tlb.scala 314:67]
      if (&_T_1609) begin // @[tlb.scala 353:8]
        r_superpage_repl_addr <= _T_1605[1:0];
      end else if (_T_1611[0]) begin // @[Mux.scala 47:69]
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_1611[1]) begin // @[Mux.scala 47:69]
        r_superpage_repl_addr <= 2'h1;
      end else begin
        r_superpage_repl_addr <= _T_1616;
      end
    end
    if (_T_1587 & tlb_miss_0 & _T_1551) begin // @[tlb.scala 314:67]
      if (&_T_1635) begin // @[tlb.scala 353:8]
        r_sectored_repl_addr <= _T_1627[0];
      end else if (_T_1637[0]) begin // @[Mux.scala 47:69]
        r_sectored_repl_addr <= 1'h0;
      end else begin
        r_sectored_repl_addr <= 1'h1;
      end
    end
    if (_T_1587 & tlb_miss_0 & _T_1551) begin // @[tlb.scala 314:67]
      r_sectored_hit_addr <= _T_1463[1]; // @[tlb.scala 320:31]
    end
    if (_T_1587 & tlb_miss_0 & _T_1551) begin // @[tlb.scala 314:67]
      r_sectored_hit <= _T_1462; // @[tlb.scala 321:31]
    end
    if (io_req_0_valid & vm_enabled_0) begin // @[tlb.scala 275:45]
      if (_T_1462) begin // @[tlb.scala 276:33]
        _T_1459 <= _T_1473[1]; // @[Replacement.scala 44:15]
      end
    end
    if (io_req_0_valid & vm_enabled_0) begin // @[tlb.scala 275:45]
      if (_T_1478) begin // @[tlb.scala 277:36]
        _T_1460 <= _T_1505[3:1]; // @[Replacement.scala 44:15]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn_0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at tlb.scala:338 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn(w))\n"
            ); // @[tlb.scala 338:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn_0 | reset)) begin
          $fatal; // @[tlb.scala 338:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_19[26:0];
  _RAND_20 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_20[33:0];
  _RAND_21 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_23[26:0];
  _RAND_24 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_24[33:0];
  _RAND_25 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_27[26:0];
  _RAND_28 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_28[33:0];
  _RAND_29 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_31[26:0];
  _RAND_32 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_32[33:0];
  _RAND_33 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  special_entry_level = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  special_entry_tag = _RAND_35[26:0];
  _RAND_36 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_36[33:0];
  _RAND_37 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  state = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  r_refill_tag = _RAND_39[26:0];
  _RAND_40 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_sectored_hit = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_1459 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_1460 = _RAND_45[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
