module Control(
  input  [6:0] io_opcode,
  output       io_itype,
  output       io_aluop,
  output       io_xsrc,
  output       io_ysrc,
  output       io_branch,
  output       io_jal,
  output       io_jalr,
  output       io_plus4,
  output       io_resultselect,
  output [1:0] io_memop,
  output       io_toreg,
  output       io_regwrite
);
  wire  _T_1 = 7'h33 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_3 = 7'h13 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_5 = 7'h3 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_7 = 7'h23 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_9 = 7'h63 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_11 = 7'h37 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_13 = 7'h17 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_15 = 7'h6f == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_17 = 7'h67 == io_opcode; // @[Lookup.scala 31:38]
  wire  _T_37 = _T_11 ? 1'h0 : _T_13 | (_T_15 | _T_17); // @[Lookup.scala 33:37]
  wire  _T_38 = _T_9 ? 1'h0 : _T_37; // @[Lookup.scala 33:37]
  wire  _T_39 = _T_7 ? 1'h0 : _T_38; // @[Lookup.scala 33:37]
  wire  _T_40 = _T_5 ? 1'h0 : _T_39; // @[Lookup.scala 33:37]
  wire  _T_41 = _T_3 ? 1'h0 : _T_40; // @[Lookup.scala 33:37]
  wire  _T_45 = _T_11 ? 1'h0 : _T_13; // @[Lookup.scala 33:37]
  wire  _T_46 = _T_9 ? 1'h0 : _T_45; // @[Lookup.scala 33:37]
  wire  _T_55 = _T_7 ? 1'h0 : _T_9; // @[Lookup.scala 33:37]
  wire  _T_56 = _T_5 ? 1'h0 : _T_55; // @[Lookup.scala 33:37]
  wire  _T_57 = _T_3 ? 1'h0 : _T_56; // @[Lookup.scala 33:37]
  wire  _T_60 = _T_13 ? 1'h0 : _T_15; // @[Lookup.scala 33:37]
  wire  _T_61 = _T_11 ? 1'h0 : _T_60; // @[Lookup.scala 33:37]
  wire  _T_62 = _T_9 ? 1'h0 : _T_61; // @[Lookup.scala 33:37]
  wire  _T_63 = _T_7 ? 1'h0 : _T_62; // @[Lookup.scala 33:37]
  wire  _T_64 = _T_5 ? 1'h0 : _T_63; // @[Lookup.scala 33:37]
  wire  _T_65 = _T_3 ? 1'h0 : _T_64; // @[Lookup.scala 33:37]
  wire  _T_67 = _T_15 ? 1'h0 : _T_17; // @[Lookup.scala 33:37]
  wire  _T_68 = _T_13 ? 1'h0 : _T_67; // @[Lookup.scala 33:37]
  wire  _T_69 = _T_11 ? 1'h0 : _T_68; // @[Lookup.scala 33:37]
  wire  _T_70 = _T_9 ? 1'h0 : _T_69; // @[Lookup.scala 33:37]
  wire  _T_71 = _T_7 ? 1'h0 : _T_70; // @[Lookup.scala 33:37]
  wire  _T_72 = _T_5 ? 1'h0 : _T_71; // @[Lookup.scala 33:37]
  wire  _T_73 = _T_3 ? 1'h0 : _T_72; // @[Lookup.scala 33:37]
  wire  _T_76 = _T_13 ? 1'h0 : _T_15 | _T_17; // @[Lookup.scala 33:37]
  wire  _T_77 = _T_11 ? 1'h0 : _T_76; // @[Lookup.scala 33:37]
  wire  _T_78 = _T_9 ? 1'h0 : _T_77; // @[Lookup.scala 33:37]
  wire  _T_79 = _T_7 ? 1'h0 : _T_78; // @[Lookup.scala 33:37]
  wire  _T_80 = _T_5 ? 1'h0 : _T_79; // @[Lookup.scala 33:37]
  wire  _T_81 = _T_3 ? 1'h0 : _T_80; // @[Lookup.scala 33:37]
  wire  _T_86 = _T_9 ? 1'h0 : _T_11; // @[Lookup.scala 33:37]
  wire  _T_87 = _T_7 ? 1'h0 : _T_86; // @[Lookup.scala 33:37]
  wire  _T_88 = _T_5 ? 1'h0 : _T_87; // @[Lookup.scala 33:37]
  wire  _T_89 = _T_3 ? 1'h0 : _T_88; // @[Lookup.scala 33:37]
  wire [1:0] _T_95 = _T_7 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_96 = _T_5 ? 2'h2 : _T_95; // @[Lookup.scala 33:37]
  wire [1:0] _T_97 = _T_3 ? 2'h0 : _T_96; // @[Lookup.scala 33:37]
  wire  _T_105 = _T_3 ? 1'h0 : _T_5; // @[Lookup.scala 33:37]
  wire  _T_110 = _T_9 ? 1'h0 : _T_11 | (_T_13 | (_T_15 | _T_17)); // @[Lookup.scala 33:37]
  wire  _T_111 = _T_7 ? 1'h0 : _T_110; // @[Lookup.scala 33:37]
  assign io_itype = _T_1 ? 1'h0 : _T_3; // @[Lookup.scala 33:37]
  assign io_aluop = _T_1 | _T_3; // @[Lookup.scala 33:37]
  assign io_xsrc = _T_1 ? 1'h0 : _T_41; // @[Lookup.scala 33:37]
  assign io_ysrc = _T_1 ? 1'h0 : _T_3 | (_T_5 | (_T_7 | _T_46)); // @[Lookup.scala 33:37]
  assign io_branch = _T_1 ? 1'h0 : _T_57; // @[Lookup.scala 33:37]
  assign io_jal = _T_1 ? 1'h0 : _T_65; // @[Lookup.scala 33:37]
  assign io_jalr = _T_1 ? 1'h0 : _T_73; // @[Lookup.scala 33:37]
  assign io_plus4 = _T_1 ? 1'h0 : _T_81; // @[Lookup.scala 33:37]
  assign io_resultselect = _T_1 ? 1'h0 : _T_89; // @[Lookup.scala 33:37]
  assign io_memop = _T_1 ? 2'h0 : _T_97; // @[Lookup.scala 33:37]
  assign io_toreg = _T_1 ? 1'h0 : _T_105; // @[Lookup.scala 33:37]
  assign io_regwrite = _T_1 | (_T_3 | (_T_5 | _T_111)); // @[Lookup.scala 33:37]
endmodule
module RegisterFile(
  input         clock,
  input  [4:0]  io_readreg1,
  input  [4:0]  io_readreg2,
  input  [4:0]  io_writereg,
  input  [31:0] io_writedata,
  input         io_wen,
  output [31:0] io_readdata1,
  output [31:0] io_readdata2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[register-file.scala 52:17]
  reg [31:0] regs_1; // @[register-file.scala 52:17]
  reg [31:0] regs_2; // @[register-file.scala 52:17]
  reg [31:0] regs_3; // @[register-file.scala 52:17]
  reg [31:0] regs_4; // @[register-file.scala 52:17]
  reg [31:0] regs_5; // @[register-file.scala 52:17]
  reg [31:0] regs_6; // @[register-file.scala 52:17]
  reg [31:0] regs_7; // @[register-file.scala 52:17]
  reg [31:0] regs_8; // @[register-file.scala 52:17]
  reg [31:0] regs_9; // @[register-file.scala 52:17]
  reg [31:0] regs_10; // @[register-file.scala 52:17]
  reg [31:0] regs_11; // @[register-file.scala 52:17]
  reg [31:0] regs_12; // @[register-file.scala 52:17]
  reg [31:0] regs_13; // @[register-file.scala 52:17]
  reg [31:0] regs_14; // @[register-file.scala 52:17]
  reg [31:0] regs_15; // @[register-file.scala 52:17]
  reg [31:0] regs_16; // @[register-file.scala 52:17]
  reg [31:0] regs_17; // @[register-file.scala 52:17]
  reg [31:0] regs_18; // @[register-file.scala 52:17]
  reg [31:0] regs_19; // @[register-file.scala 52:17]
  reg [31:0] regs_20; // @[register-file.scala 52:17]
  reg [31:0] regs_21; // @[register-file.scala 52:17]
  reg [31:0] regs_22; // @[register-file.scala 52:17]
  reg [31:0] regs_23; // @[register-file.scala 52:17]
  reg [31:0] regs_24; // @[register-file.scala 52:17]
  reg [31:0] regs_25; // @[register-file.scala 52:17]
  reg [31:0] regs_26; // @[register-file.scala 52:17]
  reg [31:0] regs_27; // @[register-file.scala 52:17]
  reg [31:0] regs_28; // @[register-file.scala 52:17]
  reg [31:0] regs_29; // @[register-file.scala 52:17]
  reg [31:0] regs_30; // @[register-file.scala 52:17]
  reg [31:0] regs_31; // @[register-file.scala 52:17]
  wire [31:0] _GEN_65 = 5'h1 == io_readreg1 ? regs_1 : regs_0; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_66 = 5'h2 == io_readreg1 ? regs_2 : _GEN_65; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_67 = 5'h3 == io_readreg1 ? regs_3 : _GEN_66; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_68 = 5'h4 == io_readreg1 ? regs_4 : _GEN_67; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_69 = 5'h5 == io_readreg1 ? regs_5 : _GEN_68; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_70 = 5'h6 == io_readreg1 ? regs_6 : _GEN_69; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_71 = 5'h7 == io_readreg1 ? regs_7 : _GEN_70; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_72 = 5'h8 == io_readreg1 ? regs_8 : _GEN_71; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_73 = 5'h9 == io_readreg1 ? regs_9 : _GEN_72; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_74 = 5'ha == io_readreg1 ? regs_10 : _GEN_73; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_75 = 5'hb == io_readreg1 ? regs_11 : _GEN_74; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_76 = 5'hc == io_readreg1 ? regs_12 : _GEN_75; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_77 = 5'hd == io_readreg1 ? regs_13 : _GEN_76; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_78 = 5'he == io_readreg1 ? regs_14 : _GEN_77; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_79 = 5'hf == io_readreg1 ? regs_15 : _GEN_78; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_80 = 5'h10 == io_readreg1 ? regs_16 : _GEN_79; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_81 = 5'h11 == io_readreg1 ? regs_17 : _GEN_80; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_82 = 5'h12 == io_readreg1 ? regs_18 : _GEN_81; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_83 = 5'h13 == io_readreg1 ? regs_19 : _GEN_82; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_84 = 5'h14 == io_readreg1 ? regs_20 : _GEN_83; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_85 = 5'h15 == io_readreg1 ? regs_21 : _GEN_84; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_86 = 5'h16 == io_readreg1 ? regs_22 : _GEN_85; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_87 = 5'h17 == io_readreg1 ? regs_23 : _GEN_86; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_88 = 5'h18 == io_readreg1 ? regs_24 : _GEN_87; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_89 = 5'h19 == io_readreg1 ? regs_25 : _GEN_88; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_90 = 5'h1a == io_readreg1 ? regs_26 : _GEN_89; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_91 = 5'h1b == io_readreg1 ? regs_27 : _GEN_90; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_92 = 5'h1c == io_readreg1 ? regs_28 : _GEN_91; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_93 = 5'h1d == io_readreg1 ? regs_29 : _GEN_92; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_94 = 5'h1e == io_readreg1 ? regs_30 : _GEN_93; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_95 = 5'h1f == io_readreg1 ? regs_31 : _GEN_94; // @[register-file.scala 61:{16,16}]
  wire [31:0] _GEN_97 = 5'h1 == io_readreg2 ? regs_1 : regs_0; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_98 = 5'h2 == io_readreg2 ? regs_2 : _GEN_97; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_99 = 5'h3 == io_readreg2 ? regs_3 : _GEN_98; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_100 = 5'h4 == io_readreg2 ? regs_4 : _GEN_99; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_101 = 5'h5 == io_readreg2 ? regs_5 : _GEN_100; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_102 = 5'h6 == io_readreg2 ? regs_6 : _GEN_101; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_103 = 5'h7 == io_readreg2 ? regs_7 : _GEN_102; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_104 = 5'h8 == io_readreg2 ? regs_8 : _GEN_103; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_105 = 5'h9 == io_readreg2 ? regs_9 : _GEN_104; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_106 = 5'ha == io_readreg2 ? regs_10 : _GEN_105; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_107 = 5'hb == io_readreg2 ? regs_11 : _GEN_106; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_108 = 5'hc == io_readreg2 ? regs_12 : _GEN_107; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_109 = 5'hd == io_readreg2 ? regs_13 : _GEN_108; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_110 = 5'he == io_readreg2 ? regs_14 : _GEN_109; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_111 = 5'hf == io_readreg2 ? regs_15 : _GEN_110; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_112 = 5'h10 == io_readreg2 ? regs_16 : _GEN_111; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_113 = 5'h11 == io_readreg2 ? regs_17 : _GEN_112; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_114 = 5'h12 == io_readreg2 ? regs_18 : _GEN_113; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_115 = 5'h13 == io_readreg2 ? regs_19 : _GEN_114; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_116 = 5'h14 == io_readreg2 ? regs_20 : _GEN_115; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_117 = 5'h15 == io_readreg2 ? regs_21 : _GEN_116; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_118 = 5'h16 == io_readreg2 ? regs_22 : _GEN_117; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_119 = 5'h17 == io_readreg2 ? regs_23 : _GEN_118; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_120 = 5'h18 == io_readreg2 ? regs_24 : _GEN_119; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_121 = 5'h19 == io_readreg2 ? regs_25 : _GEN_120; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_122 = 5'h1a == io_readreg2 ? regs_26 : _GEN_121; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_123 = 5'h1b == io_readreg2 ? regs_27 : _GEN_122; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_124 = 5'h1c == io_readreg2 ? regs_28 : _GEN_123; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_125 = 5'h1d == io_readreg2 ? regs_29 : _GEN_124; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_126 = 5'h1e == io_readreg2 ? regs_30 : _GEN_125; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_127 = 5'h1f == io_readreg2 ? regs_31 : _GEN_126; // @[register-file.scala 62:{16,16}]
  wire [31:0] _GEN_128 = io_readreg2 == io_writereg & io_wen ? io_writedata : _GEN_127; // @[register-file.scala 62:16 68:57 69:20]
  assign io_readdata1 = io_readreg1 == io_writereg & io_wen ? io_writedata : _GEN_95; // @[register-file.scala 61:16 66:50 67:20]
  assign io_readdata2 = io_readreg1 == io_writereg & io_wen ? _GEN_127 : _GEN_128; // @[register-file.scala 62:16 66:50]
  always @(posedge clock) begin
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h0 == io_writereg) begin // @[register-file.scala 56:23]
        regs_0 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1 == io_writereg) begin // @[register-file.scala 56:23]
        regs_1 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h2 == io_writereg) begin // @[register-file.scala 56:23]
        regs_2 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h3 == io_writereg) begin // @[register-file.scala 56:23]
        regs_3 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h4 == io_writereg) begin // @[register-file.scala 56:23]
        regs_4 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h5 == io_writereg) begin // @[register-file.scala 56:23]
        regs_5 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h6 == io_writereg) begin // @[register-file.scala 56:23]
        regs_6 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h7 == io_writereg) begin // @[register-file.scala 56:23]
        regs_7 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h8 == io_writereg) begin // @[register-file.scala 56:23]
        regs_8 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h9 == io_writereg) begin // @[register-file.scala 56:23]
        regs_9 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'ha == io_writereg) begin // @[register-file.scala 56:23]
        regs_10 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'hb == io_writereg) begin // @[register-file.scala 56:23]
        regs_11 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'hc == io_writereg) begin // @[register-file.scala 56:23]
        regs_12 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'hd == io_writereg) begin // @[register-file.scala 56:23]
        regs_13 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'he == io_writereg) begin // @[register-file.scala 56:23]
        regs_14 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'hf == io_writereg) begin // @[register-file.scala 56:23]
        regs_15 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h10 == io_writereg) begin // @[register-file.scala 56:23]
        regs_16 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h11 == io_writereg) begin // @[register-file.scala 56:23]
        regs_17 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h12 == io_writereg) begin // @[register-file.scala 56:23]
        regs_18 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h13 == io_writereg) begin // @[register-file.scala 56:23]
        regs_19 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h14 == io_writereg) begin // @[register-file.scala 56:23]
        regs_20 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h15 == io_writereg) begin // @[register-file.scala 56:23]
        regs_21 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h16 == io_writereg) begin // @[register-file.scala 56:23]
        regs_22 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h17 == io_writereg) begin // @[register-file.scala 56:23]
        regs_23 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h18 == io_writereg) begin // @[register-file.scala 56:23]
        regs_24 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h19 == io_writereg) begin // @[register-file.scala 56:23]
        regs_25 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1a == io_writereg) begin // @[register-file.scala 56:23]
        regs_26 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1b == io_writereg) begin // @[register-file.scala 56:23]
        regs_27 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1c == io_writereg) begin // @[register-file.scala 56:23]
        regs_28 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1d == io_writereg) begin // @[register-file.scala 56:23]
        regs_29 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1e == io_writereg) begin // @[register-file.scala 56:23]
        regs_30 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
    if (io_wen) begin // @[register-file.scala 55:17]
      if (5'h1f == io_writereg) begin // @[register-file.scala 56:23]
        regs_31 <= io_writedata; // @[register-file.scala 56:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALUControl(
  input        io_aluop,
  input        io_itype,
  input  [6:0] io_funct7,
  input  [2:0] io_funct3,
  output [3:0] io_operation
);
  wire  _T_1 = io_funct7 == 7'h0; // @[alucontrol.scala 32:35]
  wire [2:0] _GEN_0 = io_itype | io_funct7 == 7'h0 ? 3'h7 : 3'h4; // @[alucontrol.scala 32:53 33:22 35:22]
  wire [1:0] _GEN_1 = _T_1 ? 2'h2 : 2'h3; // @[alucontrol.scala 43:41 44:22 46:22]
  wire [2:0] _GEN_2 = io_funct3 == 3'h6 ? 3'h5 : 3'h6; // @[alucontrol.scala 49:{40,55} 51:20]
  wire [2:0] _GEN_3 = io_funct3 == 3'h5 ? {{1'd0}, _GEN_1} : _GEN_2; // @[alucontrol.scala 42:40]
  wire [2:0] _GEN_4 = io_funct3 == 3'h4 ? 3'h0 : _GEN_3; // @[alucontrol.scala 41:{40,55}]
  wire [2:0] _GEN_5 = io_funct3 == 3'h3 ? 3'h1 : _GEN_4; // @[alucontrol.scala 40:{40,55}]
  wire [3:0] _GEN_6 = io_funct3 == 3'h2 ? 4'h9 : {{1'd0}, _GEN_5}; // @[alucontrol.scala 39:{40,55}]
  wire [3:0] _GEN_7 = io_funct3 == 3'h1 ? 4'h8 : _GEN_6; // @[alucontrol.scala 38:{40,55}]
  wire [3:0] _GEN_8 = io_funct3 == 3'h0 ? {{1'd0}, _GEN_0} : _GEN_7; // @[alucontrol.scala 31:35]
  assign io_operation = io_aluop ? _GEN_8 : 4'h7; // @[alucontrol.scala 30:19 53:18]
endmodule
module ALU(
  input  [3:0]  io_operation,
  input  [31:0] io_inputx,
  input  [31:0] io_inputy,
  output [31:0] io_result
);
  wire [31:0] _T_1 = io_inputx & io_inputy; // @[alu.scala 26:28]
  wire [31:0] _T_3 = io_inputx | io_inputy; // @[alu.scala 29:28]
  wire [31:0] _T_6 = io_inputx + io_inputy; // @[alu.scala 32:28]
  wire [31:0] _T_9 = io_inputx - io_inputy; // @[alu.scala 35:28]
  wire [31:0] _T_11 = io_inputx; // @[alu.scala 38:29]
  wire [31:0] _T_14 = $signed(io_inputx) >>> io_inputy[4:0]; // @[alu.scala 38:55]
  wire [31:0] _T_18 = io_inputx ^ io_inputy; // @[alu.scala 44:28]
  wire [31:0] _T_21 = io_inputx >> io_inputy[4:0]; // @[alu.scala 47:28]
  wire [31:0] _T_24 = io_inputy; // @[alu.scala 50:48]
  wire [62:0] _GEN_15 = {{31'd0}, io_inputx}; // @[alu.scala 53:28]
  wire [62:0] _T_28 = _GEN_15 << io_inputy[4:0]; // @[alu.scala 53:28]
  wire [31:0] _T_31 = ~_T_3; // @[alu.scala 56:18]
  wire  _GEN_0 = io_operation == 4'he & io_inputx != io_inputy; // @[alu.scala 67:42 68:15 71:15]
  wire  _GEN_1 = io_operation == 4'hd ? io_inputx == io_inputy : _GEN_0; // @[alu.scala 64:42 65:15]
  wire  _GEN_2 = io_operation == 4'hc ? io_inputx >= io_inputy : _GEN_1; // @[alu.scala 61:42 62:15]
  wire  _GEN_3 = io_operation == 4'hb ? $signed(io_inputx) >= $signed(io_inputy) : _GEN_2; // @[alu.scala 58:42 59:15]
  wire [31:0] _GEN_4 = io_operation == 4'ha ? _T_31 : {{31'd0}, _GEN_3}; // @[alu.scala 55:42 56:15]
  wire [62:0] _GEN_5 = io_operation == 4'h8 ? _T_28 : {{31'd0}, _GEN_4}; // @[alu.scala 52:42 53:15]
  wire [62:0] _GEN_6 = io_operation == 4'h9 ? {{62'd0}, $signed(_T_11) < $signed(_T_24)} : _GEN_5; // @[alu.scala 49:42 50:15]
  wire [62:0] _GEN_7 = io_operation == 4'h2 ? {{31'd0}, _T_21} : _GEN_6; // @[alu.scala 46:42 47:15]
  wire [62:0] _GEN_8 = io_operation == 4'h0 ? {{31'd0}, _T_18} : _GEN_7; // @[alu.scala 43:42 44:15]
  wire [62:0] _GEN_9 = io_operation == 4'h1 ? {{62'd0}, io_inputx < io_inputy} : _GEN_8; // @[alu.scala 40:42 41:15]
  wire [62:0] _GEN_10 = io_operation == 4'h3 ? {{31'd0}, _T_14} : _GEN_9; // @[alu.scala 37:42 38:15]
  wire [62:0] _GEN_11 = io_operation == 4'h4 ? {{31'd0}, _T_9} : _GEN_10; // @[alu.scala 34:42 35:15]
  wire [62:0] _GEN_12 = io_operation == 4'h7 ? {{31'd0}, _T_6} : _GEN_11; // @[alu.scala 31:42 32:15]
  wire [62:0] _GEN_13 = io_operation == 4'h5 ? {{31'd0}, _T_3} : _GEN_12; // @[alu.scala 28:42 29:15]
  wire [62:0] _GEN_14 = io_operation == 4'h6 ? {{31'd0}, _T_1} : _GEN_13; // @[alu.scala 25:37 26:15]
  assign io_result = _GEN_14[31:0];
endmodule
module ImmediateGenerator(
  input  [31:0] io_instruction,
  output [31:0] io_sextImm
);
  wire [6:0] opcode = io_instruction[6:0]; // @[helpers.scala 44:30]
  wire  _T = 7'h37 == opcode; // @[Conditional.scala 37:30]
  wire [31:0] _T_3 = {io_instruction[31:12],12'h0}; // @[Cat.scala 30:58]
  wire  _T_4 = 7'h17 == opcode; // @[Conditional.scala 37:30]
  wire  _T_8 = 7'h6f == opcode; // @[Conditional.scala 37:30]
  wire [19:0] _T_15 = {io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:21]}; // @[Cat.scala 30:58]
  wire [10:0] _T_18 = _T_15[19] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_20 = {_T_18,io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:21],1'h0}; // @[Cat.scala 30:58]
  wire  _T_21 = 7'h67 == opcode; // @[Conditional.scala 37:30]
  wire [19:0] _T_25 = io_instruction[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_26 = {_T_25,io_instruction[31:20]}; // @[Cat.scala 30:58]
  wire  _T_27 = 7'h63 == opcode; // @[Conditional.scala 37:30]
  wire [11:0] _T_34 = {io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8]}; // @[Cat.scala 30:58]
  wire [18:0] _T_37 = _T_34[11] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_39 = {_T_37,io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8],1'h0}; // @[Cat.scala 30:58]
  wire  _T_40 = 7'h3 == opcode; // @[Conditional.scala 37:30]
  wire  _T_46 = 7'h23 == opcode; // @[Conditional.scala 37:30]
  wire [11:0] _T_49 = {io_instruction[31:25],io_instruction[11:7]}; // @[Cat.scala 30:58]
  wire [19:0] _T_52 = _T_49[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_53 = {_T_52,io_instruction[31:25],io_instruction[11:7]}; // @[Cat.scala 30:58]
  wire  _T_54 = 7'h13 == opcode; // @[Conditional.scala 37:30]
  wire  _T_60 = 7'h73 == opcode; // @[Conditional.scala 37:30]
  wire [31:0] _T_63 = {27'h0,io_instruction[19:15]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_0 = _T_60 ? _T_63 : 32'h0; // @[Conditional.scala 39:67 helpers.scala 42:14 81:18]
  wire [31:0] _GEN_1 = _T_54 ? _T_26 : _GEN_0; // @[Conditional.scala 39:67 helpers.scala 78:18]
  wire [31:0] _GEN_2 = _T_46 ? _T_53 : _GEN_1; // @[Conditional.scala 39:67 helpers.scala 74:18]
  wire [31:0] _GEN_3 = _T_40 ? _T_26 : _GEN_2; // @[Conditional.scala 39:67 helpers.scala 70:18]
  wire [31:0] _GEN_4 = _T_27 ? _T_39 : _GEN_3; // @[Conditional.scala 39:67 helpers.scala 66:18]
  wire [31:0] _GEN_5 = _T_21 ? _T_26 : _GEN_4; // @[Conditional.scala 39:67 helpers.scala 61:18]
  wire [31:0] _GEN_6 = _T_8 ? _T_20 : _GEN_5; // @[Conditional.scala 39:67 helpers.scala 57:18]
  wire [31:0] _GEN_7 = _T_4 ? _T_3 : _GEN_6; // @[Conditional.scala 39:67 helpers.scala 52:18]
  assign io_sextImm = _T ? _T_3 : _GEN_7; // @[Conditional.scala 40:58 helpers.scala 48:18]
endmodule
module Adder(
  input  [31:0] io_inputx,
  input  [31:0] io_inputy,
  output [31:0] io_result
);
  assign io_result = io_inputx + io_inputy; // @[helpers.scala 23:26]
endmodule
module NextPC(
  input         io_branch,
  input         io_jal,
  input         io_jalr,
  input  [31:0] io_inputx,
  input  [31:0] io_inputy,
  input  [2:0]  io_funct3,
  input  [31:0] io_pc,
  input  [31:0] io_imm,
  output [31:0] io_nextpc,
  output        io_taken
);
  wire  _GEN_0 = io_funct3 == 3'h7 & io_inputx >= io_inputy; // @[nextpc.scala 44:{40,51} 45:51]
  wire  _GEN_1 = io_funct3 == 3'h6 ? io_inputx < io_inputy : _GEN_0; // @[nextpc.scala 43:{40,51}]
  wire  _GEN_2 = io_funct3 == 3'h5 ? $signed(io_inputx) >= $signed(io_inputy) : _GEN_1; // @[nextpc.scala 42:{40,51}]
  wire  _GEN_3 = io_funct3 == 3'h4 ? $signed(io_inputx) < $signed(io_inputy) : _GEN_2; // @[nextpc.scala 41:{40,51}]
  wire  _GEN_4 = io_funct3 == 3'h1 ? io_inputx != io_inputy : _GEN_3; // @[nextpc.scala 40:{40,51}]
  wire  _GEN_5 = io_funct3 == 3'h0 ? io_inputx == io_inputy : _GEN_4; // @[nextpc.scala 39:{40,51}]
  wire [31:0] _T_17 = io_pc + io_imm; // @[nextpc.scala 48:26]
  wire [31:0] _T_19 = io_pc + 32'h4; // @[nextpc.scala 50:26]
  wire [31:0] _GEN_6 = io_taken ? _T_17 : _T_19; // @[nextpc.scala 47:21 48:17 50:17]
  wire [31:0] _T_23 = io_inputx + io_imm; // @[nextpc.scala 57:28]
  wire [31:0] _GEN_8 = io_jalr ? _T_23 : _T_19; // @[nextpc.scala 55:25 57:15 59:15]
  wire  _GEN_9 = io_jal | io_jalr; // @[nextpc.scala 52:24 53:14]
  wire [31:0] _GEN_10 = io_jal ? _T_17 : _GEN_8; // @[nextpc.scala 52:24 54:15]
  assign io_nextpc = io_branch ? _GEN_6 : _GEN_10; // @[nextpc.scala 38:20]
  assign io_taken = io_branch ? _GEN_5 : _GEN_9; // @[nextpc.scala 38:20]
endmodule
module ForwardingUnit(
  input  [4:0] io_rs1,
  input  [4:0] io_rs2,
  input  [4:0] io_exmemrd,
  input        io_exmemrw,
  input  [4:0] io_memwbrd,
  input        io_memwbrw,
  output [1:0] io_forwardA,
  output [1:0] io_forwardB
);
  wire  _T_3 = io_exmemrd != 5'h0; // @[forwarding.scala 40:70]
  wire  _T_8 = io_memwbrd != 5'h0; // @[forwarding.scala 43:75]
  wire [1:0] _GEN_0 = io_memwbrw & io_memwbrd == io_rs1 & io_memwbrd != 5'h0 ? 2'h2 : 2'h0; // @[forwarding.scala 43:84 44:17 47:17]
  wire [1:0] _GEN_2 = io_memwbrw & io_memwbrd == io_rs2 & _T_8 ? 2'h2 : 2'h0; // @[forwarding.scala 53:84 54:17 57:17]
  assign io_forwardA = io_exmemrw & io_exmemrd == io_rs1 & io_exmemrd != 5'h0 ? 2'h1 : _GEN_0; // @[forwarding.scala 40:79 41:17]
  assign io_forwardB = io_exmemrw & io_exmemrd == io_rs2 & _T_3 ? 2'h1 : _GEN_2; // @[forwarding.scala 50:79 51:17]
endmodule
module HazardUnitBP(
  input  [4:0] io_rs1,
  input  [4:0] io_rs2,
  input        io_idex_memread,
  input  [4:0] io_idex_rd,
  input        io_exmem_taken,
  output [1:0] io_pcSel,
  output       io_if_id_stall,
  output       io_if_id_flush,
  output       io_id_ex_flush,
  output       io_ex_mem_flush
);
  wire  _T_4 = io_idex_rd == io_rs1 | io_idex_rd == io_rs2; // @[hazard-bp.scala 56:32]
  wire  _T_5 = io_idex_memread & _T_4; // @[hazard-bp.scala 55:41]
  wire [1:0] _GEN_3 = _T_5 ? 2'h3 : 2'h0; // @[hazard-bp.scala 56:59 58:14]
  assign io_pcSel = io_exmem_taken ? 2'h1 : _GEN_3; // @[hazard-bp.scala 48:36 50:14]
  assign io_if_id_stall = io_exmem_taken ? 1'h0 : _T_5; // @[hazard-bp.scala 43:19 48:36]
  assign io_if_id_flush = io_exmem_taken; // @[hazard-bp.scala 48:36 51:21]
  assign io_id_ex_flush = io_exmem_taken | _T_5; // @[hazard-bp.scala 48:36 52:21]
  assign io_ex_mem_flush = io_exmem_taken; // @[hazard-bp.scala 48:36 53:21]
endmodule
module StageReg(
  input         clock,
  input         reset,
  input  [31:0] io_in_instruction,
  input  [31:0] io_in_pc,
  input         io_flush,
  input         io_valid,
  output [31:0] io_data_instruction,
  output [31:0] io_data_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_instruction; // @[stage-register.scala 43:21]
  reg [31:0] reg_pc; // @[stage-register.scala 43:21]
  assign io_data_instruction = reg_instruction; // @[stage-register.scala 45:11]
  assign io_data_pc = reg_pc; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_instruction <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_instruction <= 32'h0; // @[stage-register.scala 52:9]
    end else if (io_valid) begin // @[stage-register.scala 47:19]
      reg_instruction <= io_in_instruction; // @[stage-register.scala 48:9]
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_pc <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_pc <= 32'h0; // @[stage-register.scala 52:9]
    end else if (io_valid) begin // @[stage-register.scala 47:19]
      reg_pc <= io_in_pc; // @[stage-register.scala 48:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_instruction = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_pc = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_instruction,
  input  [31:0] io_in_sextImm,
  input  [31:0] io_in_readdata1,
  input  [31:0] io_in_readdata2,
  input         io_flush,
  output [31:0] io_data_pc,
  output [31:0] io_data_instruction,
  output [31:0] io_data_sextImm,
  output [31:0] io_data_readdata1,
  output [31:0] io_data_readdata2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[stage-register.scala 43:21]
  reg [31:0] reg_instruction; // @[stage-register.scala 43:21]
  reg [31:0] reg_sextImm; // @[stage-register.scala 43:21]
  reg [31:0] reg_readdata1; // @[stage-register.scala 43:21]
  reg [31:0] reg_readdata2; // @[stage-register.scala 43:21]
  assign io_data_pc = reg_pc; // @[stage-register.scala 45:11]
  assign io_data_instruction = reg_instruction; // @[stage-register.scala 45:11]
  assign io_data_sextImm = reg_sextImm; // @[stage-register.scala 45:11]
  assign io_data_readdata1 = reg_readdata1; // @[stage-register.scala 45:11]
  assign io_data_readdata2 = reg_readdata2; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_pc <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_pc <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_pc <= io_in_pc;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_instruction <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_instruction <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_instruction <= io_in_instruction;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_sextImm <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_sextImm <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_sextImm <= io_in_sextImm;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_readdata1 <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_readdata1 <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_readdata1 <= io_in_readdata1;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_readdata2 <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_readdata2 <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_readdata2 <= io_in_readdata2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_instruction = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_sextImm = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_readdata1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_readdata2 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_2(
  input        clock,
  input        reset,
  input        io_in_ex_ctrl_itype,
  input        io_in_ex_ctrl_aluop,
  input        io_in_ex_ctrl_resultselect,
  input        io_in_ex_ctrl_xsrc,
  input        io_in_ex_ctrl_ysrc,
  input        io_in_ex_ctrl_plus4,
  input        io_in_ex_ctrl_branch,
  input        io_in_ex_ctrl_jal,
  input        io_in_ex_ctrl_jalr,
  input  [1:0] io_in_mem_ctrl_memop,
  input        io_in_wb_ctrl_toreg,
  input        io_in_wb_ctrl_regwrite,
  input        io_flush,
  output       io_data_ex_ctrl_itype,
  output       io_data_ex_ctrl_aluop,
  output       io_data_ex_ctrl_resultselect,
  output       io_data_ex_ctrl_xsrc,
  output       io_data_ex_ctrl_ysrc,
  output       io_data_ex_ctrl_plus4,
  output       io_data_ex_ctrl_branch,
  output       io_data_ex_ctrl_jal,
  output       io_data_ex_ctrl_jalr,
  output [1:0] io_data_mem_ctrl_memop,
  output       io_data_wb_ctrl_toreg,
  output       io_data_wb_ctrl_regwrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  reg_ex_ctrl_itype; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_aluop; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_resultselect; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_xsrc; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_ysrc; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_plus4; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_branch; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_jal; // @[stage-register.scala 43:21]
  reg  reg_ex_ctrl_jalr; // @[stage-register.scala 43:21]
  reg [1:0] reg_mem_ctrl_memop; // @[stage-register.scala 43:21]
  reg  reg_wb_ctrl_toreg; // @[stage-register.scala 43:21]
  reg  reg_wb_ctrl_regwrite; // @[stage-register.scala 43:21]
  assign io_data_ex_ctrl_itype = reg_ex_ctrl_itype; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_aluop = reg_ex_ctrl_aluop; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_resultselect = reg_ex_ctrl_resultselect; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_xsrc = reg_ex_ctrl_xsrc; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_ysrc = reg_ex_ctrl_ysrc; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_plus4 = reg_ex_ctrl_plus4; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_branch = reg_ex_ctrl_branch; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_jal = reg_ex_ctrl_jal; // @[stage-register.scala 45:11]
  assign io_data_ex_ctrl_jalr = reg_ex_ctrl_jalr; // @[stage-register.scala 45:11]
  assign io_data_mem_ctrl_memop = reg_mem_ctrl_memop; // @[stage-register.scala 45:11]
  assign io_data_wb_ctrl_toreg = reg_wb_ctrl_toreg; // @[stage-register.scala 45:11]
  assign io_data_wb_ctrl_regwrite = reg_wb_ctrl_regwrite; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_itype <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_itype <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_itype <= io_in_ex_ctrl_itype;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_aluop <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_aluop <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_aluop <= io_in_ex_ctrl_aluop;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_resultselect <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_resultselect <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_resultselect <= io_in_ex_ctrl_resultselect;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_xsrc <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_xsrc <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_xsrc <= io_in_ex_ctrl_xsrc;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_ysrc <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_ysrc <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_ysrc <= io_in_ex_ctrl_ysrc;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_plus4 <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_plus4 <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_plus4 <= io_in_ex_ctrl_plus4;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_branch <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_branch <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_branch <= io_in_ex_ctrl_branch;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_jal <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_jal <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_jal <= io_in_ex_ctrl_jal;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_ctrl_jalr <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_ctrl_jalr <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_ctrl_jalr <= io_in_ex_ctrl_jalr;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_mem_ctrl_memop <= 2'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_mem_ctrl_memop <= 2'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_mem_ctrl_memop <= io_in_mem_ctrl_memop;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_toreg <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_wb_ctrl_toreg <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_wb_ctrl_toreg <= io_in_wb_ctrl_toreg;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_regwrite <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_wb_ctrl_regwrite <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_wb_ctrl_regwrite <= io_in_wb_ctrl_regwrite;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ex_ctrl_itype = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_ex_ctrl_aluop = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_ex_ctrl_resultselect = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_ex_ctrl_xsrc = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_ex_ctrl_ysrc = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_ex_ctrl_plus4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  reg_ex_ctrl_branch = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  reg_ex_ctrl_jal = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_ex_ctrl_jalr = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  reg_mem_ctrl_memop = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reg_wb_ctrl_toreg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_wb_ctrl_regwrite = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_3(
  input         clock,
  input         reset,
  input  [31:0] io_in_ex_result,
  input  [31:0] io_in_mem_writedata,
  input  [31:0] io_in_instruction,
  input  [31:0] io_in_next_pc,
  input         io_in_taken,
  input         io_flush,
  output [31:0] io_data_ex_result,
  output [31:0] io_data_mem_writedata,
  output [31:0] io_data_instruction,
  output [31:0] io_data_next_pc,
  output        io_data_taken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_ex_result; // @[stage-register.scala 43:21]
  reg [31:0] reg_mem_writedata; // @[stage-register.scala 43:21]
  reg [31:0] reg_instruction; // @[stage-register.scala 43:21]
  reg [31:0] reg_next_pc; // @[stage-register.scala 43:21]
  reg  reg_taken; // @[stage-register.scala 43:21]
  assign io_data_ex_result = reg_ex_result; // @[stage-register.scala 45:11]
  assign io_data_mem_writedata = reg_mem_writedata; // @[stage-register.scala 45:11]
  assign io_data_instruction = reg_instruction; // @[stage-register.scala 45:11]
  assign io_data_next_pc = reg_next_pc; // @[stage-register.scala 45:11]
  assign io_data_taken = reg_taken; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_result <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_ex_result <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_ex_result <= io_in_ex_result;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_mem_writedata <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_mem_writedata <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_mem_writedata <= io_in_mem_writedata;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_instruction <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_instruction <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_instruction <= io_in_instruction;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_next_pc <= 32'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_next_pc <= 32'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_next_pc <= io_in_next_pc;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_taken <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_taken <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_taken <= io_in_taken;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ex_result = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mem_writedata = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_next_pc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_taken = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_4(
  input        clock,
  input        reset,
  input  [1:0] io_in_mem_ctrl_memop,
  input        io_in_wb_ctrl_toreg,
  input        io_in_wb_ctrl_regwrite,
  input        io_flush,
  output [1:0] io_data_mem_ctrl_memop,
  output       io_data_wb_ctrl_toreg,
  output       io_data_wb_ctrl_regwrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] reg_mem_ctrl_memop; // @[stage-register.scala 43:21]
  reg  reg_wb_ctrl_toreg; // @[stage-register.scala 43:21]
  reg  reg_wb_ctrl_regwrite; // @[stage-register.scala 43:21]
  assign io_data_mem_ctrl_memop = reg_mem_ctrl_memop; // @[stage-register.scala 45:11]
  assign io_data_wb_ctrl_toreg = reg_wb_ctrl_toreg; // @[stage-register.scala 45:11]
  assign io_data_wb_ctrl_regwrite = reg_wb_ctrl_regwrite; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_mem_ctrl_memop <= 2'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_mem_ctrl_memop <= 2'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_mem_ctrl_memop <= io_in_mem_ctrl_memop;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_toreg <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_wb_ctrl_toreg <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_wb_ctrl_toreg <= io_in_wb_ctrl_toreg;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_regwrite <= 1'h0; // @[stage-register.scala 43:21]
    end else if (io_flush) begin // @[stage-register.scala 51:19]
      reg_wb_ctrl_regwrite <= 1'h0; // @[stage-register.scala 52:9]
    end else begin
      reg_wb_ctrl_regwrite <= io_in_wb_ctrl_regwrite;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mem_ctrl_memop = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reg_wb_ctrl_toreg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_wb_ctrl_regwrite = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_5(
  input         clock,
  input         reset,
  input  [31:0] io_in_instruction,
  input  [31:0] io_in_readdata,
  input  [31:0] io_in_ex_result,
  output [31:0] io_data_instruction,
  output [31:0] io_data_readdata,
  output [31:0] io_data_ex_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_instruction; // @[stage-register.scala 43:21]
  reg [31:0] reg_readdata; // @[stage-register.scala 43:21]
  reg [31:0] reg_ex_result; // @[stage-register.scala 43:21]
  assign io_data_instruction = reg_instruction; // @[stage-register.scala 45:11]
  assign io_data_readdata = reg_readdata; // @[stage-register.scala 45:11]
  assign io_data_ex_result = reg_ex_result; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_instruction <= 32'h0; // @[stage-register.scala 43:21]
    end else begin
      reg_instruction <= io_in_instruction;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_readdata <= 32'h0; // @[stage-register.scala 43:21]
    end else begin
      reg_readdata <= io_in_readdata;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_ex_result <= 32'h0; // @[stage-register.scala 43:21]
    end else begin
      reg_ex_result <= io_in_ex_result;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_instruction = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_readdata = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_ex_result = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StageReg_6(
  input   clock,
  input   reset,
  input   io_in_wb_ctrl_toreg,
  input   io_in_wb_ctrl_regwrite,
  output  io_data_wb_ctrl_toreg,
  output  io_data_wb_ctrl_regwrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  reg_wb_ctrl_toreg; // @[stage-register.scala 43:21]
  reg  reg_wb_ctrl_regwrite; // @[stage-register.scala 43:21]
  assign io_data_wb_ctrl_toreg = reg_wb_ctrl_toreg; // @[stage-register.scala 45:11]
  assign io_data_wb_ctrl_regwrite = reg_wb_ctrl_regwrite; // @[stage-register.scala 45:11]
  always @(posedge clock) begin
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_toreg <= 1'h0; // @[stage-register.scala 43:21]
    end else begin
      reg_wb_ctrl_toreg <= io_in_wb_ctrl_toreg;
    end
    if (reset) begin // @[stage-register.scala 43:21]
      reg_wb_ctrl_regwrite <= 1'h0; // @[stage-register.scala 43:21]
    end else begin
      reg_wb_ctrl_regwrite <= io_in_wb_ctrl_regwrite;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_wb_ctrl_toreg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_wb_ctrl_regwrite = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelinedCPUBP(
  input         clock,
  input         reset,
  output [31:0] io_imem_address,
  input  [31:0] io_imem_instruction,
  output [31:0] io_dmem_address,
  output        io_dmem_valid,
  output [31:0] io_dmem_writedata,
  output        io_dmem_memread,
  output        io_dmem_memwrite,
  output [1:0]  io_dmem_maskmode,
  output        io_dmem_sext,
  input  [31:0] io_dmem_readdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] control_io_opcode; // @[cpu-bp.scala 93:31]
  wire  control_io_itype; // @[cpu-bp.scala 93:31]
  wire  control_io_aluop; // @[cpu-bp.scala 93:31]
  wire  control_io_xsrc; // @[cpu-bp.scala 93:31]
  wire  control_io_ysrc; // @[cpu-bp.scala 93:31]
  wire  control_io_branch; // @[cpu-bp.scala 93:31]
  wire  control_io_jal; // @[cpu-bp.scala 93:31]
  wire  control_io_jalr; // @[cpu-bp.scala 93:31]
  wire  control_io_plus4; // @[cpu-bp.scala 93:31]
  wire  control_io_resultselect; // @[cpu-bp.scala 93:31]
  wire [1:0] control_io_memop; // @[cpu-bp.scala 93:31]
  wire  control_io_toreg; // @[cpu-bp.scala 93:31]
  wire  control_io_regwrite; // @[cpu-bp.scala 93:31]
  wire  registers_clock; // @[cpu-bp.scala 94:31]
  wire [4:0] registers_io_readreg1; // @[cpu-bp.scala 94:31]
  wire [4:0] registers_io_readreg2; // @[cpu-bp.scala 94:31]
  wire [4:0] registers_io_writereg; // @[cpu-bp.scala 94:31]
  wire [31:0] registers_io_writedata; // @[cpu-bp.scala 94:31]
  wire  registers_io_wen; // @[cpu-bp.scala 94:31]
  wire [31:0] registers_io_readdata1; // @[cpu-bp.scala 94:31]
  wire [31:0] registers_io_readdata2; // @[cpu-bp.scala 94:31]
  wire  aluControl_io_aluop; // @[cpu-bp.scala 95:31]
  wire  aluControl_io_itype; // @[cpu-bp.scala 95:31]
  wire [6:0] aluControl_io_funct7; // @[cpu-bp.scala 95:31]
  wire [2:0] aluControl_io_funct3; // @[cpu-bp.scala 95:31]
  wire [3:0] aluControl_io_operation; // @[cpu-bp.scala 95:31]
  wire [3:0] alu_io_operation; // @[cpu-bp.scala 96:31]
  wire [31:0] alu_io_inputx; // @[cpu-bp.scala 96:31]
  wire [31:0] alu_io_inputy; // @[cpu-bp.scala 96:31]
  wire [31:0] alu_io_result; // @[cpu-bp.scala 96:31]
  wire [31:0] immGen_io_instruction; // @[cpu-bp.scala 97:31]
  wire [31:0] immGen_io_sextImm; // @[cpu-bp.scala 97:31]
  wire [31:0] pcPlusFour_io_inputx; // @[cpu-bp.scala 98:31]
  wire [31:0] pcPlusFour_io_inputy; // @[cpu-bp.scala 98:31]
  wire [31:0] pcPlusFour_io_result; // @[cpu-bp.scala 98:31]
  wire  nextPCmod_io_branch; // @[cpu-bp.scala 99:31]
  wire  nextPCmod_io_jal; // @[cpu-bp.scala 99:31]
  wire  nextPCmod_io_jalr; // @[cpu-bp.scala 99:31]
  wire [31:0] nextPCmod_io_inputx; // @[cpu-bp.scala 99:31]
  wire [31:0] nextPCmod_io_inputy; // @[cpu-bp.scala 99:31]
  wire [2:0] nextPCmod_io_funct3; // @[cpu-bp.scala 99:31]
  wire [31:0] nextPCmod_io_pc; // @[cpu-bp.scala 99:31]
  wire [31:0] nextPCmod_io_imm; // @[cpu-bp.scala 99:31]
  wire [31:0] nextPCmod_io_nextpc; // @[cpu-bp.scala 99:31]
  wire  nextPCmod_io_taken; // @[cpu-bp.scala 99:31]
  wire [4:0] forwarding_io_rs1; // @[cpu-bp.scala 100:31]
  wire [4:0] forwarding_io_rs2; // @[cpu-bp.scala 100:31]
  wire [4:0] forwarding_io_exmemrd; // @[cpu-bp.scala 100:31]
  wire  forwarding_io_exmemrw; // @[cpu-bp.scala 100:31]
  wire [4:0] forwarding_io_memwbrd; // @[cpu-bp.scala 100:31]
  wire  forwarding_io_memwbrw; // @[cpu-bp.scala 100:31]
  wire [1:0] forwarding_io_forwardA; // @[cpu-bp.scala 100:31]
  wire [1:0] forwarding_io_forwardB; // @[cpu-bp.scala 100:31]
  wire [4:0] hazard_io_rs1; // @[cpu-bp.scala 101:31]
  wire [4:0] hazard_io_rs2; // @[cpu-bp.scala 101:31]
  wire  hazard_io_idex_memread; // @[cpu-bp.scala 101:31]
  wire [4:0] hazard_io_idex_rd; // @[cpu-bp.scala 101:31]
  wire  hazard_io_exmem_taken; // @[cpu-bp.scala 101:31]
  wire [1:0] hazard_io_pcSel; // @[cpu-bp.scala 101:31]
  wire  hazard_io_if_id_stall; // @[cpu-bp.scala 101:31]
  wire  hazard_io_if_id_flush; // @[cpu-bp.scala 101:31]
  wire  hazard_io_id_ex_flush; // @[cpu-bp.scala 101:31]
  wire  hazard_io_ex_mem_flush; // @[cpu-bp.scala 101:31]
  wire [31:0] branchAdd_io_inputx; // @[cpu-bp.scala 103:31]
  wire [31:0] branchAdd_io_inputy; // @[cpu-bp.scala 103:31]
  wire [31:0] branchAdd_io_result; // @[cpu-bp.scala 103:31]
  wire  if_id_clock; // @[cpu-bp.scala 107:27]
  wire  if_id_reset; // @[cpu-bp.scala 107:27]
  wire [31:0] if_id_io_in_instruction; // @[cpu-bp.scala 107:27]
  wire [31:0] if_id_io_in_pc; // @[cpu-bp.scala 107:27]
  wire  if_id_io_flush; // @[cpu-bp.scala 107:27]
  wire  if_id_io_valid; // @[cpu-bp.scala 107:27]
  wire [31:0] if_id_io_data_instruction; // @[cpu-bp.scala 107:27]
  wire [31:0] if_id_io_data_pc; // @[cpu-bp.scala 107:27]
  wire  id_ex_clock; // @[cpu-bp.scala 109:27]
  wire  id_ex_reset; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_in_pc; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_in_instruction; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_in_sextImm; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_in_readdata1; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_in_readdata2; // @[cpu-bp.scala 109:27]
  wire  id_ex_io_flush; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_data_pc; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_data_instruction; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_data_sextImm; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_data_readdata1; // @[cpu-bp.scala 109:27]
  wire [31:0] id_ex_io_data_readdata2; // @[cpu-bp.scala 109:27]
  wire  id_ex_ctrl_clock; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_reset; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_itype; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_aluop; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_resultselect; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_xsrc; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_ysrc; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_plus4; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_branch; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_jal; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_ex_ctrl_jalr; // @[cpu-bp.scala 110:27]
  wire [1:0] id_ex_ctrl_io_in_mem_ctrl_memop; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_wb_ctrl_toreg; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_in_wb_ctrl_regwrite; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_flush; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_itype; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_aluop; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_resultselect; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_xsrc; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_ysrc; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_plus4; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_branch; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_jal; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_ex_ctrl_jalr; // @[cpu-bp.scala 110:27]
  wire [1:0] id_ex_ctrl_io_data_mem_ctrl_memop; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_wb_ctrl_toreg; // @[cpu-bp.scala 110:27]
  wire  id_ex_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 110:27]
  wire  ex_mem_clock; // @[cpu-bp.scala 112:27]
  wire  ex_mem_reset; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_in_ex_result; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_in_mem_writedata; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_in_instruction; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_in_next_pc; // @[cpu-bp.scala 112:27]
  wire  ex_mem_io_in_taken; // @[cpu-bp.scala 112:27]
  wire  ex_mem_io_flush; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_data_ex_result; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_data_mem_writedata; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_data_instruction; // @[cpu-bp.scala 112:27]
  wire [31:0] ex_mem_io_data_next_pc; // @[cpu-bp.scala 112:27]
  wire  ex_mem_io_data_taken; // @[cpu-bp.scala 112:27]
  wire  ex_mem_ctrl_clock; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_reset; // @[cpu-bp.scala 113:27]
  wire [1:0] ex_mem_ctrl_io_in_mem_ctrl_memop; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_io_in_wb_ctrl_toreg; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_io_in_wb_ctrl_regwrite; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_io_flush; // @[cpu-bp.scala 113:27]
  wire [1:0] ex_mem_ctrl_io_data_mem_ctrl_memop; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_io_data_wb_ctrl_toreg; // @[cpu-bp.scala 113:27]
  wire  ex_mem_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 113:27]
  wire  mem_wb_clock; // @[cpu-bp.scala 115:27]
  wire  mem_wb_reset; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_in_instruction; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_in_readdata; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_in_ex_result; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_data_instruction; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_data_readdata; // @[cpu-bp.scala 115:27]
  wire [31:0] mem_wb_io_data_ex_result; // @[cpu-bp.scala 115:27]
  wire  mem_wb_ctrl_clock; // @[cpu-bp.scala 119:27]
  wire  mem_wb_ctrl_reset; // @[cpu-bp.scala 119:27]
  wire  mem_wb_ctrl_io_in_wb_ctrl_toreg; // @[cpu-bp.scala 119:27]
  wire  mem_wb_ctrl_io_in_wb_ctrl_regwrite; // @[cpu-bp.scala 119:27]
  wire  mem_wb_ctrl_io_data_wb_ctrl_toreg; // @[cpu-bp.scala 119:27]
  wire  mem_wb_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 119:27]
  reg [31:0] pc; // @[cpu-bp.scala 92:32]
  reg [31:0] bpCorrect; // @[cpu-bp.scala 121:28]
  reg [31:0] bpIncorrect; // @[cpu-bp.scala 122:28]
  wire  _T_5 = bpCorrect > 32'h100000; // @[cpu-bp.scala 123:19]
  wire  _T_8 = hazard_io_pcSel == 2'h0; // @[cpu-bp.scala 159:30]
  wire  _T_9 = hazard_io_pcSel == 2'h1; // @[cpu-bp.scala 160:30]
  wire  _T_10 = hazard_io_pcSel == 2'h2; // @[cpu-bp.scala 161:30]
  wire  _T_11 = hazard_io_pcSel == 2'h3; // @[cpu-bp.scala 162:30]
  wire [31:0] _T_12 = _T_11 ? pc : 32'h0; // @[Mux.scala 87:16]
  wire [31:0] id_next_pc = branchAdd_io_result; // @[cpu-bp.scala 149:24 206:14]
  wire [31:0] next_pc = ex_mem_io_data_next_pc; // @[cpu-bp.scala 148:24 400:11]
  wire [31:0] write_data = mem_wb_ctrl_io_data_wb_ctrl_toreg ? mem_wb_io_data_readdata : mem_wb_io_data_ex_result; // @[cpu-bp.scala 434:55 435:16 437:16]
  wire [31:0] _GEN_3 = forwarding_io_forwardA == 2'h1 ? ex_mem_io_data_ex_result : write_data; // @[cpu-bp.scala 284:48 285:19 287:19]
  wire [31:0] forward_a_mux = forwarding_io_forwardA == 2'h0 ? id_ex_io_data_readdata1 : _GEN_3; // @[cpu-bp.scala 282:41 283:19]
  wire [31:0] _GEN_5 = forwarding_io_forwardB == 2'h1 ? ex_mem_io_data_ex_result : write_data; // @[cpu-bp.scala 295:48 296:19 298:19]
  wire [31:0] forward_b_mux = forwarding_io_forwardB == 2'h0 ? id_ex_io_data_readdata2 : _GEN_5; // @[cpu-bp.scala 293:41 294:19]
  wire [31:0] _GEN_8 = id_ex_ctrl_io_data_ex_ctrl_ysrc ? id_ex_io_data_sextImm : forward_b_mux; // @[cpu-bp.scala 315:55 316:21 318:21]
  wire [31:0] _T_39 = bpCorrect + 32'h1; // @[cpu-bp.scala 356:32]
  wire [31:0] _T_41 = bpIncorrect + 32'h1; // @[cpu-bp.scala 359:34]
  wire  _GEN_14 = nextPCmod_io_taken; // @[cpu-bp.scala 349:71 352:25]
  Control control ( // @[cpu-bp.scala 93:31]
    .io_opcode(control_io_opcode),
    .io_itype(control_io_itype),
    .io_aluop(control_io_aluop),
    .io_xsrc(control_io_xsrc),
    .io_ysrc(control_io_ysrc),
    .io_branch(control_io_branch),
    .io_jal(control_io_jal),
    .io_jalr(control_io_jalr),
    .io_plus4(control_io_plus4),
    .io_resultselect(control_io_resultselect),
    .io_memop(control_io_memop),
    .io_toreg(control_io_toreg),
    .io_regwrite(control_io_regwrite)
  );
  RegisterFile registers ( // @[cpu-bp.scala 94:31]
    .clock(registers_clock),
    .io_readreg1(registers_io_readreg1),
    .io_readreg2(registers_io_readreg2),
    .io_writereg(registers_io_writereg),
    .io_writedata(registers_io_writedata),
    .io_wen(registers_io_wen),
    .io_readdata1(registers_io_readdata1),
    .io_readdata2(registers_io_readdata2)
  );
  ALUControl aluControl ( // @[cpu-bp.scala 95:31]
    .io_aluop(aluControl_io_aluop),
    .io_itype(aluControl_io_itype),
    .io_funct7(aluControl_io_funct7),
    .io_funct3(aluControl_io_funct3),
    .io_operation(aluControl_io_operation)
  );
  ALU alu ( // @[cpu-bp.scala 96:31]
    .io_operation(alu_io_operation),
    .io_inputx(alu_io_inputx),
    .io_inputy(alu_io_inputy),
    .io_result(alu_io_result)
  );
  ImmediateGenerator immGen ( // @[cpu-bp.scala 97:31]
    .io_instruction(immGen_io_instruction),
    .io_sextImm(immGen_io_sextImm)
  );
  Adder pcPlusFour ( // @[cpu-bp.scala 98:31]
    .io_inputx(pcPlusFour_io_inputx),
    .io_inputy(pcPlusFour_io_inputy),
    .io_result(pcPlusFour_io_result)
  );
  NextPC nextPCmod ( // @[cpu-bp.scala 99:31]
    .io_branch(nextPCmod_io_branch),
    .io_jal(nextPCmod_io_jal),
    .io_jalr(nextPCmod_io_jalr),
    .io_inputx(nextPCmod_io_inputx),
    .io_inputy(nextPCmod_io_inputy),
    .io_funct3(nextPCmod_io_funct3),
    .io_pc(nextPCmod_io_pc),
    .io_imm(nextPCmod_io_imm),
    .io_nextpc(nextPCmod_io_nextpc),
    .io_taken(nextPCmod_io_taken)
  );
  ForwardingUnit forwarding ( // @[cpu-bp.scala 100:31]
    .io_rs1(forwarding_io_rs1),
    .io_rs2(forwarding_io_rs2),
    .io_exmemrd(forwarding_io_exmemrd),
    .io_exmemrw(forwarding_io_exmemrw),
    .io_memwbrd(forwarding_io_memwbrd),
    .io_memwbrw(forwarding_io_memwbrw),
    .io_forwardA(forwarding_io_forwardA),
    .io_forwardB(forwarding_io_forwardB)
  );
  HazardUnitBP hazard ( // @[cpu-bp.scala 101:31]
    .io_rs1(hazard_io_rs1),
    .io_rs2(hazard_io_rs2),
    .io_idex_memread(hazard_io_idex_memread),
    .io_idex_rd(hazard_io_idex_rd),
    .io_exmem_taken(hazard_io_exmem_taken),
    .io_pcSel(hazard_io_pcSel),
    .io_if_id_stall(hazard_io_if_id_stall),
    .io_if_id_flush(hazard_io_if_id_flush),
    .io_id_ex_flush(hazard_io_id_ex_flush),
    .io_ex_mem_flush(hazard_io_ex_mem_flush)
  );
  Adder branchAdd ( // @[cpu-bp.scala 103:31]
    .io_inputx(branchAdd_io_inputx),
    .io_inputy(branchAdd_io_inputy),
    .io_result(branchAdd_io_result)
  );
  StageReg if_id ( // @[cpu-bp.scala 107:27]
    .clock(if_id_clock),
    .reset(if_id_reset),
    .io_in_instruction(if_id_io_in_instruction),
    .io_in_pc(if_id_io_in_pc),
    .io_flush(if_id_io_flush),
    .io_valid(if_id_io_valid),
    .io_data_instruction(if_id_io_data_instruction),
    .io_data_pc(if_id_io_data_pc)
  );
  StageReg_1 id_ex ( // @[cpu-bp.scala 109:27]
    .clock(id_ex_clock),
    .reset(id_ex_reset),
    .io_in_pc(id_ex_io_in_pc),
    .io_in_instruction(id_ex_io_in_instruction),
    .io_in_sextImm(id_ex_io_in_sextImm),
    .io_in_readdata1(id_ex_io_in_readdata1),
    .io_in_readdata2(id_ex_io_in_readdata2),
    .io_flush(id_ex_io_flush),
    .io_data_pc(id_ex_io_data_pc),
    .io_data_instruction(id_ex_io_data_instruction),
    .io_data_sextImm(id_ex_io_data_sextImm),
    .io_data_readdata1(id_ex_io_data_readdata1),
    .io_data_readdata2(id_ex_io_data_readdata2)
  );
  StageReg_2 id_ex_ctrl ( // @[cpu-bp.scala 110:27]
    .clock(id_ex_ctrl_clock),
    .reset(id_ex_ctrl_reset),
    .io_in_ex_ctrl_itype(id_ex_ctrl_io_in_ex_ctrl_itype),
    .io_in_ex_ctrl_aluop(id_ex_ctrl_io_in_ex_ctrl_aluop),
    .io_in_ex_ctrl_resultselect(id_ex_ctrl_io_in_ex_ctrl_resultselect),
    .io_in_ex_ctrl_xsrc(id_ex_ctrl_io_in_ex_ctrl_xsrc),
    .io_in_ex_ctrl_ysrc(id_ex_ctrl_io_in_ex_ctrl_ysrc),
    .io_in_ex_ctrl_plus4(id_ex_ctrl_io_in_ex_ctrl_plus4),
    .io_in_ex_ctrl_branch(id_ex_ctrl_io_in_ex_ctrl_branch),
    .io_in_ex_ctrl_jal(id_ex_ctrl_io_in_ex_ctrl_jal),
    .io_in_ex_ctrl_jalr(id_ex_ctrl_io_in_ex_ctrl_jalr),
    .io_in_mem_ctrl_memop(id_ex_ctrl_io_in_mem_ctrl_memop),
    .io_in_wb_ctrl_toreg(id_ex_ctrl_io_in_wb_ctrl_toreg),
    .io_in_wb_ctrl_regwrite(id_ex_ctrl_io_in_wb_ctrl_regwrite),
    .io_flush(id_ex_ctrl_io_flush),
    .io_data_ex_ctrl_itype(id_ex_ctrl_io_data_ex_ctrl_itype),
    .io_data_ex_ctrl_aluop(id_ex_ctrl_io_data_ex_ctrl_aluop),
    .io_data_ex_ctrl_resultselect(id_ex_ctrl_io_data_ex_ctrl_resultselect),
    .io_data_ex_ctrl_xsrc(id_ex_ctrl_io_data_ex_ctrl_xsrc),
    .io_data_ex_ctrl_ysrc(id_ex_ctrl_io_data_ex_ctrl_ysrc),
    .io_data_ex_ctrl_plus4(id_ex_ctrl_io_data_ex_ctrl_plus4),
    .io_data_ex_ctrl_branch(id_ex_ctrl_io_data_ex_ctrl_branch),
    .io_data_ex_ctrl_jal(id_ex_ctrl_io_data_ex_ctrl_jal),
    .io_data_ex_ctrl_jalr(id_ex_ctrl_io_data_ex_ctrl_jalr),
    .io_data_mem_ctrl_memop(id_ex_ctrl_io_data_mem_ctrl_memop),
    .io_data_wb_ctrl_toreg(id_ex_ctrl_io_data_wb_ctrl_toreg),
    .io_data_wb_ctrl_regwrite(id_ex_ctrl_io_data_wb_ctrl_regwrite)
  );
  StageReg_3 ex_mem ( // @[cpu-bp.scala 112:27]
    .clock(ex_mem_clock),
    .reset(ex_mem_reset),
    .io_in_ex_result(ex_mem_io_in_ex_result),
    .io_in_mem_writedata(ex_mem_io_in_mem_writedata),
    .io_in_instruction(ex_mem_io_in_instruction),
    .io_in_next_pc(ex_mem_io_in_next_pc),
    .io_in_taken(ex_mem_io_in_taken),
    .io_flush(ex_mem_io_flush),
    .io_data_ex_result(ex_mem_io_data_ex_result),
    .io_data_mem_writedata(ex_mem_io_data_mem_writedata),
    .io_data_instruction(ex_mem_io_data_instruction),
    .io_data_next_pc(ex_mem_io_data_next_pc),
    .io_data_taken(ex_mem_io_data_taken)
  );
  StageReg_4 ex_mem_ctrl ( // @[cpu-bp.scala 113:27]
    .clock(ex_mem_ctrl_clock),
    .reset(ex_mem_ctrl_reset),
    .io_in_mem_ctrl_memop(ex_mem_ctrl_io_in_mem_ctrl_memop),
    .io_in_wb_ctrl_toreg(ex_mem_ctrl_io_in_wb_ctrl_toreg),
    .io_in_wb_ctrl_regwrite(ex_mem_ctrl_io_in_wb_ctrl_regwrite),
    .io_flush(ex_mem_ctrl_io_flush),
    .io_data_mem_ctrl_memop(ex_mem_ctrl_io_data_mem_ctrl_memop),
    .io_data_wb_ctrl_toreg(ex_mem_ctrl_io_data_wb_ctrl_toreg),
    .io_data_wb_ctrl_regwrite(ex_mem_ctrl_io_data_wb_ctrl_regwrite)
  );
  StageReg_5 mem_wb ( // @[cpu-bp.scala 115:27]
    .clock(mem_wb_clock),
    .reset(mem_wb_reset),
    .io_in_instruction(mem_wb_io_in_instruction),
    .io_in_readdata(mem_wb_io_in_readdata),
    .io_in_ex_result(mem_wb_io_in_ex_result),
    .io_data_instruction(mem_wb_io_data_instruction),
    .io_data_readdata(mem_wb_io_data_readdata),
    .io_data_ex_result(mem_wb_io_data_ex_result)
  );
  StageReg_6 mem_wb_ctrl ( // @[cpu-bp.scala 119:27]
    .clock(mem_wb_ctrl_clock),
    .reset(mem_wb_ctrl_reset),
    .io_in_wb_ctrl_toreg(mem_wb_ctrl_io_in_wb_ctrl_toreg),
    .io_in_wb_ctrl_regwrite(mem_wb_ctrl_io_in_wb_ctrl_regwrite),
    .io_data_wb_ctrl_toreg(mem_wb_ctrl_io_data_wb_ctrl_toreg),
    .io_data_wb_ctrl_regwrite(mem_wb_ctrl_io_data_wb_ctrl_regwrite)
  );
  assign io_imem_address = pc; // @[cpu-bp.scala 164:19]
  assign io_dmem_address = ex_mem_io_data_ex_result; // @[cpu-bp.scala 391:21]
  assign io_dmem_valid = ex_mem_ctrl_io_data_mem_ctrl_memop[1]; // @[cpu-bp.scala 394:58]
  assign io_dmem_writedata = ex_mem_io_data_mem_writedata; // @[cpu-bp.scala 397:21]
  assign io_dmem_memread = ex_mem_ctrl_io_data_mem_ctrl_memop == 2'h2; // @[cpu-bp.scala 392:59]
  assign io_dmem_memwrite = ex_mem_ctrl_io_data_mem_ctrl_memop == 2'h3; // @[cpu-bp.scala 393:59]
  assign io_dmem_maskmode = ex_mem_io_data_instruction[13:12]; // @[cpu-bp.scala 395:50]
  assign io_dmem_sext = ~ex_mem_io_data_instruction[14]; // @[cpu-bp.scala 396:24]
  assign control_io_opcode = if_id_io_data_instruction[6:0]; // @[cpu-bp.scala 184:49]
  assign registers_clock = clock;
  assign registers_io_readreg1 = if_id_io_data_instruction[19:15]; // @[cpu-bp.scala 187:38]
  assign registers_io_readreg2 = if_id_io_data_instruction[24:20]; // @[cpu-bp.scala 188:38]
  assign registers_io_writereg = mem_wb_io_data_instruction[11:7]; // @[cpu-bp.scala 431:54]
  assign registers_io_writedata = mem_wb_ctrl_io_data_wb_ctrl_toreg ? mem_wb_io_data_readdata : mem_wb_io_data_ex_result
    ; // @[cpu-bp.scala 434:55 435:16 437:16]
  assign registers_io_wen = mem_wb_io_data_instruction[11:7] == 5'h0 ? 1'h0 : mem_wb_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 425:51 426:22 428:22]
  assign aluControl_io_aluop = id_ex_ctrl_io_data_ex_ctrl_aluop; // @[cpu-bp.scala 270:24]
  assign aluControl_io_itype = id_ex_ctrl_io_data_ex_ctrl_itype; // @[cpu-bp.scala 269:24]
  assign aluControl_io_funct7 = id_ex_io_data_instruction[31:25]; // @[cpu-bp.scala 272:52]
  assign aluControl_io_funct3 = id_ex_io_data_instruction[14:12]; // @[cpu-bp.scala 271:52]
  assign alu_io_operation = aluControl_io_operation; // @[cpu-bp.scala 302:20]
  assign alu_io_inputx = id_ex_ctrl_io_data_ex_ctrl_xsrc ? id_ex_io_data_pc : forward_a_mux; // @[cpu-bp.scala 306:53 307:19 309:19]
  assign alu_io_inputy = id_ex_ctrl_io_data_ex_ctrl_plus4 ? 32'h4 : _GEN_8; // @[cpu-bp.scala 312:54 313:19]
  assign immGen_io_instruction = if_id_io_data_instruction; // @[cpu-bp.scala 200:25]
  assign pcPlusFour_io_inputx = pc; // @[cpu-bp.scala 168:24]
  assign pcPlusFour_io_inputy = 32'h4; // @[cpu-bp.scala 169:24]
  assign nextPCmod_io_branch = id_ex_ctrl_io_data_ex_ctrl_branch; // @[cpu-bp.scala 275:23]
  assign nextPCmod_io_jal = id_ex_ctrl_io_data_ex_ctrl_jal; // @[cpu-bp.scala 276:23]
  assign nextPCmod_io_jalr = id_ex_ctrl_io_data_ex_ctrl_jalr; // @[cpu-bp.scala 277:23]
  assign nextPCmod_io_inputx = forwarding_io_forwardA == 2'h0 ? id_ex_io_data_readdata1 : _GEN_3; // @[cpu-bp.scala 282:41 283:19]
  assign nextPCmod_io_inputy = forwarding_io_forwardB == 2'h0 ? id_ex_io_data_readdata2 : _GEN_5; // @[cpu-bp.scala 293:41 294:19]
  assign nextPCmod_io_funct3 = id_ex_io_data_instruction[14:12]; // @[cpu-bp.scala 325:51]
  assign nextPCmod_io_pc = id_ex_io_data_pc; // @[cpu-bp.scala 326:23]
  assign nextPCmod_io_imm = id_ex_io_data_sextImm; // @[cpu-bp.scala 327:23]
  assign forwarding_io_rs1 = id_ex_io_data_instruction[19:15]; // @[cpu-bp.scala 263:53]
  assign forwarding_io_rs2 = id_ex_io_data_instruction[24:20]; // @[cpu-bp.scala 264:53]
  assign forwarding_io_exmemrd = ex_mem_io_data_instruction[11:7]; // @[cpu-bp.scala 265:54]
  assign forwarding_io_exmemrw = ex_mem_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 266:25]
  assign forwarding_io_memwbrd = mem_wb_io_data_instruction[11:7]; // @[cpu-bp.scala 441:54]
  assign forwarding_io_memwbrw = mem_wb_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 442:25]
  assign hazard_io_rs1 = if_id_io_data_instruction[19:15]; // @[cpu-bp.scala 187:38]
  assign hazard_io_rs2 = if_id_io_data_instruction[24:20]; // @[cpu-bp.scala 188:38]
  assign hazard_io_idex_memread = id_ex_ctrl_io_data_mem_ctrl_memop == 2'h2; // @[cpu-bp.scala 256:43]
  assign hazard_io_idex_rd = id_ex_io_data_instruction[11:7]; // @[cpu-bp.scala 254:49]
  assign hazard_io_exmem_taken = ex_mem_io_data_taken; // @[cpu-bp.scala 403:25]
  assign branchAdd_io_inputx = if_id_io_data_pc; // @[cpu-bp.scala 203:23]
  assign branchAdd_io_inputy = immGen_io_sextImm; // @[cpu-bp.scala 204:23]
  assign if_id_clock = clock;
  assign if_id_reset = reset;
  assign if_id_io_in_instruction = io_imem_instruction; // @[cpu-bp.scala 172:27]
  assign if_id_io_in_pc = pc; // @[cpu-bp.scala 173:27]
  assign if_id_io_flush = hazard_io_if_id_flush; // @[cpu-bp.scala 177:18]
  assign if_id_io_valid = ~hazard_io_if_id_stall; // @[cpu-bp.scala 176:21]
  assign id_ex_clock = clock;
  assign id_ex_reset = reset;
  assign id_ex_io_in_pc = if_id_io_data_pc; // @[cpu-bp.scala 218:27]
  assign id_ex_io_in_instruction = if_id_io_data_instruction; // @[cpu-bp.scala 220:27]
  assign id_ex_io_in_sextImm = immGen_io_sextImm; // @[cpu-bp.scala 219:27]
  assign id_ex_io_in_readdata1 = registers_io_readdata1; // @[cpu-bp.scala 221:27]
  assign id_ex_io_in_readdata2 = registers_io_readdata2; // @[cpu-bp.scala 222:27]
  assign id_ex_io_flush = hazard_io_id_ex_flush; // @[cpu-bp.scala 244:18]
  assign id_ex_ctrl_clock = clock;
  assign id_ex_ctrl_reset = reset;
  assign id_ex_ctrl_io_in_ex_ctrl_itype = control_io_itype; // @[cpu-bp.scala 226:41]
  assign id_ex_ctrl_io_in_ex_ctrl_aluop = control_io_aluop; // @[cpu-bp.scala 225:41]
  assign id_ex_ctrl_io_in_ex_ctrl_resultselect = control_io_resultselect; // @[cpu-bp.scala 227:41]
  assign id_ex_ctrl_io_in_ex_ctrl_xsrc = control_io_xsrc; // @[cpu-bp.scala 228:41]
  assign id_ex_ctrl_io_in_ex_ctrl_ysrc = control_io_ysrc; // @[cpu-bp.scala 229:41]
  assign id_ex_ctrl_io_in_ex_ctrl_plus4 = control_io_plus4; // @[cpu-bp.scala 230:41]
  assign id_ex_ctrl_io_in_ex_ctrl_branch = control_io_branch; // @[cpu-bp.scala 231:41]
  assign id_ex_ctrl_io_in_ex_ctrl_jal = control_io_jal; // @[cpu-bp.scala 232:41]
  assign id_ex_ctrl_io_in_ex_ctrl_jalr = control_io_jalr; // @[cpu-bp.scala 233:41]
  assign id_ex_ctrl_io_in_mem_ctrl_memop = control_io_memop; // @[cpu-bp.scala 237:35]
  assign id_ex_ctrl_io_in_wb_ctrl_toreg = control_io_toreg; // @[cpu-bp.scala 241:37]
  assign id_ex_ctrl_io_in_wb_ctrl_regwrite = control_io_regwrite; // @[cpu-bp.scala 240:37]
  assign id_ex_ctrl_io_flush = hazard_io_id_ex_flush; // @[cpu-bp.scala 247:23]
  assign ex_mem_clock = clock;
  assign ex_mem_reset = reset;
  assign ex_mem_io_in_ex_result = ~id_ex_ctrl_io_data_ex_ctrl_resultselect ? alu_io_result : id_ex_io_data_sextImm; // @[cpu-bp.scala 342:58 343:28 345:28]
  assign ex_mem_io_in_mem_writedata = forwarding_io_forwardB == 2'h0 ? id_ex_io_data_readdata2 : _GEN_5; // @[cpu-bp.scala 293:41 294:19]
  assign ex_mem_io_in_instruction = id_ex_io_data_instruction; // @[cpu-bp.scala 330:30]
  assign ex_mem_io_in_next_pc = nextPCmod_io_nextpc; // @[cpu-bp.scala 338:24]
  assign ex_mem_io_in_taken = id_ex_ctrl_io_data_ex_ctrl_branch ? _GEN_14 : nextPCmod_io_taken; // @[cpu-bp.scala 339:24 371:43]
  assign ex_mem_io_flush = hazard_io_ex_mem_flush; // @[cpu-bp.scala 382:24]
  assign ex_mem_ctrl_clock = clock;
  assign ex_mem_ctrl_reset = reset;
  assign ex_mem_ctrl_io_in_mem_ctrl_memop = id_ex_ctrl_io_data_mem_ctrl_memop; // @[cpu-bp.scala 333:38]
  assign ex_mem_ctrl_io_in_wb_ctrl_toreg = id_ex_ctrl_io_data_wb_ctrl_toreg; // @[cpu-bp.scala 335:38]
  assign ex_mem_ctrl_io_in_wb_ctrl_regwrite = id_ex_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 334:38]
  assign ex_mem_ctrl_io_flush = hazard_io_ex_mem_flush; // @[cpu-bp.scala 384:24]
  assign mem_wb_clock = clock;
  assign mem_wb_reset = reset;
  assign mem_wb_io_in_instruction = ex_mem_io_data_instruction; // @[cpu-bp.scala 409:28]
  assign mem_wb_io_in_readdata = io_dmem_readdata; // @[cpu-bp.scala 410:28]
  assign mem_wb_io_in_ex_result = ex_mem_io_data_ex_result; // @[cpu-bp.scala 408:28]
  assign mem_wb_ctrl_clock = clock;
  assign mem_wb_ctrl_reset = reset;
  assign mem_wb_ctrl_io_in_wb_ctrl_toreg = ex_mem_ctrl_io_data_wb_ctrl_toreg; // @[cpu-bp.scala 413:38]
  assign mem_wb_ctrl_io_in_wb_ctrl_regwrite = ex_mem_ctrl_io_data_wb_ctrl_regwrite; // @[cpu-bp.scala 412:38]
  always @(posedge clock) begin
    if (reset) begin // @[cpu-bp.scala 92:32]
      pc <= 32'h0; // @[cpu-bp.scala 92:32]
    end else if (_T_8) begin // @[Mux.scala 87:16]
      pc <= pcPlusFour_io_result;
    end else if (_T_9) begin // @[Mux.scala 87:16]
      pc <= next_pc;
    end else if (_T_10) begin // @[Mux.scala 87:16]
      pc <= id_next_pc;
    end else begin
      pc <= _T_12;
    end
    if (reset) begin // @[cpu-bp.scala 121:28]
      bpCorrect <= 32'h0; // @[cpu-bp.scala 121:28]
    end else if (id_ex_ctrl_io_data_ex_ctrl_branch & ~hazard_io_ex_mem_flush) begin // @[cpu-bp.scala 349:71]
      if (~nextPCmod_io_taken) begin // @[cpu-bp.scala 355:73]
        bpCorrect <= _T_39; // @[cpu-bp.scala 356:19]
      end
    end
    if (reset) begin // @[cpu-bp.scala 122:28]
      bpIncorrect <= 32'h0; // @[cpu-bp.scala 122:28]
    end else if (id_ex_ctrl_io_data_ex_ctrl_branch & ~hazard_io_ex_mem_flush) begin // @[cpu-bp.scala 349:71]
      if (!(~nextPCmod_io_taken)) begin // @[cpu-bp.scala 355:73]
        bpIncorrect <= _T_41; // @[cpu-bp.scala 359:19]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~reset) begin
          $fwrite(32'h80000002,"BP correct: %d; incorrect: %d\n",bpCorrect,bpIncorrect); // @[cpu-bp.scala 125:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  bpCorrect = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bpIncorrect = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortedCombinMemory(
  input         clock,
  input         reset,
  input  [31:0] io_imem_request_bits_address,
  output [31:0] io_imem_response_bits_data,
  input         io_dmem_request_valid,
  input  [31:0] io_dmem_request_bits_address,
  input  [31:0] io_dmem_request_bits_writedata,
  input  [1:0]  io_dmem_request_bits_operation,
  output        io_dmem_response_valid,
  output [31:0] io_dmem_response_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] memory [0:16383]; // @[base-memory-components.scala 39:19]
  wire  memory__T_9_en; // @[base-memory-components.scala 39:19]
  wire [13:0] memory__T_9_addr; // @[base-memory-components.scala 39:19]
  wire [31:0] memory__T_9_data; // @[base-memory-components.scala 39:19]
  wire  memory__T_20_en; // @[base-memory-components.scala 39:19]
  wire [13:0] memory__T_20_addr; // @[base-memory-components.scala 39:19]
  wire [31:0] memory__T_20_data; // @[base-memory-components.scala 39:19]
  wire [31:0] memory__T_24_data; // @[base-memory-components.scala 39:19]
  wire [13:0] memory__T_24_addr; // @[base-memory-components.scala 39:19]
  wire  memory__T_24_mask; // @[base-memory-components.scala 39:19]
  wire  memory__T_24_en; // @[base-memory-components.scala 39:19]
  wire  _T_21 = io_dmem_request_bits_operation == 2'h2; // @[memory.scala 65:29]
  assign memory__T_9_en = io_imem_request_bits_address < 32'h10000;
  assign memory__T_9_addr = io_imem_request_bits_address[15:2];
  assign memory__T_9_data = memory[memory__T_9_addr]; // @[base-memory-components.scala 39:19]
  assign memory__T_20_en = io_dmem_request_valid;
  assign memory__T_20_addr = io_dmem_request_bits_address[15:2];
  assign memory__T_20_data = memory[memory__T_20_addr]; // @[base-memory-components.scala 39:19]
  assign memory__T_24_data = io_dmem_request_bits_writedata;
  assign memory__T_24_addr = io_dmem_request_bits_address[15:2];
  assign memory__T_24_mask = 1'h1;
  assign memory__T_24_en = io_dmem_request_valid & _T_21;
  assign io_imem_response_bits_data = io_imem_request_bits_address < 32'h10000 ? memory__T_9_data : 32'h0; // @[memory.scala 35:37 base-memory-components.scala 36:20 memory.scala 37:34]
  assign io_dmem_response_valid = io_dmem_request_valid; // @[base-memory-components.scala 39:19 memory.scala 52:32 61:46]
  assign io_dmem_response_bits_data = io_dmem_request_valid ? memory__T_20_data : 32'h0; // @[base-memory-components.scala 37:20 memory.scala 52:32 61:32]
  always @(posedge clock) begin
    if (memory__T_24_en & memory__T_24_mask) begin
      memory[memory__T_24_addr] <= memory__T_24_data; // @[base-memory-components.scala 39:19]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_dmem_request_valid & ~(io_dmem_request_bits_operation != 2'h1 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at memory.scala:56 assert (request.operation =/= Write)\n"); // @[memory.scala 56:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_dmem_request_valid & ~(io_dmem_request_bits_operation != 2'h1 | reset)) begin
          $fatal; // @[memory.scala 56:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_dmem_request_valid & ~(io_dmem_request_bits_address < 32'h10000 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at memory.scala:58 assert (request.address < size.U)\n"); // @[memory.scala 58:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_dmem_request_valid & ~(io_dmem_request_bits_address < 32'h10000 | reset)) begin
          $fatal; // @[memory.scala 58:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16384; initvar = initvar+1)
    memory[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICombinMemPort(
  input  [31:0] io_pipeline_address,
  output [31:0] io_pipeline_instruction,
  output [31:0] io_bus_request_bits_address,
  input  [31:0] io_bus_response_bits_data
);
  assign io_pipeline_instruction = io_bus_response_bits_data; // @[memory-combin-ports.scala 33:27]
  assign io_bus_request_bits_address = io_pipeline_address; // @[memory-combin-ports.scala 17:23 18:23]
endmodule
module DCombinMemPort(
  input         clock,
  input         reset,
  input  [31:0] io_pipeline_address,
  input         io_pipeline_valid,
  input  [31:0] io_pipeline_writedata,
  input         io_pipeline_memread,
  input         io_pipeline_memwrite,
  input  [1:0]  io_pipeline_maskmode,
  input         io_pipeline_sext,
  output [31:0] io_pipeline_readdata,
  output        io_bus_request_valid,
  output [31:0] io_bus_request_bits_address,
  output [31:0] io_bus_request_bits_writedata,
  output [1:0]  io_bus_request_bits_operation,
  input         io_bus_response_valid,
  input  [31:0] io_bus_response_bits_data
);
  wire  _T_2 = io_pipeline_valid & (io_pipeline_memread | io_pipeline_memwrite); // @[memory-combin-ports.scala 44:27]
  wire  _T_12 = io_pipeline_maskmode == 2'h0; // @[memory-combin-ports.scala 85:36]
  wire  _T_13 = io_pipeline_address[1:0] == 2'h0; // @[memory-combin-ports.scala 86:23]
  wire [31:0] _T_16 = {io_bus_response_bits_data[31:8],io_pipeline_writedata[7:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_22 = {io_bus_response_bits_data[31:16],io_pipeline_writedata[15:8],io_bus_response_bits_data[7:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_28 = {io_bus_response_bits_data[31:24],io_pipeline_writedata[23:16],io_bus_response_bits_data[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_31 = {io_pipeline_writedata[31:24],io_bus_response_bits_data[23:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_4 = io_pipeline_address[1:0] == 2'h2 ? _T_28 : _T_31; // @[memory-combin-ports.scala 90:38 91:23 93:23]
  wire [31:0] _GEN_5 = io_pipeline_address[1:0] == 2'h1 ? _T_22 : _GEN_4; // @[memory-combin-ports.scala 88:38 89:23]
  wire [31:0] _GEN_6 = io_pipeline_address[1:0] == 2'h0 ? _T_16 : _GEN_5; // @[memory-combin-ports.scala 86:32 87:23]
  wire [31:0] _T_35 = {io_bus_response_bits_data[31:16],io_pipeline_writedata[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_38 = {io_pipeline_writedata[31:16],io_bus_response_bits_data[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_7 = _T_13 ? _T_35 : _T_38; // @[memory-combin-ports.scala 96:33 97:23 99:23]
  wire [31:0] _GEN_8 = io_pipeline_maskmode == 2'h0 ? _GEN_6 : _GEN_7; // @[memory-combin-ports.scala 85:45]
  wire [5:0] _T_43 = io_pipeline_address[1:0] * 4'h8; // @[memory-combin-ports.scala 116:64]
  wire [31:0] _T_44 = io_bus_response_bits_data >> _T_43; // @[memory-combin-ports.scala 116:53]
  wire [31:0] _T_45 = _T_44 & 32'hff; // @[memory-combin-ports.scala 116:72]
  wire  _T_46 = io_pipeline_maskmode == 2'h1; // @[memory-combin-ports.scala 117:41]
  wire [31:0] _T_49 = _T_44 & 32'hffff; // @[memory-combin-ports.scala 119:72]
  wire [31:0] _GEN_10 = io_pipeline_maskmode == 2'h1 ? _T_49 : io_bus_response_bits_data; // @[memory-combin-ports.scala 117:50 119:23 121:23]
  wire [31:0] _GEN_11 = _T_12 ? _T_45 : _GEN_10; // @[memory-combin-ports.scala 114:43 116:23]
  wire [23:0] _T_53 = _GEN_11[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_55 = {_T_53,_GEN_11[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_59 = _GEN_11[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_61 = {_T_59,_GEN_11[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_12 = _T_46 ? _T_61 : _GEN_11; // @[memory-combin-ports.scala 128:52 130:30 133:30]
  wire [31:0] _GEN_13 = _T_12 ? _T_55 : _GEN_12; // @[memory-combin-ports.scala 125:45 127:30]
  wire [31:0] _GEN_14 = io_pipeline_sext ? _GEN_13 : _GEN_11; // @[memory-combin-ports.scala 124:31 136:28]
  wire [31:0] _GEN_15 = io_pipeline_memread ? _GEN_14 : 32'h0; // @[memory-combin-ports.scala 108:39 139:28 base-memory-components.scala 69:15]
  wire [31:0] _GEN_17 = io_pipeline_memwrite ? 32'h0 : _GEN_15; // @[base-memory-components.scala 69:15 memory-combin-ports.scala 72:33]
  assign io_pipeline_readdata = io_bus_response_valid ? _GEN_17 : 32'h0; // @[base-memory-components.scala 69:15 memory-combin-ports.scala 71:32]
  assign io_bus_request_valid = io_pipeline_valid & (io_pipeline_memread | io_pipeline_memwrite); // @[memory-combin-ports.scala 44:27]
  assign io_bus_request_bits_address = io_pipeline_address; // @[memory-combin-ports.scala 44:77 48:33]
  assign io_bus_request_bits_writedata = io_pipeline_maskmode != 2'h2 ? _GEN_8 : io_pipeline_writedata; // @[memory-combin-ports.scala 104:19 77:43]
  assign io_bus_request_bits_operation = io_pipeline_memwrite ? 2'h2 : 2'h0; // @[memory-combin-ports.scala 51:33 60:37 63:37]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~(io_pipeline_memread & io_pipeline_memwrite) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at memory-combin-ports.scala:46 assert(!(io.pipeline.memread && io.pipeline.memwrite))\n"
            ); // @[memory-combin-ports.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~(io_pipeline_memread & io_pipeline_memwrite) | reset)) begin
          $fatal; // @[memory-combin-ports.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Dino128Core(
  input   clock,
  input   reset,
  output  io_success
);
  wire  cpu0_clock; // @[top.scala 12:20]
  wire  cpu0_reset; // @[top.scala 12:20]
  wire [31:0] cpu0_io_imem_address; // @[top.scala 12:20]
  wire [31:0] cpu0_io_imem_instruction; // @[top.scala 12:20]
  wire [31:0] cpu0_io_dmem_address; // @[top.scala 12:20]
  wire  cpu0_io_dmem_valid; // @[top.scala 12:20]
  wire [31:0] cpu0_io_dmem_writedata; // @[top.scala 12:20]
  wire  cpu0_io_dmem_memread; // @[top.scala 12:20]
  wire  cpu0_io_dmem_memwrite; // @[top.scala 12:20]
  wire [1:0] cpu0_io_dmem_maskmode; // @[top.scala 12:20]
  wire  cpu0_io_dmem_sext; // @[top.scala 12:20]
  wire [31:0] cpu0_io_dmem_readdata; // @[top.scala 12:20]
  wire  mem0_clock; // @[top.scala 13:20]
  wire  mem0_reset; // @[top.scala 13:20]
  wire [31:0] mem0_io_imem_request_bits_address; // @[top.scala 13:20]
  wire [31:0] mem0_io_imem_response_bits_data; // @[top.scala 13:20]
  wire  mem0_io_dmem_request_valid; // @[top.scala 13:20]
  wire [31:0] mem0_io_dmem_request_bits_address; // @[top.scala 13:20]
  wire [31:0] mem0_io_dmem_request_bits_writedata; // @[top.scala 13:20]
  wire [1:0] mem0_io_dmem_request_bits_operation; // @[top.scala 13:20]
  wire  mem0_io_dmem_response_valid; // @[top.scala 13:20]
  wire [31:0] mem0_io_dmem_response_bits_data; // @[top.scala 13:20]
  wire [31:0] imem0_io_pipeline_address; // @[top.scala 14:21]
  wire [31:0] imem0_io_pipeline_instruction; // @[top.scala 14:21]
  wire [31:0] imem0_io_bus_request_bits_address; // @[top.scala 14:21]
  wire [31:0] imem0_io_bus_response_bits_data; // @[top.scala 14:21]
  wire  dmem0_clock; // @[top.scala 15:21]
  wire  dmem0_reset; // @[top.scala 15:21]
  wire [31:0] dmem0_io_pipeline_address; // @[top.scala 15:21]
  wire  dmem0_io_pipeline_valid; // @[top.scala 15:21]
  wire [31:0] dmem0_io_pipeline_writedata; // @[top.scala 15:21]
  wire  dmem0_io_pipeline_memread; // @[top.scala 15:21]
  wire  dmem0_io_pipeline_memwrite; // @[top.scala 15:21]
  wire [1:0] dmem0_io_pipeline_maskmode; // @[top.scala 15:21]
  wire  dmem0_io_pipeline_sext; // @[top.scala 15:21]
  wire [31:0] dmem0_io_pipeline_readdata; // @[top.scala 15:21]
  wire  dmem0_io_bus_request_valid; // @[top.scala 15:21]
  wire [31:0] dmem0_io_bus_request_bits_address; // @[top.scala 15:21]
  wire [31:0] dmem0_io_bus_request_bits_writedata; // @[top.scala 15:21]
  wire [1:0] dmem0_io_bus_request_bits_operation; // @[top.scala 15:21]
  wire  dmem0_io_bus_response_valid; // @[top.scala 15:21]
  wire [31:0] dmem0_io_bus_response_bits_data; // @[top.scala 15:21]
  wire  cpu1_clock; // @[top.scala 19:20]
  wire  cpu1_reset; // @[top.scala 19:20]
  wire [31:0] cpu1_io_imem_address; // @[top.scala 19:20]
  wire [31:0] cpu1_io_imem_instruction; // @[top.scala 19:20]
  wire [31:0] cpu1_io_dmem_address; // @[top.scala 19:20]
  wire  cpu1_io_dmem_valid; // @[top.scala 19:20]
  wire [31:0] cpu1_io_dmem_writedata; // @[top.scala 19:20]
  wire  cpu1_io_dmem_memread; // @[top.scala 19:20]
  wire  cpu1_io_dmem_memwrite; // @[top.scala 19:20]
  wire [1:0] cpu1_io_dmem_maskmode; // @[top.scala 19:20]
  wire  cpu1_io_dmem_sext; // @[top.scala 19:20]
  wire [31:0] cpu1_io_dmem_readdata; // @[top.scala 19:20]
  wire  mem1_clock; // @[top.scala 20:20]
  wire  mem1_reset; // @[top.scala 20:20]
  wire [31:0] mem1_io_imem_request_bits_address; // @[top.scala 20:20]
  wire [31:0] mem1_io_imem_response_bits_data; // @[top.scala 20:20]
  wire  mem1_io_dmem_request_valid; // @[top.scala 20:20]
  wire [31:0] mem1_io_dmem_request_bits_address; // @[top.scala 20:20]
  wire [31:0] mem1_io_dmem_request_bits_writedata; // @[top.scala 20:20]
  wire [1:0] mem1_io_dmem_request_bits_operation; // @[top.scala 20:20]
  wire  mem1_io_dmem_response_valid; // @[top.scala 20:20]
  wire [31:0] mem1_io_dmem_response_bits_data; // @[top.scala 20:20]
  wire [31:0] imem1_io_pipeline_address; // @[top.scala 21:21]
  wire [31:0] imem1_io_pipeline_instruction; // @[top.scala 21:21]
  wire [31:0] imem1_io_bus_request_bits_address; // @[top.scala 21:21]
  wire [31:0] imem1_io_bus_response_bits_data; // @[top.scala 21:21]
  wire  dmem1_clock; // @[top.scala 22:21]
  wire  dmem1_reset; // @[top.scala 22:21]
  wire [31:0] dmem1_io_pipeline_address; // @[top.scala 22:21]
  wire  dmem1_io_pipeline_valid; // @[top.scala 22:21]
  wire [31:0] dmem1_io_pipeline_writedata; // @[top.scala 22:21]
  wire  dmem1_io_pipeline_memread; // @[top.scala 22:21]
  wire  dmem1_io_pipeline_memwrite; // @[top.scala 22:21]
  wire [1:0] dmem1_io_pipeline_maskmode; // @[top.scala 22:21]
  wire  dmem1_io_pipeline_sext; // @[top.scala 22:21]
  wire [31:0] dmem1_io_pipeline_readdata; // @[top.scala 22:21]
  wire  dmem1_io_bus_request_valid; // @[top.scala 22:21]
  wire [31:0] dmem1_io_bus_request_bits_address; // @[top.scala 22:21]
  wire [31:0] dmem1_io_bus_request_bits_writedata; // @[top.scala 22:21]
  wire [1:0] dmem1_io_bus_request_bits_operation; // @[top.scala 22:21]
  wire  dmem1_io_bus_response_valid; // @[top.scala 22:21]
  wire [31:0] dmem1_io_bus_response_bits_data; // @[top.scala 22:21]
  wire  cpu2_clock; // @[top.scala 26:20]
  wire  cpu2_reset; // @[top.scala 26:20]
  wire [31:0] cpu2_io_imem_address; // @[top.scala 26:20]
  wire [31:0] cpu2_io_imem_instruction; // @[top.scala 26:20]
  wire [31:0] cpu2_io_dmem_address; // @[top.scala 26:20]
  wire  cpu2_io_dmem_valid; // @[top.scala 26:20]
  wire [31:0] cpu2_io_dmem_writedata; // @[top.scala 26:20]
  wire  cpu2_io_dmem_memread; // @[top.scala 26:20]
  wire  cpu2_io_dmem_memwrite; // @[top.scala 26:20]
  wire [1:0] cpu2_io_dmem_maskmode; // @[top.scala 26:20]
  wire  cpu2_io_dmem_sext; // @[top.scala 26:20]
  wire [31:0] cpu2_io_dmem_readdata; // @[top.scala 26:20]
  wire  mem2_clock; // @[top.scala 27:20]
  wire  mem2_reset; // @[top.scala 27:20]
  wire [31:0] mem2_io_imem_request_bits_address; // @[top.scala 27:20]
  wire [31:0] mem2_io_imem_response_bits_data; // @[top.scala 27:20]
  wire  mem2_io_dmem_request_valid; // @[top.scala 27:20]
  wire [31:0] mem2_io_dmem_request_bits_address; // @[top.scala 27:20]
  wire [31:0] mem2_io_dmem_request_bits_writedata; // @[top.scala 27:20]
  wire [1:0] mem2_io_dmem_request_bits_operation; // @[top.scala 27:20]
  wire  mem2_io_dmem_response_valid; // @[top.scala 27:20]
  wire [31:0] mem2_io_dmem_response_bits_data; // @[top.scala 27:20]
  wire [31:0] imem2_io_pipeline_address; // @[top.scala 28:21]
  wire [31:0] imem2_io_pipeline_instruction; // @[top.scala 28:21]
  wire [31:0] imem2_io_bus_request_bits_address; // @[top.scala 28:21]
  wire [31:0] imem2_io_bus_response_bits_data; // @[top.scala 28:21]
  wire  dmem2_clock; // @[top.scala 29:21]
  wire  dmem2_reset; // @[top.scala 29:21]
  wire [31:0] dmem2_io_pipeline_address; // @[top.scala 29:21]
  wire  dmem2_io_pipeline_valid; // @[top.scala 29:21]
  wire [31:0] dmem2_io_pipeline_writedata; // @[top.scala 29:21]
  wire  dmem2_io_pipeline_memread; // @[top.scala 29:21]
  wire  dmem2_io_pipeline_memwrite; // @[top.scala 29:21]
  wire [1:0] dmem2_io_pipeline_maskmode; // @[top.scala 29:21]
  wire  dmem2_io_pipeline_sext; // @[top.scala 29:21]
  wire [31:0] dmem2_io_pipeline_readdata; // @[top.scala 29:21]
  wire  dmem2_io_bus_request_valid; // @[top.scala 29:21]
  wire [31:0] dmem2_io_bus_request_bits_address; // @[top.scala 29:21]
  wire [31:0] dmem2_io_bus_request_bits_writedata; // @[top.scala 29:21]
  wire [1:0] dmem2_io_bus_request_bits_operation; // @[top.scala 29:21]
  wire  dmem2_io_bus_response_valid; // @[top.scala 29:21]
  wire [31:0] dmem2_io_bus_response_bits_data; // @[top.scala 29:21]
  wire  cpu3_clock; // @[top.scala 33:20]
  wire  cpu3_reset; // @[top.scala 33:20]
  wire [31:0] cpu3_io_imem_address; // @[top.scala 33:20]
  wire [31:0] cpu3_io_imem_instruction; // @[top.scala 33:20]
  wire [31:0] cpu3_io_dmem_address; // @[top.scala 33:20]
  wire  cpu3_io_dmem_valid; // @[top.scala 33:20]
  wire [31:0] cpu3_io_dmem_writedata; // @[top.scala 33:20]
  wire  cpu3_io_dmem_memread; // @[top.scala 33:20]
  wire  cpu3_io_dmem_memwrite; // @[top.scala 33:20]
  wire [1:0] cpu3_io_dmem_maskmode; // @[top.scala 33:20]
  wire  cpu3_io_dmem_sext; // @[top.scala 33:20]
  wire [31:0] cpu3_io_dmem_readdata; // @[top.scala 33:20]
  wire  mem3_clock; // @[top.scala 34:20]
  wire  mem3_reset; // @[top.scala 34:20]
  wire [31:0] mem3_io_imem_request_bits_address; // @[top.scala 34:20]
  wire [31:0] mem3_io_imem_response_bits_data; // @[top.scala 34:20]
  wire  mem3_io_dmem_request_valid; // @[top.scala 34:20]
  wire [31:0] mem3_io_dmem_request_bits_address; // @[top.scala 34:20]
  wire [31:0] mem3_io_dmem_request_bits_writedata; // @[top.scala 34:20]
  wire [1:0] mem3_io_dmem_request_bits_operation; // @[top.scala 34:20]
  wire  mem3_io_dmem_response_valid; // @[top.scala 34:20]
  wire [31:0] mem3_io_dmem_response_bits_data; // @[top.scala 34:20]
  wire [31:0] imem3_io_pipeline_address; // @[top.scala 35:21]
  wire [31:0] imem3_io_pipeline_instruction; // @[top.scala 35:21]
  wire [31:0] imem3_io_bus_request_bits_address; // @[top.scala 35:21]
  wire [31:0] imem3_io_bus_response_bits_data; // @[top.scala 35:21]
  wire  dmem3_clock; // @[top.scala 36:21]
  wire  dmem3_reset; // @[top.scala 36:21]
  wire [31:0] dmem3_io_pipeline_address; // @[top.scala 36:21]
  wire  dmem3_io_pipeline_valid; // @[top.scala 36:21]
  wire [31:0] dmem3_io_pipeline_writedata; // @[top.scala 36:21]
  wire  dmem3_io_pipeline_memread; // @[top.scala 36:21]
  wire  dmem3_io_pipeline_memwrite; // @[top.scala 36:21]
  wire [1:0] dmem3_io_pipeline_maskmode; // @[top.scala 36:21]
  wire  dmem3_io_pipeline_sext; // @[top.scala 36:21]
  wire [31:0] dmem3_io_pipeline_readdata; // @[top.scala 36:21]
  wire  dmem3_io_bus_request_valid; // @[top.scala 36:21]
  wire [31:0] dmem3_io_bus_request_bits_address; // @[top.scala 36:21]
  wire [31:0] dmem3_io_bus_request_bits_writedata; // @[top.scala 36:21]
  wire [1:0] dmem3_io_bus_request_bits_operation; // @[top.scala 36:21]
  wire  dmem3_io_bus_response_valid; // @[top.scala 36:21]
  wire [31:0] dmem3_io_bus_response_bits_data; // @[top.scala 36:21]
  wire  cpu4_clock; // @[top.scala 40:20]
  wire  cpu4_reset; // @[top.scala 40:20]
  wire [31:0] cpu4_io_imem_address; // @[top.scala 40:20]
  wire [31:0] cpu4_io_imem_instruction; // @[top.scala 40:20]
  wire [31:0] cpu4_io_dmem_address; // @[top.scala 40:20]
  wire  cpu4_io_dmem_valid; // @[top.scala 40:20]
  wire [31:0] cpu4_io_dmem_writedata; // @[top.scala 40:20]
  wire  cpu4_io_dmem_memread; // @[top.scala 40:20]
  wire  cpu4_io_dmem_memwrite; // @[top.scala 40:20]
  wire [1:0] cpu4_io_dmem_maskmode; // @[top.scala 40:20]
  wire  cpu4_io_dmem_sext; // @[top.scala 40:20]
  wire [31:0] cpu4_io_dmem_readdata; // @[top.scala 40:20]
  wire  mem4_clock; // @[top.scala 41:20]
  wire  mem4_reset; // @[top.scala 41:20]
  wire [31:0] mem4_io_imem_request_bits_address; // @[top.scala 41:20]
  wire [31:0] mem4_io_imem_response_bits_data; // @[top.scala 41:20]
  wire  mem4_io_dmem_request_valid; // @[top.scala 41:20]
  wire [31:0] mem4_io_dmem_request_bits_address; // @[top.scala 41:20]
  wire [31:0] mem4_io_dmem_request_bits_writedata; // @[top.scala 41:20]
  wire [1:0] mem4_io_dmem_request_bits_operation; // @[top.scala 41:20]
  wire  mem4_io_dmem_response_valid; // @[top.scala 41:20]
  wire [31:0] mem4_io_dmem_response_bits_data; // @[top.scala 41:20]
  wire [31:0] imem4_io_pipeline_address; // @[top.scala 42:21]
  wire [31:0] imem4_io_pipeline_instruction; // @[top.scala 42:21]
  wire [31:0] imem4_io_bus_request_bits_address; // @[top.scala 42:21]
  wire [31:0] imem4_io_bus_response_bits_data; // @[top.scala 42:21]
  wire  dmem4_clock; // @[top.scala 43:21]
  wire  dmem4_reset; // @[top.scala 43:21]
  wire [31:0] dmem4_io_pipeline_address; // @[top.scala 43:21]
  wire  dmem4_io_pipeline_valid; // @[top.scala 43:21]
  wire [31:0] dmem4_io_pipeline_writedata; // @[top.scala 43:21]
  wire  dmem4_io_pipeline_memread; // @[top.scala 43:21]
  wire  dmem4_io_pipeline_memwrite; // @[top.scala 43:21]
  wire [1:0] dmem4_io_pipeline_maskmode; // @[top.scala 43:21]
  wire  dmem4_io_pipeline_sext; // @[top.scala 43:21]
  wire [31:0] dmem4_io_pipeline_readdata; // @[top.scala 43:21]
  wire  dmem4_io_bus_request_valid; // @[top.scala 43:21]
  wire [31:0] dmem4_io_bus_request_bits_address; // @[top.scala 43:21]
  wire [31:0] dmem4_io_bus_request_bits_writedata; // @[top.scala 43:21]
  wire [1:0] dmem4_io_bus_request_bits_operation; // @[top.scala 43:21]
  wire  dmem4_io_bus_response_valid; // @[top.scala 43:21]
  wire [31:0] dmem4_io_bus_response_bits_data; // @[top.scala 43:21]
  wire  cpu5_clock; // @[top.scala 47:20]
  wire  cpu5_reset; // @[top.scala 47:20]
  wire [31:0] cpu5_io_imem_address; // @[top.scala 47:20]
  wire [31:0] cpu5_io_imem_instruction; // @[top.scala 47:20]
  wire [31:0] cpu5_io_dmem_address; // @[top.scala 47:20]
  wire  cpu5_io_dmem_valid; // @[top.scala 47:20]
  wire [31:0] cpu5_io_dmem_writedata; // @[top.scala 47:20]
  wire  cpu5_io_dmem_memread; // @[top.scala 47:20]
  wire  cpu5_io_dmem_memwrite; // @[top.scala 47:20]
  wire [1:0] cpu5_io_dmem_maskmode; // @[top.scala 47:20]
  wire  cpu5_io_dmem_sext; // @[top.scala 47:20]
  wire [31:0] cpu5_io_dmem_readdata; // @[top.scala 47:20]
  wire  mem5_clock; // @[top.scala 48:20]
  wire  mem5_reset; // @[top.scala 48:20]
  wire [31:0] mem5_io_imem_request_bits_address; // @[top.scala 48:20]
  wire [31:0] mem5_io_imem_response_bits_data; // @[top.scala 48:20]
  wire  mem5_io_dmem_request_valid; // @[top.scala 48:20]
  wire [31:0] mem5_io_dmem_request_bits_address; // @[top.scala 48:20]
  wire [31:0] mem5_io_dmem_request_bits_writedata; // @[top.scala 48:20]
  wire [1:0] mem5_io_dmem_request_bits_operation; // @[top.scala 48:20]
  wire  mem5_io_dmem_response_valid; // @[top.scala 48:20]
  wire [31:0] mem5_io_dmem_response_bits_data; // @[top.scala 48:20]
  wire [31:0] imem5_io_pipeline_address; // @[top.scala 49:21]
  wire [31:0] imem5_io_pipeline_instruction; // @[top.scala 49:21]
  wire [31:0] imem5_io_bus_request_bits_address; // @[top.scala 49:21]
  wire [31:0] imem5_io_bus_response_bits_data; // @[top.scala 49:21]
  wire  dmem5_clock; // @[top.scala 50:21]
  wire  dmem5_reset; // @[top.scala 50:21]
  wire [31:0] dmem5_io_pipeline_address; // @[top.scala 50:21]
  wire  dmem5_io_pipeline_valid; // @[top.scala 50:21]
  wire [31:0] dmem5_io_pipeline_writedata; // @[top.scala 50:21]
  wire  dmem5_io_pipeline_memread; // @[top.scala 50:21]
  wire  dmem5_io_pipeline_memwrite; // @[top.scala 50:21]
  wire [1:0] dmem5_io_pipeline_maskmode; // @[top.scala 50:21]
  wire  dmem5_io_pipeline_sext; // @[top.scala 50:21]
  wire [31:0] dmem5_io_pipeline_readdata; // @[top.scala 50:21]
  wire  dmem5_io_bus_request_valid; // @[top.scala 50:21]
  wire [31:0] dmem5_io_bus_request_bits_address; // @[top.scala 50:21]
  wire [31:0] dmem5_io_bus_request_bits_writedata; // @[top.scala 50:21]
  wire [1:0] dmem5_io_bus_request_bits_operation; // @[top.scala 50:21]
  wire  dmem5_io_bus_response_valid; // @[top.scala 50:21]
  wire [31:0] dmem5_io_bus_response_bits_data; // @[top.scala 50:21]
  wire  cpu6_clock; // @[top.scala 54:20]
  wire  cpu6_reset; // @[top.scala 54:20]
  wire [31:0] cpu6_io_imem_address; // @[top.scala 54:20]
  wire [31:0] cpu6_io_imem_instruction; // @[top.scala 54:20]
  wire [31:0] cpu6_io_dmem_address; // @[top.scala 54:20]
  wire  cpu6_io_dmem_valid; // @[top.scala 54:20]
  wire [31:0] cpu6_io_dmem_writedata; // @[top.scala 54:20]
  wire  cpu6_io_dmem_memread; // @[top.scala 54:20]
  wire  cpu6_io_dmem_memwrite; // @[top.scala 54:20]
  wire [1:0] cpu6_io_dmem_maskmode; // @[top.scala 54:20]
  wire  cpu6_io_dmem_sext; // @[top.scala 54:20]
  wire [31:0] cpu6_io_dmem_readdata; // @[top.scala 54:20]
  wire  mem6_clock; // @[top.scala 55:20]
  wire  mem6_reset; // @[top.scala 55:20]
  wire [31:0] mem6_io_imem_request_bits_address; // @[top.scala 55:20]
  wire [31:0] mem6_io_imem_response_bits_data; // @[top.scala 55:20]
  wire  mem6_io_dmem_request_valid; // @[top.scala 55:20]
  wire [31:0] mem6_io_dmem_request_bits_address; // @[top.scala 55:20]
  wire [31:0] mem6_io_dmem_request_bits_writedata; // @[top.scala 55:20]
  wire [1:0] mem6_io_dmem_request_bits_operation; // @[top.scala 55:20]
  wire  mem6_io_dmem_response_valid; // @[top.scala 55:20]
  wire [31:0] mem6_io_dmem_response_bits_data; // @[top.scala 55:20]
  wire [31:0] imem6_io_pipeline_address; // @[top.scala 56:21]
  wire [31:0] imem6_io_pipeline_instruction; // @[top.scala 56:21]
  wire [31:0] imem6_io_bus_request_bits_address; // @[top.scala 56:21]
  wire [31:0] imem6_io_bus_response_bits_data; // @[top.scala 56:21]
  wire  dmem6_clock; // @[top.scala 57:21]
  wire  dmem6_reset; // @[top.scala 57:21]
  wire [31:0] dmem6_io_pipeline_address; // @[top.scala 57:21]
  wire  dmem6_io_pipeline_valid; // @[top.scala 57:21]
  wire [31:0] dmem6_io_pipeline_writedata; // @[top.scala 57:21]
  wire  dmem6_io_pipeline_memread; // @[top.scala 57:21]
  wire  dmem6_io_pipeline_memwrite; // @[top.scala 57:21]
  wire [1:0] dmem6_io_pipeline_maskmode; // @[top.scala 57:21]
  wire  dmem6_io_pipeline_sext; // @[top.scala 57:21]
  wire [31:0] dmem6_io_pipeline_readdata; // @[top.scala 57:21]
  wire  dmem6_io_bus_request_valid; // @[top.scala 57:21]
  wire [31:0] dmem6_io_bus_request_bits_address; // @[top.scala 57:21]
  wire [31:0] dmem6_io_bus_request_bits_writedata; // @[top.scala 57:21]
  wire [1:0] dmem6_io_bus_request_bits_operation; // @[top.scala 57:21]
  wire  dmem6_io_bus_response_valid; // @[top.scala 57:21]
  wire [31:0] dmem6_io_bus_response_bits_data; // @[top.scala 57:21]
  wire  cpu7_clock; // @[top.scala 61:20]
  wire  cpu7_reset; // @[top.scala 61:20]
  wire [31:0] cpu7_io_imem_address; // @[top.scala 61:20]
  wire [31:0] cpu7_io_imem_instruction; // @[top.scala 61:20]
  wire [31:0] cpu7_io_dmem_address; // @[top.scala 61:20]
  wire  cpu7_io_dmem_valid; // @[top.scala 61:20]
  wire [31:0] cpu7_io_dmem_writedata; // @[top.scala 61:20]
  wire  cpu7_io_dmem_memread; // @[top.scala 61:20]
  wire  cpu7_io_dmem_memwrite; // @[top.scala 61:20]
  wire [1:0] cpu7_io_dmem_maskmode; // @[top.scala 61:20]
  wire  cpu7_io_dmem_sext; // @[top.scala 61:20]
  wire [31:0] cpu7_io_dmem_readdata; // @[top.scala 61:20]
  wire  mem7_clock; // @[top.scala 62:20]
  wire  mem7_reset; // @[top.scala 62:20]
  wire [31:0] mem7_io_imem_request_bits_address; // @[top.scala 62:20]
  wire [31:0] mem7_io_imem_response_bits_data; // @[top.scala 62:20]
  wire  mem7_io_dmem_request_valid; // @[top.scala 62:20]
  wire [31:0] mem7_io_dmem_request_bits_address; // @[top.scala 62:20]
  wire [31:0] mem7_io_dmem_request_bits_writedata; // @[top.scala 62:20]
  wire [1:0] mem7_io_dmem_request_bits_operation; // @[top.scala 62:20]
  wire  mem7_io_dmem_response_valid; // @[top.scala 62:20]
  wire [31:0] mem7_io_dmem_response_bits_data; // @[top.scala 62:20]
  wire [31:0] imem7_io_pipeline_address; // @[top.scala 63:21]
  wire [31:0] imem7_io_pipeline_instruction; // @[top.scala 63:21]
  wire [31:0] imem7_io_bus_request_bits_address; // @[top.scala 63:21]
  wire [31:0] imem7_io_bus_response_bits_data; // @[top.scala 63:21]
  wire  dmem7_clock; // @[top.scala 64:21]
  wire  dmem7_reset; // @[top.scala 64:21]
  wire [31:0] dmem7_io_pipeline_address; // @[top.scala 64:21]
  wire  dmem7_io_pipeline_valid; // @[top.scala 64:21]
  wire [31:0] dmem7_io_pipeline_writedata; // @[top.scala 64:21]
  wire  dmem7_io_pipeline_memread; // @[top.scala 64:21]
  wire  dmem7_io_pipeline_memwrite; // @[top.scala 64:21]
  wire [1:0] dmem7_io_pipeline_maskmode; // @[top.scala 64:21]
  wire  dmem7_io_pipeline_sext; // @[top.scala 64:21]
  wire [31:0] dmem7_io_pipeline_readdata; // @[top.scala 64:21]
  wire  dmem7_io_bus_request_valid; // @[top.scala 64:21]
  wire [31:0] dmem7_io_bus_request_bits_address; // @[top.scala 64:21]
  wire [31:0] dmem7_io_bus_request_bits_writedata; // @[top.scala 64:21]
  wire [1:0] dmem7_io_bus_request_bits_operation; // @[top.scala 64:21]
  wire  dmem7_io_bus_response_valid; // @[top.scala 64:21]
  wire [31:0] dmem7_io_bus_response_bits_data; // @[top.scala 64:21]
  wire  cpu8_clock; // @[top.scala 68:20]
  wire  cpu8_reset; // @[top.scala 68:20]
  wire [31:0] cpu8_io_imem_address; // @[top.scala 68:20]
  wire [31:0] cpu8_io_imem_instruction; // @[top.scala 68:20]
  wire [31:0] cpu8_io_dmem_address; // @[top.scala 68:20]
  wire  cpu8_io_dmem_valid; // @[top.scala 68:20]
  wire [31:0] cpu8_io_dmem_writedata; // @[top.scala 68:20]
  wire  cpu8_io_dmem_memread; // @[top.scala 68:20]
  wire  cpu8_io_dmem_memwrite; // @[top.scala 68:20]
  wire [1:0] cpu8_io_dmem_maskmode; // @[top.scala 68:20]
  wire  cpu8_io_dmem_sext; // @[top.scala 68:20]
  wire [31:0] cpu8_io_dmem_readdata; // @[top.scala 68:20]
  wire  mem8_clock; // @[top.scala 69:20]
  wire  mem8_reset; // @[top.scala 69:20]
  wire [31:0] mem8_io_imem_request_bits_address; // @[top.scala 69:20]
  wire [31:0] mem8_io_imem_response_bits_data; // @[top.scala 69:20]
  wire  mem8_io_dmem_request_valid; // @[top.scala 69:20]
  wire [31:0] mem8_io_dmem_request_bits_address; // @[top.scala 69:20]
  wire [31:0] mem8_io_dmem_request_bits_writedata; // @[top.scala 69:20]
  wire [1:0] mem8_io_dmem_request_bits_operation; // @[top.scala 69:20]
  wire  mem8_io_dmem_response_valid; // @[top.scala 69:20]
  wire [31:0] mem8_io_dmem_response_bits_data; // @[top.scala 69:20]
  wire [31:0] imem8_io_pipeline_address; // @[top.scala 70:21]
  wire [31:0] imem8_io_pipeline_instruction; // @[top.scala 70:21]
  wire [31:0] imem8_io_bus_request_bits_address; // @[top.scala 70:21]
  wire [31:0] imem8_io_bus_response_bits_data; // @[top.scala 70:21]
  wire  dmem8_clock; // @[top.scala 71:21]
  wire  dmem8_reset; // @[top.scala 71:21]
  wire [31:0] dmem8_io_pipeline_address; // @[top.scala 71:21]
  wire  dmem8_io_pipeline_valid; // @[top.scala 71:21]
  wire [31:0] dmem8_io_pipeline_writedata; // @[top.scala 71:21]
  wire  dmem8_io_pipeline_memread; // @[top.scala 71:21]
  wire  dmem8_io_pipeline_memwrite; // @[top.scala 71:21]
  wire [1:0] dmem8_io_pipeline_maskmode; // @[top.scala 71:21]
  wire  dmem8_io_pipeline_sext; // @[top.scala 71:21]
  wire [31:0] dmem8_io_pipeline_readdata; // @[top.scala 71:21]
  wire  dmem8_io_bus_request_valid; // @[top.scala 71:21]
  wire [31:0] dmem8_io_bus_request_bits_address; // @[top.scala 71:21]
  wire [31:0] dmem8_io_bus_request_bits_writedata; // @[top.scala 71:21]
  wire [1:0] dmem8_io_bus_request_bits_operation; // @[top.scala 71:21]
  wire  dmem8_io_bus_response_valid; // @[top.scala 71:21]
  wire [31:0] dmem8_io_bus_response_bits_data; // @[top.scala 71:21]
  wire  cpu9_clock; // @[top.scala 75:20]
  wire  cpu9_reset; // @[top.scala 75:20]
  wire [31:0] cpu9_io_imem_address; // @[top.scala 75:20]
  wire [31:0] cpu9_io_imem_instruction; // @[top.scala 75:20]
  wire [31:0] cpu9_io_dmem_address; // @[top.scala 75:20]
  wire  cpu9_io_dmem_valid; // @[top.scala 75:20]
  wire [31:0] cpu9_io_dmem_writedata; // @[top.scala 75:20]
  wire  cpu9_io_dmem_memread; // @[top.scala 75:20]
  wire  cpu9_io_dmem_memwrite; // @[top.scala 75:20]
  wire [1:0] cpu9_io_dmem_maskmode; // @[top.scala 75:20]
  wire  cpu9_io_dmem_sext; // @[top.scala 75:20]
  wire [31:0] cpu9_io_dmem_readdata; // @[top.scala 75:20]
  wire  mem9_clock; // @[top.scala 76:20]
  wire  mem9_reset; // @[top.scala 76:20]
  wire [31:0] mem9_io_imem_request_bits_address; // @[top.scala 76:20]
  wire [31:0] mem9_io_imem_response_bits_data; // @[top.scala 76:20]
  wire  mem9_io_dmem_request_valid; // @[top.scala 76:20]
  wire [31:0] mem9_io_dmem_request_bits_address; // @[top.scala 76:20]
  wire [31:0] mem9_io_dmem_request_bits_writedata; // @[top.scala 76:20]
  wire [1:0] mem9_io_dmem_request_bits_operation; // @[top.scala 76:20]
  wire  mem9_io_dmem_response_valid; // @[top.scala 76:20]
  wire [31:0] mem9_io_dmem_response_bits_data; // @[top.scala 76:20]
  wire [31:0] imem9_io_pipeline_address; // @[top.scala 77:21]
  wire [31:0] imem9_io_pipeline_instruction; // @[top.scala 77:21]
  wire [31:0] imem9_io_bus_request_bits_address; // @[top.scala 77:21]
  wire [31:0] imem9_io_bus_response_bits_data; // @[top.scala 77:21]
  wire  dmem9_clock; // @[top.scala 78:21]
  wire  dmem9_reset; // @[top.scala 78:21]
  wire [31:0] dmem9_io_pipeline_address; // @[top.scala 78:21]
  wire  dmem9_io_pipeline_valid; // @[top.scala 78:21]
  wire [31:0] dmem9_io_pipeline_writedata; // @[top.scala 78:21]
  wire  dmem9_io_pipeline_memread; // @[top.scala 78:21]
  wire  dmem9_io_pipeline_memwrite; // @[top.scala 78:21]
  wire [1:0] dmem9_io_pipeline_maskmode; // @[top.scala 78:21]
  wire  dmem9_io_pipeline_sext; // @[top.scala 78:21]
  wire [31:0] dmem9_io_pipeline_readdata; // @[top.scala 78:21]
  wire  dmem9_io_bus_request_valid; // @[top.scala 78:21]
  wire [31:0] dmem9_io_bus_request_bits_address; // @[top.scala 78:21]
  wire [31:0] dmem9_io_bus_request_bits_writedata; // @[top.scala 78:21]
  wire [1:0] dmem9_io_bus_request_bits_operation; // @[top.scala 78:21]
  wire  dmem9_io_bus_response_valid; // @[top.scala 78:21]
  wire [31:0] dmem9_io_bus_response_bits_data; // @[top.scala 78:21]
  wire  cpu10_clock; // @[top.scala 82:21]
  wire  cpu10_reset; // @[top.scala 82:21]
  wire [31:0] cpu10_io_imem_address; // @[top.scala 82:21]
  wire [31:0] cpu10_io_imem_instruction; // @[top.scala 82:21]
  wire [31:0] cpu10_io_dmem_address; // @[top.scala 82:21]
  wire  cpu10_io_dmem_valid; // @[top.scala 82:21]
  wire [31:0] cpu10_io_dmem_writedata; // @[top.scala 82:21]
  wire  cpu10_io_dmem_memread; // @[top.scala 82:21]
  wire  cpu10_io_dmem_memwrite; // @[top.scala 82:21]
  wire [1:0] cpu10_io_dmem_maskmode; // @[top.scala 82:21]
  wire  cpu10_io_dmem_sext; // @[top.scala 82:21]
  wire [31:0] cpu10_io_dmem_readdata; // @[top.scala 82:21]
  wire  mem10_clock; // @[top.scala 83:21]
  wire  mem10_reset; // @[top.scala 83:21]
  wire [31:0] mem10_io_imem_request_bits_address; // @[top.scala 83:21]
  wire [31:0] mem10_io_imem_response_bits_data; // @[top.scala 83:21]
  wire  mem10_io_dmem_request_valid; // @[top.scala 83:21]
  wire [31:0] mem10_io_dmem_request_bits_address; // @[top.scala 83:21]
  wire [31:0] mem10_io_dmem_request_bits_writedata; // @[top.scala 83:21]
  wire [1:0] mem10_io_dmem_request_bits_operation; // @[top.scala 83:21]
  wire  mem10_io_dmem_response_valid; // @[top.scala 83:21]
  wire [31:0] mem10_io_dmem_response_bits_data; // @[top.scala 83:21]
  wire [31:0] imem10_io_pipeline_address; // @[top.scala 84:22]
  wire [31:0] imem10_io_pipeline_instruction; // @[top.scala 84:22]
  wire [31:0] imem10_io_bus_request_bits_address; // @[top.scala 84:22]
  wire [31:0] imem10_io_bus_response_bits_data; // @[top.scala 84:22]
  wire  dmem10_clock; // @[top.scala 85:22]
  wire  dmem10_reset; // @[top.scala 85:22]
  wire [31:0] dmem10_io_pipeline_address; // @[top.scala 85:22]
  wire  dmem10_io_pipeline_valid; // @[top.scala 85:22]
  wire [31:0] dmem10_io_pipeline_writedata; // @[top.scala 85:22]
  wire  dmem10_io_pipeline_memread; // @[top.scala 85:22]
  wire  dmem10_io_pipeline_memwrite; // @[top.scala 85:22]
  wire [1:0] dmem10_io_pipeline_maskmode; // @[top.scala 85:22]
  wire  dmem10_io_pipeline_sext; // @[top.scala 85:22]
  wire [31:0] dmem10_io_pipeline_readdata; // @[top.scala 85:22]
  wire  dmem10_io_bus_request_valid; // @[top.scala 85:22]
  wire [31:0] dmem10_io_bus_request_bits_address; // @[top.scala 85:22]
  wire [31:0] dmem10_io_bus_request_bits_writedata; // @[top.scala 85:22]
  wire [1:0] dmem10_io_bus_request_bits_operation; // @[top.scala 85:22]
  wire  dmem10_io_bus_response_valid; // @[top.scala 85:22]
  wire [31:0] dmem10_io_bus_response_bits_data; // @[top.scala 85:22]
  wire  cpu11_clock; // @[top.scala 89:21]
  wire  cpu11_reset; // @[top.scala 89:21]
  wire [31:0] cpu11_io_imem_address; // @[top.scala 89:21]
  wire [31:0] cpu11_io_imem_instruction; // @[top.scala 89:21]
  wire [31:0] cpu11_io_dmem_address; // @[top.scala 89:21]
  wire  cpu11_io_dmem_valid; // @[top.scala 89:21]
  wire [31:0] cpu11_io_dmem_writedata; // @[top.scala 89:21]
  wire  cpu11_io_dmem_memread; // @[top.scala 89:21]
  wire  cpu11_io_dmem_memwrite; // @[top.scala 89:21]
  wire [1:0] cpu11_io_dmem_maskmode; // @[top.scala 89:21]
  wire  cpu11_io_dmem_sext; // @[top.scala 89:21]
  wire [31:0] cpu11_io_dmem_readdata; // @[top.scala 89:21]
  wire  mem11_clock; // @[top.scala 90:21]
  wire  mem11_reset; // @[top.scala 90:21]
  wire [31:0] mem11_io_imem_request_bits_address; // @[top.scala 90:21]
  wire [31:0] mem11_io_imem_response_bits_data; // @[top.scala 90:21]
  wire  mem11_io_dmem_request_valid; // @[top.scala 90:21]
  wire [31:0] mem11_io_dmem_request_bits_address; // @[top.scala 90:21]
  wire [31:0] mem11_io_dmem_request_bits_writedata; // @[top.scala 90:21]
  wire [1:0] mem11_io_dmem_request_bits_operation; // @[top.scala 90:21]
  wire  mem11_io_dmem_response_valid; // @[top.scala 90:21]
  wire [31:0] mem11_io_dmem_response_bits_data; // @[top.scala 90:21]
  wire [31:0] imem11_io_pipeline_address; // @[top.scala 91:22]
  wire [31:0] imem11_io_pipeline_instruction; // @[top.scala 91:22]
  wire [31:0] imem11_io_bus_request_bits_address; // @[top.scala 91:22]
  wire [31:0] imem11_io_bus_response_bits_data; // @[top.scala 91:22]
  wire  dmem11_clock; // @[top.scala 92:22]
  wire  dmem11_reset; // @[top.scala 92:22]
  wire [31:0] dmem11_io_pipeline_address; // @[top.scala 92:22]
  wire  dmem11_io_pipeline_valid; // @[top.scala 92:22]
  wire [31:0] dmem11_io_pipeline_writedata; // @[top.scala 92:22]
  wire  dmem11_io_pipeline_memread; // @[top.scala 92:22]
  wire  dmem11_io_pipeline_memwrite; // @[top.scala 92:22]
  wire [1:0] dmem11_io_pipeline_maskmode; // @[top.scala 92:22]
  wire  dmem11_io_pipeline_sext; // @[top.scala 92:22]
  wire [31:0] dmem11_io_pipeline_readdata; // @[top.scala 92:22]
  wire  dmem11_io_bus_request_valid; // @[top.scala 92:22]
  wire [31:0] dmem11_io_bus_request_bits_address; // @[top.scala 92:22]
  wire [31:0] dmem11_io_bus_request_bits_writedata; // @[top.scala 92:22]
  wire [1:0] dmem11_io_bus_request_bits_operation; // @[top.scala 92:22]
  wire  dmem11_io_bus_response_valid; // @[top.scala 92:22]
  wire [31:0] dmem11_io_bus_response_bits_data; // @[top.scala 92:22]
  wire  cpu12_clock; // @[top.scala 96:21]
  wire  cpu12_reset; // @[top.scala 96:21]
  wire [31:0] cpu12_io_imem_address; // @[top.scala 96:21]
  wire [31:0] cpu12_io_imem_instruction; // @[top.scala 96:21]
  wire [31:0] cpu12_io_dmem_address; // @[top.scala 96:21]
  wire  cpu12_io_dmem_valid; // @[top.scala 96:21]
  wire [31:0] cpu12_io_dmem_writedata; // @[top.scala 96:21]
  wire  cpu12_io_dmem_memread; // @[top.scala 96:21]
  wire  cpu12_io_dmem_memwrite; // @[top.scala 96:21]
  wire [1:0] cpu12_io_dmem_maskmode; // @[top.scala 96:21]
  wire  cpu12_io_dmem_sext; // @[top.scala 96:21]
  wire [31:0] cpu12_io_dmem_readdata; // @[top.scala 96:21]
  wire  mem12_clock; // @[top.scala 97:21]
  wire  mem12_reset; // @[top.scala 97:21]
  wire [31:0] mem12_io_imem_request_bits_address; // @[top.scala 97:21]
  wire [31:0] mem12_io_imem_response_bits_data; // @[top.scala 97:21]
  wire  mem12_io_dmem_request_valid; // @[top.scala 97:21]
  wire [31:0] mem12_io_dmem_request_bits_address; // @[top.scala 97:21]
  wire [31:0] mem12_io_dmem_request_bits_writedata; // @[top.scala 97:21]
  wire [1:0] mem12_io_dmem_request_bits_operation; // @[top.scala 97:21]
  wire  mem12_io_dmem_response_valid; // @[top.scala 97:21]
  wire [31:0] mem12_io_dmem_response_bits_data; // @[top.scala 97:21]
  wire [31:0] imem12_io_pipeline_address; // @[top.scala 98:22]
  wire [31:0] imem12_io_pipeline_instruction; // @[top.scala 98:22]
  wire [31:0] imem12_io_bus_request_bits_address; // @[top.scala 98:22]
  wire [31:0] imem12_io_bus_response_bits_data; // @[top.scala 98:22]
  wire  dmem12_clock; // @[top.scala 99:22]
  wire  dmem12_reset; // @[top.scala 99:22]
  wire [31:0] dmem12_io_pipeline_address; // @[top.scala 99:22]
  wire  dmem12_io_pipeline_valid; // @[top.scala 99:22]
  wire [31:0] dmem12_io_pipeline_writedata; // @[top.scala 99:22]
  wire  dmem12_io_pipeline_memread; // @[top.scala 99:22]
  wire  dmem12_io_pipeline_memwrite; // @[top.scala 99:22]
  wire [1:0] dmem12_io_pipeline_maskmode; // @[top.scala 99:22]
  wire  dmem12_io_pipeline_sext; // @[top.scala 99:22]
  wire [31:0] dmem12_io_pipeline_readdata; // @[top.scala 99:22]
  wire  dmem12_io_bus_request_valid; // @[top.scala 99:22]
  wire [31:0] dmem12_io_bus_request_bits_address; // @[top.scala 99:22]
  wire [31:0] dmem12_io_bus_request_bits_writedata; // @[top.scala 99:22]
  wire [1:0] dmem12_io_bus_request_bits_operation; // @[top.scala 99:22]
  wire  dmem12_io_bus_response_valid; // @[top.scala 99:22]
  wire [31:0] dmem12_io_bus_response_bits_data; // @[top.scala 99:22]
  wire  cpu13_clock; // @[top.scala 103:21]
  wire  cpu13_reset; // @[top.scala 103:21]
  wire [31:0] cpu13_io_imem_address; // @[top.scala 103:21]
  wire [31:0] cpu13_io_imem_instruction; // @[top.scala 103:21]
  wire [31:0] cpu13_io_dmem_address; // @[top.scala 103:21]
  wire  cpu13_io_dmem_valid; // @[top.scala 103:21]
  wire [31:0] cpu13_io_dmem_writedata; // @[top.scala 103:21]
  wire  cpu13_io_dmem_memread; // @[top.scala 103:21]
  wire  cpu13_io_dmem_memwrite; // @[top.scala 103:21]
  wire [1:0] cpu13_io_dmem_maskmode; // @[top.scala 103:21]
  wire  cpu13_io_dmem_sext; // @[top.scala 103:21]
  wire [31:0] cpu13_io_dmem_readdata; // @[top.scala 103:21]
  wire  mem13_clock; // @[top.scala 104:21]
  wire  mem13_reset; // @[top.scala 104:21]
  wire [31:0] mem13_io_imem_request_bits_address; // @[top.scala 104:21]
  wire [31:0] mem13_io_imem_response_bits_data; // @[top.scala 104:21]
  wire  mem13_io_dmem_request_valid; // @[top.scala 104:21]
  wire [31:0] mem13_io_dmem_request_bits_address; // @[top.scala 104:21]
  wire [31:0] mem13_io_dmem_request_bits_writedata; // @[top.scala 104:21]
  wire [1:0] mem13_io_dmem_request_bits_operation; // @[top.scala 104:21]
  wire  mem13_io_dmem_response_valid; // @[top.scala 104:21]
  wire [31:0] mem13_io_dmem_response_bits_data; // @[top.scala 104:21]
  wire [31:0] imem13_io_pipeline_address; // @[top.scala 105:22]
  wire [31:0] imem13_io_pipeline_instruction; // @[top.scala 105:22]
  wire [31:0] imem13_io_bus_request_bits_address; // @[top.scala 105:22]
  wire [31:0] imem13_io_bus_response_bits_data; // @[top.scala 105:22]
  wire  dmem13_clock; // @[top.scala 106:22]
  wire  dmem13_reset; // @[top.scala 106:22]
  wire [31:0] dmem13_io_pipeline_address; // @[top.scala 106:22]
  wire  dmem13_io_pipeline_valid; // @[top.scala 106:22]
  wire [31:0] dmem13_io_pipeline_writedata; // @[top.scala 106:22]
  wire  dmem13_io_pipeline_memread; // @[top.scala 106:22]
  wire  dmem13_io_pipeline_memwrite; // @[top.scala 106:22]
  wire [1:0] dmem13_io_pipeline_maskmode; // @[top.scala 106:22]
  wire  dmem13_io_pipeline_sext; // @[top.scala 106:22]
  wire [31:0] dmem13_io_pipeline_readdata; // @[top.scala 106:22]
  wire  dmem13_io_bus_request_valid; // @[top.scala 106:22]
  wire [31:0] dmem13_io_bus_request_bits_address; // @[top.scala 106:22]
  wire [31:0] dmem13_io_bus_request_bits_writedata; // @[top.scala 106:22]
  wire [1:0] dmem13_io_bus_request_bits_operation; // @[top.scala 106:22]
  wire  dmem13_io_bus_response_valid; // @[top.scala 106:22]
  wire [31:0] dmem13_io_bus_response_bits_data; // @[top.scala 106:22]
  wire  cpu14_clock; // @[top.scala 110:21]
  wire  cpu14_reset; // @[top.scala 110:21]
  wire [31:0] cpu14_io_imem_address; // @[top.scala 110:21]
  wire [31:0] cpu14_io_imem_instruction; // @[top.scala 110:21]
  wire [31:0] cpu14_io_dmem_address; // @[top.scala 110:21]
  wire  cpu14_io_dmem_valid; // @[top.scala 110:21]
  wire [31:0] cpu14_io_dmem_writedata; // @[top.scala 110:21]
  wire  cpu14_io_dmem_memread; // @[top.scala 110:21]
  wire  cpu14_io_dmem_memwrite; // @[top.scala 110:21]
  wire [1:0] cpu14_io_dmem_maskmode; // @[top.scala 110:21]
  wire  cpu14_io_dmem_sext; // @[top.scala 110:21]
  wire [31:0] cpu14_io_dmem_readdata; // @[top.scala 110:21]
  wire  mem14_clock; // @[top.scala 111:21]
  wire  mem14_reset; // @[top.scala 111:21]
  wire [31:0] mem14_io_imem_request_bits_address; // @[top.scala 111:21]
  wire [31:0] mem14_io_imem_response_bits_data; // @[top.scala 111:21]
  wire  mem14_io_dmem_request_valid; // @[top.scala 111:21]
  wire [31:0] mem14_io_dmem_request_bits_address; // @[top.scala 111:21]
  wire [31:0] mem14_io_dmem_request_bits_writedata; // @[top.scala 111:21]
  wire [1:0] mem14_io_dmem_request_bits_operation; // @[top.scala 111:21]
  wire  mem14_io_dmem_response_valid; // @[top.scala 111:21]
  wire [31:0] mem14_io_dmem_response_bits_data; // @[top.scala 111:21]
  wire [31:0] imem14_io_pipeline_address; // @[top.scala 112:22]
  wire [31:0] imem14_io_pipeline_instruction; // @[top.scala 112:22]
  wire [31:0] imem14_io_bus_request_bits_address; // @[top.scala 112:22]
  wire [31:0] imem14_io_bus_response_bits_data; // @[top.scala 112:22]
  wire  dmem14_clock; // @[top.scala 113:22]
  wire  dmem14_reset; // @[top.scala 113:22]
  wire [31:0] dmem14_io_pipeline_address; // @[top.scala 113:22]
  wire  dmem14_io_pipeline_valid; // @[top.scala 113:22]
  wire [31:0] dmem14_io_pipeline_writedata; // @[top.scala 113:22]
  wire  dmem14_io_pipeline_memread; // @[top.scala 113:22]
  wire  dmem14_io_pipeline_memwrite; // @[top.scala 113:22]
  wire [1:0] dmem14_io_pipeline_maskmode; // @[top.scala 113:22]
  wire  dmem14_io_pipeline_sext; // @[top.scala 113:22]
  wire [31:0] dmem14_io_pipeline_readdata; // @[top.scala 113:22]
  wire  dmem14_io_bus_request_valid; // @[top.scala 113:22]
  wire [31:0] dmem14_io_bus_request_bits_address; // @[top.scala 113:22]
  wire [31:0] dmem14_io_bus_request_bits_writedata; // @[top.scala 113:22]
  wire [1:0] dmem14_io_bus_request_bits_operation; // @[top.scala 113:22]
  wire  dmem14_io_bus_response_valid; // @[top.scala 113:22]
  wire [31:0] dmem14_io_bus_response_bits_data; // @[top.scala 113:22]
  wire  cpu15_clock; // @[top.scala 117:21]
  wire  cpu15_reset; // @[top.scala 117:21]
  wire [31:0] cpu15_io_imem_address; // @[top.scala 117:21]
  wire [31:0] cpu15_io_imem_instruction; // @[top.scala 117:21]
  wire [31:0] cpu15_io_dmem_address; // @[top.scala 117:21]
  wire  cpu15_io_dmem_valid; // @[top.scala 117:21]
  wire [31:0] cpu15_io_dmem_writedata; // @[top.scala 117:21]
  wire  cpu15_io_dmem_memread; // @[top.scala 117:21]
  wire  cpu15_io_dmem_memwrite; // @[top.scala 117:21]
  wire [1:0] cpu15_io_dmem_maskmode; // @[top.scala 117:21]
  wire  cpu15_io_dmem_sext; // @[top.scala 117:21]
  wire [31:0] cpu15_io_dmem_readdata; // @[top.scala 117:21]
  wire  mem15_clock; // @[top.scala 118:21]
  wire  mem15_reset; // @[top.scala 118:21]
  wire [31:0] mem15_io_imem_request_bits_address; // @[top.scala 118:21]
  wire [31:0] mem15_io_imem_response_bits_data; // @[top.scala 118:21]
  wire  mem15_io_dmem_request_valid; // @[top.scala 118:21]
  wire [31:0] mem15_io_dmem_request_bits_address; // @[top.scala 118:21]
  wire [31:0] mem15_io_dmem_request_bits_writedata; // @[top.scala 118:21]
  wire [1:0] mem15_io_dmem_request_bits_operation; // @[top.scala 118:21]
  wire  mem15_io_dmem_response_valid; // @[top.scala 118:21]
  wire [31:0] mem15_io_dmem_response_bits_data; // @[top.scala 118:21]
  wire [31:0] imem15_io_pipeline_address; // @[top.scala 119:22]
  wire [31:0] imem15_io_pipeline_instruction; // @[top.scala 119:22]
  wire [31:0] imem15_io_bus_request_bits_address; // @[top.scala 119:22]
  wire [31:0] imem15_io_bus_response_bits_data; // @[top.scala 119:22]
  wire  dmem15_clock; // @[top.scala 120:22]
  wire  dmem15_reset; // @[top.scala 120:22]
  wire [31:0] dmem15_io_pipeline_address; // @[top.scala 120:22]
  wire  dmem15_io_pipeline_valid; // @[top.scala 120:22]
  wire [31:0] dmem15_io_pipeline_writedata; // @[top.scala 120:22]
  wire  dmem15_io_pipeline_memread; // @[top.scala 120:22]
  wire  dmem15_io_pipeline_memwrite; // @[top.scala 120:22]
  wire [1:0] dmem15_io_pipeline_maskmode; // @[top.scala 120:22]
  wire  dmem15_io_pipeline_sext; // @[top.scala 120:22]
  wire [31:0] dmem15_io_pipeline_readdata; // @[top.scala 120:22]
  wire  dmem15_io_bus_request_valid; // @[top.scala 120:22]
  wire [31:0] dmem15_io_bus_request_bits_address; // @[top.scala 120:22]
  wire [31:0] dmem15_io_bus_request_bits_writedata; // @[top.scala 120:22]
  wire [1:0] dmem15_io_bus_request_bits_operation; // @[top.scala 120:22]
  wire  dmem15_io_bus_response_valid; // @[top.scala 120:22]
  wire [31:0] dmem15_io_bus_response_bits_data; // @[top.scala 120:22]
  wire  cpu16_clock; // @[top.scala 124:21]
  wire  cpu16_reset; // @[top.scala 124:21]
  wire [31:0] cpu16_io_imem_address; // @[top.scala 124:21]
  wire [31:0] cpu16_io_imem_instruction; // @[top.scala 124:21]
  wire [31:0] cpu16_io_dmem_address; // @[top.scala 124:21]
  wire  cpu16_io_dmem_valid; // @[top.scala 124:21]
  wire [31:0] cpu16_io_dmem_writedata; // @[top.scala 124:21]
  wire  cpu16_io_dmem_memread; // @[top.scala 124:21]
  wire  cpu16_io_dmem_memwrite; // @[top.scala 124:21]
  wire [1:0] cpu16_io_dmem_maskmode; // @[top.scala 124:21]
  wire  cpu16_io_dmem_sext; // @[top.scala 124:21]
  wire [31:0] cpu16_io_dmem_readdata; // @[top.scala 124:21]
  wire  mem16_clock; // @[top.scala 125:21]
  wire  mem16_reset; // @[top.scala 125:21]
  wire [31:0] mem16_io_imem_request_bits_address; // @[top.scala 125:21]
  wire [31:0] mem16_io_imem_response_bits_data; // @[top.scala 125:21]
  wire  mem16_io_dmem_request_valid; // @[top.scala 125:21]
  wire [31:0] mem16_io_dmem_request_bits_address; // @[top.scala 125:21]
  wire [31:0] mem16_io_dmem_request_bits_writedata; // @[top.scala 125:21]
  wire [1:0] mem16_io_dmem_request_bits_operation; // @[top.scala 125:21]
  wire  mem16_io_dmem_response_valid; // @[top.scala 125:21]
  wire [31:0] mem16_io_dmem_response_bits_data; // @[top.scala 125:21]
  wire [31:0] imem16_io_pipeline_address; // @[top.scala 126:22]
  wire [31:0] imem16_io_pipeline_instruction; // @[top.scala 126:22]
  wire [31:0] imem16_io_bus_request_bits_address; // @[top.scala 126:22]
  wire [31:0] imem16_io_bus_response_bits_data; // @[top.scala 126:22]
  wire  dmem16_clock; // @[top.scala 127:22]
  wire  dmem16_reset; // @[top.scala 127:22]
  wire [31:0] dmem16_io_pipeline_address; // @[top.scala 127:22]
  wire  dmem16_io_pipeline_valid; // @[top.scala 127:22]
  wire [31:0] dmem16_io_pipeline_writedata; // @[top.scala 127:22]
  wire  dmem16_io_pipeline_memread; // @[top.scala 127:22]
  wire  dmem16_io_pipeline_memwrite; // @[top.scala 127:22]
  wire [1:0] dmem16_io_pipeline_maskmode; // @[top.scala 127:22]
  wire  dmem16_io_pipeline_sext; // @[top.scala 127:22]
  wire [31:0] dmem16_io_pipeline_readdata; // @[top.scala 127:22]
  wire  dmem16_io_bus_request_valid; // @[top.scala 127:22]
  wire [31:0] dmem16_io_bus_request_bits_address; // @[top.scala 127:22]
  wire [31:0] dmem16_io_bus_request_bits_writedata; // @[top.scala 127:22]
  wire [1:0] dmem16_io_bus_request_bits_operation; // @[top.scala 127:22]
  wire  dmem16_io_bus_response_valid; // @[top.scala 127:22]
  wire [31:0] dmem16_io_bus_response_bits_data; // @[top.scala 127:22]
  wire  cpu17_clock; // @[top.scala 131:21]
  wire  cpu17_reset; // @[top.scala 131:21]
  wire [31:0] cpu17_io_imem_address; // @[top.scala 131:21]
  wire [31:0] cpu17_io_imem_instruction; // @[top.scala 131:21]
  wire [31:0] cpu17_io_dmem_address; // @[top.scala 131:21]
  wire  cpu17_io_dmem_valid; // @[top.scala 131:21]
  wire [31:0] cpu17_io_dmem_writedata; // @[top.scala 131:21]
  wire  cpu17_io_dmem_memread; // @[top.scala 131:21]
  wire  cpu17_io_dmem_memwrite; // @[top.scala 131:21]
  wire [1:0] cpu17_io_dmem_maskmode; // @[top.scala 131:21]
  wire  cpu17_io_dmem_sext; // @[top.scala 131:21]
  wire [31:0] cpu17_io_dmem_readdata; // @[top.scala 131:21]
  wire  mem17_clock; // @[top.scala 132:21]
  wire  mem17_reset; // @[top.scala 132:21]
  wire [31:0] mem17_io_imem_request_bits_address; // @[top.scala 132:21]
  wire [31:0] mem17_io_imem_response_bits_data; // @[top.scala 132:21]
  wire  mem17_io_dmem_request_valid; // @[top.scala 132:21]
  wire [31:0] mem17_io_dmem_request_bits_address; // @[top.scala 132:21]
  wire [31:0] mem17_io_dmem_request_bits_writedata; // @[top.scala 132:21]
  wire [1:0] mem17_io_dmem_request_bits_operation; // @[top.scala 132:21]
  wire  mem17_io_dmem_response_valid; // @[top.scala 132:21]
  wire [31:0] mem17_io_dmem_response_bits_data; // @[top.scala 132:21]
  wire [31:0] imem17_io_pipeline_address; // @[top.scala 133:22]
  wire [31:0] imem17_io_pipeline_instruction; // @[top.scala 133:22]
  wire [31:0] imem17_io_bus_request_bits_address; // @[top.scala 133:22]
  wire [31:0] imem17_io_bus_response_bits_data; // @[top.scala 133:22]
  wire  dmem17_clock; // @[top.scala 134:22]
  wire  dmem17_reset; // @[top.scala 134:22]
  wire [31:0] dmem17_io_pipeline_address; // @[top.scala 134:22]
  wire  dmem17_io_pipeline_valid; // @[top.scala 134:22]
  wire [31:0] dmem17_io_pipeline_writedata; // @[top.scala 134:22]
  wire  dmem17_io_pipeline_memread; // @[top.scala 134:22]
  wire  dmem17_io_pipeline_memwrite; // @[top.scala 134:22]
  wire [1:0] dmem17_io_pipeline_maskmode; // @[top.scala 134:22]
  wire  dmem17_io_pipeline_sext; // @[top.scala 134:22]
  wire [31:0] dmem17_io_pipeline_readdata; // @[top.scala 134:22]
  wire  dmem17_io_bus_request_valid; // @[top.scala 134:22]
  wire [31:0] dmem17_io_bus_request_bits_address; // @[top.scala 134:22]
  wire [31:0] dmem17_io_bus_request_bits_writedata; // @[top.scala 134:22]
  wire [1:0] dmem17_io_bus_request_bits_operation; // @[top.scala 134:22]
  wire  dmem17_io_bus_response_valid; // @[top.scala 134:22]
  wire [31:0] dmem17_io_bus_response_bits_data; // @[top.scala 134:22]
  wire  cpu18_clock; // @[top.scala 138:21]
  wire  cpu18_reset; // @[top.scala 138:21]
  wire [31:0] cpu18_io_imem_address; // @[top.scala 138:21]
  wire [31:0] cpu18_io_imem_instruction; // @[top.scala 138:21]
  wire [31:0] cpu18_io_dmem_address; // @[top.scala 138:21]
  wire  cpu18_io_dmem_valid; // @[top.scala 138:21]
  wire [31:0] cpu18_io_dmem_writedata; // @[top.scala 138:21]
  wire  cpu18_io_dmem_memread; // @[top.scala 138:21]
  wire  cpu18_io_dmem_memwrite; // @[top.scala 138:21]
  wire [1:0] cpu18_io_dmem_maskmode; // @[top.scala 138:21]
  wire  cpu18_io_dmem_sext; // @[top.scala 138:21]
  wire [31:0] cpu18_io_dmem_readdata; // @[top.scala 138:21]
  wire  mem18_clock; // @[top.scala 139:21]
  wire  mem18_reset; // @[top.scala 139:21]
  wire [31:0] mem18_io_imem_request_bits_address; // @[top.scala 139:21]
  wire [31:0] mem18_io_imem_response_bits_data; // @[top.scala 139:21]
  wire  mem18_io_dmem_request_valid; // @[top.scala 139:21]
  wire [31:0] mem18_io_dmem_request_bits_address; // @[top.scala 139:21]
  wire [31:0] mem18_io_dmem_request_bits_writedata; // @[top.scala 139:21]
  wire [1:0] mem18_io_dmem_request_bits_operation; // @[top.scala 139:21]
  wire  mem18_io_dmem_response_valid; // @[top.scala 139:21]
  wire [31:0] mem18_io_dmem_response_bits_data; // @[top.scala 139:21]
  wire [31:0] imem18_io_pipeline_address; // @[top.scala 140:22]
  wire [31:0] imem18_io_pipeline_instruction; // @[top.scala 140:22]
  wire [31:0] imem18_io_bus_request_bits_address; // @[top.scala 140:22]
  wire [31:0] imem18_io_bus_response_bits_data; // @[top.scala 140:22]
  wire  dmem18_clock; // @[top.scala 141:22]
  wire  dmem18_reset; // @[top.scala 141:22]
  wire [31:0] dmem18_io_pipeline_address; // @[top.scala 141:22]
  wire  dmem18_io_pipeline_valid; // @[top.scala 141:22]
  wire [31:0] dmem18_io_pipeline_writedata; // @[top.scala 141:22]
  wire  dmem18_io_pipeline_memread; // @[top.scala 141:22]
  wire  dmem18_io_pipeline_memwrite; // @[top.scala 141:22]
  wire [1:0] dmem18_io_pipeline_maskmode; // @[top.scala 141:22]
  wire  dmem18_io_pipeline_sext; // @[top.scala 141:22]
  wire [31:0] dmem18_io_pipeline_readdata; // @[top.scala 141:22]
  wire  dmem18_io_bus_request_valid; // @[top.scala 141:22]
  wire [31:0] dmem18_io_bus_request_bits_address; // @[top.scala 141:22]
  wire [31:0] dmem18_io_bus_request_bits_writedata; // @[top.scala 141:22]
  wire [1:0] dmem18_io_bus_request_bits_operation; // @[top.scala 141:22]
  wire  dmem18_io_bus_response_valid; // @[top.scala 141:22]
  wire [31:0] dmem18_io_bus_response_bits_data; // @[top.scala 141:22]
  wire  cpu19_clock; // @[top.scala 145:21]
  wire  cpu19_reset; // @[top.scala 145:21]
  wire [31:0] cpu19_io_imem_address; // @[top.scala 145:21]
  wire [31:0] cpu19_io_imem_instruction; // @[top.scala 145:21]
  wire [31:0] cpu19_io_dmem_address; // @[top.scala 145:21]
  wire  cpu19_io_dmem_valid; // @[top.scala 145:21]
  wire [31:0] cpu19_io_dmem_writedata; // @[top.scala 145:21]
  wire  cpu19_io_dmem_memread; // @[top.scala 145:21]
  wire  cpu19_io_dmem_memwrite; // @[top.scala 145:21]
  wire [1:0] cpu19_io_dmem_maskmode; // @[top.scala 145:21]
  wire  cpu19_io_dmem_sext; // @[top.scala 145:21]
  wire [31:0] cpu19_io_dmem_readdata; // @[top.scala 145:21]
  wire  mem19_clock; // @[top.scala 146:21]
  wire  mem19_reset; // @[top.scala 146:21]
  wire [31:0] mem19_io_imem_request_bits_address; // @[top.scala 146:21]
  wire [31:0] mem19_io_imem_response_bits_data; // @[top.scala 146:21]
  wire  mem19_io_dmem_request_valid; // @[top.scala 146:21]
  wire [31:0] mem19_io_dmem_request_bits_address; // @[top.scala 146:21]
  wire [31:0] mem19_io_dmem_request_bits_writedata; // @[top.scala 146:21]
  wire [1:0] mem19_io_dmem_request_bits_operation; // @[top.scala 146:21]
  wire  mem19_io_dmem_response_valid; // @[top.scala 146:21]
  wire [31:0] mem19_io_dmem_response_bits_data; // @[top.scala 146:21]
  wire [31:0] imem19_io_pipeline_address; // @[top.scala 147:22]
  wire [31:0] imem19_io_pipeline_instruction; // @[top.scala 147:22]
  wire [31:0] imem19_io_bus_request_bits_address; // @[top.scala 147:22]
  wire [31:0] imem19_io_bus_response_bits_data; // @[top.scala 147:22]
  wire  dmem19_clock; // @[top.scala 148:22]
  wire  dmem19_reset; // @[top.scala 148:22]
  wire [31:0] dmem19_io_pipeline_address; // @[top.scala 148:22]
  wire  dmem19_io_pipeline_valid; // @[top.scala 148:22]
  wire [31:0] dmem19_io_pipeline_writedata; // @[top.scala 148:22]
  wire  dmem19_io_pipeline_memread; // @[top.scala 148:22]
  wire  dmem19_io_pipeline_memwrite; // @[top.scala 148:22]
  wire [1:0] dmem19_io_pipeline_maskmode; // @[top.scala 148:22]
  wire  dmem19_io_pipeline_sext; // @[top.scala 148:22]
  wire [31:0] dmem19_io_pipeline_readdata; // @[top.scala 148:22]
  wire  dmem19_io_bus_request_valid; // @[top.scala 148:22]
  wire [31:0] dmem19_io_bus_request_bits_address; // @[top.scala 148:22]
  wire [31:0] dmem19_io_bus_request_bits_writedata; // @[top.scala 148:22]
  wire [1:0] dmem19_io_bus_request_bits_operation; // @[top.scala 148:22]
  wire  dmem19_io_bus_response_valid; // @[top.scala 148:22]
  wire [31:0] dmem19_io_bus_response_bits_data; // @[top.scala 148:22]
  wire  cpu20_clock; // @[top.scala 152:21]
  wire  cpu20_reset; // @[top.scala 152:21]
  wire [31:0] cpu20_io_imem_address; // @[top.scala 152:21]
  wire [31:0] cpu20_io_imem_instruction; // @[top.scala 152:21]
  wire [31:0] cpu20_io_dmem_address; // @[top.scala 152:21]
  wire  cpu20_io_dmem_valid; // @[top.scala 152:21]
  wire [31:0] cpu20_io_dmem_writedata; // @[top.scala 152:21]
  wire  cpu20_io_dmem_memread; // @[top.scala 152:21]
  wire  cpu20_io_dmem_memwrite; // @[top.scala 152:21]
  wire [1:0] cpu20_io_dmem_maskmode; // @[top.scala 152:21]
  wire  cpu20_io_dmem_sext; // @[top.scala 152:21]
  wire [31:0] cpu20_io_dmem_readdata; // @[top.scala 152:21]
  wire  mem20_clock; // @[top.scala 153:21]
  wire  mem20_reset; // @[top.scala 153:21]
  wire [31:0] mem20_io_imem_request_bits_address; // @[top.scala 153:21]
  wire [31:0] mem20_io_imem_response_bits_data; // @[top.scala 153:21]
  wire  mem20_io_dmem_request_valid; // @[top.scala 153:21]
  wire [31:0] mem20_io_dmem_request_bits_address; // @[top.scala 153:21]
  wire [31:0] mem20_io_dmem_request_bits_writedata; // @[top.scala 153:21]
  wire [1:0] mem20_io_dmem_request_bits_operation; // @[top.scala 153:21]
  wire  mem20_io_dmem_response_valid; // @[top.scala 153:21]
  wire [31:0] mem20_io_dmem_response_bits_data; // @[top.scala 153:21]
  wire [31:0] imem20_io_pipeline_address; // @[top.scala 154:22]
  wire [31:0] imem20_io_pipeline_instruction; // @[top.scala 154:22]
  wire [31:0] imem20_io_bus_request_bits_address; // @[top.scala 154:22]
  wire [31:0] imem20_io_bus_response_bits_data; // @[top.scala 154:22]
  wire  dmem20_clock; // @[top.scala 155:22]
  wire  dmem20_reset; // @[top.scala 155:22]
  wire [31:0] dmem20_io_pipeline_address; // @[top.scala 155:22]
  wire  dmem20_io_pipeline_valid; // @[top.scala 155:22]
  wire [31:0] dmem20_io_pipeline_writedata; // @[top.scala 155:22]
  wire  dmem20_io_pipeline_memread; // @[top.scala 155:22]
  wire  dmem20_io_pipeline_memwrite; // @[top.scala 155:22]
  wire [1:0] dmem20_io_pipeline_maskmode; // @[top.scala 155:22]
  wire  dmem20_io_pipeline_sext; // @[top.scala 155:22]
  wire [31:0] dmem20_io_pipeline_readdata; // @[top.scala 155:22]
  wire  dmem20_io_bus_request_valid; // @[top.scala 155:22]
  wire [31:0] dmem20_io_bus_request_bits_address; // @[top.scala 155:22]
  wire [31:0] dmem20_io_bus_request_bits_writedata; // @[top.scala 155:22]
  wire [1:0] dmem20_io_bus_request_bits_operation; // @[top.scala 155:22]
  wire  dmem20_io_bus_response_valid; // @[top.scala 155:22]
  wire [31:0] dmem20_io_bus_response_bits_data; // @[top.scala 155:22]
  wire  cpu21_clock; // @[top.scala 159:21]
  wire  cpu21_reset; // @[top.scala 159:21]
  wire [31:0] cpu21_io_imem_address; // @[top.scala 159:21]
  wire [31:0] cpu21_io_imem_instruction; // @[top.scala 159:21]
  wire [31:0] cpu21_io_dmem_address; // @[top.scala 159:21]
  wire  cpu21_io_dmem_valid; // @[top.scala 159:21]
  wire [31:0] cpu21_io_dmem_writedata; // @[top.scala 159:21]
  wire  cpu21_io_dmem_memread; // @[top.scala 159:21]
  wire  cpu21_io_dmem_memwrite; // @[top.scala 159:21]
  wire [1:0] cpu21_io_dmem_maskmode; // @[top.scala 159:21]
  wire  cpu21_io_dmem_sext; // @[top.scala 159:21]
  wire [31:0] cpu21_io_dmem_readdata; // @[top.scala 159:21]
  wire  mem21_clock; // @[top.scala 160:21]
  wire  mem21_reset; // @[top.scala 160:21]
  wire [31:0] mem21_io_imem_request_bits_address; // @[top.scala 160:21]
  wire [31:0] mem21_io_imem_response_bits_data; // @[top.scala 160:21]
  wire  mem21_io_dmem_request_valid; // @[top.scala 160:21]
  wire [31:0] mem21_io_dmem_request_bits_address; // @[top.scala 160:21]
  wire [31:0] mem21_io_dmem_request_bits_writedata; // @[top.scala 160:21]
  wire [1:0] mem21_io_dmem_request_bits_operation; // @[top.scala 160:21]
  wire  mem21_io_dmem_response_valid; // @[top.scala 160:21]
  wire [31:0] mem21_io_dmem_response_bits_data; // @[top.scala 160:21]
  wire [31:0] imem21_io_pipeline_address; // @[top.scala 161:22]
  wire [31:0] imem21_io_pipeline_instruction; // @[top.scala 161:22]
  wire [31:0] imem21_io_bus_request_bits_address; // @[top.scala 161:22]
  wire [31:0] imem21_io_bus_response_bits_data; // @[top.scala 161:22]
  wire  dmem21_clock; // @[top.scala 162:22]
  wire  dmem21_reset; // @[top.scala 162:22]
  wire [31:0] dmem21_io_pipeline_address; // @[top.scala 162:22]
  wire  dmem21_io_pipeline_valid; // @[top.scala 162:22]
  wire [31:0] dmem21_io_pipeline_writedata; // @[top.scala 162:22]
  wire  dmem21_io_pipeline_memread; // @[top.scala 162:22]
  wire  dmem21_io_pipeline_memwrite; // @[top.scala 162:22]
  wire [1:0] dmem21_io_pipeline_maskmode; // @[top.scala 162:22]
  wire  dmem21_io_pipeline_sext; // @[top.scala 162:22]
  wire [31:0] dmem21_io_pipeline_readdata; // @[top.scala 162:22]
  wire  dmem21_io_bus_request_valid; // @[top.scala 162:22]
  wire [31:0] dmem21_io_bus_request_bits_address; // @[top.scala 162:22]
  wire [31:0] dmem21_io_bus_request_bits_writedata; // @[top.scala 162:22]
  wire [1:0] dmem21_io_bus_request_bits_operation; // @[top.scala 162:22]
  wire  dmem21_io_bus_response_valid; // @[top.scala 162:22]
  wire [31:0] dmem21_io_bus_response_bits_data; // @[top.scala 162:22]
  wire  cpu22_clock; // @[top.scala 166:21]
  wire  cpu22_reset; // @[top.scala 166:21]
  wire [31:0] cpu22_io_imem_address; // @[top.scala 166:21]
  wire [31:0] cpu22_io_imem_instruction; // @[top.scala 166:21]
  wire [31:0] cpu22_io_dmem_address; // @[top.scala 166:21]
  wire  cpu22_io_dmem_valid; // @[top.scala 166:21]
  wire [31:0] cpu22_io_dmem_writedata; // @[top.scala 166:21]
  wire  cpu22_io_dmem_memread; // @[top.scala 166:21]
  wire  cpu22_io_dmem_memwrite; // @[top.scala 166:21]
  wire [1:0] cpu22_io_dmem_maskmode; // @[top.scala 166:21]
  wire  cpu22_io_dmem_sext; // @[top.scala 166:21]
  wire [31:0] cpu22_io_dmem_readdata; // @[top.scala 166:21]
  wire  mem22_clock; // @[top.scala 167:21]
  wire  mem22_reset; // @[top.scala 167:21]
  wire [31:0] mem22_io_imem_request_bits_address; // @[top.scala 167:21]
  wire [31:0] mem22_io_imem_response_bits_data; // @[top.scala 167:21]
  wire  mem22_io_dmem_request_valid; // @[top.scala 167:21]
  wire [31:0] mem22_io_dmem_request_bits_address; // @[top.scala 167:21]
  wire [31:0] mem22_io_dmem_request_bits_writedata; // @[top.scala 167:21]
  wire [1:0] mem22_io_dmem_request_bits_operation; // @[top.scala 167:21]
  wire  mem22_io_dmem_response_valid; // @[top.scala 167:21]
  wire [31:0] mem22_io_dmem_response_bits_data; // @[top.scala 167:21]
  wire [31:0] imem22_io_pipeline_address; // @[top.scala 168:22]
  wire [31:0] imem22_io_pipeline_instruction; // @[top.scala 168:22]
  wire [31:0] imem22_io_bus_request_bits_address; // @[top.scala 168:22]
  wire [31:0] imem22_io_bus_response_bits_data; // @[top.scala 168:22]
  wire  dmem22_clock; // @[top.scala 169:22]
  wire  dmem22_reset; // @[top.scala 169:22]
  wire [31:0] dmem22_io_pipeline_address; // @[top.scala 169:22]
  wire  dmem22_io_pipeline_valid; // @[top.scala 169:22]
  wire [31:0] dmem22_io_pipeline_writedata; // @[top.scala 169:22]
  wire  dmem22_io_pipeline_memread; // @[top.scala 169:22]
  wire  dmem22_io_pipeline_memwrite; // @[top.scala 169:22]
  wire [1:0] dmem22_io_pipeline_maskmode; // @[top.scala 169:22]
  wire  dmem22_io_pipeline_sext; // @[top.scala 169:22]
  wire [31:0] dmem22_io_pipeline_readdata; // @[top.scala 169:22]
  wire  dmem22_io_bus_request_valid; // @[top.scala 169:22]
  wire [31:0] dmem22_io_bus_request_bits_address; // @[top.scala 169:22]
  wire [31:0] dmem22_io_bus_request_bits_writedata; // @[top.scala 169:22]
  wire [1:0] dmem22_io_bus_request_bits_operation; // @[top.scala 169:22]
  wire  dmem22_io_bus_response_valid; // @[top.scala 169:22]
  wire [31:0] dmem22_io_bus_response_bits_data; // @[top.scala 169:22]
  wire  cpu23_clock; // @[top.scala 173:21]
  wire  cpu23_reset; // @[top.scala 173:21]
  wire [31:0] cpu23_io_imem_address; // @[top.scala 173:21]
  wire [31:0] cpu23_io_imem_instruction; // @[top.scala 173:21]
  wire [31:0] cpu23_io_dmem_address; // @[top.scala 173:21]
  wire  cpu23_io_dmem_valid; // @[top.scala 173:21]
  wire [31:0] cpu23_io_dmem_writedata; // @[top.scala 173:21]
  wire  cpu23_io_dmem_memread; // @[top.scala 173:21]
  wire  cpu23_io_dmem_memwrite; // @[top.scala 173:21]
  wire [1:0] cpu23_io_dmem_maskmode; // @[top.scala 173:21]
  wire  cpu23_io_dmem_sext; // @[top.scala 173:21]
  wire [31:0] cpu23_io_dmem_readdata; // @[top.scala 173:21]
  wire  mem23_clock; // @[top.scala 174:21]
  wire  mem23_reset; // @[top.scala 174:21]
  wire [31:0] mem23_io_imem_request_bits_address; // @[top.scala 174:21]
  wire [31:0] mem23_io_imem_response_bits_data; // @[top.scala 174:21]
  wire  mem23_io_dmem_request_valid; // @[top.scala 174:21]
  wire [31:0] mem23_io_dmem_request_bits_address; // @[top.scala 174:21]
  wire [31:0] mem23_io_dmem_request_bits_writedata; // @[top.scala 174:21]
  wire [1:0] mem23_io_dmem_request_bits_operation; // @[top.scala 174:21]
  wire  mem23_io_dmem_response_valid; // @[top.scala 174:21]
  wire [31:0] mem23_io_dmem_response_bits_data; // @[top.scala 174:21]
  wire [31:0] imem23_io_pipeline_address; // @[top.scala 175:22]
  wire [31:0] imem23_io_pipeline_instruction; // @[top.scala 175:22]
  wire [31:0] imem23_io_bus_request_bits_address; // @[top.scala 175:22]
  wire [31:0] imem23_io_bus_response_bits_data; // @[top.scala 175:22]
  wire  dmem23_clock; // @[top.scala 176:22]
  wire  dmem23_reset; // @[top.scala 176:22]
  wire [31:0] dmem23_io_pipeline_address; // @[top.scala 176:22]
  wire  dmem23_io_pipeline_valid; // @[top.scala 176:22]
  wire [31:0] dmem23_io_pipeline_writedata; // @[top.scala 176:22]
  wire  dmem23_io_pipeline_memread; // @[top.scala 176:22]
  wire  dmem23_io_pipeline_memwrite; // @[top.scala 176:22]
  wire [1:0] dmem23_io_pipeline_maskmode; // @[top.scala 176:22]
  wire  dmem23_io_pipeline_sext; // @[top.scala 176:22]
  wire [31:0] dmem23_io_pipeline_readdata; // @[top.scala 176:22]
  wire  dmem23_io_bus_request_valid; // @[top.scala 176:22]
  wire [31:0] dmem23_io_bus_request_bits_address; // @[top.scala 176:22]
  wire [31:0] dmem23_io_bus_request_bits_writedata; // @[top.scala 176:22]
  wire [1:0] dmem23_io_bus_request_bits_operation; // @[top.scala 176:22]
  wire  dmem23_io_bus_response_valid; // @[top.scala 176:22]
  wire [31:0] dmem23_io_bus_response_bits_data; // @[top.scala 176:22]
  wire  cpu24_clock; // @[top.scala 180:21]
  wire  cpu24_reset; // @[top.scala 180:21]
  wire [31:0] cpu24_io_imem_address; // @[top.scala 180:21]
  wire [31:0] cpu24_io_imem_instruction; // @[top.scala 180:21]
  wire [31:0] cpu24_io_dmem_address; // @[top.scala 180:21]
  wire  cpu24_io_dmem_valid; // @[top.scala 180:21]
  wire [31:0] cpu24_io_dmem_writedata; // @[top.scala 180:21]
  wire  cpu24_io_dmem_memread; // @[top.scala 180:21]
  wire  cpu24_io_dmem_memwrite; // @[top.scala 180:21]
  wire [1:0] cpu24_io_dmem_maskmode; // @[top.scala 180:21]
  wire  cpu24_io_dmem_sext; // @[top.scala 180:21]
  wire [31:0] cpu24_io_dmem_readdata; // @[top.scala 180:21]
  wire  mem24_clock; // @[top.scala 181:21]
  wire  mem24_reset; // @[top.scala 181:21]
  wire [31:0] mem24_io_imem_request_bits_address; // @[top.scala 181:21]
  wire [31:0] mem24_io_imem_response_bits_data; // @[top.scala 181:21]
  wire  mem24_io_dmem_request_valid; // @[top.scala 181:21]
  wire [31:0] mem24_io_dmem_request_bits_address; // @[top.scala 181:21]
  wire [31:0] mem24_io_dmem_request_bits_writedata; // @[top.scala 181:21]
  wire [1:0] mem24_io_dmem_request_bits_operation; // @[top.scala 181:21]
  wire  mem24_io_dmem_response_valid; // @[top.scala 181:21]
  wire [31:0] mem24_io_dmem_response_bits_data; // @[top.scala 181:21]
  wire [31:0] imem24_io_pipeline_address; // @[top.scala 182:22]
  wire [31:0] imem24_io_pipeline_instruction; // @[top.scala 182:22]
  wire [31:0] imem24_io_bus_request_bits_address; // @[top.scala 182:22]
  wire [31:0] imem24_io_bus_response_bits_data; // @[top.scala 182:22]
  wire  dmem24_clock; // @[top.scala 183:22]
  wire  dmem24_reset; // @[top.scala 183:22]
  wire [31:0] dmem24_io_pipeline_address; // @[top.scala 183:22]
  wire  dmem24_io_pipeline_valid; // @[top.scala 183:22]
  wire [31:0] dmem24_io_pipeline_writedata; // @[top.scala 183:22]
  wire  dmem24_io_pipeline_memread; // @[top.scala 183:22]
  wire  dmem24_io_pipeline_memwrite; // @[top.scala 183:22]
  wire [1:0] dmem24_io_pipeline_maskmode; // @[top.scala 183:22]
  wire  dmem24_io_pipeline_sext; // @[top.scala 183:22]
  wire [31:0] dmem24_io_pipeline_readdata; // @[top.scala 183:22]
  wire  dmem24_io_bus_request_valid; // @[top.scala 183:22]
  wire [31:0] dmem24_io_bus_request_bits_address; // @[top.scala 183:22]
  wire [31:0] dmem24_io_bus_request_bits_writedata; // @[top.scala 183:22]
  wire [1:0] dmem24_io_bus_request_bits_operation; // @[top.scala 183:22]
  wire  dmem24_io_bus_response_valid; // @[top.scala 183:22]
  wire [31:0] dmem24_io_bus_response_bits_data; // @[top.scala 183:22]
  wire  cpu25_clock; // @[top.scala 187:21]
  wire  cpu25_reset; // @[top.scala 187:21]
  wire [31:0] cpu25_io_imem_address; // @[top.scala 187:21]
  wire [31:0] cpu25_io_imem_instruction; // @[top.scala 187:21]
  wire [31:0] cpu25_io_dmem_address; // @[top.scala 187:21]
  wire  cpu25_io_dmem_valid; // @[top.scala 187:21]
  wire [31:0] cpu25_io_dmem_writedata; // @[top.scala 187:21]
  wire  cpu25_io_dmem_memread; // @[top.scala 187:21]
  wire  cpu25_io_dmem_memwrite; // @[top.scala 187:21]
  wire [1:0] cpu25_io_dmem_maskmode; // @[top.scala 187:21]
  wire  cpu25_io_dmem_sext; // @[top.scala 187:21]
  wire [31:0] cpu25_io_dmem_readdata; // @[top.scala 187:21]
  wire  mem25_clock; // @[top.scala 188:21]
  wire  mem25_reset; // @[top.scala 188:21]
  wire [31:0] mem25_io_imem_request_bits_address; // @[top.scala 188:21]
  wire [31:0] mem25_io_imem_response_bits_data; // @[top.scala 188:21]
  wire  mem25_io_dmem_request_valid; // @[top.scala 188:21]
  wire [31:0] mem25_io_dmem_request_bits_address; // @[top.scala 188:21]
  wire [31:0] mem25_io_dmem_request_bits_writedata; // @[top.scala 188:21]
  wire [1:0] mem25_io_dmem_request_bits_operation; // @[top.scala 188:21]
  wire  mem25_io_dmem_response_valid; // @[top.scala 188:21]
  wire [31:0] mem25_io_dmem_response_bits_data; // @[top.scala 188:21]
  wire [31:0] imem25_io_pipeline_address; // @[top.scala 189:22]
  wire [31:0] imem25_io_pipeline_instruction; // @[top.scala 189:22]
  wire [31:0] imem25_io_bus_request_bits_address; // @[top.scala 189:22]
  wire [31:0] imem25_io_bus_response_bits_data; // @[top.scala 189:22]
  wire  dmem25_clock; // @[top.scala 190:22]
  wire  dmem25_reset; // @[top.scala 190:22]
  wire [31:0] dmem25_io_pipeline_address; // @[top.scala 190:22]
  wire  dmem25_io_pipeline_valid; // @[top.scala 190:22]
  wire [31:0] dmem25_io_pipeline_writedata; // @[top.scala 190:22]
  wire  dmem25_io_pipeline_memread; // @[top.scala 190:22]
  wire  dmem25_io_pipeline_memwrite; // @[top.scala 190:22]
  wire [1:0] dmem25_io_pipeline_maskmode; // @[top.scala 190:22]
  wire  dmem25_io_pipeline_sext; // @[top.scala 190:22]
  wire [31:0] dmem25_io_pipeline_readdata; // @[top.scala 190:22]
  wire  dmem25_io_bus_request_valid; // @[top.scala 190:22]
  wire [31:0] dmem25_io_bus_request_bits_address; // @[top.scala 190:22]
  wire [31:0] dmem25_io_bus_request_bits_writedata; // @[top.scala 190:22]
  wire [1:0] dmem25_io_bus_request_bits_operation; // @[top.scala 190:22]
  wire  dmem25_io_bus_response_valid; // @[top.scala 190:22]
  wire [31:0] dmem25_io_bus_response_bits_data; // @[top.scala 190:22]
  wire  cpu26_clock; // @[top.scala 194:21]
  wire  cpu26_reset; // @[top.scala 194:21]
  wire [31:0] cpu26_io_imem_address; // @[top.scala 194:21]
  wire [31:0] cpu26_io_imem_instruction; // @[top.scala 194:21]
  wire [31:0] cpu26_io_dmem_address; // @[top.scala 194:21]
  wire  cpu26_io_dmem_valid; // @[top.scala 194:21]
  wire [31:0] cpu26_io_dmem_writedata; // @[top.scala 194:21]
  wire  cpu26_io_dmem_memread; // @[top.scala 194:21]
  wire  cpu26_io_dmem_memwrite; // @[top.scala 194:21]
  wire [1:0] cpu26_io_dmem_maskmode; // @[top.scala 194:21]
  wire  cpu26_io_dmem_sext; // @[top.scala 194:21]
  wire [31:0] cpu26_io_dmem_readdata; // @[top.scala 194:21]
  wire  mem26_clock; // @[top.scala 195:21]
  wire  mem26_reset; // @[top.scala 195:21]
  wire [31:0] mem26_io_imem_request_bits_address; // @[top.scala 195:21]
  wire [31:0] mem26_io_imem_response_bits_data; // @[top.scala 195:21]
  wire  mem26_io_dmem_request_valid; // @[top.scala 195:21]
  wire [31:0] mem26_io_dmem_request_bits_address; // @[top.scala 195:21]
  wire [31:0] mem26_io_dmem_request_bits_writedata; // @[top.scala 195:21]
  wire [1:0] mem26_io_dmem_request_bits_operation; // @[top.scala 195:21]
  wire  mem26_io_dmem_response_valid; // @[top.scala 195:21]
  wire [31:0] mem26_io_dmem_response_bits_data; // @[top.scala 195:21]
  wire [31:0] imem26_io_pipeline_address; // @[top.scala 196:22]
  wire [31:0] imem26_io_pipeline_instruction; // @[top.scala 196:22]
  wire [31:0] imem26_io_bus_request_bits_address; // @[top.scala 196:22]
  wire [31:0] imem26_io_bus_response_bits_data; // @[top.scala 196:22]
  wire  dmem26_clock; // @[top.scala 197:22]
  wire  dmem26_reset; // @[top.scala 197:22]
  wire [31:0] dmem26_io_pipeline_address; // @[top.scala 197:22]
  wire  dmem26_io_pipeline_valid; // @[top.scala 197:22]
  wire [31:0] dmem26_io_pipeline_writedata; // @[top.scala 197:22]
  wire  dmem26_io_pipeline_memread; // @[top.scala 197:22]
  wire  dmem26_io_pipeline_memwrite; // @[top.scala 197:22]
  wire [1:0] dmem26_io_pipeline_maskmode; // @[top.scala 197:22]
  wire  dmem26_io_pipeline_sext; // @[top.scala 197:22]
  wire [31:0] dmem26_io_pipeline_readdata; // @[top.scala 197:22]
  wire  dmem26_io_bus_request_valid; // @[top.scala 197:22]
  wire [31:0] dmem26_io_bus_request_bits_address; // @[top.scala 197:22]
  wire [31:0] dmem26_io_bus_request_bits_writedata; // @[top.scala 197:22]
  wire [1:0] dmem26_io_bus_request_bits_operation; // @[top.scala 197:22]
  wire  dmem26_io_bus_response_valid; // @[top.scala 197:22]
  wire [31:0] dmem26_io_bus_response_bits_data; // @[top.scala 197:22]
  wire  cpu27_clock; // @[top.scala 201:21]
  wire  cpu27_reset; // @[top.scala 201:21]
  wire [31:0] cpu27_io_imem_address; // @[top.scala 201:21]
  wire [31:0] cpu27_io_imem_instruction; // @[top.scala 201:21]
  wire [31:0] cpu27_io_dmem_address; // @[top.scala 201:21]
  wire  cpu27_io_dmem_valid; // @[top.scala 201:21]
  wire [31:0] cpu27_io_dmem_writedata; // @[top.scala 201:21]
  wire  cpu27_io_dmem_memread; // @[top.scala 201:21]
  wire  cpu27_io_dmem_memwrite; // @[top.scala 201:21]
  wire [1:0] cpu27_io_dmem_maskmode; // @[top.scala 201:21]
  wire  cpu27_io_dmem_sext; // @[top.scala 201:21]
  wire [31:0] cpu27_io_dmem_readdata; // @[top.scala 201:21]
  wire  mem27_clock; // @[top.scala 202:21]
  wire  mem27_reset; // @[top.scala 202:21]
  wire [31:0] mem27_io_imem_request_bits_address; // @[top.scala 202:21]
  wire [31:0] mem27_io_imem_response_bits_data; // @[top.scala 202:21]
  wire  mem27_io_dmem_request_valid; // @[top.scala 202:21]
  wire [31:0] mem27_io_dmem_request_bits_address; // @[top.scala 202:21]
  wire [31:0] mem27_io_dmem_request_bits_writedata; // @[top.scala 202:21]
  wire [1:0] mem27_io_dmem_request_bits_operation; // @[top.scala 202:21]
  wire  mem27_io_dmem_response_valid; // @[top.scala 202:21]
  wire [31:0] mem27_io_dmem_response_bits_data; // @[top.scala 202:21]
  wire [31:0] imem27_io_pipeline_address; // @[top.scala 203:22]
  wire [31:0] imem27_io_pipeline_instruction; // @[top.scala 203:22]
  wire [31:0] imem27_io_bus_request_bits_address; // @[top.scala 203:22]
  wire [31:0] imem27_io_bus_response_bits_data; // @[top.scala 203:22]
  wire  dmem27_clock; // @[top.scala 204:22]
  wire  dmem27_reset; // @[top.scala 204:22]
  wire [31:0] dmem27_io_pipeline_address; // @[top.scala 204:22]
  wire  dmem27_io_pipeline_valid; // @[top.scala 204:22]
  wire [31:0] dmem27_io_pipeline_writedata; // @[top.scala 204:22]
  wire  dmem27_io_pipeline_memread; // @[top.scala 204:22]
  wire  dmem27_io_pipeline_memwrite; // @[top.scala 204:22]
  wire [1:0] dmem27_io_pipeline_maskmode; // @[top.scala 204:22]
  wire  dmem27_io_pipeline_sext; // @[top.scala 204:22]
  wire [31:0] dmem27_io_pipeline_readdata; // @[top.scala 204:22]
  wire  dmem27_io_bus_request_valid; // @[top.scala 204:22]
  wire [31:0] dmem27_io_bus_request_bits_address; // @[top.scala 204:22]
  wire [31:0] dmem27_io_bus_request_bits_writedata; // @[top.scala 204:22]
  wire [1:0] dmem27_io_bus_request_bits_operation; // @[top.scala 204:22]
  wire  dmem27_io_bus_response_valid; // @[top.scala 204:22]
  wire [31:0] dmem27_io_bus_response_bits_data; // @[top.scala 204:22]
  wire  cpu28_clock; // @[top.scala 208:21]
  wire  cpu28_reset; // @[top.scala 208:21]
  wire [31:0] cpu28_io_imem_address; // @[top.scala 208:21]
  wire [31:0] cpu28_io_imem_instruction; // @[top.scala 208:21]
  wire [31:0] cpu28_io_dmem_address; // @[top.scala 208:21]
  wire  cpu28_io_dmem_valid; // @[top.scala 208:21]
  wire [31:0] cpu28_io_dmem_writedata; // @[top.scala 208:21]
  wire  cpu28_io_dmem_memread; // @[top.scala 208:21]
  wire  cpu28_io_dmem_memwrite; // @[top.scala 208:21]
  wire [1:0] cpu28_io_dmem_maskmode; // @[top.scala 208:21]
  wire  cpu28_io_dmem_sext; // @[top.scala 208:21]
  wire [31:0] cpu28_io_dmem_readdata; // @[top.scala 208:21]
  wire  mem28_clock; // @[top.scala 209:21]
  wire  mem28_reset; // @[top.scala 209:21]
  wire [31:0] mem28_io_imem_request_bits_address; // @[top.scala 209:21]
  wire [31:0] mem28_io_imem_response_bits_data; // @[top.scala 209:21]
  wire  mem28_io_dmem_request_valid; // @[top.scala 209:21]
  wire [31:0] mem28_io_dmem_request_bits_address; // @[top.scala 209:21]
  wire [31:0] mem28_io_dmem_request_bits_writedata; // @[top.scala 209:21]
  wire [1:0] mem28_io_dmem_request_bits_operation; // @[top.scala 209:21]
  wire  mem28_io_dmem_response_valid; // @[top.scala 209:21]
  wire [31:0] mem28_io_dmem_response_bits_data; // @[top.scala 209:21]
  wire [31:0] imem28_io_pipeline_address; // @[top.scala 210:22]
  wire [31:0] imem28_io_pipeline_instruction; // @[top.scala 210:22]
  wire [31:0] imem28_io_bus_request_bits_address; // @[top.scala 210:22]
  wire [31:0] imem28_io_bus_response_bits_data; // @[top.scala 210:22]
  wire  dmem28_clock; // @[top.scala 211:22]
  wire  dmem28_reset; // @[top.scala 211:22]
  wire [31:0] dmem28_io_pipeline_address; // @[top.scala 211:22]
  wire  dmem28_io_pipeline_valid; // @[top.scala 211:22]
  wire [31:0] dmem28_io_pipeline_writedata; // @[top.scala 211:22]
  wire  dmem28_io_pipeline_memread; // @[top.scala 211:22]
  wire  dmem28_io_pipeline_memwrite; // @[top.scala 211:22]
  wire [1:0] dmem28_io_pipeline_maskmode; // @[top.scala 211:22]
  wire  dmem28_io_pipeline_sext; // @[top.scala 211:22]
  wire [31:0] dmem28_io_pipeline_readdata; // @[top.scala 211:22]
  wire  dmem28_io_bus_request_valid; // @[top.scala 211:22]
  wire [31:0] dmem28_io_bus_request_bits_address; // @[top.scala 211:22]
  wire [31:0] dmem28_io_bus_request_bits_writedata; // @[top.scala 211:22]
  wire [1:0] dmem28_io_bus_request_bits_operation; // @[top.scala 211:22]
  wire  dmem28_io_bus_response_valid; // @[top.scala 211:22]
  wire [31:0] dmem28_io_bus_response_bits_data; // @[top.scala 211:22]
  wire  cpu29_clock; // @[top.scala 215:21]
  wire  cpu29_reset; // @[top.scala 215:21]
  wire [31:0] cpu29_io_imem_address; // @[top.scala 215:21]
  wire [31:0] cpu29_io_imem_instruction; // @[top.scala 215:21]
  wire [31:0] cpu29_io_dmem_address; // @[top.scala 215:21]
  wire  cpu29_io_dmem_valid; // @[top.scala 215:21]
  wire [31:0] cpu29_io_dmem_writedata; // @[top.scala 215:21]
  wire  cpu29_io_dmem_memread; // @[top.scala 215:21]
  wire  cpu29_io_dmem_memwrite; // @[top.scala 215:21]
  wire [1:0] cpu29_io_dmem_maskmode; // @[top.scala 215:21]
  wire  cpu29_io_dmem_sext; // @[top.scala 215:21]
  wire [31:0] cpu29_io_dmem_readdata; // @[top.scala 215:21]
  wire  mem29_clock; // @[top.scala 216:21]
  wire  mem29_reset; // @[top.scala 216:21]
  wire [31:0] mem29_io_imem_request_bits_address; // @[top.scala 216:21]
  wire [31:0] mem29_io_imem_response_bits_data; // @[top.scala 216:21]
  wire  mem29_io_dmem_request_valid; // @[top.scala 216:21]
  wire [31:0] mem29_io_dmem_request_bits_address; // @[top.scala 216:21]
  wire [31:0] mem29_io_dmem_request_bits_writedata; // @[top.scala 216:21]
  wire [1:0] mem29_io_dmem_request_bits_operation; // @[top.scala 216:21]
  wire  mem29_io_dmem_response_valid; // @[top.scala 216:21]
  wire [31:0] mem29_io_dmem_response_bits_data; // @[top.scala 216:21]
  wire [31:0] imem29_io_pipeline_address; // @[top.scala 217:22]
  wire [31:0] imem29_io_pipeline_instruction; // @[top.scala 217:22]
  wire [31:0] imem29_io_bus_request_bits_address; // @[top.scala 217:22]
  wire [31:0] imem29_io_bus_response_bits_data; // @[top.scala 217:22]
  wire  dmem29_clock; // @[top.scala 218:22]
  wire  dmem29_reset; // @[top.scala 218:22]
  wire [31:0] dmem29_io_pipeline_address; // @[top.scala 218:22]
  wire  dmem29_io_pipeline_valid; // @[top.scala 218:22]
  wire [31:0] dmem29_io_pipeline_writedata; // @[top.scala 218:22]
  wire  dmem29_io_pipeline_memread; // @[top.scala 218:22]
  wire  dmem29_io_pipeline_memwrite; // @[top.scala 218:22]
  wire [1:0] dmem29_io_pipeline_maskmode; // @[top.scala 218:22]
  wire  dmem29_io_pipeline_sext; // @[top.scala 218:22]
  wire [31:0] dmem29_io_pipeline_readdata; // @[top.scala 218:22]
  wire  dmem29_io_bus_request_valid; // @[top.scala 218:22]
  wire [31:0] dmem29_io_bus_request_bits_address; // @[top.scala 218:22]
  wire [31:0] dmem29_io_bus_request_bits_writedata; // @[top.scala 218:22]
  wire [1:0] dmem29_io_bus_request_bits_operation; // @[top.scala 218:22]
  wire  dmem29_io_bus_response_valid; // @[top.scala 218:22]
  wire [31:0] dmem29_io_bus_response_bits_data; // @[top.scala 218:22]
  wire  cpu30_clock; // @[top.scala 222:21]
  wire  cpu30_reset; // @[top.scala 222:21]
  wire [31:0] cpu30_io_imem_address; // @[top.scala 222:21]
  wire [31:0] cpu30_io_imem_instruction; // @[top.scala 222:21]
  wire [31:0] cpu30_io_dmem_address; // @[top.scala 222:21]
  wire  cpu30_io_dmem_valid; // @[top.scala 222:21]
  wire [31:0] cpu30_io_dmem_writedata; // @[top.scala 222:21]
  wire  cpu30_io_dmem_memread; // @[top.scala 222:21]
  wire  cpu30_io_dmem_memwrite; // @[top.scala 222:21]
  wire [1:0] cpu30_io_dmem_maskmode; // @[top.scala 222:21]
  wire  cpu30_io_dmem_sext; // @[top.scala 222:21]
  wire [31:0] cpu30_io_dmem_readdata; // @[top.scala 222:21]
  wire  mem30_clock; // @[top.scala 223:21]
  wire  mem30_reset; // @[top.scala 223:21]
  wire [31:0] mem30_io_imem_request_bits_address; // @[top.scala 223:21]
  wire [31:0] mem30_io_imem_response_bits_data; // @[top.scala 223:21]
  wire  mem30_io_dmem_request_valid; // @[top.scala 223:21]
  wire [31:0] mem30_io_dmem_request_bits_address; // @[top.scala 223:21]
  wire [31:0] mem30_io_dmem_request_bits_writedata; // @[top.scala 223:21]
  wire [1:0] mem30_io_dmem_request_bits_operation; // @[top.scala 223:21]
  wire  mem30_io_dmem_response_valid; // @[top.scala 223:21]
  wire [31:0] mem30_io_dmem_response_bits_data; // @[top.scala 223:21]
  wire [31:0] imem30_io_pipeline_address; // @[top.scala 224:22]
  wire [31:0] imem30_io_pipeline_instruction; // @[top.scala 224:22]
  wire [31:0] imem30_io_bus_request_bits_address; // @[top.scala 224:22]
  wire [31:0] imem30_io_bus_response_bits_data; // @[top.scala 224:22]
  wire  dmem30_clock; // @[top.scala 225:22]
  wire  dmem30_reset; // @[top.scala 225:22]
  wire [31:0] dmem30_io_pipeline_address; // @[top.scala 225:22]
  wire  dmem30_io_pipeline_valid; // @[top.scala 225:22]
  wire [31:0] dmem30_io_pipeline_writedata; // @[top.scala 225:22]
  wire  dmem30_io_pipeline_memread; // @[top.scala 225:22]
  wire  dmem30_io_pipeline_memwrite; // @[top.scala 225:22]
  wire [1:0] dmem30_io_pipeline_maskmode; // @[top.scala 225:22]
  wire  dmem30_io_pipeline_sext; // @[top.scala 225:22]
  wire [31:0] dmem30_io_pipeline_readdata; // @[top.scala 225:22]
  wire  dmem30_io_bus_request_valid; // @[top.scala 225:22]
  wire [31:0] dmem30_io_bus_request_bits_address; // @[top.scala 225:22]
  wire [31:0] dmem30_io_bus_request_bits_writedata; // @[top.scala 225:22]
  wire [1:0] dmem30_io_bus_request_bits_operation; // @[top.scala 225:22]
  wire  dmem30_io_bus_response_valid; // @[top.scala 225:22]
  wire [31:0] dmem30_io_bus_response_bits_data; // @[top.scala 225:22]
  wire  cpu31_clock; // @[top.scala 229:21]
  wire  cpu31_reset; // @[top.scala 229:21]
  wire [31:0] cpu31_io_imem_address; // @[top.scala 229:21]
  wire [31:0] cpu31_io_imem_instruction; // @[top.scala 229:21]
  wire [31:0] cpu31_io_dmem_address; // @[top.scala 229:21]
  wire  cpu31_io_dmem_valid; // @[top.scala 229:21]
  wire [31:0] cpu31_io_dmem_writedata; // @[top.scala 229:21]
  wire  cpu31_io_dmem_memread; // @[top.scala 229:21]
  wire  cpu31_io_dmem_memwrite; // @[top.scala 229:21]
  wire [1:0] cpu31_io_dmem_maskmode; // @[top.scala 229:21]
  wire  cpu31_io_dmem_sext; // @[top.scala 229:21]
  wire [31:0] cpu31_io_dmem_readdata; // @[top.scala 229:21]
  wire  mem31_clock; // @[top.scala 230:21]
  wire  mem31_reset; // @[top.scala 230:21]
  wire [31:0] mem31_io_imem_request_bits_address; // @[top.scala 230:21]
  wire [31:0] mem31_io_imem_response_bits_data; // @[top.scala 230:21]
  wire  mem31_io_dmem_request_valid; // @[top.scala 230:21]
  wire [31:0] mem31_io_dmem_request_bits_address; // @[top.scala 230:21]
  wire [31:0] mem31_io_dmem_request_bits_writedata; // @[top.scala 230:21]
  wire [1:0] mem31_io_dmem_request_bits_operation; // @[top.scala 230:21]
  wire  mem31_io_dmem_response_valid; // @[top.scala 230:21]
  wire [31:0] mem31_io_dmem_response_bits_data; // @[top.scala 230:21]
  wire [31:0] imem31_io_pipeline_address; // @[top.scala 231:22]
  wire [31:0] imem31_io_pipeline_instruction; // @[top.scala 231:22]
  wire [31:0] imem31_io_bus_request_bits_address; // @[top.scala 231:22]
  wire [31:0] imem31_io_bus_response_bits_data; // @[top.scala 231:22]
  wire  dmem31_clock; // @[top.scala 232:22]
  wire  dmem31_reset; // @[top.scala 232:22]
  wire [31:0] dmem31_io_pipeline_address; // @[top.scala 232:22]
  wire  dmem31_io_pipeline_valid; // @[top.scala 232:22]
  wire [31:0] dmem31_io_pipeline_writedata; // @[top.scala 232:22]
  wire  dmem31_io_pipeline_memread; // @[top.scala 232:22]
  wire  dmem31_io_pipeline_memwrite; // @[top.scala 232:22]
  wire [1:0] dmem31_io_pipeline_maskmode; // @[top.scala 232:22]
  wire  dmem31_io_pipeline_sext; // @[top.scala 232:22]
  wire [31:0] dmem31_io_pipeline_readdata; // @[top.scala 232:22]
  wire  dmem31_io_bus_request_valid; // @[top.scala 232:22]
  wire [31:0] dmem31_io_bus_request_bits_address; // @[top.scala 232:22]
  wire [31:0] dmem31_io_bus_request_bits_writedata; // @[top.scala 232:22]
  wire [1:0] dmem31_io_bus_request_bits_operation; // @[top.scala 232:22]
  wire  dmem31_io_bus_response_valid; // @[top.scala 232:22]
  wire [31:0] dmem31_io_bus_response_bits_data; // @[top.scala 232:22]
  wire  cpu32_clock; // @[top.scala 236:21]
  wire  cpu32_reset; // @[top.scala 236:21]
  wire [31:0] cpu32_io_imem_address; // @[top.scala 236:21]
  wire [31:0] cpu32_io_imem_instruction; // @[top.scala 236:21]
  wire [31:0] cpu32_io_dmem_address; // @[top.scala 236:21]
  wire  cpu32_io_dmem_valid; // @[top.scala 236:21]
  wire [31:0] cpu32_io_dmem_writedata; // @[top.scala 236:21]
  wire  cpu32_io_dmem_memread; // @[top.scala 236:21]
  wire  cpu32_io_dmem_memwrite; // @[top.scala 236:21]
  wire [1:0] cpu32_io_dmem_maskmode; // @[top.scala 236:21]
  wire  cpu32_io_dmem_sext; // @[top.scala 236:21]
  wire [31:0] cpu32_io_dmem_readdata; // @[top.scala 236:21]
  wire  mem32_clock; // @[top.scala 237:21]
  wire  mem32_reset; // @[top.scala 237:21]
  wire [31:0] mem32_io_imem_request_bits_address; // @[top.scala 237:21]
  wire [31:0] mem32_io_imem_response_bits_data; // @[top.scala 237:21]
  wire  mem32_io_dmem_request_valid; // @[top.scala 237:21]
  wire [31:0] mem32_io_dmem_request_bits_address; // @[top.scala 237:21]
  wire [31:0] mem32_io_dmem_request_bits_writedata; // @[top.scala 237:21]
  wire [1:0] mem32_io_dmem_request_bits_operation; // @[top.scala 237:21]
  wire  mem32_io_dmem_response_valid; // @[top.scala 237:21]
  wire [31:0] mem32_io_dmem_response_bits_data; // @[top.scala 237:21]
  wire [31:0] imem32_io_pipeline_address; // @[top.scala 238:22]
  wire [31:0] imem32_io_pipeline_instruction; // @[top.scala 238:22]
  wire [31:0] imem32_io_bus_request_bits_address; // @[top.scala 238:22]
  wire [31:0] imem32_io_bus_response_bits_data; // @[top.scala 238:22]
  wire  dmem32_clock; // @[top.scala 239:22]
  wire  dmem32_reset; // @[top.scala 239:22]
  wire [31:0] dmem32_io_pipeline_address; // @[top.scala 239:22]
  wire  dmem32_io_pipeline_valid; // @[top.scala 239:22]
  wire [31:0] dmem32_io_pipeline_writedata; // @[top.scala 239:22]
  wire  dmem32_io_pipeline_memread; // @[top.scala 239:22]
  wire  dmem32_io_pipeline_memwrite; // @[top.scala 239:22]
  wire [1:0] dmem32_io_pipeline_maskmode; // @[top.scala 239:22]
  wire  dmem32_io_pipeline_sext; // @[top.scala 239:22]
  wire [31:0] dmem32_io_pipeline_readdata; // @[top.scala 239:22]
  wire  dmem32_io_bus_request_valid; // @[top.scala 239:22]
  wire [31:0] dmem32_io_bus_request_bits_address; // @[top.scala 239:22]
  wire [31:0] dmem32_io_bus_request_bits_writedata; // @[top.scala 239:22]
  wire [1:0] dmem32_io_bus_request_bits_operation; // @[top.scala 239:22]
  wire  dmem32_io_bus_response_valid; // @[top.scala 239:22]
  wire [31:0] dmem32_io_bus_response_bits_data; // @[top.scala 239:22]
  wire  cpu33_clock; // @[top.scala 243:21]
  wire  cpu33_reset; // @[top.scala 243:21]
  wire [31:0] cpu33_io_imem_address; // @[top.scala 243:21]
  wire [31:0] cpu33_io_imem_instruction; // @[top.scala 243:21]
  wire [31:0] cpu33_io_dmem_address; // @[top.scala 243:21]
  wire  cpu33_io_dmem_valid; // @[top.scala 243:21]
  wire [31:0] cpu33_io_dmem_writedata; // @[top.scala 243:21]
  wire  cpu33_io_dmem_memread; // @[top.scala 243:21]
  wire  cpu33_io_dmem_memwrite; // @[top.scala 243:21]
  wire [1:0] cpu33_io_dmem_maskmode; // @[top.scala 243:21]
  wire  cpu33_io_dmem_sext; // @[top.scala 243:21]
  wire [31:0] cpu33_io_dmem_readdata; // @[top.scala 243:21]
  wire  mem33_clock; // @[top.scala 244:21]
  wire  mem33_reset; // @[top.scala 244:21]
  wire [31:0] mem33_io_imem_request_bits_address; // @[top.scala 244:21]
  wire [31:0] mem33_io_imem_response_bits_data; // @[top.scala 244:21]
  wire  mem33_io_dmem_request_valid; // @[top.scala 244:21]
  wire [31:0] mem33_io_dmem_request_bits_address; // @[top.scala 244:21]
  wire [31:0] mem33_io_dmem_request_bits_writedata; // @[top.scala 244:21]
  wire [1:0] mem33_io_dmem_request_bits_operation; // @[top.scala 244:21]
  wire  mem33_io_dmem_response_valid; // @[top.scala 244:21]
  wire [31:0] mem33_io_dmem_response_bits_data; // @[top.scala 244:21]
  wire [31:0] imem33_io_pipeline_address; // @[top.scala 245:22]
  wire [31:0] imem33_io_pipeline_instruction; // @[top.scala 245:22]
  wire [31:0] imem33_io_bus_request_bits_address; // @[top.scala 245:22]
  wire [31:0] imem33_io_bus_response_bits_data; // @[top.scala 245:22]
  wire  dmem33_clock; // @[top.scala 246:22]
  wire  dmem33_reset; // @[top.scala 246:22]
  wire [31:0] dmem33_io_pipeline_address; // @[top.scala 246:22]
  wire  dmem33_io_pipeline_valid; // @[top.scala 246:22]
  wire [31:0] dmem33_io_pipeline_writedata; // @[top.scala 246:22]
  wire  dmem33_io_pipeline_memread; // @[top.scala 246:22]
  wire  dmem33_io_pipeline_memwrite; // @[top.scala 246:22]
  wire [1:0] dmem33_io_pipeline_maskmode; // @[top.scala 246:22]
  wire  dmem33_io_pipeline_sext; // @[top.scala 246:22]
  wire [31:0] dmem33_io_pipeline_readdata; // @[top.scala 246:22]
  wire  dmem33_io_bus_request_valid; // @[top.scala 246:22]
  wire [31:0] dmem33_io_bus_request_bits_address; // @[top.scala 246:22]
  wire [31:0] dmem33_io_bus_request_bits_writedata; // @[top.scala 246:22]
  wire [1:0] dmem33_io_bus_request_bits_operation; // @[top.scala 246:22]
  wire  dmem33_io_bus_response_valid; // @[top.scala 246:22]
  wire [31:0] dmem33_io_bus_response_bits_data; // @[top.scala 246:22]
  wire  cpu34_clock; // @[top.scala 250:21]
  wire  cpu34_reset; // @[top.scala 250:21]
  wire [31:0] cpu34_io_imem_address; // @[top.scala 250:21]
  wire [31:0] cpu34_io_imem_instruction; // @[top.scala 250:21]
  wire [31:0] cpu34_io_dmem_address; // @[top.scala 250:21]
  wire  cpu34_io_dmem_valid; // @[top.scala 250:21]
  wire [31:0] cpu34_io_dmem_writedata; // @[top.scala 250:21]
  wire  cpu34_io_dmem_memread; // @[top.scala 250:21]
  wire  cpu34_io_dmem_memwrite; // @[top.scala 250:21]
  wire [1:0] cpu34_io_dmem_maskmode; // @[top.scala 250:21]
  wire  cpu34_io_dmem_sext; // @[top.scala 250:21]
  wire [31:0] cpu34_io_dmem_readdata; // @[top.scala 250:21]
  wire  mem34_clock; // @[top.scala 251:21]
  wire  mem34_reset; // @[top.scala 251:21]
  wire [31:0] mem34_io_imem_request_bits_address; // @[top.scala 251:21]
  wire [31:0] mem34_io_imem_response_bits_data; // @[top.scala 251:21]
  wire  mem34_io_dmem_request_valid; // @[top.scala 251:21]
  wire [31:0] mem34_io_dmem_request_bits_address; // @[top.scala 251:21]
  wire [31:0] mem34_io_dmem_request_bits_writedata; // @[top.scala 251:21]
  wire [1:0] mem34_io_dmem_request_bits_operation; // @[top.scala 251:21]
  wire  mem34_io_dmem_response_valid; // @[top.scala 251:21]
  wire [31:0] mem34_io_dmem_response_bits_data; // @[top.scala 251:21]
  wire [31:0] imem34_io_pipeline_address; // @[top.scala 252:22]
  wire [31:0] imem34_io_pipeline_instruction; // @[top.scala 252:22]
  wire [31:0] imem34_io_bus_request_bits_address; // @[top.scala 252:22]
  wire [31:0] imem34_io_bus_response_bits_data; // @[top.scala 252:22]
  wire  dmem34_clock; // @[top.scala 253:22]
  wire  dmem34_reset; // @[top.scala 253:22]
  wire [31:0] dmem34_io_pipeline_address; // @[top.scala 253:22]
  wire  dmem34_io_pipeline_valid; // @[top.scala 253:22]
  wire [31:0] dmem34_io_pipeline_writedata; // @[top.scala 253:22]
  wire  dmem34_io_pipeline_memread; // @[top.scala 253:22]
  wire  dmem34_io_pipeline_memwrite; // @[top.scala 253:22]
  wire [1:0] dmem34_io_pipeline_maskmode; // @[top.scala 253:22]
  wire  dmem34_io_pipeline_sext; // @[top.scala 253:22]
  wire [31:0] dmem34_io_pipeline_readdata; // @[top.scala 253:22]
  wire  dmem34_io_bus_request_valid; // @[top.scala 253:22]
  wire [31:0] dmem34_io_bus_request_bits_address; // @[top.scala 253:22]
  wire [31:0] dmem34_io_bus_request_bits_writedata; // @[top.scala 253:22]
  wire [1:0] dmem34_io_bus_request_bits_operation; // @[top.scala 253:22]
  wire  dmem34_io_bus_response_valid; // @[top.scala 253:22]
  wire [31:0] dmem34_io_bus_response_bits_data; // @[top.scala 253:22]
  wire  cpu35_clock; // @[top.scala 257:21]
  wire  cpu35_reset; // @[top.scala 257:21]
  wire [31:0] cpu35_io_imem_address; // @[top.scala 257:21]
  wire [31:0] cpu35_io_imem_instruction; // @[top.scala 257:21]
  wire [31:0] cpu35_io_dmem_address; // @[top.scala 257:21]
  wire  cpu35_io_dmem_valid; // @[top.scala 257:21]
  wire [31:0] cpu35_io_dmem_writedata; // @[top.scala 257:21]
  wire  cpu35_io_dmem_memread; // @[top.scala 257:21]
  wire  cpu35_io_dmem_memwrite; // @[top.scala 257:21]
  wire [1:0] cpu35_io_dmem_maskmode; // @[top.scala 257:21]
  wire  cpu35_io_dmem_sext; // @[top.scala 257:21]
  wire [31:0] cpu35_io_dmem_readdata; // @[top.scala 257:21]
  wire  mem35_clock; // @[top.scala 258:21]
  wire  mem35_reset; // @[top.scala 258:21]
  wire [31:0] mem35_io_imem_request_bits_address; // @[top.scala 258:21]
  wire [31:0] mem35_io_imem_response_bits_data; // @[top.scala 258:21]
  wire  mem35_io_dmem_request_valid; // @[top.scala 258:21]
  wire [31:0] mem35_io_dmem_request_bits_address; // @[top.scala 258:21]
  wire [31:0] mem35_io_dmem_request_bits_writedata; // @[top.scala 258:21]
  wire [1:0] mem35_io_dmem_request_bits_operation; // @[top.scala 258:21]
  wire  mem35_io_dmem_response_valid; // @[top.scala 258:21]
  wire [31:0] mem35_io_dmem_response_bits_data; // @[top.scala 258:21]
  wire [31:0] imem35_io_pipeline_address; // @[top.scala 259:22]
  wire [31:0] imem35_io_pipeline_instruction; // @[top.scala 259:22]
  wire [31:0] imem35_io_bus_request_bits_address; // @[top.scala 259:22]
  wire [31:0] imem35_io_bus_response_bits_data; // @[top.scala 259:22]
  wire  dmem35_clock; // @[top.scala 260:22]
  wire  dmem35_reset; // @[top.scala 260:22]
  wire [31:0] dmem35_io_pipeline_address; // @[top.scala 260:22]
  wire  dmem35_io_pipeline_valid; // @[top.scala 260:22]
  wire [31:0] dmem35_io_pipeline_writedata; // @[top.scala 260:22]
  wire  dmem35_io_pipeline_memread; // @[top.scala 260:22]
  wire  dmem35_io_pipeline_memwrite; // @[top.scala 260:22]
  wire [1:0] dmem35_io_pipeline_maskmode; // @[top.scala 260:22]
  wire  dmem35_io_pipeline_sext; // @[top.scala 260:22]
  wire [31:0] dmem35_io_pipeline_readdata; // @[top.scala 260:22]
  wire  dmem35_io_bus_request_valid; // @[top.scala 260:22]
  wire [31:0] dmem35_io_bus_request_bits_address; // @[top.scala 260:22]
  wire [31:0] dmem35_io_bus_request_bits_writedata; // @[top.scala 260:22]
  wire [1:0] dmem35_io_bus_request_bits_operation; // @[top.scala 260:22]
  wire  dmem35_io_bus_response_valid; // @[top.scala 260:22]
  wire [31:0] dmem35_io_bus_response_bits_data; // @[top.scala 260:22]
  wire  cpu36_clock; // @[top.scala 264:21]
  wire  cpu36_reset; // @[top.scala 264:21]
  wire [31:0] cpu36_io_imem_address; // @[top.scala 264:21]
  wire [31:0] cpu36_io_imem_instruction; // @[top.scala 264:21]
  wire [31:0] cpu36_io_dmem_address; // @[top.scala 264:21]
  wire  cpu36_io_dmem_valid; // @[top.scala 264:21]
  wire [31:0] cpu36_io_dmem_writedata; // @[top.scala 264:21]
  wire  cpu36_io_dmem_memread; // @[top.scala 264:21]
  wire  cpu36_io_dmem_memwrite; // @[top.scala 264:21]
  wire [1:0] cpu36_io_dmem_maskmode; // @[top.scala 264:21]
  wire  cpu36_io_dmem_sext; // @[top.scala 264:21]
  wire [31:0] cpu36_io_dmem_readdata; // @[top.scala 264:21]
  wire  mem36_clock; // @[top.scala 265:21]
  wire  mem36_reset; // @[top.scala 265:21]
  wire [31:0] mem36_io_imem_request_bits_address; // @[top.scala 265:21]
  wire [31:0] mem36_io_imem_response_bits_data; // @[top.scala 265:21]
  wire  mem36_io_dmem_request_valid; // @[top.scala 265:21]
  wire [31:0] mem36_io_dmem_request_bits_address; // @[top.scala 265:21]
  wire [31:0] mem36_io_dmem_request_bits_writedata; // @[top.scala 265:21]
  wire [1:0] mem36_io_dmem_request_bits_operation; // @[top.scala 265:21]
  wire  mem36_io_dmem_response_valid; // @[top.scala 265:21]
  wire [31:0] mem36_io_dmem_response_bits_data; // @[top.scala 265:21]
  wire [31:0] imem36_io_pipeline_address; // @[top.scala 266:22]
  wire [31:0] imem36_io_pipeline_instruction; // @[top.scala 266:22]
  wire [31:0] imem36_io_bus_request_bits_address; // @[top.scala 266:22]
  wire [31:0] imem36_io_bus_response_bits_data; // @[top.scala 266:22]
  wire  dmem36_clock; // @[top.scala 267:22]
  wire  dmem36_reset; // @[top.scala 267:22]
  wire [31:0] dmem36_io_pipeline_address; // @[top.scala 267:22]
  wire  dmem36_io_pipeline_valid; // @[top.scala 267:22]
  wire [31:0] dmem36_io_pipeline_writedata; // @[top.scala 267:22]
  wire  dmem36_io_pipeline_memread; // @[top.scala 267:22]
  wire  dmem36_io_pipeline_memwrite; // @[top.scala 267:22]
  wire [1:0] dmem36_io_pipeline_maskmode; // @[top.scala 267:22]
  wire  dmem36_io_pipeline_sext; // @[top.scala 267:22]
  wire [31:0] dmem36_io_pipeline_readdata; // @[top.scala 267:22]
  wire  dmem36_io_bus_request_valid; // @[top.scala 267:22]
  wire [31:0] dmem36_io_bus_request_bits_address; // @[top.scala 267:22]
  wire [31:0] dmem36_io_bus_request_bits_writedata; // @[top.scala 267:22]
  wire [1:0] dmem36_io_bus_request_bits_operation; // @[top.scala 267:22]
  wire  dmem36_io_bus_response_valid; // @[top.scala 267:22]
  wire [31:0] dmem36_io_bus_response_bits_data; // @[top.scala 267:22]
  wire  cpu37_clock; // @[top.scala 271:21]
  wire  cpu37_reset; // @[top.scala 271:21]
  wire [31:0] cpu37_io_imem_address; // @[top.scala 271:21]
  wire [31:0] cpu37_io_imem_instruction; // @[top.scala 271:21]
  wire [31:0] cpu37_io_dmem_address; // @[top.scala 271:21]
  wire  cpu37_io_dmem_valid; // @[top.scala 271:21]
  wire [31:0] cpu37_io_dmem_writedata; // @[top.scala 271:21]
  wire  cpu37_io_dmem_memread; // @[top.scala 271:21]
  wire  cpu37_io_dmem_memwrite; // @[top.scala 271:21]
  wire [1:0] cpu37_io_dmem_maskmode; // @[top.scala 271:21]
  wire  cpu37_io_dmem_sext; // @[top.scala 271:21]
  wire [31:0] cpu37_io_dmem_readdata; // @[top.scala 271:21]
  wire  mem37_clock; // @[top.scala 272:21]
  wire  mem37_reset; // @[top.scala 272:21]
  wire [31:0] mem37_io_imem_request_bits_address; // @[top.scala 272:21]
  wire [31:0] mem37_io_imem_response_bits_data; // @[top.scala 272:21]
  wire  mem37_io_dmem_request_valid; // @[top.scala 272:21]
  wire [31:0] mem37_io_dmem_request_bits_address; // @[top.scala 272:21]
  wire [31:0] mem37_io_dmem_request_bits_writedata; // @[top.scala 272:21]
  wire [1:0] mem37_io_dmem_request_bits_operation; // @[top.scala 272:21]
  wire  mem37_io_dmem_response_valid; // @[top.scala 272:21]
  wire [31:0] mem37_io_dmem_response_bits_data; // @[top.scala 272:21]
  wire [31:0] imem37_io_pipeline_address; // @[top.scala 273:22]
  wire [31:0] imem37_io_pipeline_instruction; // @[top.scala 273:22]
  wire [31:0] imem37_io_bus_request_bits_address; // @[top.scala 273:22]
  wire [31:0] imem37_io_bus_response_bits_data; // @[top.scala 273:22]
  wire  dmem37_clock; // @[top.scala 274:22]
  wire  dmem37_reset; // @[top.scala 274:22]
  wire [31:0] dmem37_io_pipeline_address; // @[top.scala 274:22]
  wire  dmem37_io_pipeline_valid; // @[top.scala 274:22]
  wire [31:0] dmem37_io_pipeline_writedata; // @[top.scala 274:22]
  wire  dmem37_io_pipeline_memread; // @[top.scala 274:22]
  wire  dmem37_io_pipeline_memwrite; // @[top.scala 274:22]
  wire [1:0] dmem37_io_pipeline_maskmode; // @[top.scala 274:22]
  wire  dmem37_io_pipeline_sext; // @[top.scala 274:22]
  wire [31:0] dmem37_io_pipeline_readdata; // @[top.scala 274:22]
  wire  dmem37_io_bus_request_valid; // @[top.scala 274:22]
  wire [31:0] dmem37_io_bus_request_bits_address; // @[top.scala 274:22]
  wire [31:0] dmem37_io_bus_request_bits_writedata; // @[top.scala 274:22]
  wire [1:0] dmem37_io_bus_request_bits_operation; // @[top.scala 274:22]
  wire  dmem37_io_bus_response_valid; // @[top.scala 274:22]
  wire [31:0] dmem37_io_bus_response_bits_data; // @[top.scala 274:22]
  wire  cpu38_clock; // @[top.scala 278:21]
  wire  cpu38_reset; // @[top.scala 278:21]
  wire [31:0] cpu38_io_imem_address; // @[top.scala 278:21]
  wire [31:0] cpu38_io_imem_instruction; // @[top.scala 278:21]
  wire [31:0] cpu38_io_dmem_address; // @[top.scala 278:21]
  wire  cpu38_io_dmem_valid; // @[top.scala 278:21]
  wire [31:0] cpu38_io_dmem_writedata; // @[top.scala 278:21]
  wire  cpu38_io_dmem_memread; // @[top.scala 278:21]
  wire  cpu38_io_dmem_memwrite; // @[top.scala 278:21]
  wire [1:0] cpu38_io_dmem_maskmode; // @[top.scala 278:21]
  wire  cpu38_io_dmem_sext; // @[top.scala 278:21]
  wire [31:0] cpu38_io_dmem_readdata; // @[top.scala 278:21]
  wire  mem38_clock; // @[top.scala 279:21]
  wire  mem38_reset; // @[top.scala 279:21]
  wire [31:0] mem38_io_imem_request_bits_address; // @[top.scala 279:21]
  wire [31:0] mem38_io_imem_response_bits_data; // @[top.scala 279:21]
  wire  mem38_io_dmem_request_valid; // @[top.scala 279:21]
  wire [31:0] mem38_io_dmem_request_bits_address; // @[top.scala 279:21]
  wire [31:0] mem38_io_dmem_request_bits_writedata; // @[top.scala 279:21]
  wire [1:0] mem38_io_dmem_request_bits_operation; // @[top.scala 279:21]
  wire  mem38_io_dmem_response_valid; // @[top.scala 279:21]
  wire [31:0] mem38_io_dmem_response_bits_data; // @[top.scala 279:21]
  wire [31:0] imem38_io_pipeline_address; // @[top.scala 280:22]
  wire [31:0] imem38_io_pipeline_instruction; // @[top.scala 280:22]
  wire [31:0] imem38_io_bus_request_bits_address; // @[top.scala 280:22]
  wire [31:0] imem38_io_bus_response_bits_data; // @[top.scala 280:22]
  wire  dmem38_clock; // @[top.scala 281:22]
  wire  dmem38_reset; // @[top.scala 281:22]
  wire [31:0] dmem38_io_pipeline_address; // @[top.scala 281:22]
  wire  dmem38_io_pipeline_valid; // @[top.scala 281:22]
  wire [31:0] dmem38_io_pipeline_writedata; // @[top.scala 281:22]
  wire  dmem38_io_pipeline_memread; // @[top.scala 281:22]
  wire  dmem38_io_pipeline_memwrite; // @[top.scala 281:22]
  wire [1:0] dmem38_io_pipeline_maskmode; // @[top.scala 281:22]
  wire  dmem38_io_pipeline_sext; // @[top.scala 281:22]
  wire [31:0] dmem38_io_pipeline_readdata; // @[top.scala 281:22]
  wire  dmem38_io_bus_request_valid; // @[top.scala 281:22]
  wire [31:0] dmem38_io_bus_request_bits_address; // @[top.scala 281:22]
  wire [31:0] dmem38_io_bus_request_bits_writedata; // @[top.scala 281:22]
  wire [1:0] dmem38_io_bus_request_bits_operation; // @[top.scala 281:22]
  wire  dmem38_io_bus_response_valid; // @[top.scala 281:22]
  wire [31:0] dmem38_io_bus_response_bits_data; // @[top.scala 281:22]
  wire  cpu39_clock; // @[top.scala 285:21]
  wire  cpu39_reset; // @[top.scala 285:21]
  wire [31:0] cpu39_io_imem_address; // @[top.scala 285:21]
  wire [31:0] cpu39_io_imem_instruction; // @[top.scala 285:21]
  wire [31:0] cpu39_io_dmem_address; // @[top.scala 285:21]
  wire  cpu39_io_dmem_valid; // @[top.scala 285:21]
  wire [31:0] cpu39_io_dmem_writedata; // @[top.scala 285:21]
  wire  cpu39_io_dmem_memread; // @[top.scala 285:21]
  wire  cpu39_io_dmem_memwrite; // @[top.scala 285:21]
  wire [1:0] cpu39_io_dmem_maskmode; // @[top.scala 285:21]
  wire  cpu39_io_dmem_sext; // @[top.scala 285:21]
  wire [31:0] cpu39_io_dmem_readdata; // @[top.scala 285:21]
  wire  mem39_clock; // @[top.scala 286:21]
  wire  mem39_reset; // @[top.scala 286:21]
  wire [31:0] mem39_io_imem_request_bits_address; // @[top.scala 286:21]
  wire [31:0] mem39_io_imem_response_bits_data; // @[top.scala 286:21]
  wire  mem39_io_dmem_request_valid; // @[top.scala 286:21]
  wire [31:0] mem39_io_dmem_request_bits_address; // @[top.scala 286:21]
  wire [31:0] mem39_io_dmem_request_bits_writedata; // @[top.scala 286:21]
  wire [1:0] mem39_io_dmem_request_bits_operation; // @[top.scala 286:21]
  wire  mem39_io_dmem_response_valid; // @[top.scala 286:21]
  wire [31:0] mem39_io_dmem_response_bits_data; // @[top.scala 286:21]
  wire [31:0] imem39_io_pipeline_address; // @[top.scala 287:22]
  wire [31:0] imem39_io_pipeline_instruction; // @[top.scala 287:22]
  wire [31:0] imem39_io_bus_request_bits_address; // @[top.scala 287:22]
  wire [31:0] imem39_io_bus_response_bits_data; // @[top.scala 287:22]
  wire  dmem39_clock; // @[top.scala 288:22]
  wire  dmem39_reset; // @[top.scala 288:22]
  wire [31:0] dmem39_io_pipeline_address; // @[top.scala 288:22]
  wire  dmem39_io_pipeline_valid; // @[top.scala 288:22]
  wire [31:0] dmem39_io_pipeline_writedata; // @[top.scala 288:22]
  wire  dmem39_io_pipeline_memread; // @[top.scala 288:22]
  wire  dmem39_io_pipeline_memwrite; // @[top.scala 288:22]
  wire [1:0] dmem39_io_pipeline_maskmode; // @[top.scala 288:22]
  wire  dmem39_io_pipeline_sext; // @[top.scala 288:22]
  wire [31:0] dmem39_io_pipeline_readdata; // @[top.scala 288:22]
  wire  dmem39_io_bus_request_valid; // @[top.scala 288:22]
  wire [31:0] dmem39_io_bus_request_bits_address; // @[top.scala 288:22]
  wire [31:0] dmem39_io_bus_request_bits_writedata; // @[top.scala 288:22]
  wire [1:0] dmem39_io_bus_request_bits_operation; // @[top.scala 288:22]
  wire  dmem39_io_bus_response_valid; // @[top.scala 288:22]
  wire [31:0] dmem39_io_bus_response_bits_data; // @[top.scala 288:22]
  wire  cpu40_clock; // @[top.scala 292:21]
  wire  cpu40_reset; // @[top.scala 292:21]
  wire [31:0] cpu40_io_imem_address; // @[top.scala 292:21]
  wire [31:0] cpu40_io_imem_instruction; // @[top.scala 292:21]
  wire [31:0] cpu40_io_dmem_address; // @[top.scala 292:21]
  wire  cpu40_io_dmem_valid; // @[top.scala 292:21]
  wire [31:0] cpu40_io_dmem_writedata; // @[top.scala 292:21]
  wire  cpu40_io_dmem_memread; // @[top.scala 292:21]
  wire  cpu40_io_dmem_memwrite; // @[top.scala 292:21]
  wire [1:0] cpu40_io_dmem_maskmode; // @[top.scala 292:21]
  wire  cpu40_io_dmem_sext; // @[top.scala 292:21]
  wire [31:0] cpu40_io_dmem_readdata; // @[top.scala 292:21]
  wire  mem40_clock; // @[top.scala 293:21]
  wire  mem40_reset; // @[top.scala 293:21]
  wire [31:0] mem40_io_imem_request_bits_address; // @[top.scala 293:21]
  wire [31:0] mem40_io_imem_response_bits_data; // @[top.scala 293:21]
  wire  mem40_io_dmem_request_valid; // @[top.scala 293:21]
  wire [31:0] mem40_io_dmem_request_bits_address; // @[top.scala 293:21]
  wire [31:0] mem40_io_dmem_request_bits_writedata; // @[top.scala 293:21]
  wire [1:0] mem40_io_dmem_request_bits_operation; // @[top.scala 293:21]
  wire  mem40_io_dmem_response_valid; // @[top.scala 293:21]
  wire [31:0] mem40_io_dmem_response_bits_data; // @[top.scala 293:21]
  wire [31:0] imem40_io_pipeline_address; // @[top.scala 294:22]
  wire [31:0] imem40_io_pipeline_instruction; // @[top.scala 294:22]
  wire [31:0] imem40_io_bus_request_bits_address; // @[top.scala 294:22]
  wire [31:0] imem40_io_bus_response_bits_data; // @[top.scala 294:22]
  wire  dmem40_clock; // @[top.scala 295:22]
  wire  dmem40_reset; // @[top.scala 295:22]
  wire [31:0] dmem40_io_pipeline_address; // @[top.scala 295:22]
  wire  dmem40_io_pipeline_valid; // @[top.scala 295:22]
  wire [31:0] dmem40_io_pipeline_writedata; // @[top.scala 295:22]
  wire  dmem40_io_pipeline_memread; // @[top.scala 295:22]
  wire  dmem40_io_pipeline_memwrite; // @[top.scala 295:22]
  wire [1:0] dmem40_io_pipeline_maskmode; // @[top.scala 295:22]
  wire  dmem40_io_pipeline_sext; // @[top.scala 295:22]
  wire [31:0] dmem40_io_pipeline_readdata; // @[top.scala 295:22]
  wire  dmem40_io_bus_request_valid; // @[top.scala 295:22]
  wire [31:0] dmem40_io_bus_request_bits_address; // @[top.scala 295:22]
  wire [31:0] dmem40_io_bus_request_bits_writedata; // @[top.scala 295:22]
  wire [1:0] dmem40_io_bus_request_bits_operation; // @[top.scala 295:22]
  wire  dmem40_io_bus_response_valid; // @[top.scala 295:22]
  wire [31:0] dmem40_io_bus_response_bits_data; // @[top.scala 295:22]
  wire  cpu41_clock; // @[top.scala 299:21]
  wire  cpu41_reset; // @[top.scala 299:21]
  wire [31:0] cpu41_io_imem_address; // @[top.scala 299:21]
  wire [31:0] cpu41_io_imem_instruction; // @[top.scala 299:21]
  wire [31:0] cpu41_io_dmem_address; // @[top.scala 299:21]
  wire  cpu41_io_dmem_valid; // @[top.scala 299:21]
  wire [31:0] cpu41_io_dmem_writedata; // @[top.scala 299:21]
  wire  cpu41_io_dmem_memread; // @[top.scala 299:21]
  wire  cpu41_io_dmem_memwrite; // @[top.scala 299:21]
  wire [1:0] cpu41_io_dmem_maskmode; // @[top.scala 299:21]
  wire  cpu41_io_dmem_sext; // @[top.scala 299:21]
  wire [31:0] cpu41_io_dmem_readdata; // @[top.scala 299:21]
  wire  mem41_clock; // @[top.scala 300:21]
  wire  mem41_reset; // @[top.scala 300:21]
  wire [31:0] mem41_io_imem_request_bits_address; // @[top.scala 300:21]
  wire [31:0] mem41_io_imem_response_bits_data; // @[top.scala 300:21]
  wire  mem41_io_dmem_request_valid; // @[top.scala 300:21]
  wire [31:0] mem41_io_dmem_request_bits_address; // @[top.scala 300:21]
  wire [31:0] mem41_io_dmem_request_bits_writedata; // @[top.scala 300:21]
  wire [1:0] mem41_io_dmem_request_bits_operation; // @[top.scala 300:21]
  wire  mem41_io_dmem_response_valid; // @[top.scala 300:21]
  wire [31:0] mem41_io_dmem_response_bits_data; // @[top.scala 300:21]
  wire [31:0] imem41_io_pipeline_address; // @[top.scala 301:22]
  wire [31:0] imem41_io_pipeline_instruction; // @[top.scala 301:22]
  wire [31:0] imem41_io_bus_request_bits_address; // @[top.scala 301:22]
  wire [31:0] imem41_io_bus_response_bits_data; // @[top.scala 301:22]
  wire  dmem41_clock; // @[top.scala 302:22]
  wire  dmem41_reset; // @[top.scala 302:22]
  wire [31:0] dmem41_io_pipeline_address; // @[top.scala 302:22]
  wire  dmem41_io_pipeline_valid; // @[top.scala 302:22]
  wire [31:0] dmem41_io_pipeline_writedata; // @[top.scala 302:22]
  wire  dmem41_io_pipeline_memread; // @[top.scala 302:22]
  wire  dmem41_io_pipeline_memwrite; // @[top.scala 302:22]
  wire [1:0] dmem41_io_pipeline_maskmode; // @[top.scala 302:22]
  wire  dmem41_io_pipeline_sext; // @[top.scala 302:22]
  wire [31:0] dmem41_io_pipeline_readdata; // @[top.scala 302:22]
  wire  dmem41_io_bus_request_valid; // @[top.scala 302:22]
  wire [31:0] dmem41_io_bus_request_bits_address; // @[top.scala 302:22]
  wire [31:0] dmem41_io_bus_request_bits_writedata; // @[top.scala 302:22]
  wire [1:0] dmem41_io_bus_request_bits_operation; // @[top.scala 302:22]
  wire  dmem41_io_bus_response_valid; // @[top.scala 302:22]
  wire [31:0] dmem41_io_bus_response_bits_data; // @[top.scala 302:22]
  wire  cpu42_clock; // @[top.scala 306:21]
  wire  cpu42_reset; // @[top.scala 306:21]
  wire [31:0] cpu42_io_imem_address; // @[top.scala 306:21]
  wire [31:0] cpu42_io_imem_instruction; // @[top.scala 306:21]
  wire [31:0] cpu42_io_dmem_address; // @[top.scala 306:21]
  wire  cpu42_io_dmem_valid; // @[top.scala 306:21]
  wire [31:0] cpu42_io_dmem_writedata; // @[top.scala 306:21]
  wire  cpu42_io_dmem_memread; // @[top.scala 306:21]
  wire  cpu42_io_dmem_memwrite; // @[top.scala 306:21]
  wire [1:0] cpu42_io_dmem_maskmode; // @[top.scala 306:21]
  wire  cpu42_io_dmem_sext; // @[top.scala 306:21]
  wire [31:0] cpu42_io_dmem_readdata; // @[top.scala 306:21]
  wire  mem42_clock; // @[top.scala 307:21]
  wire  mem42_reset; // @[top.scala 307:21]
  wire [31:0] mem42_io_imem_request_bits_address; // @[top.scala 307:21]
  wire [31:0] mem42_io_imem_response_bits_data; // @[top.scala 307:21]
  wire  mem42_io_dmem_request_valid; // @[top.scala 307:21]
  wire [31:0] mem42_io_dmem_request_bits_address; // @[top.scala 307:21]
  wire [31:0] mem42_io_dmem_request_bits_writedata; // @[top.scala 307:21]
  wire [1:0] mem42_io_dmem_request_bits_operation; // @[top.scala 307:21]
  wire  mem42_io_dmem_response_valid; // @[top.scala 307:21]
  wire [31:0] mem42_io_dmem_response_bits_data; // @[top.scala 307:21]
  wire [31:0] imem42_io_pipeline_address; // @[top.scala 308:22]
  wire [31:0] imem42_io_pipeline_instruction; // @[top.scala 308:22]
  wire [31:0] imem42_io_bus_request_bits_address; // @[top.scala 308:22]
  wire [31:0] imem42_io_bus_response_bits_data; // @[top.scala 308:22]
  wire  dmem42_clock; // @[top.scala 309:22]
  wire  dmem42_reset; // @[top.scala 309:22]
  wire [31:0] dmem42_io_pipeline_address; // @[top.scala 309:22]
  wire  dmem42_io_pipeline_valid; // @[top.scala 309:22]
  wire [31:0] dmem42_io_pipeline_writedata; // @[top.scala 309:22]
  wire  dmem42_io_pipeline_memread; // @[top.scala 309:22]
  wire  dmem42_io_pipeline_memwrite; // @[top.scala 309:22]
  wire [1:0] dmem42_io_pipeline_maskmode; // @[top.scala 309:22]
  wire  dmem42_io_pipeline_sext; // @[top.scala 309:22]
  wire [31:0] dmem42_io_pipeline_readdata; // @[top.scala 309:22]
  wire  dmem42_io_bus_request_valid; // @[top.scala 309:22]
  wire [31:0] dmem42_io_bus_request_bits_address; // @[top.scala 309:22]
  wire [31:0] dmem42_io_bus_request_bits_writedata; // @[top.scala 309:22]
  wire [1:0] dmem42_io_bus_request_bits_operation; // @[top.scala 309:22]
  wire  dmem42_io_bus_response_valid; // @[top.scala 309:22]
  wire [31:0] dmem42_io_bus_response_bits_data; // @[top.scala 309:22]
  wire  cpu43_clock; // @[top.scala 313:21]
  wire  cpu43_reset; // @[top.scala 313:21]
  wire [31:0] cpu43_io_imem_address; // @[top.scala 313:21]
  wire [31:0] cpu43_io_imem_instruction; // @[top.scala 313:21]
  wire [31:0] cpu43_io_dmem_address; // @[top.scala 313:21]
  wire  cpu43_io_dmem_valid; // @[top.scala 313:21]
  wire [31:0] cpu43_io_dmem_writedata; // @[top.scala 313:21]
  wire  cpu43_io_dmem_memread; // @[top.scala 313:21]
  wire  cpu43_io_dmem_memwrite; // @[top.scala 313:21]
  wire [1:0] cpu43_io_dmem_maskmode; // @[top.scala 313:21]
  wire  cpu43_io_dmem_sext; // @[top.scala 313:21]
  wire [31:0] cpu43_io_dmem_readdata; // @[top.scala 313:21]
  wire  mem43_clock; // @[top.scala 314:21]
  wire  mem43_reset; // @[top.scala 314:21]
  wire [31:0] mem43_io_imem_request_bits_address; // @[top.scala 314:21]
  wire [31:0] mem43_io_imem_response_bits_data; // @[top.scala 314:21]
  wire  mem43_io_dmem_request_valid; // @[top.scala 314:21]
  wire [31:0] mem43_io_dmem_request_bits_address; // @[top.scala 314:21]
  wire [31:0] mem43_io_dmem_request_bits_writedata; // @[top.scala 314:21]
  wire [1:0] mem43_io_dmem_request_bits_operation; // @[top.scala 314:21]
  wire  mem43_io_dmem_response_valid; // @[top.scala 314:21]
  wire [31:0] mem43_io_dmem_response_bits_data; // @[top.scala 314:21]
  wire [31:0] imem43_io_pipeline_address; // @[top.scala 315:22]
  wire [31:0] imem43_io_pipeline_instruction; // @[top.scala 315:22]
  wire [31:0] imem43_io_bus_request_bits_address; // @[top.scala 315:22]
  wire [31:0] imem43_io_bus_response_bits_data; // @[top.scala 315:22]
  wire  dmem43_clock; // @[top.scala 316:22]
  wire  dmem43_reset; // @[top.scala 316:22]
  wire [31:0] dmem43_io_pipeline_address; // @[top.scala 316:22]
  wire  dmem43_io_pipeline_valid; // @[top.scala 316:22]
  wire [31:0] dmem43_io_pipeline_writedata; // @[top.scala 316:22]
  wire  dmem43_io_pipeline_memread; // @[top.scala 316:22]
  wire  dmem43_io_pipeline_memwrite; // @[top.scala 316:22]
  wire [1:0] dmem43_io_pipeline_maskmode; // @[top.scala 316:22]
  wire  dmem43_io_pipeline_sext; // @[top.scala 316:22]
  wire [31:0] dmem43_io_pipeline_readdata; // @[top.scala 316:22]
  wire  dmem43_io_bus_request_valid; // @[top.scala 316:22]
  wire [31:0] dmem43_io_bus_request_bits_address; // @[top.scala 316:22]
  wire [31:0] dmem43_io_bus_request_bits_writedata; // @[top.scala 316:22]
  wire [1:0] dmem43_io_bus_request_bits_operation; // @[top.scala 316:22]
  wire  dmem43_io_bus_response_valid; // @[top.scala 316:22]
  wire [31:0] dmem43_io_bus_response_bits_data; // @[top.scala 316:22]
  wire  cpu44_clock; // @[top.scala 320:21]
  wire  cpu44_reset; // @[top.scala 320:21]
  wire [31:0] cpu44_io_imem_address; // @[top.scala 320:21]
  wire [31:0] cpu44_io_imem_instruction; // @[top.scala 320:21]
  wire [31:0] cpu44_io_dmem_address; // @[top.scala 320:21]
  wire  cpu44_io_dmem_valid; // @[top.scala 320:21]
  wire [31:0] cpu44_io_dmem_writedata; // @[top.scala 320:21]
  wire  cpu44_io_dmem_memread; // @[top.scala 320:21]
  wire  cpu44_io_dmem_memwrite; // @[top.scala 320:21]
  wire [1:0] cpu44_io_dmem_maskmode; // @[top.scala 320:21]
  wire  cpu44_io_dmem_sext; // @[top.scala 320:21]
  wire [31:0] cpu44_io_dmem_readdata; // @[top.scala 320:21]
  wire  mem44_clock; // @[top.scala 321:21]
  wire  mem44_reset; // @[top.scala 321:21]
  wire [31:0] mem44_io_imem_request_bits_address; // @[top.scala 321:21]
  wire [31:0] mem44_io_imem_response_bits_data; // @[top.scala 321:21]
  wire  mem44_io_dmem_request_valid; // @[top.scala 321:21]
  wire [31:0] mem44_io_dmem_request_bits_address; // @[top.scala 321:21]
  wire [31:0] mem44_io_dmem_request_bits_writedata; // @[top.scala 321:21]
  wire [1:0] mem44_io_dmem_request_bits_operation; // @[top.scala 321:21]
  wire  mem44_io_dmem_response_valid; // @[top.scala 321:21]
  wire [31:0] mem44_io_dmem_response_bits_data; // @[top.scala 321:21]
  wire [31:0] imem44_io_pipeline_address; // @[top.scala 322:22]
  wire [31:0] imem44_io_pipeline_instruction; // @[top.scala 322:22]
  wire [31:0] imem44_io_bus_request_bits_address; // @[top.scala 322:22]
  wire [31:0] imem44_io_bus_response_bits_data; // @[top.scala 322:22]
  wire  dmem44_clock; // @[top.scala 323:22]
  wire  dmem44_reset; // @[top.scala 323:22]
  wire [31:0] dmem44_io_pipeline_address; // @[top.scala 323:22]
  wire  dmem44_io_pipeline_valid; // @[top.scala 323:22]
  wire [31:0] dmem44_io_pipeline_writedata; // @[top.scala 323:22]
  wire  dmem44_io_pipeline_memread; // @[top.scala 323:22]
  wire  dmem44_io_pipeline_memwrite; // @[top.scala 323:22]
  wire [1:0] dmem44_io_pipeline_maskmode; // @[top.scala 323:22]
  wire  dmem44_io_pipeline_sext; // @[top.scala 323:22]
  wire [31:0] dmem44_io_pipeline_readdata; // @[top.scala 323:22]
  wire  dmem44_io_bus_request_valid; // @[top.scala 323:22]
  wire [31:0] dmem44_io_bus_request_bits_address; // @[top.scala 323:22]
  wire [31:0] dmem44_io_bus_request_bits_writedata; // @[top.scala 323:22]
  wire [1:0] dmem44_io_bus_request_bits_operation; // @[top.scala 323:22]
  wire  dmem44_io_bus_response_valid; // @[top.scala 323:22]
  wire [31:0] dmem44_io_bus_response_bits_data; // @[top.scala 323:22]
  wire  cpu45_clock; // @[top.scala 327:21]
  wire  cpu45_reset; // @[top.scala 327:21]
  wire [31:0] cpu45_io_imem_address; // @[top.scala 327:21]
  wire [31:0] cpu45_io_imem_instruction; // @[top.scala 327:21]
  wire [31:0] cpu45_io_dmem_address; // @[top.scala 327:21]
  wire  cpu45_io_dmem_valid; // @[top.scala 327:21]
  wire [31:0] cpu45_io_dmem_writedata; // @[top.scala 327:21]
  wire  cpu45_io_dmem_memread; // @[top.scala 327:21]
  wire  cpu45_io_dmem_memwrite; // @[top.scala 327:21]
  wire [1:0] cpu45_io_dmem_maskmode; // @[top.scala 327:21]
  wire  cpu45_io_dmem_sext; // @[top.scala 327:21]
  wire [31:0] cpu45_io_dmem_readdata; // @[top.scala 327:21]
  wire  mem45_clock; // @[top.scala 328:21]
  wire  mem45_reset; // @[top.scala 328:21]
  wire [31:0] mem45_io_imem_request_bits_address; // @[top.scala 328:21]
  wire [31:0] mem45_io_imem_response_bits_data; // @[top.scala 328:21]
  wire  mem45_io_dmem_request_valid; // @[top.scala 328:21]
  wire [31:0] mem45_io_dmem_request_bits_address; // @[top.scala 328:21]
  wire [31:0] mem45_io_dmem_request_bits_writedata; // @[top.scala 328:21]
  wire [1:0] mem45_io_dmem_request_bits_operation; // @[top.scala 328:21]
  wire  mem45_io_dmem_response_valid; // @[top.scala 328:21]
  wire [31:0] mem45_io_dmem_response_bits_data; // @[top.scala 328:21]
  wire [31:0] imem45_io_pipeline_address; // @[top.scala 329:22]
  wire [31:0] imem45_io_pipeline_instruction; // @[top.scala 329:22]
  wire [31:0] imem45_io_bus_request_bits_address; // @[top.scala 329:22]
  wire [31:0] imem45_io_bus_response_bits_data; // @[top.scala 329:22]
  wire  dmem45_clock; // @[top.scala 330:22]
  wire  dmem45_reset; // @[top.scala 330:22]
  wire [31:0] dmem45_io_pipeline_address; // @[top.scala 330:22]
  wire  dmem45_io_pipeline_valid; // @[top.scala 330:22]
  wire [31:0] dmem45_io_pipeline_writedata; // @[top.scala 330:22]
  wire  dmem45_io_pipeline_memread; // @[top.scala 330:22]
  wire  dmem45_io_pipeline_memwrite; // @[top.scala 330:22]
  wire [1:0] dmem45_io_pipeline_maskmode; // @[top.scala 330:22]
  wire  dmem45_io_pipeline_sext; // @[top.scala 330:22]
  wire [31:0] dmem45_io_pipeline_readdata; // @[top.scala 330:22]
  wire  dmem45_io_bus_request_valid; // @[top.scala 330:22]
  wire [31:0] dmem45_io_bus_request_bits_address; // @[top.scala 330:22]
  wire [31:0] dmem45_io_bus_request_bits_writedata; // @[top.scala 330:22]
  wire [1:0] dmem45_io_bus_request_bits_operation; // @[top.scala 330:22]
  wire  dmem45_io_bus_response_valid; // @[top.scala 330:22]
  wire [31:0] dmem45_io_bus_response_bits_data; // @[top.scala 330:22]
  wire  cpu46_clock; // @[top.scala 334:21]
  wire  cpu46_reset; // @[top.scala 334:21]
  wire [31:0] cpu46_io_imem_address; // @[top.scala 334:21]
  wire [31:0] cpu46_io_imem_instruction; // @[top.scala 334:21]
  wire [31:0] cpu46_io_dmem_address; // @[top.scala 334:21]
  wire  cpu46_io_dmem_valid; // @[top.scala 334:21]
  wire [31:0] cpu46_io_dmem_writedata; // @[top.scala 334:21]
  wire  cpu46_io_dmem_memread; // @[top.scala 334:21]
  wire  cpu46_io_dmem_memwrite; // @[top.scala 334:21]
  wire [1:0] cpu46_io_dmem_maskmode; // @[top.scala 334:21]
  wire  cpu46_io_dmem_sext; // @[top.scala 334:21]
  wire [31:0] cpu46_io_dmem_readdata; // @[top.scala 334:21]
  wire  mem46_clock; // @[top.scala 335:21]
  wire  mem46_reset; // @[top.scala 335:21]
  wire [31:0] mem46_io_imem_request_bits_address; // @[top.scala 335:21]
  wire [31:0] mem46_io_imem_response_bits_data; // @[top.scala 335:21]
  wire  mem46_io_dmem_request_valid; // @[top.scala 335:21]
  wire [31:0] mem46_io_dmem_request_bits_address; // @[top.scala 335:21]
  wire [31:0] mem46_io_dmem_request_bits_writedata; // @[top.scala 335:21]
  wire [1:0] mem46_io_dmem_request_bits_operation; // @[top.scala 335:21]
  wire  mem46_io_dmem_response_valid; // @[top.scala 335:21]
  wire [31:0] mem46_io_dmem_response_bits_data; // @[top.scala 335:21]
  wire [31:0] imem46_io_pipeline_address; // @[top.scala 336:22]
  wire [31:0] imem46_io_pipeline_instruction; // @[top.scala 336:22]
  wire [31:0] imem46_io_bus_request_bits_address; // @[top.scala 336:22]
  wire [31:0] imem46_io_bus_response_bits_data; // @[top.scala 336:22]
  wire  dmem46_clock; // @[top.scala 337:22]
  wire  dmem46_reset; // @[top.scala 337:22]
  wire [31:0] dmem46_io_pipeline_address; // @[top.scala 337:22]
  wire  dmem46_io_pipeline_valid; // @[top.scala 337:22]
  wire [31:0] dmem46_io_pipeline_writedata; // @[top.scala 337:22]
  wire  dmem46_io_pipeline_memread; // @[top.scala 337:22]
  wire  dmem46_io_pipeline_memwrite; // @[top.scala 337:22]
  wire [1:0] dmem46_io_pipeline_maskmode; // @[top.scala 337:22]
  wire  dmem46_io_pipeline_sext; // @[top.scala 337:22]
  wire [31:0] dmem46_io_pipeline_readdata; // @[top.scala 337:22]
  wire  dmem46_io_bus_request_valid; // @[top.scala 337:22]
  wire [31:0] dmem46_io_bus_request_bits_address; // @[top.scala 337:22]
  wire [31:0] dmem46_io_bus_request_bits_writedata; // @[top.scala 337:22]
  wire [1:0] dmem46_io_bus_request_bits_operation; // @[top.scala 337:22]
  wire  dmem46_io_bus_response_valid; // @[top.scala 337:22]
  wire [31:0] dmem46_io_bus_response_bits_data; // @[top.scala 337:22]
  wire  cpu47_clock; // @[top.scala 341:21]
  wire  cpu47_reset; // @[top.scala 341:21]
  wire [31:0] cpu47_io_imem_address; // @[top.scala 341:21]
  wire [31:0] cpu47_io_imem_instruction; // @[top.scala 341:21]
  wire [31:0] cpu47_io_dmem_address; // @[top.scala 341:21]
  wire  cpu47_io_dmem_valid; // @[top.scala 341:21]
  wire [31:0] cpu47_io_dmem_writedata; // @[top.scala 341:21]
  wire  cpu47_io_dmem_memread; // @[top.scala 341:21]
  wire  cpu47_io_dmem_memwrite; // @[top.scala 341:21]
  wire [1:0] cpu47_io_dmem_maskmode; // @[top.scala 341:21]
  wire  cpu47_io_dmem_sext; // @[top.scala 341:21]
  wire [31:0] cpu47_io_dmem_readdata; // @[top.scala 341:21]
  wire  mem47_clock; // @[top.scala 342:21]
  wire  mem47_reset; // @[top.scala 342:21]
  wire [31:0] mem47_io_imem_request_bits_address; // @[top.scala 342:21]
  wire [31:0] mem47_io_imem_response_bits_data; // @[top.scala 342:21]
  wire  mem47_io_dmem_request_valid; // @[top.scala 342:21]
  wire [31:0] mem47_io_dmem_request_bits_address; // @[top.scala 342:21]
  wire [31:0] mem47_io_dmem_request_bits_writedata; // @[top.scala 342:21]
  wire [1:0] mem47_io_dmem_request_bits_operation; // @[top.scala 342:21]
  wire  mem47_io_dmem_response_valid; // @[top.scala 342:21]
  wire [31:0] mem47_io_dmem_response_bits_data; // @[top.scala 342:21]
  wire [31:0] imem47_io_pipeline_address; // @[top.scala 343:22]
  wire [31:0] imem47_io_pipeline_instruction; // @[top.scala 343:22]
  wire [31:0] imem47_io_bus_request_bits_address; // @[top.scala 343:22]
  wire [31:0] imem47_io_bus_response_bits_data; // @[top.scala 343:22]
  wire  dmem47_clock; // @[top.scala 344:22]
  wire  dmem47_reset; // @[top.scala 344:22]
  wire [31:0] dmem47_io_pipeline_address; // @[top.scala 344:22]
  wire  dmem47_io_pipeline_valid; // @[top.scala 344:22]
  wire [31:0] dmem47_io_pipeline_writedata; // @[top.scala 344:22]
  wire  dmem47_io_pipeline_memread; // @[top.scala 344:22]
  wire  dmem47_io_pipeline_memwrite; // @[top.scala 344:22]
  wire [1:0] dmem47_io_pipeline_maskmode; // @[top.scala 344:22]
  wire  dmem47_io_pipeline_sext; // @[top.scala 344:22]
  wire [31:0] dmem47_io_pipeline_readdata; // @[top.scala 344:22]
  wire  dmem47_io_bus_request_valid; // @[top.scala 344:22]
  wire [31:0] dmem47_io_bus_request_bits_address; // @[top.scala 344:22]
  wire [31:0] dmem47_io_bus_request_bits_writedata; // @[top.scala 344:22]
  wire [1:0] dmem47_io_bus_request_bits_operation; // @[top.scala 344:22]
  wire  dmem47_io_bus_response_valid; // @[top.scala 344:22]
  wire [31:0] dmem47_io_bus_response_bits_data; // @[top.scala 344:22]
  wire  cpu48_clock; // @[top.scala 348:21]
  wire  cpu48_reset; // @[top.scala 348:21]
  wire [31:0] cpu48_io_imem_address; // @[top.scala 348:21]
  wire [31:0] cpu48_io_imem_instruction; // @[top.scala 348:21]
  wire [31:0] cpu48_io_dmem_address; // @[top.scala 348:21]
  wire  cpu48_io_dmem_valid; // @[top.scala 348:21]
  wire [31:0] cpu48_io_dmem_writedata; // @[top.scala 348:21]
  wire  cpu48_io_dmem_memread; // @[top.scala 348:21]
  wire  cpu48_io_dmem_memwrite; // @[top.scala 348:21]
  wire [1:0] cpu48_io_dmem_maskmode; // @[top.scala 348:21]
  wire  cpu48_io_dmem_sext; // @[top.scala 348:21]
  wire [31:0] cpu48_io_dmem_readdata; // @[top.scala 348:21]
  wire  mem48_clock; // @[top.scala 349:21]
  wire  mem48_reset; // @[top.scala 349:21]
  wire [31:0] mem48_io_imem_request_bits_address; // @[top.scala 349:21]
  wire [31:0] mem48_io_imem_response_bits_data; // @[top.scala 349:21]
  wire  mem48_io_dmem_request_valid; // @[top.scala 349:21]
  wire [31:0] mem48_io_dmem_request_bits_address; // @[top.scala 349:21]
  wire [31:0] mem48_io_dmem_request_bits_writedata; // @[top.scala 349:21]
  wire [1:0] mem48_io_dmem_request_bits_operation; // @[top.scala 349:21]
  wire  mem48_io_dmem_response_valid; // @[top.scala 349:21]
  wire [31:0] mem48_io_dmem_response_bits_data; // @[top.scala 349:21]
  wire [31:0] imem48_io_pipeline_address; // @[top.scala 350:22]
  wire [31:0] imem48_io_pipeline_instruction; // @[top.scala 350:22]
  wire [31:0] imem48_io_bus_request_bits_address; // @[top.scala 350:22]
  wire [31:0] imem48_io_bus_response_bits_data; // @[top.scala 350:22]
  wire  dmem48_clock; // @[top.scala 351:22]
  wire  dmem48_reset; // @[top.scala 351:22]
  wire [31:0] dmem48_io_pipeline_address; // @[top.scala 351:22]
  wire  dmem48_io_pipeline_valid; // @[top.scala 351:22]
  wire [31:0] dmem48_io_pipeline_writedata; // @[top.scala 351:22]
  wire  dmem48_io_pipeline_memread; // @[top.scala 351:22]
  wire  dmem48_io_pipeline_memwrite; // @[top.scala 351:22]
  wire [1:0] dmem48_io_pipeline_maskmode; // @[top.scala 351:22]
  wire  dmem48_io_pipeline_sext; // @[top.scala 351:22]
  wire [31:0] dmem48_io_pipeline_readdata; // @[top.scala 351:22]
  wire  dmem48_io_bus_request_valid; // @[top.scala 351:22]
  wire [31:0] dmem48_io_bus_request_bits_address; // @[top.scala 351:22]
  wire [31:0] dmem48_io_bus_request_bits_writedata; // @[top.scala 351:22]
  wire [1:0] dmem48_io_bus_request_bits_operation; // @[top.scala 351:22]
  wire  dmem48_io_bus_response_valid; // @[top.scala 351:22]
  wire [31:0] dmem48_io_bus_response_bits_data; // @[top.scala 351:22]
  wire  cpu49_clock; // @[top.scala 355:21]
  wire  cpu49_reset; // @[top.scala 355:21]
  wire [31:0] cpu49_io_imem_address; // @[top.scala 355:21]
  wire [31:0] cpu49_io_imem_instruction; // @[top.scala 355:21]
  wire [31:0] cpu49_io_dmem_address; // @[top.scala 355:21]
  wire  cpu49_io_dmem_valid; // @[top.scala 355:21]
  wire [31:0] cpu49_io_dmem_writedata; // @[top.scala 355:21]
  wire  cpu49_io_dmem_memread; // @[top.scala 355:21]
  wire  cpu49_io_dmem_memwrite; // @[top.scala 355:21]
  wire [1:0] cpu49_io_dmem_maskmode; // @[top.scala 355:21]
  wire  cpu49_io_dmem_sext; // @[top.scala 355:21]
  wire [31:0] cpu49_io_dmem_readdata; // @[top.scala 355:21]
  wire  mem49_clock; // @[top.scala 356:21]
  wire  mem49_reset; // @[top.scala 356:21]
  wire [31:0] mem49_io_imem_request_bits_address; // @[top.scala 356:21]
  wire [31:0] mem49_io_imem_response_bits_data; // @[top.scala 356:21]
  wire  mem49_io_dmem_request_valid; // @[top.scala 356:21]
  wire [31:0] mem49_io_dmem_request_bits_address; // @[top.scala 356:21]
  wire [31:0] mem49_io_dmem_request_bits_writedata; // @[top.scala 356:21]
  wire [1:0] mem49_io_dmem_request_bits_operation; // @[top.scala 356:21]
  wire  mem49_io_dmem_response_valid; // @[top.scala 356:21]
  wire [31:0] mem49_io_dmem_response_bits_data; // @[top.scala 356:21]
  wire [31:0] imem49_io_pipeline_address; // @[top.scala 357:22]
  wire [31:0] imem49_io_pipeline_instruction; // @[top.scala 357:22]
  wire [31:0] imem49_io_bus_request_bits_address; // @[top.scala 357:22]
  wire [31:0] imem49_io_bus_response_bits_data; // @[top.scala 357:22]
  wire  dmem49_clock; // @[top.scala 358:22]
  wire  dmem49_reset; // @[top.scala 358:22]
  wire [31:0] dmem49_io_pipeline_address; // @[top.scala 358:22]
  wire  dmem49_io_pipeline_valid; // @[top.scala 358:22]
  wire [31:0] dmem49_io_pipeline_writedata; // @[top.scala 358:22]
  wire  dmem49_io_pipeline_memread; // @[top.scala 358:22]
  wire  dmem49_io_pipeline_memwrite; // @[top.scala 358:22]
  wire [1:0] dmem49_io_pipeline_maskmode; // @[top.scala 358:22]
  wire  dmem49_io_pipeline_sext; // @[top.scala 358:22]
  wire [31:0] dmem49_io_pipeline_readdata; // @[top.scala 358:22]
  wire  dmem49_io_bus_request_valid; // @[top.scala 358:22]
  wire [31:0] dmem49_io_bus_request_bits_address; // @[top.scala 358:22]
  wire [31:0] dmem49_io_bus_request_bits_writedata; // @[top.scala 358:22]
  wire [1:0] dmem49_io_bus_request_bits_operation; // @[top.scala 358:22]
  wire  dmem49_io_bus_response_valid; // @[top.scala 358:22]
  wire [31:0] dmem49_io_bus_response_bits_data; // @[top.scala 358:22]
  wire  cpu50_clock; // @[top.scala 362:21]
  wire  cpu50_reset; // @[top.scala 362:21]
  wire [31:0] cpu50_io_imem_address; // @[top.scala 362:21]
  wire [31:0] cpu50_io_imem_instruction; // @[top.scala 362:21]
  wire [31:0] cpu50_io_dmem_address; // @[top.scala 362:21]
  wire  cpu50_io_dmem_valid; // @[top.scala 362:21]
  wire [31:0] cpu50_io_dmem_writedata; // @[top.scala 362:21]
  wire  cpu50_io_dmem_memread; // @[top.scala 362:21]
  wire  cpu50_io_dmem_memwrite; // @[top.scala 362:21]
  wire [1:0] cpu50_io_dmem_maskmode; // @[top.scala 362:21]
  wire  cpu50_io_dmem_sext; // @[top.scala 362:21]
  wire [31:0] cpu50_io_dmem_readdata; // @[top.scala 362:21]
  wire  mem50_clock; // @[top.scala 363:21]
  wire  mem50_reset; // @[top.scala 363:21]
  wire [31:0] mem50_io_imem_request_bits_address; // @[top.scala 363:21]
  wire [31:0] mem50_io_imem_response_bits_data; // @[top.scala 363:21]
  wire  mem50_io_dmem_request_valid; // @[top.scala 363:21]
  wire [31:0] mem50_io_dmem_request_bits_address; // @[top.scala 363:21]
  wire [31:0] mem50_io_dmem_request_bits_writedata; // @[top.scala 363:21]
  wire [1:0] mem50_io_dmem_request_bits_operation; // @[top.scala 363:21]
  wire  mem50_io_dmem_response_valid; // @[top.scala 363:21]
  wire [31:0] mem50_io_dmem_response_bits_data; // @[top.scala 363:21]
  wire [31:0] imem50_io_pipeline_address; // @[top.scala 364:22]
  wire [31:0] imem50_io_pipeline_instruction; // @[top.scala 364:22]
  wire [31:0] imem50_io_bus_request_bits_address; // @[top.scala 364:22]
  wire [31:0] imem50_io_bus_response_bits_data; // @[top.scala 364:22]
  wire  dmem50_clock; // @[top.scala 365:22]
  wire  dmem50_reset; // @[top.scala 365:22]
  wire [31:0] dmem50_io_pipeline_address; // @[top.scala 365:22]
  wire  dmem50_io_pipeline_valid; // @[top.scala 365:22]
  wire [31:0] dmem50_io_pipeline_writedata; // @[top.scala 365:22]
  wire  dmem50_io_pipeline_memread; // @[top.scala 365:22]
  wire  dmem50_io_pipeline_memwrite; // @[top.scala 365:22]
  wire [1:0] dmem50_io_pipeline_maskmode; // @[top.scala 365:22]
  wire  dmem50_io_pipeline_sext; // @[top.scala 365:22]
  wire [31:0] dmem50_io_pipeline_readdata; // @[top.scala 365:22]
  wire  dmem50_io_bus_request_valid; // @[top.scala 365:22]
  wire [31:0] dmem50_io_bus_request_bits_address; // @[top.scala 365:22]
  wire [31:0] dmem50_io_bus_request_bits_writedata; // @[top.scala 365:22]
  wire [1:0] dmem50_io_bus_request_bits_operation; // @[top.scala 365:22]
  wire  dmem50_io_bus_response_valid; // @[top.scala 365:22]
  wire [31:0] dmem50_io_bus_response_bits_data; // @[top.scala 365:22]
  wire  cpu51_clock; // @[top.scala 369:21]
  wire  cpu51_reset; // @[top.scala 369:21]
  wire [31:0] cpu51_io_imem_address; // @[top.scala 369:21]
  wire [31:0] cpu51_io_imem_instruction; // @[top.scala 369:21]
  wire [31:0] cpu51_io_dmem_address; // @[top.scala 369:21]
  wire  cpu51_io_dmem_valid; // @[top.scala 369:21]
  wire [31:0] cpu51_io_dmem_writedata; // @[top.scala 369:21]
  wire  cpu51_io_dmem_memread; // @[top.scala 369:21]
  wire  cpu51_io_dmem_memwrite; // @[top.scala 369:21]
  wire [1:0] cpu51_io_dmem_maskmode; // @[top.scala 369:21]
  wire  cpu51_io_dmem_sext; // @[top.scala 369:21]
  wire [31:0] cpu51_io_dmem_readdata; // @[top.scala 369:21]
  wire  mem51_clock; // @[top.scala 370:21]
  wire  mem51_reset; // @[top.scala 370:21]
  wire [31:0] mem51_io_imem_request_bits_address; // @[top.scala 370:21]
  wire [31:0] mem51_io_imem_response_bits_data; // @[top.scala 370:21]
  wire  mem51_io_dmem_request_valid; // @[top.scala 370:21]
  wire [31:0] mem51_io_dmem_request_bits_address; // @[top.scala 370:21]
  wire [31:0] mem51_io_dmem_request_bits_writedata; // @[top.scala 370:21]
  wire [1:0] mem51_io_dmem_request_bits_operation; // @[top.scala 370:21]
  wire  mem51_io_dmem_response_valid; // @[top.scala 370:21]
  wire [31:0] mem51_io_dmem_response_bits_data; // @[top.scala 370:21]
  wire [31:0] imem51_io_pipeline_address; // @[top.scala 371:22]
  wire [31:0] imem51_io_pipeline_instruction; // @[top.scala 371:22]
  wire [31:0] imem51_io_bus_request_bits_address; // @[top.scala 371:22]
  wire [31:0] imem51_io_bus_response_bits_data; // @[top.scala 371:22]
  wire  dmem51_clock; // @[top.scala 372:22]
  wire  dmem51_reset; // @[top.scala 372:22]
  wire [31:0] dmem51_io_pipeline_address; // @[top.scala 372:22]
  wire  dmem51_io_pipeline_valid; // @[top.scala 372:22]
  wire [31:0] dmem51_io_pipeline_writedata; // @[top.scala 372:22]
  wire  dmem51_io_pipeline_memread; // @[top.scala 372:22]
  wire  dmem51_io_pipeline_memwrite; // @[top.scala 372:22]
  wire [1:0] dmem51_io_pipeline_maskmode; // @[top.scala 372:22]
  wire  dmem51_io_pipeline_sext; // @[top.scala 372:22]
  wire [31:0] dmem51_io_pipeline_readdata; // @[top.scala 372:22]
  wire  dmem51_io_bus_request_valid; // @[top.scala 372:22]
  wire [31:0] dmem51_io_bus_request_bits_address; // @[top.scala 372:22]
  wire [31:0] dmem51_io_bus_request_bits_writedata; // @[top.scala 372:22]
  wire [1:0] dmem51_io_bus_request_bits_operation; // @[top.scala 372:22]
  wire  dmem51_io_bus_response_valid; // @[top.scala 372:22]
  wire [31:0] dmem51_io_bus_response_bits_data; // @[top.scala 372:22]
  wire  cpu52_clock; // @[top.scala 376:21]
  wire  cpu52_reset; // @[top.scala 376:21]
  wire [31:0] cpu52_io_imem_address; // @[top.scala 376:21]
  wire [31:0] cpu52_io_imem_instruction; // @[top.scala 376:21]
  wire [31:0] cpu52_io_dmem_address; // @[top.scala 376:21]
  wire  cpu52_io_dmem_valid; // @[top.scala 376:21]
  wire [31:0] cpu52_io_dmem_writedata; // @[top.scala 376:21]
  wire  cpu52_io_dmem_memread; // @[top.scala 376:21]
  wire  cpu52_io_dmem_memwrite; // @[top.scala 376:21]
  wire [1:0] cpu52_io_dmem_maskmode; // @[top.scala 376:21]
  wire  cpu52_io_dmem_sext; // @[top.scala 376:21]
  wire [31:0] cpu52_io_dmem_readdata; // @[top.scala 376:21]
  wire  mem52_clock; // @[top.scala 377:21]
  wire  mem52_reset; // @[top.scala 377:21]
  wire [31:0] mem52_io_imem_request_bits_address; // @[top.scala 377:21]
  wire [31:0] mem52_io_imem_response_bits_data; // @[top.scala 377:21]
  wire  mem52_io_dmem_request_valid; // @[top.scala 377:21]
  wire [31:0] mem52_io_dmem_request_bits_address; // @[top.scala 377:21]
  wire [31:0] mem52_io_dmem_request_bits_writedata; // @[top.scala 377:21]
  wire [1:0] mem52_io_dmem_request_bits_operation; // @[top.scala 377:21]
  wire  mem52_io_dmem_response_valid; // @[top.scala 377:21]
  wire [31:0] mem52_io_dmem_response_bits_data; // @[top.scala 377:21]
  wire [31:0] imem52_io_pipeline_address; // @[top.scala 378:22]
  wire [31:0] imem52_io_pipeline_instruction; // @[top.scala 378:22]
  wire [31:0] imem52_io_bus_request_bits_address; // @[top.scala 378:22]
  wire [31:0] imem52_io_bus_response_bits_data; // @[top.scala 378:22]
  wire  dmem52_clock; // @[top.scala 379:22]
  wire  dmem52_reset; // @[top.scala 379:22]
  wire [31:0] dmem52_io_pipeline_address; // @[top.scala 379:22]
  wire  dmem52_io_pipeline_valid; // @[top.scala 379:22]
  wire [31:0] dmem52_io_pipeline_writedata; // @[top.scala 379:22]
  wire  dmem52_io_pipeline_memread; // @[top.scala 379:22]
  wire  dmem52_io_pipeline_memwrite; // @[top.scala 379:22]
  wire [1:0] dmem52_io_pipeline_maskmode; // @[top.scala 379:22]
  wire  dmem52_io_pipeline_sext; // @[top.scala 379:22]
  wire [31:0] dmem52_io_pipeline_readdata; // @[top.scala 379:22]
  wire  dmem52_io_bus_request_valid; // @[top.scala 379:22]
  wire [31:0] dmem52_io_bus_request_bits_address; // @[top.scala 379:22]
  wire [31:0] dmem52_io_bus_request_bits_writedata; // @[top.scala 379:22]
  wire [1:0] dmem52_io_bus_request_bits_operation; // @[top.scala 379:22]
  wire  dmem52_io_bus_response_valid; // @[top.scala 379:22]
  wire [31:0] dmem52_io_bus_response_bits_data; // @[top.scala 379:22]
  wire  cpu53_clock; // @[top.scala 383:21]
  wire  cpu53_reset; // @[top.scala 383:21]
  wire [31:0] cpu53_io_imem_address; // @[top.scala 383:21]
  wire [31:0] cpu53_io_imem_instruction; // @[top.scala 383:21]
  wire [31:0] cpu53_io_dmem_address; // @[top.scala 383:21]
  wire  cpu53_io_dmem_valid; // @[top.scala 383:21]
  wire [31:0] cpu53_io_dmem_writedata; // @[top.scala 383:21]
  wire  cpu53_io_dmem_memread; // @[top.scala 383:21]
  wire  cpu53_io_dmem_memwrite; // @[top.scala 383:21]
  wire [1:0] cpu53_io_dmem_maskmode; // @[top.scala 383:21]
  wire  cpu53_io_dmem_sext; // @[top.scala 383:21]
  wire [31:0] cpu53_io_dmem_readdata; // @[top.scala 383:21]
  wire  mem53_clock; // @[top.scala 384:21]
  wire  mem53_reset; // @[top.scala 384:21]
  wire [31:0] mem53_io_imem_request_bits_address; // @[top.scala 384:21]
  wire [31:0] mem53_io_imem_response_bits_data; // @[top.scala 384:21]
  wire  mem53_io_dmem_request_valid; // @[top.scala 384:21]
  wire [31:0] mem53_io_dmem_request_bits_address; // @[top.scala 384:21]
  wire [31:0] mem53_io_dmem_request_bits_writedata; // @[top.scala 384:21]
  wire [1:0] mem53_io_dmem_request_bits_operation; // @[top.scala 384:21]
  wire  mem53_io_dmem_response_valid; // @[top.scala 384:21]
  wire [31:0] mem53_io_dmem_response_bits_data; // @[top.scala 384:21]
  wire [31:0] imem53_io_pipeline_address; // @[top.scala 385:22]
  wire [31:0] imem53_io_pipeline_instruction; // @[top.scala 385:22]
  wire [31:0] imem53_io_bus_request_bits_address; // @[top.scala 385:22]
  wire [31:0] imem53_io_bus_response_bits_data; // @[top.scala 385:22]
  wire  dmem53_clock; // @[top.scala 386:22]
  wire  dmem53_reset; // @[top.scala 386:22]
  wire [31:0] dmem53_io_pipeline_address; // @[top.scala 386:22]
  wire  dmem53_io_pipeline_valid; // @[top.scala 386:22]
  wire [31:0] dmem53_io_pipeline_writedata; // @[top.scala 386:22]
  wire  dmem53_io_pipeline_memread; // @[top.scala 386:22]
  wire  dmem53_io_pipeline_memwrite; // @[top.scala 386:22]
  wire [1:0] dmem53_io_pipeline_maskmode; // @[top.scala 386:22]
  wire  dmem53_io_pipeline_sext; // @[top.scala 386:22]
  wire [31:0] dmem53_io_pipeline_readdata; // @[top.scala 386:22]
  wire  dmem53_io_bus_request_valid; // @[top.scala 386:22]
  wire [31:0] dmem53_io_bus_request_bits_address; // @[top.scala 386:22]
  wire [31:0] dmem53_io_bus_request_bits_writedata; // @[top.scala 386:22]
  wire [1:0] dmem53_io_bus_request_bits_operation; // @[top.scala 386:22]
  wire  dmem53_io_bus_response_valid; // @[top.scala 386:22]
  wire [31:0] dmem53_io_bus_response_bits_data; // @[top.scala 386:22]
  wire  cpu54_clock; // @[top.scala 390:21]
  wire  cpu54_reset; // @[top.scala 390:21]
  wire [31:0] cpu54_io_imem_address; // @[top.scala 390:21]
  wire [31:0] cpu54_io_imem_instruction; // @[top.scala 390:21]
  wire [31:0] cpu54_io_dmem_address; // @[top.scala 390:21]
  wire  cpu54_io_dmem_valid; // @[top.scala 390:21]
  wire [31:0] cpu54_io_dmem_writedata; // @[top.scala 390:21]
  wire  cpu54_io_dmem_memread; // @[top.scala 390:21]
  wire  cpu54_io_dmem_memwrite; // @[top.scala 390:21]
  wire [1:0] cpu54_io_dmem_maskmode; // @[top.scala 390:21]
  wire  cpu54_io_dmem_sext; // @[top.scala 390:21]
  wire [31:0] cpu54_io_dmem_readdata; // @[top.scala 390:21]
  wire  mem54_clock; // @[top.scala 391:21]
  wire  mem54_reset; // @[top.scala 391:21]
  wire [31:0] mem54_io_imem_request_bits_address; // @[top.scala 391:21]
  wire [31:0] mem54_io_imem_response_bits_data; // @[top.scala 391:21]
  wire  mem54_io_dmem_request_valid; // @[top.scala 391:21]
  wire [31:0] mem54_io_dmem_request_bits_address; // @[top.scala 391:21]
  wire [31:0] mem54_io_dmem_request_bits_writedata; // @[top.scala 391:21]
  wire [1:0] mem54_io_dmem_request_bits_operation; // @[top.scala 391:21]
  wire  mem54_io_dmem_response_valid; // @[top.scala 391:21]
  wire [31:0] mem54_io_dmem_response_bits_data; // @[top.scala 391:21]
  wire [31:0] imem54_io_pipeline_address; // @[top.scala 392:22]
  wire [31:0] imem54_io_pipeline_instruction; // @[top.scala 392:22]
  wire [31:0] imem54_io_bus_request_bits_address; // @[top.scala 392:22]
  wire [31:0] imem54_io_bus_response_bits_data; // @[top.scala 392:22]
  wire  dmem54_clock; // @[top.scala 393:22]
  wire  dmem54_reset; // @[top.scala 393:22]
  wire [31:0] dmem54_io_pipeline_address; // @[top.scala 393:22]
  wire  dmem54_io_pipeline_valid; // @[top.scala 393:22]
  wire [31:0] dmem54_io_pipeline_writedata; // @[top.scala 393:22]
  wire  dmem54_io_pipeline_memread; // @[top.scala 393:22]
  wire  dmem54_io_pipeline_memwrite; // @[top.scala 393:22]
  wire [1:0] dmem54_io_pipeline_maskmode; // @[top.scala 393:22]
  wire  dmem54_io_pipeline_sext; // @[top.scala 393:22]
  wire [31:0] dmem54_io_pipeline_readdata; // @[top.scala 393:22]
  wire  dmem54_io_bus_request_valid; // @[top.scala 393:22]
  wire [31:0] dmem54_io_bus_request_bits_address; // @[top.scala 393:22]
  wire [31:0] dmem54_io_bus_request_bits_writedata; // @[top.scala 393:22]
  wire [1:0] dmem54_io_bus_request_bits_operation; // @[top.scala 393:22]
  wire  dmem54_io_bus_response_valid; // @[top.scala 393:22]
  wire [31:0] dmem54_io_bus_response_bits_data; // @[top.scala 393:22]
  wire  cpu55_clock; // @[top.scala 397:21]
  wire  cpu55_reset; // @[top.scala 397:21]
  wire [31:0] cpu55_io_imem_address; // @[top.scala 397:21]
  wire [31:0] cpu55_io_imem_instruction; // @[top.scala 397:21]
  wire [31:0] cpu55_io_dmem_address; // @[top.scala 397:21]
  wire  cpu55_io_dmem_valid; // @[top.scala 397:21]
  wire [31:0] cpu55_io_dmem_writedata; // @[top.scala 397:21]
  wire  cpu55_io_dmem_memread; // @[top.scala 397:21]
  wire  cpu55_io_dmem_memwrite; // @[top.scala 397:21]
  wire [1:0] cpu55_io_dmem_maskmode; // @[top.scala 397:21]
  wire  cpu55_io_dmem_sext; // @[top.scala 397:21]
  wire [31:0] cpu55_io_dmem_readdata; // @[top.scala 397:21]
  wire  mem55_clock; // @[top.scala 398:21]
  wire  mem55_reset; // @[top.scala 398:21]
  wire [31:0] mem55_io_imem_request_bits_address; // @[top.scala 398:21]
  wire [31:0] mem55_io_imem_response_bits_data; // @[top.scala 398:21]
  wire  mem55_io_dmem_request_valid; // @[top.scala 398:21]
  wire [31:0] mem55_io_dmem_request_bits_address; // @[top.scala 398:21]
  wire [31:0] mem55_io_dmem_request_bits_writedata; // @[top.scala 398:21]
  wire [1:0] mem55_io_dmem_request_bits_operation; // @[top.scala 398:21]
  wire  mem55_io_dmem_response_valid; // @[top.scala 398:21]
  wire [31:0] mem55_io_dmem_response_bits_data; // @[top.scala 398:21]
  wire [31:0] imem55_io_pipeline_address; // @[top.scala 399:22]
  wire [31:0] imem55_io_pipeline_instruction; // @[top.scala 399:22]
  wire [31:0] imem55_io_bus_request_bits_address; // @[top.scala 399:22]
  wire [31:0] imem55_io_bus_response_bits_data; // @[top.scala 399:22]
  wire  dmem55_clock; // @[top.scala 400:22]
  wire  dmem55_reset; // @[top.scala 400:22]
  wire [31:0] dmem55_io_pipeline_address; // @[top.scala 400:22]
  wire  dmem55_io_pipeline_valid; // @[top.scala 400:22]
  wire [31:0] dmem55_io_pipeline_writedata; // @[top.scala 400:22]
  wire  dmem55_io_pipeline_memread; // @[top.scala 400:22]
  wire  dmem55_io_pipeline_memwrite; // @[top.scala 400:22]
  wire [1:0] dmem55_io_pipeline_maskmode; // @[top.scala 400:22]
  wire  dmem55_io_pipeline_sext; // @[top.scala 400:22]
  wire [31:0] dmem55_io_pipeline_readdata; // @[top.scala 400:22]
  wire  dmem55_io_bus_request_valid; // @[top.scala 400:22]
  wire [31:0] dmem55_io_bus_request_bits_address; // @[top.scala 400:22]
  wire [31:0] dmem55_io_bus_request_bits_writedata; // @[top.scala 400:22]
  wire [1:0] dmem55_io_bus_request_bits_operation; // @[top.scala 400:22]
  wire  dmem55_io_bus_response_valid; // @[top.scala 400:22]
  wire [31:0] dmem55_io_bus_response_bits_data; // @[top.scala 400:22]
  wire  cpu56_clock; // @[top.scala 404:21]
  wire  cpu56_reset; // @[top.scala 404:21]
  wire [31:0] cpu56_io_imem_address; // @[top.scala 404:21]
  wire [31:0] cpu56_io_imem_instruction; // @[top.scala 404:21]
  wire [31:0] cpu56_io_dmem_address; // @[top.scala 404:21]
  wire  cpu56_io_dmem_valid; // @[top.scala 404:21]
  wire [31:0] cpu56_io_dmem_writedata; // @[top.scala 404:21]
  wire  cpu56_io_dmem_memread; // @[top.scala 404:21]
  wire  cpu56_io_dmem_memwrite; // @[top.scala 404:21]
  wire [1:0] cpu56_io_dmem_maskmode; // @[top.scala 404:21]
  wire  cpu56_io_dmem_sext; // @[top.scala 404:21]
  wire [31:0] cpu56_io_dmem_readdata; // @[top.scala 404:21]
  wire  mem56_clock; // @[top.scala 405:21]
  wire  mem56_reset; // @[top.scala 405:21]
  wire [31:0] mem56_io_imem_request_bits_address; // @[top.scala 405:21]
  wire [31:0] mem56_io_imem_response_bits_data; // @[top.scala 405:21]
  wire  mem56_io_dmem_request_valid; // @[top.scala 405:21]
  wire [31:0] mem56_io_dmem_request_bits_address; // @[top.scala 405:21]
  wire [31:0] mem56_io_dmem_request_bits_writedata; // @[top.scala 405:21]
  wire [1:0] mem56_io_dmem_request_bits_operation; // @[top.scala 405:21]
  wire  mem56_io_dmem_response_valid; // @[top.scala 405:21]
  wire [31:0] mem56_io_dmem_response_bits_data; // @[top.scala 405:21]
  wire [31:0] imem56_io_pipeline_address; // @[top.scala 406:22]
  wire [31:0] imem56_io_pipeline_instruction; // @[top.scala 406:22]
  wire [31:0] imem56_io_bus_request_bits_address; // @[top.scala 406:22]
  wire [31:0] imem56_io_bus_response_bits_data; // @[top.scala 406:22]
  wire  dmem56_clock; // @[top.scala 407:22]
  wire  dmem56_reset; // @[top.scala 407:22]
  wire [31:0] dmem56_io_pipeline_address; // @[top.scala 407:22]
  wire  dmem56_io_pipeline_valid; // @[top.scala 407:22]
  wire [31:0] dmem56_io_pipeline_writedata; // @[top.scala 407:22]
  wire  dmem56_io_pipeline_memread; // @[top.scala 407:22]
  wire  dmem56_io_pipeline_memwrite; // @[top.scala 407:22]
  wire [1:0] dmem56_io_pipeline_maskmode; // @[top.scala 407:22]
  wire  dmem56_io_pipeline_sext; // @[top.scala 407:22]
  wire [31:0] dmem56_io_pipeline_readdata; // @[top.scala 407:22]
  wire  dmem56_io_bus_request_valid; // @[top.scala 407:22]
  wire [31:0] dmem56_io_bus_request_bits_address; // @[top.scala 407:22]
  wire [31:0] dmem56_io_bus_request_bits_writedata; // @[top.scala 407:22]
  wire [1:0] dmem56_io_bus_request_bits_operation; // @[top.scala 407:22]
  wire  dmem56_io_bus_response_valid; // @[top.scala 407:22]
  wire [31:0] dmem56_io_bus_response_bits_data; // @[top.scala 407:22]
  wire  cpu57_clock; // @[top.scala 411:21]
  wire  cpu57_reset; // @[top.scala 411:21]
  wire [31:0] cpu57_io_imem_address; // @[top.scala 411:21]
  wire [31:0] cpu57_io_imem_instruction; // @[top.scala 411:21]
  wire [31:0] cpu57_io_dmem_address; // @[top.scala 411:21]
  wire  cpu57_io_dmem_valid; // @[top.scala 411:21]
  wire [31:0] cpu57_io_dmem_writedata; // @[top.scala 411:21]
  wire  cpu57_io_dmem_memread; // @[top.scala 411:21]
  wire  cpu57_io_dmem_memwrite; // @[top.scala 411:21]
  wire [1:0] cpu57_io_dmem_maskmode; // @[top.scala 411:21]
  wire  cpu57_io_dmem_sext; // @[top.scala 411:21]
  wire [31:0] cpu57_io_dmem_readdata; // @[top.scala 411:21]
  wire  mem57_clock; // @[top.scala 412:21]
  wire  mem57_reset; // @[top.scala 412:21]
  wire [31:0] mem57_io_imem_request_bits_address; // @[top.scala 412:21]
  wire [31:0] mem57_io_imem_response_bits_data; // @[top.scala 412:21]
  wire  mem57_io_dmem_request_valid; // @[top.scala 412:21]
  wire [31:0] mem57_io_dmem_request_bits_address; // @[top.scala 412:21]
  wire [31:0] mem57_io_dmem_request_bits_writedata; // @[top.scala 412:21]
  wire [1:0] mem57_io_dmem_request_bits_operation; // @[top.scala 412:21]
  wire  mem57_io_dmem_response_valid; // @[top.scala 412:21]
  wire [31:0] mem57_io_dmem_response_bits_data; // @[top.scala 412:21]
  wire [31:0] imem57_io_pipeline_address; // @[top.scala 413:22]
  wire [31:0] imem57_io_pipeline_instruction; // @[top.scala 413:22]
  wire [31:0] imem57_io_bus_request_bits_address; // @[top.scala 413:22]
  wire [31:0] imem57_io_bus_response_bits_data; // @[top.scala 413:22]
  wire  dmem57_clock; // @[top.scala 414:22]
  wire  dmem57_reset; // @[top.scala 414:22]
  wire [31:0] dmem57_io_pipeline_address; // @[top.scala 414:22]
  wire  dmem57_io_pipeline_valid; // @[top.scala 414:22]
  wire [31:0] dmem57_io_pipeline_writedata; // @[top.scala 414:22]
  wire  dmem57_io_pipeline_memread; // @[top.scala 414:22]
  wire  dmem57_io_pipeline_memwrite; // @[top.scala 414:22]
  wire [1:0] dmem57_io_pipeline_maskmode; // @[top.scala 414:22]
  wire  dmem57_io_pipeline_sext; // @[top.scala 414:22]
  wire [31:0] dmem57_io_pipeline_readdata; // @[top.scala 414:22]
  wire  dmem57_io_bus_request_valid; // @[top.scala 414:22]
  wire [31:0] dmem57_io_bus_request_bits_address; // @[top.scala 414:22]
  wire [31:0] dmem57_io_bus_request_bits_writedata; // @[top.scala 414:22]
  wire [1:0] dmem57_io_bus_request_bits_operation; // @[top.scala 414:22]
  wire  dmem57_io_bus_response_valid; // @[top.scala 414:22]
  wire [31:0] dmem57_io_bus_response_bits_data; // @[top.scala 414:22]
  wire  cpu58_clock; // @[top.scala 418:21]
  wire  cpu58_reset; // @[top.scala 418:21]
  wire [31:0] cpu58_io_imem_address; // @[top.scala 418:21]
  wire [31:0] cpu58_io_imem_instruction; // @[top.scala 418:21]
  wire [31:0] cpu58_io_dmem_address; // @[top.scala 418:21]
  wire  cpu58_io_dmem_valid; // @[top.scala 418:21]
  wire [31:0] cpu58_io_dmem_writedata; // @[top.scala 418:21]
  wire  cpu58_io_dmem_memread; // @[top.scala 418:21]
  wire  cpu58_io_dmem_memwrite; // @[top.scala 418:21]
  wire [1:0] cpu58_io_dmem_maskmode; // @[top.scala 418:21]
  wire  cpu58_io_dmem_sext; // @[top.scala 418:21]
  wire [31:0] cpu58_io_dmem_readdata; // @[top.scala 418:21]
  wire  mem58_clock; // @[top.scala 419:21]
  wire  mem58_reset; // @[top.scala 419:21]
  wire [31:0] mem58_io_imem_request_bits_address; // @[top.scala 419:21]
  wire [31:0] mem58_io_imem_response_bits_data; // @[top.scala 419:21]
  wire  mem58_io_dmem_request_valid; // @[top.scala 419:21]
  wire [31:0] mem58_io_dmem_request_bits_address; // @[top.scala 419:21]
  wire [31:0] mem58_io_dmem_request_bits_writedata; // @[top.scala 419:21]
  wire [1:0] mem58_io_dmem_request_bits_operation; // @[top.scala 419:21]
  wire  mem58_io_dmem_response_valid; // @[top.scala 419:21]
  wire [31:0] mem58_io_dmem_response_bits_data; // @[top.scala 419:21]
  wire [31:0] imem58_io_pipeline_address; // @[top.scala 420:22]
  wire [31:0] imem58_io_pipeline_instruction; // @[top.scala 420:22]
  wire [31:0] imem58_io_bus_request_bits_address; // @[top.scala 420:22]
  wire [31:0] imem58_io_bus_response_bits_data; // @[top.scala 420:22]
  wire  dmem58_clock; // @[top.scala 421:22]
  wire  dmem58_reset; // @[top.scala 421:22]
  wire [31:0] dmem58_io_pipeline_address; // @[top.scala 421:22]
  wire  dmem58_io_pipeline_valid; // @[top.scala 421:22]
  wire [31:0] dmem58_io_pipeline_writedata; // @[top.scala 421:22]
  wire  dmem58_io_pipeline_memread; // @[top.scala 421:22]
  wire  dmem58_io_pipeline_memwrite; // @[top.scala 421:22]
  wire [1:0] dmem58_io_pipeline_maskmode; // @[top.scala 421:22]
  wire  dmem58_io_pipeline_sext; // @[top.scala 421:22]
  wire [31:0] dmem58_io_pipeline_readdata; // @[top.scala 421:22]
  wire  dmem58_io_bus_request_valid; // @[top.scala 421:22]
  wire [31:0] dmem58_io_bus_request_bits_address; // @[top.scala 421:22]
  wire [31:0] dmem58_io_bus_request_bits_writedata; // @[top.scala 421:22]
  wire [1:0] dmem58_io_bus_request_bits_operation; // @[top.scala 421:22]
  wire  dmem58_io_bus_response_valid; // @[top.scala 421:22]
  wire [31:0] dmem58_io_bus_response_bits_data; // @[top.scala 421:22]
  wire  cpu59_clock; // @[top.scala 425:21]
  wire  cpu59_reset; // @[top.scala 425:21]
  wire [31:0] cpu59_io_imem_address; // @[top.scala 425:21]
  wire [31:0] cpu59_io_imem_instruction; // @[top.scala 425:21]
  wire [31:0] cpu59_io_dmem_address; // @[top.scala 425:21]
  wire  cpu59_io_dmem_valid; // @[top.scala 425:21]
  wire [31:0] cpu59_io_dmem_writedata; // @[top.scala 425:21]
  wire  cpu59_io_dmem_memread; // @[top.scala 425:21]
  wire  cpu59_io_dmem_memwrite; // @[top.scala 425:21]
  wire [1:0] cpu59_io_dmem_maskmode; // @[top.scala 425:21]
  wire  cpu59_io_dmem_sext; // @[top.scala 425:21]
  wire [31:0] cpu59_io_dmem_readdata; // @[top.scala 425:21]
  wire  mem59_clock; // @[top.scala 426:21]
  wire  mem59_reset; // @[top.scala 426:21]
  wire [31:0] mem59_io_imem_request_bits_address; // @[top.scala 426:21]
  wire [31:0] mem59_io_imem_response_bits_data; // @[top.scala 426:21]
  wire  mem59_io_dmem_request_valid; // @[top.scala 426:21]
  wire [31:0] mem59_io_dmem_request_bits_address; // @[top.scala 426:21]
  wire [31:0] mem59_io_dmem_request_bits_writedata; // @[top.scala 426:21]
  wire [1:0] mem59_io_dmem_request_bits_operation; // @[top.scala 426:21]
  wire  mem59_io_dmem_response_valid; // @[top.scala 426:21]
  wire [31:0] mem59_io_dmem_response_bits_data; // @[top.scala 426:21]
  wire [31:0] imem59_io_pipeline_address; // @[top.scala 427:22]
  wire [31:0] imem59_io_pipeline_instruction; // @[top.scala 427:22]
  wire [31:0] imem59_io_bus_request_bits_address; // @[top.scala 427:22]
  wire [31:0] imem59_io_bus_response_bits_data; // @[top.scala 427:22]
  wire  dmem59_clock; // @[top.scala 428:22]
  wire  dmem59_reset; // @[top.scala 428:22]
  wire [31:0] dmem59_io_pipeline_address; // @[top.scala 428:22]
  wire  dmem59_io_pipeline_valid; // @[top.scala 428:22]
  wire [31:0] dmem59_io_pipeline_writedata; // @[top.scala 428:22]
  wire  dmem59_io_pipeline_memread; // @[top.scala 428:22]
  wire  dmem59_io_pipeline_memwrite; // @[top.scala 428:22]
  wire [1:0] dmem59_io_pipeline_maskmode; // @[top.scala 428:22]
  wire  dmem59_io_pipeline_sext; // @[top.scala 428:22]
  wire [31:0] dmem59_io_pipeline_readdata; // @[top.scala 428:22]
  wire  dmem59_io_bus_request_valid; // @[top.scala 428:22]
  wire [31:0] dmem59_io_bus_request_bits_address; // @[top.scala 428:22]
  wire [31:0] dmem59_io_bus_request_bits_writedata; // @[top.scala 428:22]
  wire [1:0] dmem59_io_bus_request_bits_operation; // @[top.scala 428:22]
  wire  dmem59_io_bus_response_valid; // @[top.scala 428:22]
  wire [31:0] dmem59_io_bus_response_bits_data; // @[top.scala 428:22]
  wire  cpu60_clock; // @[top.scala 432:21]
  wire  cpu60_reset; // @[top.scala 432:21]
  wire [31:0] cpu60_io_imem_address; // @[top.scala 432:21]
  wire [31:0] cpu60_io_imem_instruction; // @[top.scala 432:21]
  wire [31:0] cpu60_io_dmem_address; // @[top.scala 432:21]
  wire  cpu60_io_dmem_valid; // @[top.scala 432:21]
  wire [31:0] cpu60_io_dmem_writedata; // @[top.scala 432:21]
  wire  cpu60_io_dmem_memread; // @[top.scala 432:21]
  wire  cpu60_io_dmem_memwrite; // @[top.scala 432:21]
  wire [1:0] cpu60_io_dmem_maskmode; // @[top.scala 432:21]
  wire  cpu60_io_dmem_sext; // @[top.scala 432:21]
  wire [31:0] cpu60_io_dmem_readdata; // @[top.scala 432:21]
  wire  mem60_clock; // @[top.scala 433:21]
  wire  mem60_reset; // @[top.scala 433:21]
  wire [31:0] mem60_io_imem_request_bits_address; // @[top.scala 433:21]
  wire [31:0] mem60_io_imem_response_bits_data; // @[top.scala 433:21]
  wire  mem60_io_dmem_request_valid; // @[top.scala 433:21]
  wire [31:0] mem60_io_dmem_request_bits_address; // @[top.scala 433:21]
  wire [31:0] mem60_io_dmem_request_bits_writedata; // @[top.scala 433:21]
  wire [1:0] mem60_io_dmem_request_bits_operation; // @[top.scala 433:21]
  wire  mem60_io_dmem_response_valid; // @[top.scala 433:21]
  wire [31:0] mem60_io_dmem_response_bits_data; // @[top.scala 433:21]
  wire [31:0] imem60_io_pipeline_address; // @[top.scala 434:22]
  wire [31:0] imem60_io_pipeline_instruction; // @[top.scala 434:22]
  wire [31:0] imem60_io_bus_request_bits_address; // @[top.scala 434:22]
  wire [31:0] imem60_io_bus_response_bits_data; // @[top.scala 434:22]
  wire  dmem60_clock; // @[top.scala 435:22]
  wire  dmem60_reset; // @[top.scala 435:22]
  wire [31:0] dmem60_io_pipeline_address; // @[top.scala 435:22]
  wire  dmem60_io_pipeline_valid; // @[top.scala 435:22]
  wire [31:0] dmem60_io_pipeline_writedata; // @[top.scala 435:22]
  wire  dmem60_io_pipeline_memread; // @[top.scala 435:22]
  wire  dmem60_io_pipeline_memwrite; // @[top.scala 435:22]
  wire [1:0] dmem60_io_pipeline_maskmode; // @[top.scala 435:22]
  wire  dmem60_io_pipeline_sext; // @[top.scala 435:22]
  wire [31:0] dmem60_io_pipeline_readdata; // @[top.scala 435:22]
  wire  dmem60_io_bus_request_valid; // @[top.scala 435:22]
  wire [31:0] dmem60_io_bus_request_bits_address; // @[top.scala 435:22]
  wire [31:0] dmem60_io_bus_request_bits_writedata; // @[top.scala 435:22]
  wire [1:0] dmem60_io_bus_request_bits_operation; // @[top.scala 435:22]
  wire  dmem60_io_bus_response_valid; // @[top.scala 435:22]
  wire [31:0] dmem60_io_bus_response_bits_data; // @[top.scala 435:22]
  wire  cpu61_clock; // @[top.scala 439:21]
  wire  cpu61_reset; // @[top.scala 439:21]
  wire [31:0] cpu61_io_imem_address; // @[top.scala 439:21]
  wire [31:0] cpu61_io_imem_instruction; // @[top.scala 439:21]
  wire [31:0] cpu61_io_dmem_address; // @[top.scala 439:21]
  wire  cpu61_io_dmem_valid; // @[top.scala 439:21]
  wire [31:0] cpu61_io_dmem_writedata; // @[top.scala 439:21]
  wire  cpu61_io_dmem_memread; // @[top.scala 439:21]
  wire  cpu61_io_dmem_memwrite; // @[top.scala 439:21]
  wire [1:0] cpu61_io_dmem_maskmode; // @[top.scala 439:21]
  wire  cpu61_io_dmem_sext; // @[top.scala 439:21]
  wire [31:0] cpu61_io_dmem_readdata; // @[top.scala 439:21]
  wire  mem61_clock; // @[top.scala 440:21]
  wire  mem61_reset; // @[top.scala 440:21]
  wire [31:0] mem61_io_imem_request_bits_address; // @[top.scala 440:21]
  wire [31:0] mem61_io_imem_response_bits_data; // @[top.scala 440:21]
  wire  mem61_io_dmem_request_valid; // @[top.scala 440:21]
  wire [31:0] mem61_io_dmem_request_bits_address; // @[top.scala 440:21]
  wire [31:0] mem61_io_dmem_request_bits_writedata; // @[top.scala 440:21]
  wire [1:0] mem61_io_dmem_request_bits_operation; // @[top.scala 440:21]
  wire  mem61_io_dmem_response_valid; // @[top.scala 440:21]
  wire [31:0] mem61_io_dmem_response_bits_data; // @[top.scala 440:21]
  wire [31:0] imem61_io_pipeline_address; // @[top.scala 441:22]
  wire [31:0] imem61_io_pipeline_instruction; // @[top.scala 441:22]
  wire [31:0] imem61_io_bus_request_bits_address; // @[top.scala 441:22]
  wire [31:0] imem61_io_bus_response_bits_data; // @[top.scala 441:22]
  wire  dmem61_clock; // @[top.scala 442:22]
  wire  dmem61_reset; // @[top.scala 442:22]
  wire [31:0] dmem61_io_pipeline_address; // @[top.scala 442:22]
  wire  dmem61_io_pipeline_valid; // @[top.scala 442:22]
  wire [31:0] dmem61_io_pipeline_writedata; // @[top.scala 442:22]
  wire  dmem61_io_pipeline_memread; // @[top.scala 442:22]
  wire  dmem61_io_pipeline_memwrite; // @[top.scala 442:22]
  wire [1:0] dmem61_io_pipeline_maskmode; // @[top.scala 442:22]
  wire  dmem61_io_pipeline_sext; // @[top.scala 442:22]
  wire [31:0] dmem61_io_pipeline_readdata; // @[top.scala 442:22]
  wire  dmem61_io_bus_request_valid; // @[top.scala 442:22]
  wire [31:0] dmem61_io_bus_request_bits_address; // @[top.scala 442:22]
  wire [31:0] dmem61_io_bus_request_bits_writedata; // @[top.scala 442:22]
  wire [1:0] dmem61_io_bus_request_bits_operation; // @[top.scala 442:22]
  wire  dmem61_io_bus_response_valid; // @[top.scala 442:22]
  wire [31:0] dmem61_io_bus_response_bits_data; // @[top.scala 442:22]
  wire  cpu62_clock; // @[top.scala 446:21]
  wire  cpu62_reset; // @[top.scala 446:21]
  wire [31:0] cpu62_io_imem_address; // @[top.scala 446:21]
  wire [31:0] cpu62_io_imem_instruction; // @[top.scala 446:21]
  wire [31:0] cpu62_io_dmem_address; // @[top.scala 446:21]
  wire  cpu62_io_dmem_valid; // @[top.scala 446:21]
  wire [31:0] cpu62_io_dmem_writedata; // @[top.scala 446:21]
  wire  cpu62_io_dmem_memread; // @[top.scala 446:21]
  wire  cpu62_io_dmem_memwrite; // @[top.scala 446:21]
  wire [1:0] cpu62_io_dmem_maskmode; // @[top.scala 446:21]
  wire  cpu62_io_dmem_sext; // @[top.scala 446:21]
  wire [31:0] cpu62_io_dmem_readdata; // @[top.scala 446:21]
  wire  mem62_clock; // @[top.scala 447:21]
  wire  mem62_reset; // @[top.scala 447:21]
  wire [31:0] mem62_io_imem_request_bits_address; // @[top.scala 447:21]
  wire [31:0] mem62_io_imem_response_bits_data; // @[top.scala 447:21]
  wire  mem62_io_dmem_request_valid; // @[top.scala 447:21]
  wire [31:0] mem62_io_dmem_request_bits_address; // @[top.scala 447:21]
  wire [31:0] mem62_io_dmem_request_bits_writedata; // @[top.scala 447:21]
  wire [1:0] mem62_io_dmem_request_bits_operation; // @[top.scala 447:21]
  wire  mem62_io_dmem_response_valid; // @[top.scala 447:21]
  wire [31:0] mem62_io_dmem_response_bits_data; // @[top.scala 447:21]
  wire [31:0] imem62_io_pipeline_address; // @[top.scala 448:22]
  wire [31:0] imem62_io_pipeline_instruction; // @[top.scala 448:22]
  wire [31:0] imem62_io_bus_request_bits_address; // @[top.scala 448:22]
  wire [31:0] imem62_io_bus_response_bits_data; // @[top.scala 448:22]
  wire  dmem62_clock; // @[top.scala 449:22]
  wire  dmem62_reset; // @[top.scala 449:22]
  wire [31:0] dmem62_io_pipeline_address; // @[top.scala 449:22]
  wire  dmem62_io_pipeline_valid; // @[top.scala 449:22]
  wire [31:0] dmem62_io_pipeline_writedata; // @[top.scala 449:22]
  wire  dmem62_io_pipeline_memread; // @[top.scala 449:22]
  wire  dmem62_io_pipeline_memwrite; // @[top.scala 449:22]
  wire [1:0] dmem62_io_pipeline_maskmode; // @[top.scala 449:22]
  wire  dmem62_io_pipeline_sext; // @[top.scala 449:22]
  wire [31:0] dmem62_io_pipeline_readdata; // @[top.scala 449:22]
  wire  dmem62_io_bus_request_valid; // @[top.scala 449:22]
  wire [31:0] dmem62_io_bus_request_bits_address; // @[top.scala 449:22]
  wire [31:0] dmem62_io_bus_request_bits_writedata; // @[top.scala 449:22]
  wire [1:0] dmem62_io_bus_request_bits_operation; // @[top.scala 449:22]
  wire  dmem62_io_bus_response_valid; // @[top.scala 449:22]
  wire [31:0] dmem62_io_bus_response_bits_data; // @[top.scala 449:22]
  wire  cpu63_clock; // @[top.scala 453:21]
  wire  cpu63_reset; // @[top.scala 453:21]
  wire [31:0] cpu63_io_imem_address; // @[top.scala 453:21]
  wire [31:0] cpu63_io_imem_instruction; // @[top.scala 453:21]
  wire [31:0] cpu63_io_dmem_address; // @[top.scala 453:21]
  wire  cpu63_io_dmem_valid; // @[top.scala 453:21]
  wire [31:0] cpu63_io_dmem_writedata; // @[top.scala 453:21]
  wire  cpu63_io_dmem_memread; // @[top.scala 453:21]
  wire  cpu63_io_dmem_memwrite; // @[top.scala 453:21]
  wire [1:0] cpu63_io_dmem_maskmode; // @[top.scala 453:21]
  wire  cpu63_io_dmem_sext; // @[top.scala 453:21]
  wire [31:0] cpu63_io_dmem_readdata; // @[top.scala 453:21]
  wire  mem63_clock; // @[top.scala 454:21]
  wire  mem63_reset; // @[top.scala 454:21]
  wire [31:0] mem63_io_imem_request_bits_address; // @[top.scala 454:21]
  wire [31:0] mem63_io_imem_response_bits_data; // @[top.scala 454:21]
  wire  mem63_io_dmem_request_valid; // @[top.scala 454:21]
  wire [31:0] mem63_io_dmem_request_bits_address; // @[top.scala 454:21]
  wire [31:0] mem63_io_dmem_request_bits_writedata; // @[top.scala 454:21]
  wire [1:0] mem63_io_dmem_request_bits_operation; // @[top.scala 454:21]
  wire  mem63_io_dmem_response_valid; // @[top.scala 454:21]
  wire [31:0] mem63_io_dmem_response_bits_data; // @[top.scala 454:21]
  wire [31:0] imem63_io_pipeline_address; // @[top.scala 455:22]
  wire [31:0] imem63_io_pipeline_instruction; // @[top.scala 455:22]
  wire [31:0] imem63_io_bus_request_bits_address; // @[top.scala 455:22]
  wire [31:0] imem63_io_bus_response_bits_data; // @[top.scala 455:22]
  wire  dmem63_clock; // @[top.scala 456:22]
  wire  dmem63_reset; // @[top.scala 456:22]
  wire [31:0] dmem63_io_pipeline_address; // @[top.scala 456:22]
  wire  dmem63_io_pipeline_valid; // @[top.scala 456:22]
  wire [31:0] dmem63_io_pipeline_writedata; // @[top.scala 456:22]
  wire  dmem63_io_pipeline_memread; // @[top.scala 456:22]
  wire  dmem63_io_pipeline_memwrite; // @[top.scala 456:22]
  wire [1:0] dmem63_io_pipeline_maskmode; // @[top.scala 456:22]
  wire  dmem63_io_pipeline_sext; // @[top.scala 456:22]
  wire [31:0] dmem63_io_pipeline_readdata; // @[top.scala 456:22]
  wire  dmem63_io_bus_request_valid; // @[top.scala 456:22]
  wire [31:0] dmem63_io_bus_request_bits_address; // @[top.scala 456:22]
  wire [31:0] dmem63_io_bus_request_bits_writedata; // @[top.scala 456:22]
  wire [1:0] dmem63_io_bus_request_bits_operation; // @[top.scala 456:22]
  wire  dmem63_io_bus_response_valid; // @[top.scala 456:22]
  wire [31:0] dmem63_io_bus_response_bits_data; // @[top.scala 456:22]
  wire  cpu64_clock; // @[top.scala 460:21]
  wire  cpu64_reset; // @[top.scala 460:21]
  wire [31:0] cpu64_io_imem_address; // @[top.scala 460:21]
  wire [31:0] cpu64_io_imem_instruction; // @[top.scala 460:21]
  wire [31:0] cpu64_io_dmem_address; // @[top.scala 460:21]
  wire  cpu64_io_dmem_valid; // @[top.scala 460:21]
  wire [31:0] cpu64_io_dmem_writedata; // @[top.scala 460:21]
  wire  cpu64_io_dmem_memread; // @[top.scala 460:21]
  wire  cpu64_io_dmem_memwrite; // @[top.scala 460:21]
  wire [1:0] cpu64_io_dmem_maskmode; // @[top.scala 460:21]
  wire  cpu64_io_dmem_sext; // @[top.scala 460:21]
  wire [31:0] cpu64_io_dmem_readdata; // @[top.scala 460:21]
  wire  mem64_clock; // @[top.scala 461:21]
  wire  mem64_reset; // @[top.scala 461:21]
  wire [31:0] mem64_io_imem_request_bits_address; // @[top.scala 461:21]
  wire [31:0] mem64_io_imem_response_bits_data; // @[top.scala 461:21]
  wire  mem64_io_dmem_request_valid; // @[top.scala 461:21]
  wire [31:0] mem64_io_dmem_request_bits_address; // @[top.scala 461:21]
  wire [31:0] mem64_io_dmem_request_bits_writedata; // @[top.scala 461:21]
  wire [1:0] mem64_io_dmem_request_bits_operation; // @[top.scala 461:21]
  wire  mem64_io_dmem_response_valid; // @[top.scala 461:21]
  wire [31:0] mem64_io_dmem_response_bits_data; // @[top.scala 461:21]
  wire [31:0] imem64_io_pipeline_address; // @[top.scala 462:22]
  wire [31:0] imem64_io_pipeline_instruction; // @[top.scala 462:22]
  wire [31:0] imem64_io_bus_request_bits_address; // @[top.scala 462:22]
  wire [31:0] imem64_io_bus_response_bits_data; // @[top.scala 462:22]
  wire  dmem64_clock; // @[top.scala 463:22]
  wire  dmem64_reset; // @[top.scala 463:22]
  wire [31:0] dmem64_io_pipeline_address; // @[top.scala 463:22]
  wire  dmem64_io_pipeline_valid; // @[top.scala 463:22]
  wire [31:0] dmem64_io_pipeline_writedata; // @[top.scala 463:22]
  wire  dmem64_io_pipeline_memread; // @[top.scala 463:22]
  wire  dmem64_io_pipeline_memwrite; // @[top.scala 463:22]
  wire [1:0] dmem64_io_pipeline_maskmode; // @[top.scala 463:22]
  wire  dmem64_io_pipeline_sext; // @[top.scala 463:22]
  wire [31:0] dmem64_io_pipeline_readdata; // @[top.scala 463:22]
  wire  dmem64_io_bus_request_valid; // @[top.scala 463:22]
  wire [31:0] dmem64_io_bus_request_bits_address; // @[top.scala 463:22]
  wire [31:0] dmem64_io_bus_request_bits_writedata; // @[top.scala 463:22]
  wire [1:0] dmem64_io_bus_request_bits_operation; // @[top.scala 463:22]
  wire  dmem64_io_bus_response_valid; // @[top.scala 463:22]
  wire [31:0] dmem64_io_bus_response_bits_data; // @[top.scala 463:22]
  wire  cpu65_clock; // @[top.scala 467:21]
  wire  cpu65_reset; // @[top.scala 467:21]
  wire [31:0] cpu65_io_imem_address; // @[top.scala 467:21]
  wire [31:0] cpu65_io_imem_instruction; // @[top.scala 467:21]
  wire [31:0] cpu65_io_dmem_address; // @[top.scala 467:21]
  wire  cpu65_io_dmem_valid; // @[top.scala 467:21]
  wire [31:0] cpu65_io_dmem_writedata; // @[top.scala 467:21]
  wire  cpu65_io_dmem_memread; // @[top.scala 467:21]
  wire  cpu65_io_dmem_memwrite; // @[top.scala 467:21]
  wire [1:0] cpu65_io_dmem_maskmode; // @[top.scala 467:21]
  wire  cpu65_io_dmem_sext; // @[top.scala 467:21]
  wire [31:0] cpu65_io_dmem_readdata; // @[top.scala 467:21]
  wire  mem65_clock; // @[top.scala 468:21]
  wire  mem65_reset; // @[top.scala 468:21]
  wire [31:0] mem65_io_imem_request_bits_address; // @[top.scala 468:21]
  wire [31:0] mem65_io_imem_response_bits_data; // @[top.scala 468:21]
  wire  mem65_io_dmem_request_valid; // @[top.scala 468:21]
  wire [31:0] mem65_io_dmem_request_bits_address; // @[top.scala 468:21]
  wire [31:0] mem65_io_dmem_request_bits_writedata; // @[top.scala 468:21]
  wire [1:0] mem65_io_dmem_request_bits_operation; // @[top.scala 468:21]
  wire  mem65_io_dmem_response_valid; // @[top.scala 468:21]
  wire [31:0] mem65_io_dmem_response_bits_data; // @[top.scala 468:21]
  wire [31:0] imem65_io_pipeline_address; // @[top.scala 469:22]
  wire [31:0] imem65_io_pipeline_instruction; // @[top.scala 469:22]
  wire [31:0] imem65_io_bus_request_bits_address; // @[top.scala 469:22]
  wire [31:0] imem65_io_bus_response_bits_data; // @[top.scala 469:22]
  wire  dmem65_clock; // @[top.scala 470:22]
  wire  dmem65_reset; // @[top.scala 470:22]
  wire [31:0] dmem65_io_pipeline_address; // @[top.scala 470:22]
  wire  dmem65_io_pipeline_valid; // @[top.scala 470:22]
  wire [31:0] dmem65_io_pipeline_writedata; // @[top.scala 470:22]
  wire  dmem65_io_pipeline_memread; // @[top.scala 470:22]
  wire  dmem65_io_pipeline_memwrite; // @[top.scala 470:22]
  wire [1:0] dmem65_io_pipeline_maskmode; // @[top.scala 470:22]
  wire  dmem65_io_pipeline_sext; // @[top.scala 470:22]
  wire [31:0] dmem65_io_pipeline_readdata; // @[top.scala 470:22]
  wire  dmem65_io_bus_request_valid; // @[top.scala 470:22]
  wire [31:0] dmem65_io_bus_request_bits_address; // @[top.scala 470:22]
  wire [31:0] dmem65_io_bus_request_bits_writedata; // @[top.scala 470:22]
  wire [1:0] dmem65_io_bus_request_bits_operation; // @[top.scala 470:22]
  wire  dmem65_io_bus_response_valid; // @[top.scala 470:22]
  wire [31:0] dmem65_io_bus_response_bits_data; // @[top.scala 470:22]
  wire  cpu66_clock; // @[top.scala 474:21]
  wire  cpu66_reset; // @[top.scala 474:21]
  wire [31:0] cpu66_io_imem_address; // @[top.scala 474:21]
  wire [31:0] cpu66_io_imem_instruction; // @[top.scala 474:21]
  wire [31:0] cpu66_io_dmem_address; // @[top.scala 474:21]
  wire  cpu66_io_dmem_valid; // @[top.scala 474:21]
  wire [31:0] cpu66_io_dmem_writedata; // @[top.scala 474:21]
  wire  cpu66_io_dmem_memread; // @[top.scala 474:21]
  wire  cpu66_io_dmem_memwrite; // @[top.scala 474:21]
  wire [1:0] cpu66_io_dmem_maskmode; // @[top.scala 474:21]
  wire  cpu66_io_dmem_sext; // @[top.scala 474:21]
  wire [31:0] cpu66_io_dmem_readdata; // @[top.scala 474:21]
  wire  mem66_clock; // @[top.scala 475:21]
  wire  mem66_reset; // @[top.scala 475:21]
  wire [31:0] mem66_io_imem_request_bits_address; // @[top.scala 475:21]
  wire [31:0] mem66_io_imem_response_bits_data; // @[top.scala 475:21]
  wire  mem66_io_dmem_request_valid; // @[top.scala 475:21]
  wire [31:0] mem66_io_dmem_request_bits_address; // @[top.scala 475:21]
  wire [31:0] mem66_io_dmem_request_bits_writedata; // @[top.scala 475:21]
  wire [1:0] mem66_io_dmem_request_bits_operation; // @[top.scala 475:21]
  wire  mem66_io_dmem_response_valid; // @[top.scala 475:21]
  wire [31:0] mem66_io_dmem_response_bits_data; // @[top.scala 475:21]
  wire [31:0] imem66_io_pipeline_address; // @[top.scala 476:22]
  wire [31:0] imem66_io_pipeline_instruction; // @[top.scala 476:22]
  wire [31:0] imem66_io_bus_request_bits_address; // @[top.scala 476:22]
  wire [31:0] imem66_io_bus_response_bits_data; // @[top.scala 476:22]
  wire  dmem66_clock; // @[top.scala 477:22]
  wire  dmem66_reset; // @[top.scala 477:22]
  wire [31:0] dmem66_io_pipeline_address; // @[top.scala 477:22]
  wire  dmem66_io_pipeline_valid; // @[top.scala 477:22]
  wire [31:0] dmem66_io_pipeline_writedata; // @[top.scala 477:22]
  wire  dmem66_io_pipeline_memread; // @[top.scala 477:22]
  wire  dmem66_io_pipeline_memwrite; // @[top.scala 477:22]
  wire [1:0] dmem66_io_pipeline_maskmode; // @[top.scala 477:22]
  wire  dmem66_io_pipeline_sext; // @[top.scala 477:22]
  wire [31:0] dmem66_io_pipeline_readdata; // @[top.scala 477:22]
  wire  dmem66_io_bus_request_valid; // @[top.scala 477:22]
  wire [31:0] dmem66_io_bus_request_bits_address; // @[top.scala 477:22]
  wire [31:0] dmem66_io_bus_request_bits_writedata; // @[top.scala 477:22]
  wire [1:0] dmem66_io_bus_request_bits_operation; // @[top.scala 477:22]
  wire  dmem66_io_bus_response_valid; // @[top.scala 477:22]
  wire [31:0] dmem66_io_bus_response_bits_data; // @[top.scala 477:22]
  wire  cpu67_clock; // @[top.scala 481:21]
  wire  cpu67_reset; // @[top.scala 481:21]
  wire [31:0] cpu67_io_imem_address; // @[top.scala 481:21]
  wire [31:0] cpu67_io_imem_instruction; // @[top.scala 481:21]
  wire [31:0] cpu67_io_dmem_address; // @[top.scala 481:21]
  wire  cpu67_io_dmem_valid; // @[top.scala 481:21]
  wire [31:0] cpu67_io_dmem_writedata; // @[top.scala 481:21]
  wire  cpu67_io_dmem_memread; // @[top.scala 481:21]
  wire  cpu67_io_dmem_memwrite; // @[top.scala 481:21]
  wire [1:0] cpu67_io_dmem_maskmode; // @[top.scala 481:21]
  wire  cpu67_io_dmem_sext; // @[top.scala 481:21]
  wire [31:0] cpu67_io_dmem_readdata; // @[top.scala 481:21]
  wire  mem67_clock; // @[top.scala 482:21]
  wire  mem67_reset; // @[top.scala 482:21]
  wire [31:0] mem67_io_imem_request_bits_address; // @[top.scala 482:21]
  wire [31:0] mem67_io_imem_response_bits_data; // @[top.scala 482:21]
  wire  mem67_io_dmem_request_valid; // @[top.scala 482:21]
  wire [31:0] mem67_io_dmem_request_bits_address; // @[top.scala 482:21]
  wire [31:0] mem67_io_dmem_request_bits_writedata; // @[top.scala 482:21]
  wire [1:0] mem67_io_dmem_request_bits_operation; // @[top.scala 482:21]
  wire  mem67_io_dmem_response_valid; // @[top.scala 482:21]
  wire [31:0] mem67_io_dmem_response_bits_data; // @[top.scala 482:21]
  wire [31:0] imem67_io_pipeline_address; // @[top.scala 483:22]
  wire [31:0] imem67_io_pipeline_instruction; // @[top.scala 483:22]
  wire [31:0] imem67_io_bus_request_bits_address; // @[top.scala 483:22]
  wire [31:0] imem67_io_bus_response_bits_data; // @[top.scala 483:22]
  wire  dmem67_clock; // @[top.scala 484:22]
  wire  dmem67_reset; // @[top.scala 484:22]
  wire [31:0] dmem67_io_pipeline_address; // @[top.scala 484:22]
  wire  dmem67_io_pipeline_valid; // @[top.scala 484:22]
  wire [31:0] dmem67_io_pipeline_writedata; // @[top.scala 484:22]
  wire  dmem67_io_pipeline_memread; // @[top.scala 484:22]
  wire  dmem67_io_pipeline_memwrite; // @[top.scala 484:22]
  wire [1:0] dmem67_io_pipeline_maskmode; // @[top.scala 484:22]
  wire  dmem67_io_pipeline_sext; // @[top.scala 484:22]
  wire [31:0] dmem67_io_pipeline_readdata; // @[top.scala 484:22]
  wire  dmem67_io_bus_request_valid; // @[top.scala 484:22]
  wire [31:0] dmem67_io_bus_request_bits_address; // @[top.scala 484:22]
  wire [31:0] dmem67_io_bus_request_bits_writedata; // @[top.scala 484:22]
  wire [1:0] dmem67_io_bus_request_bits_operation; // @[top.scala 484:22]
  wire  dmem67_io_bus_response_valid; // @[top.scala 484:22]
  wire [31:0] dmem67_io_bus_response_bits_data; // @[top.scala 484:22]
  wire  cpu68_clock; // @[top.scala 488:21]
  wire  cpu68_reset; // @[top.scala 488:21]
  wire [31:0] cpu68_io_imem_address; // @[top.scala 488:21]
  wire [31:0] cpu68_io_imem_instruction; // @[top.scala 488:21]
  wire [31:0] cpu68_io_dmem_address; // @[top.scala 488:21]
  wire  cpu68_io_dmem_valid; // @[top.scala 488:21]
  wire [31:0] cpu68_io_dmem_writedata; // @[top.scala 488:21]
  wire  cpu68_io_dmem_memread; // @[top.scala 488:21]
  wire  cpu68_io_dmem_memwrite; // @[top.scala 488:21]
  wire [1:0] cpu68_io_dmem_maskmode; // @[top.scala 488:21]
  wire  cpu68_io_dmem_sext; // @[top.scala 488:21]
  wire [31:0] cpu68_io_dmem_readdata; // @[top.scala 488:21]
  wire  mem68_clock; // @[top.scala 489:21]
  wire  mem68_reset; // @[top.scala 489:21]
  wire [31:0] mem68_io_imem_request_bits_address; // @[top.scala 489:21]
  wire [31:0] mem68_io_imem_response_bits_data; // @[top.scala 489:21]
  wire  mem68_io_dmem_request_valid; // @[top.scala 489:21]
  wire [31:0] mem68_io_dmem_request_bits_address; // @[top.scala 489:21]
  wire [31:0] mem68_io_dmem_request_bits_writedata; // @[top.scala 489:21]
  wire [1:0] mem68_io_dmem_request_bits_operation; // @[top.scala 489:21]
  wire  mem68_io_dmem_response_valid; // @[top.scala 489:21]
  wire [31:0] mem68_io_dmem_response_bits_data; // @[top.scala 489:21]
  wire [31:0] imem68_io_pipeline_address; // @[top.scala 490:22]
  wire [31:0] imem68_io_pipeline_instruction; // @[top.scala 490:22]
  wire [31:0] imem68_io_bus_request_bits_address; // @[top.scala 490:22]
  wire [31:0] imem68_io_bus_response_bits_data; // @[top.scala 490:22]
  wire  dmem68_clock; // @[top.scala 491:22]
  wire  dmem68_reset; // @[top.scala 491:22]
  wire [31:0] dmem68_io_pipeline_address; // @[top.scala 491:22]
  wire  dmem68_io_pipeline_valid; // @[top.scala 491:22]
  wire [31:0] dmem68_io_pipeline_writedata; // @[top.scala 491:22]
  wire  dmem68_io_pipeline_memread; // @[top.scala 491:22]
  wire  dmem68_io_pipeline_memwrite; // @[top.scala 491:22]
  wire [1:0] dmem68_io_pipeline_maskmode; // @[top.scala 491:22]
  wire  dmem68_io_pipeline_sext; // @[top.scala 491:22]
  wire [31:0] dmem68_io_pipeline_readdata; // @[top.scala 491:22]
  wire  dmem68_io_bus_request_valid; // @[top.scala 491:22]
  wire [31:0] dmem68_io_bus_request_bits_address; // @[top.scala 491:22]
  wire [31:0] dmem68_io_bus_request_bits_writedata; // @[top.scala 491:22]
  wire [1:0] dmem68_io_bus_request_bits_operation; // @[top.scala 491:22]
  wire  dmem68_io_bus_response_valid; // @[top.scala 491:22]
  wire [31:0] dmem68_io_bus_response_bits_data; // @[top.scala 491:22]
  wire  cpu69_clock; // @[top.scala 495:21]
  wire  cpu69_reset; // @[top.scala 495:21]
  wire [31:0] cpu69_io_imem_address; // @[top.scala 495:21]
  wire [31:0] cpu69_io_imem_instruction; // @[top.scala 495:21]
  wire [31:0] cpu69_io_dmem_address; // @[top.scala 495:21]
  wire  cpu69_io_dmem_valid; // @[top.scala 495:21]
  wire [31:0] cpu69_io_dmem_writedata; // @[top.scala 495:21]
  wire  cpu69_io_dmem_memread; // @[top.scala 495:21]
  wire  cpu69_io_dmem_memwrite; // @[top.scala 495:21]
  wire [1:0] cpu69_io_dmem_maskmode; // @[top.scala 495:21]
  wire  cpu69_io_dmem_sext; // @[top.scala 495:21]
  wire [31:0] cpu69_io_dmem_readdata; // @[top.scala 495:21]
  wire  mem69_clock; // @[top.scala 496:21]
  wire  mem69_reset; // @[top.scala 496:21]
  wire [31:0] mem69_io_imem_request_bits_address; // @[top.scala 496:21]
  wire [31:0] mem69_io_imem_response_bits_data; // @[top.scala 496:21]
  wire  mem69_io_dmem_request_valid; // @[top.scala 496:21]
  wire [31:0] mem69_io_dmem_request_bits_address; // @[top.scala 496:21]
  wire [31:0] mem69_io_dmem_request_bits_writedata; // @[top.scala 496:21]
  wire [1:0] mem69_io_dmem_request_bits_operation; // @[top.scala 496:21]
  wire  mem69_io_dmem_response_valid; // @[top.scala 496:21]
  wire [31:0] mem69_io_dmem_response_bits_data; // @[top.scala 496:21]
  wire [31:0] imem69_io_pipeline_address; // @[top.scala 497:22]
  wire [31:0] imem69_io_pipeline_instruction; // @[top.scala 497:22]
  wire [31:0] imem69_io_bus_request_bits_address; // @[top.scala 497:22]
  wire [31:0] imem69_io_bus_response_bits_data; // @[top.scala 497:22]
  wire  dmem69_clock; // @[top.scala 498:22]
  wire  dmem69_reset; // @[top.scala 498:22]
  wire [31:0] dmem69_io_pipeline_address; // @[top.scala 498:22]
  wire  dmem69_io_pipeline_valid; // @[top.scala 498:22]
  wire [31:0] dmem69_io_pipeline_writedata; // @[top.scala 498:22]
  wire  dmem69_io_pipeline_memread; // @[top.scala 498:22]
  wire  dmem69_io_pipeline_memwrite; // @[top.scala 498:22]
  wire [1:0] dmem69_io_pipeline_maskmode; // @[top.scala 498:22]
  wire  dmem69_io_pipeline_sext; // @[top.scala 498:22]
  wire [31:0] dmem69_io_pipeline_readdata; // @[top.scala 498:22]
  wire  dmem69_io_bus_request_valid; // @[top.scala 498:22]
  wire [31:0] dmem69_io_bus_request_bits_address; // @[top.scala 498:22]
  wire [31:0] dmem69_io_bus_request_bits_writedata; // @[top.scala 498:22]
  wire [1:0] dmem69_io_bus_request_bits_operation; // @[top.scala 498:22]
  wire  dmem69_io_bus_response_valid; // @[top.scala 498:22]
  wire [31:0] dmem69_io_bus_response_bits_data; // @[top.scala 498:22]
  wire  cpu70_clock; // @[top.scala 502:21]
  wire  cpu70_reset; // @[top.scala 502:21]
  wire [31:0] cpu70_io_imem_address; // @[top.scala 502:21]
  wire [31:0] cpu70_io_imem_instruction; // @[top.scala 502:21]
  wire [31:0] cpu70_io_dmem_address; // @[top.scala 502:21]
  wire  cpu70_io_dmem_valid; // @[top.scala 502:21]
  wire [31:0] cpu70_io_dmem_writedata; // @[top.scala 502:21]
  wire  cpu70_io_dmem_memread; // @[top.scala 502:21]
  wire  cpu70_io_dmem_memwrite; // @[top.scala 502:21]
  wire [1:0] cpu70_io_dmem_maskmode; // @[top.scala 502:21]
  wire  cpu70_io_dmem_sext; // @[top.scala 502:21]
  wire [31:0] cpu70_io_dmem_readdata; // @[top.scala 502:21]
  wire  mem70_clock; // @[top.scala 503:21]
  wire  mem70_reset; // @[top.scala 503:21]
  wire [31:0] mem70_io_imem_request_bits_address; // @[top.scala 503:21]
  wire [31:0] mem70_io_imem_response_bits_data; // @[top.scala 503:21]
  wire  mem70_io_dmem_request_valid; // @[top.scala 503:21]
  wire [31:0] mem70_io_dmem_request_bits_address; // @[top.scala 503:21]
  wire [31:0] mem70_io_dmem_request_bits_writedata; // @[top.scala 503:21]
  wire [1:0] mem70_io_dmem_request_bits_operation; // @[top.scala 503:21]
  wire  mem70_io_dmem_response_valid; // @[top.scala 503:21]
  wire [31:0] mem70_io_dmem_response_bits_data; // @[top.scala 503:21]
  wire [31:0] imem70_io_pipeline_address; // @[top.scala 504:22]
  wire [31:0] imem70_io_pipeline_instruction; // @[top.scala 504:22]
  wire [31:0] imem70_io_bus_request_bits_address; // @[top.scala 504:22]
  wire [31:0] imem70_io_bus_response_bits_data; // @[top.scala 504:22]
  wire  dmem70_clock; // @[top.scala 505:22]
  wire  dmem70_reset; // @[top.scala 505:22]
  wire [31:0] dmem70_io_pipeline_address; // @[top.scala 505:22]
  wire  dmem70_io_pipeline_valid; // @[top.scala 505:22]
  wire [31:0] dmem70_io_pipeline_writedata; // @[top.scala 505:22]
  wire  dmem70_io_pipeline_memread; // @[top.scala 505:22]
  wire  dmem70_io_pipeline_memwrite; // @[top.scala 505:22]
  wire [1:0] dmem70_io_pipeline_maskmode; // @[top.scala 505:22]
  wire  dmem70_io_pipeline_sext; // @[top.scala 505:22]
  wire [31:0] dmem70_io_pipeline_readdata; // @[top.scala 505:22]
  wire  dmem70_io_bus_request_valid; // @[top.scala 505:22]
  wire [31:0] dmem70_io_bus_request_bits_address; // @[top.scala 505:22]
  wire [31:0] dmem70_io_bus_request_bits_writedata; // @[top.scala 505:22]
  wire [1:0] dmem70_io_bus_request_bits_operation; // @[top.scala 505:22]
  wire  dmem70_io_bus_response_valid; // @[top.scala 505:22]
  wire [31:0] dmem70_io_bus_response_bits_data; // @[top.scala 505:22]
  wire  cpu71_clock; // @[top.scala 509:21]
  wire  cpu71_reset; // @[top.scala 509:21]
  wire [31:0] cpu71_io_imem_address; // @[top.scala 509:21]
  wire [31:0] cpu71_io_imem_instruction; // @[top.scala 509:21]
  wire [31:0] cpu71_io_dmem_address; // @[top.scala 509:21]
  wire  cpu71_io_dmem_valid; // @[top.scala 509:21]
  wire [31:0] cpu71_io_dmem_writedata; // @[top.scala 509:21]
  wire  cpu71_io_dmem_memread; // @[top.scala 509:21]
  wire  cpu71_io_dmem_memwrite; // @[top.scala 509:21]
  wire [1:0] cpu71_io_dmem_maskmode; // @[top.scala 509:21]
  wire  cpu71_io_dmem_sext; // @[top.scala 509:21]
  wire [31:0] cpu71_io_dmem_readdata; // @[top.scala 509:21]
  wire  mem71_clock; // @[top.scala 510:21]
  wire  mem71_reset; // @[top.scala 510:21]
  wire [31:0] mem71_io_imem_request_bits_address; // @[top.scala 510:21]
  wire [31:0] mem71_io_imem_response_bits_data; // @[top.scala 510:21]
  wire  mem71_io_dmem_request_valid; // @[top.scala 510:21]
  wire [31:0] mem71_io_dmem_request_bits_address; // @[top.scala 510:21]
  wire [31:0] mem71_io_dmem_request_bits_writedata; // @[top.scala 510:21]
  wire [1:0] mem71_io_dmem_request_bits_operation; // @[top.scala 510:21]
  wire  mem71_io_dmem_response_valid; // @[top.scala 510:21]
  wire [31:0] mem71_io_dmem_response_bits_data; // @[top.scala 510:21]
  wire [31:0] imem71_io_pipeline_address; // @[top.scala 511:22]
  wire [31:0] imem71_io_pipeline_instruction; // @[top.scala 511:22]
  wire [31:0] imem71_io_bus_request_bits_address; // @[top.scala 511:22]
  wire [31:0] imem71_io_bus_response_bits_data; // @[top.scala 511:22]
  wire  dmem71_clock; // @[top.scala 512:22]
  wire  dmem71_reset; // @[top.scala 512:22]
  wire [31:0] dmem71_io_pipeline_address; // @[top.scala 512:22]
  wire  dmem71_io_pipeline_valid; // @[top.scala 512:22]
  wire [31:0] dmem71_io_pipeline_writedata; // @[top.scala 512:22]
  wire  dmem71_io_pipeline_memread; // @[top.scala 512:22]
  wire  dmem71_io_pipeline_memwrite; // @[top.scala 512:22]
  wire [1:0] dmem71_io_pipeline_maskmode; // @[top.scala 512:22]
  wire  dmem71_io_pipeline_sext; // @[top.scala 512:22]
  wire [31:0] dmem71_io_pipeline_readdata; // @[top.scala 512:22]
  wire  dmem71_io_bus_request_valid; // @[top.scala 512:22]
  wire [31:0] dmem71_io_bus_request_bits_address; // @[top.scala 512:22]
  wire [31:0] dmem71_io_bus_request_bits_writedata; // @[top.scala 512:22]
  wire [1:0] dmem71_io_bus_request_bits_operation; // @[top.scala 512:22]
  wire  dmem71_io_bus_response_valid; // @[top.scala 512:22]
  wire [31:0] dmem71_io_bus_response_bits_data; // @[top.scala 512:22]
  wire  cpu72_clock; // @[top.scala 516:21]
  wire  cpu72_reset; // @[top.scala 516:21]
  wire [31:0] cpu72_io_imem_address; // @[top.scala 516:21]
  wire [31:0] cpu72_io_imem_instruction; // @[top.scala 516:21]
  wire [31:0] cpu72_io_dmem_address; // @[top.scala 516:21]
  wire  cpu72_io_dmem_valid; // @[top.scala 516:21]
  wire [31:0] cpu72_io_dmem_writedata; // @[top.scala 516:21]
  wire  cpu72_io_dmem_memread; // @[top.scala 516:21]
  wire  cpu72_io_dmem_memwrite; // @[top.scala 516:21]
  wire [1:0] cpu72_io_dmem_maskmode; // @[top.scala 516:21]
  wire  cpu72_io_dmem_sext; // @[top.scala 516:21]
  wire [31:0] cpu72_io_dmem_readdata; // @[top.scala 516:21]
  wire  mem72_clock; // @[top.scala 517:21]
  wire  mem72_reset; // @[top.scala 517:21]
  wire [31:0] mem72_io_imem_request_bits_address; // @[top.scala 517:21]
  wire [31:0] mem72_io_imem_response_bits_data; // @[top.scala 517:21]
  wire  mem72_io_dmem_request_valid; // @[top.scala 517:21]
  wire [31:0] mem72_io_dmem_request_bits_address; // @[top.scala 517:21]
  wire [31:0] mem72_io_dmem_request_bits_writedata; // @[top.scala 517:21]
  wire [1:0] mem72_io_dmem_request_bits_operation; // @[top.scala 517:21]
  wire  mem72_io_dmem_response_valid; // @[top.scala 517:21]
  wire [31:0] mem72_io_dmem_response_bits_data; // @[top.scala 517:21]
  wire [31:0] imem72_io_pipeline_address; // @[top.scala 518:22]
  wire [31:0] imem72_io_pipeline_instruction; // @[top.scala 518:22]
  wire [31:0] imem72_io_bus_request_bits_address; // @[top.scala 518:22]
  wire [31:0] imem72_io_bus_response_bits_data; // @[top.scala 518:22]
  wire  dmem72_clock; // @[top.scala 519:22]
  wire  dmem72_reset; // @[top.scala 519:22]
  wire [31:0] dmem72_io_pipeline_address; // @[top.scala 519:22]
  wire  dmem72_io_pipeline_valid; // @[top.scala 519:22]
  wire [31:0] dmem72_io_pipeline_writedata; // @[top.scala 519:22]
  wire  dmem72_io_pipeline_memread; // @[top.scala 519:22]
  wire  dmem72_io_pipeline_memwrite; // @[top.scala 519:22]
  wire [1:0] dmem72_io_pipeline_maskmode; // @[top.scala 519:22]
  wire  dmem72_io_pipeline_sext; // @[top.scala 519:22]
  wire [31:0] dmem72_io_pipeline_readdata; // @[top.scala 519:22]
  wire  dmem72_io_bus_request_valid; // @[top.scala 519:22]
  wire [31:0] dmem72_io_bus_request_bits_address; // @[top.scala 519:22]
  wire [31:0] dmem72_io_bus_request_bits_writedata; // @[top.scala 519:22]
  wire [1:0] dmem72_io_bus_request_bits_operation; // @[top.scala 519:22]
  wire  dmem72_io_bus_response_valid; // @[top.scala 519:22]
  wire [31:0] dmem72_io_bus_response_bits_data; // @[top.scala 519:22]
  wire  cpu73_clock; // @[top.scala 523:21]
  wire  cpu73_reset; // @[top.scala 523:21]
  wire [31:0] cpu73_io_imem_address; // @[top.scala 523:21]
  wire [31:0] cpu73_io_imem_instruction; // @[top.scala 523:21]
  wire [31:0] cpu73_io_dmem_address; // @[top.scala 523:21]
  wire  cpu73_io_dmem_valid; // @[top.scala 523:21]
  wire [31:0] cpu73_io_dmem_writedata; // @[top.scala 523:21]
  wire  cpu73_io_dmem_memread; // @[top.scala 523:21]
  wire  cpu73_io_dmem_memwrite; // @[top.scala 523:21]
  wire [1:0] cpu73_io_dmem_maskmode; // @[top.scala 523:21]
  wire  cpu73_io_dmem_sext; // @[top.scala 523:21]
  wire [31:0] cpu73_io_dmem_readdata; // @[top.scala 523:21]
  wire  mem73_clock; // @[top.scala 524:21]
  wire  mem73_reset; // @[top.scala 524:21]
  wire [31:0] mem73_io_imem_request_bits_address; // @[top.scala 524:21]
  wire [31:0] mem73_io_imem_response_bits_data; // @[top.scala 524:21]
  wire  mem73_io_dmem_request_valid; // @[top.scala 524:21]
  wire [31:0] mem73_io_dmem_request_bits_address; // @[top.scala 524:21]
  wire [31:0] mem73_io_dmem_request_bits_writedata; // @[top.scala 524:21]
  wire [1:0] mem73_io_dmem_request_bits_operation; // @[top.scala 524:21]
  wire  mem73_io_dmem_response_valid; // @[top.scala 524:21]
  wire [31:0] mem73_io_dmem_response_bits_data; // @[top.scala 524:21]
  wire [31:0] imem73_io_pipeline_address; // @[top.scala 525:22]
  wire [31:0] imem73_io_pipeline_instruction; // @[top.scala 525:22]
  wire [31:0] imem73_io_bus_request_bits_address; // @[top.scala 525:22]
  wire [31:0] imem73_io_bus_response_bits_data; // @[top.scala 525:22]
  wire  dmem73_clock; // @[top.scala 526:22]
  wire  dmem73_reset; // @[top.scala 526:22]
  wire [31:0] dmem73_io_pipeline_address; // @[top.scala 526:22]
  wire  dmem73_io_pipeline_valid; // @[top.scala 526:22]
  wire [31:0] dmem73_io_pipeline_writedata; // @[top.scala 526:22]
  wire  dmem73_io_pipeline_memread; // @[top.scala 526:22]
  wire  dmem73_io_pipeline_memwrite; // @[top.scala 526:22]
  wire [1:0] dmem73_io_pipeline_maskmode; // @[top.scala 526:22]
  wire  dmem73_io_pipeline_sext; // @[top.scala 526:22]
  wire [31:0] dmem73_io_pipeline_readdata; // @[top.scala 526:22]
  wire  dmem73_io_bus_request_valid; // @[top.scala 526:22]
  wire [31:0] dmem73_io_bus_request_bits_address; // @[top.scala 526:22]
  wire [31:0] dmem73_io_bus_request_bits_writedata; // @[top.scala 526:22]
  wire [1:0] dmem73_io_bus_request_bits_operation; // @[top.scala 526:22]
  wire  dmem73_io_bus_response_valid; // @[top.scala 526:22]
  wire [31:0] dmem73_io_bus_response_bits_data; // @[top.scala 526:22]
  wire  cpu74_clock; // @[top.scala 530:21]
  wire  cpu74_reset; // @[top.scala 530:21]
  wire [31:0] cpu74_io_imem_address; // @[top.scala 530:21]
  wire [31:0] cpu74_io_imem_instruction; // @[top.scala 530:21]
  wire [31:0] cpu74_io_dmem_address; // @[top.scala 530:21]
  wire  cpu74_io_dmem_valid; // @[top.scala 530:21]
  wire [31:0] cpu74_io_dmem_writedata; // @[top.scala 530:21]
  wire  cpu74_io_dmem_memread; // @[top.scala 530:21]
  wire  cpu74_io_dmem_memwrite; // @[top.scala 530:21]
  wire [1:0] cpu74_io_dmem_maskmode; // @[top.scala 530:21]
  wire  cpu74_io_dmem_sext; // @[top.scala 530:21]
  wire [31:0] cpu74_io_dmem_readdata; // @[top.scala 530:21]
  wire  mem74_clock; // @[top.scala 531:21]
  wire  mem74_reset; // @[top.scala 531:21]
  wire [31:0] mem74_io_imem_request_bits_address; // @[top.scala 531:21]
  wire [31:0] mem74_io_imem_response_bits_data; // @[top.scala 531:21]
  wire  mem74_io_dmem_request_valid; // @[top.scala 531:21]
  wire [31:0] mem74_io_dmem_request_bits_address; // @[top.scala 531:21]
  wire [31:0] mem74_io_dmem_request_bits_writedata; // @[top.scala 531:21]
  wire [1:0] mem74_io_dmem_request_bits_operation; // @[top.scala 531:21]
  wire  mem74_io_dmem_response_valid; // @[top.scala 531:21]
  wire [31:0] mem74_io_dmem_response_bits_data; // @[top.scala 531:21]
  wire [31:0] imem74_io_pipeline_address; // @[top.scala 532:22]
  wire [31:0] imem74_io_pipeline_instruction; // @[top.scala 532:22]
  wire [31:0] imem74_io_bus_request_bits_address; // @[top.scala 532:22]
  wire [31:0] imem74_io_bus_response_bits_data; // @[top.scala 532:22]
  wire  dmem74_clock; // @[top.scala 533:22]
  wire  dmem74_reset; // @[top.scala 533:22]
  wire [31:0] dmem74_io_pipeline_address; // @[top.scala 533:22]
  wire  dmem74_io_pipeline_valid; // @[top.scala 533:22]
  wire [31:0] dmem74_io_pipeline_writedata; // @[top.scala 533:22]
  wire  dmem74_io_pipeline_memread; // @[top.scala 533:22]
  wire  dmem74_io_pipeline_memwrite; // @[top.scala 533:22]
  wire [1:0] dmem74_io_pipeline_maskmode; // @[top.scala 533:22]
  wire  dmem74_io_pipeline_sext; // @[top.scala 533:22]
  wire [31:0] dmem74_io_pipeline_readdata; // @[top.scala 533:22]
  wire  dmem74_io_bus_request_valid; // @[top.scala 533:22]
  wire [31:0] dmem74_io_bus_request_bits_address; // @[top.scala 533:22]
  wire [31:0] dmem74_io_bus_request_bits_writedata; // @[top.scala 533:22]
  wire [1:0] dmem74_io_bus_request_bits_operation; // @[top.scala 533:22]
  wire  dmem74_io_bus_response_valid; // @[top.scala 533:22]
  wire [31:0] dmem74_io_bus_response_bits_data; // @[top.scala 533:22]
  wire  cpu75_clock; // @[top.scala 537:21]
  wire  cpu75_reset; // @[top.scala 537:21]
  wire [31:0] cpu75_io_imem_address; // @[top.scala 537:21]
  wire [31:0] cpu75_io_imem_instruction; // @[top.scala 537:21]
  wire [31:0] cpu75_io_dmem_address; // @[top.scala 537:21]
  wire  cpu75_io_dmem_valid; // @[top.scala 537:21]
  wire [31:0] cpu75_io_dmem_writedata; // @[top.scala 537:21]
  wire  cpu75_io_dmem_memread; // @[top.scala 537:21]
  wire  cpu75_io_dmem_memwrite; // @[top.scala 537:21]
  wire [1:0] cpu75_io_dmem_maskmode; // @[top.scala 537:21]
  wire  cpu75_io_dmem_sext; // @[top.scala 537:21]
  wire [31:0] cpu75_io_dmem_readdata; // @[top.scala 537:21]
  wire  mem75_clock; // @[top.scala 538:21]
  wire  mem75_reset; // @[top.scala 538:21]
  wire [31:0] mem75_io_imem_request_bits_address; // @[top.scala 538:21]
  wire [31:0] mem75_io_imem_response_bits_data; // @[top.scala 538:21]
  wire  mem75_io_dmem_request_valid; // @[top.scala 538:21]
  wire [31:0] mem75_io_dmem_request_bits_address; // @[top.scala 538:21]
  wire [31:0] mem75_io_dmem_request_bits_writedata; // @[top.scala 538:21]
  wire [1:0] mem75_io_dmem_request_bits_operation; // @[top.scala 538:21]
  wire  mem75_io_dmem_response_valid; // @[top.scala 538:21]
  wire [31:0] mem75_io_dmem_response_bits_data; // @[top.scala 538:21]
  wire [31:0] imem75_io_pipeline_address; // @[top.scala 539:22]
  wire [31:0] imem75_io_pipeline_instruction; // @[top.scala 539:22]
  wire [31:0] imem75_io_bus_request_bits_address; // @[top.scala 539:22]
  wire [31:0] imem75_io_bus_response_bits_data; // @[top.scala 539:22]
  wire  dmem75_clock; // @[top.scala 540:22]
  wire  dmem75_reset; // @[top.scala 540:22]
  wire [31:0] dmem75_io_pipeline_address; // @[top.scala 540:22]
  wire  dmem75_io_pipeline_valid; // @[top.scala 540:22]
  wire [31:0] dmem75_io_pipeline_writedata; // @[top.scala 540:22]
  wire  dmem75_io_pipeline_memread; // @[top.scala 540:22]
  wire  dmem75_io_pipeline_memwrite; // @[top.scala 540:22]
  wire [1:0] dmem75_io_pipeline_maskmode; // @[top.scala 540:22]
  wire  dmem75_io_pipeline_sext; // @[top.scala 540:22]
  wire [31:0] dmem75_io_pipeline_readdata; // @[top.scala 540:22]
  wire  dmem75_io_bus_request_valid; // @[top.scala 540:22]
  wire [31:0] dmem75_io_bus_request_bits_address; // @[top.scala 540:22]
  wire [31:0] dmem75_io_bus_request_bits_writedata; // @[top.scala 540:22]
  wire [1:0] dmem75_io_bus_request_bits_operation; // @[top.scala 540:22]
  wire  dmem75_io_bus_response_valid; // @[top.scala 540:22]
  wire [31:0] dmem75_io_bus_response_bits_data; // @[top.scala 540:22]
  wire  cpu76_clock; // @[top.scala 544:21]
  wire  cpu76_reset; // @[top.scala 544:21]
  wire [31:0] cpu76_io_imem_address; // @[top.scala 544:21]
  wire [31:0] cpu76_io_imem_instruction; // @[top.scala 544:21]
  wire [31:0] cpu76_io_dmem_address; // @[top.scala 544:21]
  wire  cpu76_io_dmem_valid; // @[top.scala 544:21]
  wire [31:0] cpu76_io_dmem_writedata; // @[top.scala 544:21]
  wire  cpu76_io_dmem_memread; // @[top.scala 544:21]
  wire  cpu76_io_dmem_memwrite; // @[top.scala 544:21]
  wire [1:0] cpu76_io_dmem_maskmode; // @[top.scala 544:21]
  wire  cpu76_io_dmem_sext; // @[top.scala 544:21]
  wire [31:0] cpu76_io_dmem_readdata; // @[top.scala 544:21]
  wire  mem76_clock; // @[top.scala 545:21]
  wire  mem76_reset; // @[top.scala 545:21]
  wire [31:0] mem76_io_imem_request_bits_address; // @[top.scala 545:21]
  wire [31:0] mem76_io_imem_response_bits_data; // @[top.scala 545:21]
  wire  mem76_io_dmem_request_valid; // @[top.scala 545:21]
  wire [31:0] mem76_io_dmem_request_bits_address; // @[top.scala 545:21]
  wire [31:0] mem76_io_dmem_request_bits_writedata; // @[top.scala 545:21]
  wire [1:0] mem76_io_dmem_request_bits_operation; // @[top.scala 545:21]
  wire  mem76_io_dmem_response_valid; // @[top.scala 545:21]
  wire [31:0] mem76_io_dmem_response_bits_data; // @[top.scala 545:21]
  wire [31:0] imem76_io_pipeline_address; // @[top.scala 546:22]
  wire [31:0] imem76_io_pipeline_instruction; // @[top.scala 546:22]
  wire [31:0] imem76_io_bus_request_bits_address; // @[top.scala 546:22]
  wire [31:0] imem76_io_bus_response_bits_data; // @[top.scala 546:22]
  wire  dmem76_clock; // @[top.scala 547:22]
  wire  dmem76_reset; // @[top.scala 547:22]
  wire [31:0] dmem76_io_pipeline_address; // @[top.scala 547:22]
  wire  dmem76_io_pipeline_valid; // @[top.scala 547:22]
  wire [31:0] dmem76_io_pipeline_writedata; // @[top.scala 547:22]
  wire  dmem76_io_pipeline_memread; // @[top.scala 547:22]
  wire  dmem76_io_pipeline_memwrite; // @[top.scala 547:22]
  wire [1:0] dmem76_io_pipeline_maskmode; // @[top.scala 547:22]
  wire  dmem76_io_pipeline_sext; // @[top.scala 547:22]
  wire [31:0] dmem76_io_pipeline_readdata; // @[top.scala 547:22]
  wire  dmem76_io_bus_request_valid; // @[top.scala 547:22]
  wire [31:0] dmem76_io_bus_request_bits_address; // @[top.scala 547:22]
  wire [31:0] dmem76_io_bus_request_bits_writedata; // @[top.scala 547:22]
  wire [1:0] dmem76_io_bus_request_bits_operation; // @[top.scala 547:22]
  wire  dmem76_io_bus_response_valid; // @[top.scala 547:22]
  wire [31:0] dmem76_io_bus_response_bits_data; // @[top.scala 547:22]
  wire  cpu77_clock; // @[top.scala 551:21]
  wire  cpu77_reset; // @[top.scala 551:21]
  wire [31:0] cpu77_io_imem_address; // @[top.scala 551:21]
  wire [31:0] cpu77_io_imem_instruction; // @[top.scala 551:21]
  wire [31:0] cpu77_io_dmem_address; // @[top.scala 551:21]
  wire  cpu77_io_dmem_valid; // @[top.scala 551:21]
  wire [31:0] cpu77_io_dmem_writedata; // @[top.scala 551:21]
  wire  cpu77_io_dmem_memread; // @[top.scala 551:21]
  wire  cpu77_io_dmem_memwrite; // @[top.scala 551:21]
  wire [1:0] cpu77_io_dmem_maskmode; // @[top.scala 551:21]
  wire  cpu77_io_dmem_sext; // @[top.scala 551:21]
  wire [31:0] cpu77_io_dmem_readdata; // @[top.scala 551:21]
  wire  mem77_clock; // @[top.scala 552:21]
  wire  mem77_reset; // @[top.scala 552:21]
  wire [31:0] mem77_io_imem_request_bits_address; // @[top.scala 552:21]
  wire [31:0] mem77_io_imem_response_bits_data; // @[top.scala 552:21]
  wire  mem77_io_dmem_request_valid; // @[top.scala 552:21]
  wire [31:0] mem77_io_dmem_request_bits_address; // @[top.scala 552:21]
  wire [31:0] mem77_io_dmem_request_bits_writedata; // @[top.scala 552:21]
  wire [1:0] mem77_io_dmem_request_bits_operation; // @[top.scala 552:21]
  wire  mem77_io_dmem_response_valid; // @[top.scala 552:21]
  wire [31:0] mem77_io_dmem_response_bits_data; // @[top.scala 552:21]
  wire [31:0] imem77_io_pipeline_address; // @[top.scala 553:22]
  wire [31:0] imem77_io_pipeline_instruction; // @[top.scala 553:22]
  wire [31:0] imem77_io_bus_request_bits_address; // @[top.scala 553:22]
  wire [31:0] imem77_io_bus_response_bits_data; // @[top.scala 553:22]
  wire  dmem77_clock; // @[top.scala 554:22]
  wire  dmem77_reset; // @[top.scala 554:22]
  wire [31:0] dmem77_io_pipeline_address; // @[top.scala 554:22]
  wire  dmem77_io_pipeline_valid; // @[top.scala 554:22]
  wire [31:0] dmem77_io_pipeline_writedata; // @[top.scala 554:22]
  wire  dmem77_io_pipeline_memread; // @[top.scala 554:22]
  wire  dmem77_io_pipeline_memwrite; // @[top.scala 554:22]
  wire [1:0] dmem77_io_pipeline_maskmode; // @[top.scala 554:22]
  wire  dmem77_io_pipeline_sext; // @[top.scala 554:22]
  wire [31:0] dmem77_io_pipeline_readdata; // @[top.scala 554:22]
  wire  dmem77_io_bus_request_valid; // @[top.scala 554:22]
  wire [31:0] dmem77_io_bus_request_bits_address; // @[top.scala 554:22]
  wire [31:0] dmem77_io_bus_request_bits_writedata; // @[top.scala 554:22]
  wire [1:0] dmem77_io_bus_request_bits_operation; // @[top.scala 554:22]
  wire  dmem77_io_bus_response_valid; // @[top.scala 554:22]
  wire [31:0] dmem77_io_bus_response_bits_data; // @[top.scala 554:22]
  wire  cpu78_clock; // @[top.scala 558:21]
  wire  cpu78_reset; // @[top.scala 558:21]
  wire [31:0] cpu78_io_imem_address; // @[top.scala 558:21]
  wire [31:0] cpu78_io_imem_instruction; // @[top.scala 558:21]
  wire [31:0] cpu78_io_dmem_address; // @[top.scala 558:21]
  wire  cpu78_io_dmem_valid; // @[top.scala 558:21]
  wire [31:0] cpu78_io_dmem_writedata; // @[top.scala 558:21]
  wire  cpu78_io_dmem_memread; // @[top.scala 558:21]
  wire  cpu78_io_dmem_memwrite; // @[top.scala 558:21]
  wire [1:0] cpu78_io_dmem_maskmode; // @[top.scala 558:21]
  wire  cpu78_io_dmem_sext; // @[top.scala 558:21]
  wire [31:0] cpu78_io_dmem_readdata; // @[top.scala 558:21]
  wire  mem78_clock; // @[top.scala 559:21]
  wire  mem78_reset; // @[top.scala 559:21]
  wire [31:0] mem78_io_imem_request_bits_address; // @[top.scala 559:21]
  wire [31:0] mem78_io_imem_response_bits_data; // @[top.scala 559:21]
  wire  mem78_io_dmem_request_valid; // @[top.scala 559:21]
  wire [31:0] mem78_io_dmem_request_bits_address; // @[top.scala 559:21]
  wire [31:0] mem78_io_dmem_request_bits_writedata; // @[top.scala 559:21]
  wire [1:0] mem78_io_dmem_request_bits_operation; // @[top.scala 559:21]
  wire  mem78_io_dmem_response_valid; // @[top.scala 559:21]
  wire [31:0] mem78_io_dmem_response_bits_data; // @[top.scala 559:21]
  wire [31:0] imem78_io_pipeline_address; // @[top.scala 560:22]
  wire [31:0] imem78_io_pipeline_instruction; // @[top.scala 560:22]
  wire [31:0] imem78_io_bus_request_bits_address; // @[top.scala 560:22]
  wire [31:0] imem78_io_bus_response_bits_data; // @[top.scala 560:22]
  wire  dmem78_clock; // @[top.scala 561:22]
  wire  dmem78_reset; // @[top.scala 561:22]
  wire [31:0] dmem78_io_pipeline_address; // @[top.scala 561:22]
  wire  dmem78_io_pipeline_valid; // @[top.scala 561:22]
  wire [31:0] dmem78_io_pipeline_writedata; // @[top.scala 561:22]
  wire  dmem78_io_pipeline_memread; // @[top.scala 561:22]
  wire  dmem78_io_pipeline_memwrite; // @[top.scala 561:22]
  wire [1:0] dmem78_io_pipeline_maskmode; // @[top.scala 561:22]
  wire  dmem78_io_pipeline_sext; // @[top.scala 561:22]
  wire [31:0] dmem78_io_pipeline_readdata; // @[top.scala 561:22]
  wire  dmem78_io_bus_request_valid; // @[top.scala 561:22]
  wire [31:0] dmem78_io_bus_request_bits_address; // @[top.scala 561:22]
  wire [31:0] dmem78_io_bus_request_bits_writedata; // @[top.scala 561:22]
  wire [1:0] dmem78_io_bus_request_bits_operation; // @[top.scala 561:22]
  wire  dmem78_io_bus_response_valid; // @[top.scala 561:22]
  wire [31:0] dmem78_io_bus_response_bits_data; // @[top.scala 561:22]
  wire  cpu79_clock; // @[top.scala 565:21]
  wire  cpu79_reset; // @[top.scala 565:21]
  wire [31:0] cpu79_io_imem_address; // @[top.scala 565:21]
  wire [31:0] cpu79_io_imem_instruction; // @[top.scala 565:21]
  wire [31:0] cpu79_io_dmem_address; // @[top.scala 565:21]
  wire  cpu79_io_dmem_valid; // @[top.scala 565:21]
  wire [31:0] cpu79_io_dmem_writedata; // @[top.scala 565:21]
  wire  cpu79_io_dmem_memread; // @[top.scala 565:21]
  wire  cpu79_io_dmem_memwrite; // @[top.scala 565:21]
  wire [1:0] cpu79_io_dmem_maskmode; // @[top.scala 565:21]
  wire  cpu79_io_dmem_sext; // @[top.scala 565:21]
  wire [31:0] cpu79_io_dmem_readdata; // @[top.scala 565:21]
  wire  mem79_clock; // @[top.scala 566:21]
  wire  mem79_reset; // @[top.scala 566:21]
  wire [31:0] mem79_io_imem_request_bits_address; // @[top.scala 566:21]
  wire [31:0] mem79_io_imem_response_bits_data; // @[top.scala 566:21]
  wire  mem79_io_dmem_request_valid; // @[top.scala 566:21]
  wire [31:0] mem79_io_dmem_request_bits_address; // @[top.scala 566:21]
  wire [31:0] mem79_io_dmem_request_bits_writedata; // @[top.scala 566:21]
  wire [1:0] mem79_io_dmem_request_bits_operation; // @[top.scala 566:21]
  wire  mem79_io_dmem_response_valid; // @[top.scala 566:21]
  wire [31:0] mem79_io_dmem_response_bits_data; // @[top.scala 566:21]
  wire [31:0] imem79_io_pipeline_address; // @[top.scala 567:22]
  wire [31:0] imem79_io_pipeline_instruction; // @[top.scala 567:22]
  wire [31:0] imem79_io_bus_request_bits_address; // @[top.scala 567:22]
  wire [31:0] imem79_io_bus_response_bits_data; // @[top.scala 567:22]
  wire  dmem79_clock; // @[top.scala 568:22]
  wire  dmem79_reset; // @[top.scala 568:22]
  wire [31:0] dmem79_io_pipeline_address; // @[top.scala 568:22]
  wire  dmem79_io_pipeline_valid; // @[top.scala 568:22]
  wire [31:0] dmem79_io_pipeline_writedata; // @[top.scala 568:22]
  wire  dmem79_io_pipeline_memread; // @[top.scala 568:22]
  wire  dmem79_io_pipeline_memwrite; // @[top.scala 568:22]
  wire [1:0] dmem79_io_pipeline_maskmode; // @[top.scala 568:22]
  wire  dmem79_io_pipeline_sext; // @[top.scala 568:22]
  wire [31:0] dmem79_io_pipeline_readdata; // @[top.scala 568:22]
  wire  dmem79_io_bus_request_valid; // @[top.scala 568:22]
  wire [31:0] dmem79_io_bus_request_bits_address; // @[top.scala 568:22]
  wire [31:0] dmem79_io_bus_request_bits_writedata; // @[top.scala 568:22]
  wire [1:0] dmem79_io_bus_request_bits_operation; // @[top.scala 568:22]
  wire  dmem79_io_bus_response_valid; // @[top.scala 568:22]
  wire [31:0] dmem79_io_bus_response_bits_data; // @[top.scala 568:22]
  wire  cpu80_clock; // @[top.scala 572:21]
  wire  cpu80_reset; // @[top.scala 572:21]
  wire [31:0] cpu80_io_imem_address; // @[top.scala 572:21]
  wire [31:0] cpu80_io_imem_instruction; // @[top.scala 572:21]
  wire [31:0] cpu80_io_dmem_address; // @[top.scala 572:21]
  wire  cpu80_io_dmem_valid; // @[top.scala 572:21]
  wire [31:0] cpu80_io_dmem_writedata; // @[top.scala 572:21]
  wire  cpu80_io_dmem_memread; // @[top.scala 572:21]
  wire  cpu80_io_dmem_memwrite; // @[top.scala 572:21]
  wire [1:0] cpu80_io_dmem_maskmode; // @[top.scala 572:21]
  wire  cpu80_io_dmem_sext; // @[top.scala 572:21]
  wire [31:0] cpu80_io_dmem_readdata; // @[top.scala 572:21]
  wire  mem80_clock; // @[top.scala 573:21]
  wire  mem80_reset; // @[top.scala 573:21]
  wire [31:0] mem80_io_imem_request_bits_address; // @[top.scala 573:21]
  wire [31:0] mem80_io_imem_response_bits_data; // @[top.scala 573:21]
  wire  mem80_io_dmem_request_valid; // @[top.scala 573:21]
  wire [31:0] mem80_io_dmem_request_bits_address; // @[top.scala 573:21]
  wire [31:0] mem80_io_dmem_request_bits_writedata; // @[top.scala 573:21]
  wire [1:0] mem80_io_dmem_request_bits_operation; // @[top.scala 573:21]
  wire  mem80_io_dmem_response_valid; // @[top.scala 573:21]
  wire [31:0] mem80_io_dmem_response_bits_data; // @[top.scala 573:21]
  wire [31:0] imem80_io_pipeline_address; // @[top.scala 574:22]
  wire [31:0] imem80_io_pipeline_instruction; // @[top.scala 574:22]
  wire [31:0] imem80_io_bus_request_bits_address; // @[top.scala 574:22]
  wire [31:0] imem80_io_bus_response_bits_data; // @[top.scala 574:22]
  wire  dmem80_clock; // @[top.scala 575:22]
  wire  dmem80_reset; // @[top.scala 575:22]
  wire [31:0] dmem80_io_pipeline_address; // @[top.scala 575:22]
  wire  dmem80_io_pipeline_valid; // @[top.scala 575:22]
  wire [31:0] dmem80_io_pipeline_writedata; // @[top.scala 575:22]
  wire  dmem80_io_pipeline_memread; // @[top.scala 575:22]
  wire  dmem80_io_pipeline_memwrite; // @[top.scala 575:22]
  wire [1:0] dmem80_io_pipeline_maskmode; // @[top.scala 575:22]
  wire  dmem80_io_pipeline_sext; // @[top.scala 575:22]
  wire [31:0] dmem80_io_pipeline_readdata; // @[top.scala 575:22]
  wire  dmem80_io_bus_request_valid; // @[top.scala 575:22]
  wire [31:0] dmem80_io_bus_request_bits_address; // @[top.scala 575:22]
  wire [31:0] dmem80_io_bus_request_bits_writedata; // @[top.scala 575:22]
  wire [1:0] dmem80_io_bus_request_bits_operation; // @[top.scala 575:22]
  wire  dmem80_io_bus_response_valid; // @[top.scala 575:22]
  wire [31:0] dmem80_io_bus_response_bits_data; // @[top.scala 575:22]
  wire  cpu81_clock; // @[top.scala 579:21]
  wire  cpu81_reset; // @[top.scala 579:21]
  wire [31:0] cpu81_io_imem_address; // @[top.scala 579:21]
  wire [31:0] cpu81_io_imem_instruction; // @[top.scala 579:21]
  wire [31:0] cpu81_io_dmem_address; // @[top.scala 579:21]
  wire  cpu81_io_dmem_valid; // @[top.scala 579:21]
  wire [31:0] cpu81_io_dmem_writedata; // @[top.scala 579:21]
  wire  cpu81_io_dmem_memread; // @[top.scala 579:21]
  wire  cpu81_io_dmem_memwrite; // @[top.scala 579:21]
  wire [1:0] cpu81_io_dmem_maskmode; // @[top.scala 579:21]
  wire  cpu81_io_dmem_sext; // @[top.scala 579:21]
  wire [31:0] cpu81_io_dmem_readdata; // @[top.scala 579:21]
  wire  mem81_clock; // @[top.scala 580:21]
  wire  mem81_reset; // @[top.scala 580:21]
  wire [31:0] mem81_io_imem_request_bits_address; // @[top.scala 580:21]
  wire [31:0] mem81_io_imem_response_bits_data; // @[top.scala 580:21]
  wire  mem81_io_dmem_request_valid; // @[top.scala 580:21]
  wire [31:0] mem81_io_dmem_request_bits_address; // @[top.scala 580:21]
  wire [31:0] mem81_io_dmem_request_bits_writedata; // @[top.scala 580:21]
  wire [1:0] mem81_io_dmem_request_bits_operation; // @[top.scala 580:21]
  wire  mem81_io_dmem_response_valid; // @[top.scala 580:21]
  wire [31:0] mem81_io_dmem_response_bits_data; // @[top.scala 580:21]
  wire [31:0] imem81_io_pipeline_address; // @[top.scala 581:22]
  wire [31:0] imem81_io_pipeline_instruction; // @[top.scala 581:22]
  wire [31:0] imem81_io_bus_request_bits_address; // @[top.scala 581:22]
  wire [31:0] imem81_io_bus_response_bits_data; // @[top.scala 581:22]
  wire  dmem81_clock; // @[top.scala 582:22]
  wire  dmem81_reset; // @[top.scala 582:22]
  wire [31:0] dmem81_io_pipeline_address; // @[top.scala 582:22]
  wire  dmem81_io_pipeline_valid; // @[top.scala 582:22]
  wire [31:0] dmem81_io_pipeline_writedata; // @[top.scala 582:22]
  wire  dmem81_io_pipeline_memread; // @[top.scala 582:22]
  wire  dmem81_io_pipeline_memwrite; // @[top.scala 582:22]
  wire [1:0] dmem81_io_pipeline_maskmode; // @[top.scala 582:22]
  wire  dmem81_io_pipeline_sext; // @[top.scala 582:22]
  wire [31:0] dmem81_io_pipeline_readdata; // @[top.scala 582:22]
  wire  dmem81_io_bus_request_valid; // @[top.scala 582:22]
  wire [31:0] dmem81_io_bus_request_bits_address; // @[top.scala 582:22]
  wire [31:0] dmem81_io_bus_request_bits_writedata; // @[top.scala 582:22]
  wire [1:0] dmem81_io_bus_request_bits_operation; // @[top.scala 582:22]
  wire  dmem81_io_bus_response_valid; // @[top.scala 582:22]
  wire [31:0] dmem81_io_bus_response_bits_data; // @[top.scala 582:22]
  wire  cpu82_clock; // @[top.scala 586:21]
  wire  cpu82_reset; // @[top.scala 586:21]
  wire [31:0] cpu82_io_imem_address; // @[top.scala 586:21]
  wire [31:0] cpu82_io_imem_instruction; // @[top.scala 586:21]
  wire [31:0] cpu82_io_dmem_address; // @[top.scala 586:21]
  wire  cpu82_io_dmem_valid; // @[top.scala 586:21]
  wire [31:0] cpu82_io_dmem_writedata; // @[top.scala 586:21]
  wire  cpu82_io_dmem_memread; // @[top.scala 586:21]
  wire  cpu82_io_dmem_memwrite; // @[top.scala 586:21]
  wire [1:0] cpu82_io_dmem_maskmode; // @[top.scala 586:21]
  wire  cpu82_io_dmem_sext; // @[top.scala 586:21]
  wire [31:0] cpu82_io_dmem_readdata; // @[top.scala 586:21]
  wire  mem82_clock; // @[top.scala 587:21]
  wire  mem82_reset; // @[top.scala 587:21]
  wire [31:0] mem82_io_imem_request_bits_address; // @[top.scala 587:21]
  wire [31:0] mem82_io_imem_response_bits_data; // @[top.scala 587:21]
  wire  mem82_io_dmem_request_valid; // @[top.scala 587:21]
  wire [31:0] mem82_io_dmem_request_bits_address; // @[top.scala 587:21]
  wire [31:0] mem82_io_dmem_request_bits_writedata; // @[top.scala 587:21]
  wire [1:0] mem82_io_dmem_request_bits_operation; // @[top.scala 587:21]
  wire  mem82_io_dmem_response_valid; // @[top.scala 587:21]
  wire [31:0] mem82_io_dmem_response_bits_data; // @[top.scala 587:21]
  wire [31:0] imem82_io_pipeline_address; // @[top.scala 588:22]
  wire [31:0] imem82_io_pipeline_instruction; // @[top.scala 588:22]
  wire [31:0] imem82_io_bus_request_bits_address; // @[top.scala 588:22]
  wire [31:0] imem82_io_bus_response_bits_data; // @[top.scala 588:22]
  wire  dmem82_clock; // @[top.scala 589:22]
  wire  dmem82_reset; // @[top.scala 589:22]
  wire [31:0] dmem82_io_pipeline_address; // @[top.scala 589:22]
  wire  dmem82_io_pipeline_valid; // @[top.scala 589:22]
  wire [31:0] dmem82_io_pipeline_writedata; // @[top.scala 589:22]
  wire  dmem82_io_pipeline_memread; // @[top.scala 589:22]
  wire  dmem82_io_pipeline_memwrite; // @[top.scala 589:22]
  wire [1:0] dmem82_io_pipeline_maskmode; // @[top.scala 589:22]
  wire  dmem82_io_pipeline_sext; // @[top.scala 589:22]
  wire [31:0] dmem82_io_pipeline_readdata; // @[top.scala 589:22]
  wire  dmem82_io_bus_request_valid; // @[top.scala 589:22]
  wire [31:0] dmem82_io_bus_request_bits_address; // @[top.scala 589:22]
  wire [31:0] dmem82_io_bus_request_bits_writedata; // @[top.scala 589:22]
  wire [1:0] dmem82_io_bus_request_bits_operation; // @[top.scala 589:22]
  wire  dmem82_io_bus_response_valid; // @[top.scala 589:22]
  wire [31:0] dmem82_io_bus_response_bits_data; // @[top.scala 589:22]
  wire  cpu83_clock; // @[top.scala 593:21]
  wire  cpu83_reset; // @[top.scala 593:21]
  wire [31:0] cpu83_io_imem_address; // @[top.scala 593:21]
  wire [31:0] cpu83_io_imem_instruction; // @[top.scala 593:21]
  wire [31:0] cpu83_io_dmem_address; // @[top.scala 593:21]
  wire  cpu83_io_dmem_valid; // @[top.scala 593:21]
  wire [31:0] cpu83_io_dmem_writedata; // @[top.scala 593:21]
  wire  cpu83_io_dmem_memread; // @[top.scala 593:21]
  wire  cpu83_io_dmem_memwrite; // @[top.scala 593:21]
  wire [1:0] cpu83_io_dmem_maskmode; // @[top.scala 593:21]
  wire  cpu83_io_dmem_sext; // @[top.scala 593:21]
  wire [31:0] cpu83_io_dmem_readdata; // @[top.scala 593:21]
  wire  mem83_clock; // @[top.scala 594:21]
  wire  mem83_reset; // @[top.scala 594:21]
  wire [31:0] mem83_io_imem_request_bits_address; // @[top.scala 594:21]
  wire [31:0] mem83_io_imem_response_bits_data; // @[top.scala 594:21]
  wire  mem83_io_dmem_request_valid; // @[top.scala 594:21]
  wire [31:0] mem83_io_dmem_request_bits_address; // @[top.scala 594:21]
  wire [31:0] mem83_io_dmem_request_bits_writedata; // @[top.scala 594:21]
  wire [1:0] mem83_io_dmem_request_bits_operation; // @[top.scala 594:21]
  wire  mem83_io_dmem_response_valid; // @[top.scala 594:21]
  wire [31:0] mem83_io_dmem_response_bits_data; // @[top.scala 594:21]
  wire [31:0] imem83_io_pipeline_address; // @[top.scala 595:22]
  wire [31:0] imem83_io_pipeline_instruction; // @[top.scala 595:22]
  wire [31:0] imem83_io_bus_request_bits_address; // @[top.scala 595:22]
  wire [31:0] imem83_io_bus_response_bits_data; // @[top.scala 595:22]
  wire  dmem83_clock; // @[top.scala 596:22]
  wire  dmem83_reset; // @[top.scala 596:22]
  wire [31:0] dmem83_io_pipeline_address; // @[top.scala 596:22]
  wire  dmem83_io_pipeline_valid; // @[top.scala 596:22]
  wire [31:0] dmem83_io_pipeline_writedata; // @[top.scala 596:22]
  wire  dmem83_io_pipeline_memread; // @[top.scala 596:22]
  wire  dmem83_io_pipeline_memwrite; // @[top.scala 596:22]
  wire [1:0] dmem83_io_pipeline_maskmode; // @[top.scala 596:22]
  wire  dmem83_io_pipeline_sext; // @[top.scala 596:22]
  wire [31:0] dmem83_io_pipeline_readdata; // @[top.scala 596:22]
  wire  dmem83_io_bus_request_valid; // @[top.scala 596:22]
  wire [31:0] dmem83_io_bus_request_bits_address; // @[top.scala 596:22]
  wire [31:0] dmem83_io_bus_request_bits_writedata; // @[top.scala 596:22]
  wire [1:0] dmem83_io_bus_request_bits_operation; // @[top.scala 596:22]
  wire  dmem83_io_bus_response_valid; // @[top.scala 596:22]
  wire [31:0] dmem83_io_bus_response_bits_data; // @[top.scala 596:22]
  wire  cpu84_clock; // @[top.scala 600:21]
  wire  cpu84_reset; // @[top.scala 600:21]
  wire [31:0] cpu84_io_imem_address; // @[top.scala 600:21]
  wire [31:0] cpu84_io_imem_instruction; // @[top.scala 600:21]
  wire [31:0] cpu84_io_dmem_address; // @[top.scala 600:21]
  wire  cpu84_io_dmem_valid; // @[top.scala 600:21]
  wire [31:0] cpu84_io_dmem_writedata; // @[top.scala 600:21]
  wire  cpu84_io_dmem_memread; // @[top.scala 600:21]
  wire  cpu84_io_dmem_memwrite; // @[top.scala 600:21]
  wire [1:0] cpu84_io_dmem_maskmode; // @[top.scala 600:21]
  wire  cpu84_io_dmem_sext; // @[top.scala 600:21]
  wire [31:0] cpu84_io_dmem_readdata; // @[top.scala 600:21]
  wire  mem84_clock; // @[top.scala 601:21]
  wire  mem84_reset; // @[top.scala 601:21]
  wire [31:0] mem84_io_imem_request_bits_address; // @[top.scala 601:21]
  wire [31:0] mem84_io_imem_response_bits_data; // @[top.scala 601:21]
  wire  mem84_io_dmem_request_valid; // @[top.scala 601:21]
  wire [31:0] mem84_io_dmem_request_bits_address; // @[top.scala 601:21]
  wire [31:0] mem84_io_dmem_request_bits_writedata; // @[top.scala 601:21]
  wire [1:0] mem84_io_dmem_request_bits_operation; // @[top.scala 601:21]
  wire  mem84_io_dmem_response_valid; // @[top.scala 601:21]
  wire [31:0] mem84_io_dmem_response_bits_data; // @[top.scala 601:21]
  wire [31:0] imem84_io_pipeline_address; // @[top.scala 602:22]
  wire [31:0] imem84_io_pipeline_instruction; // @[top.scala 602:22]
  wire [31:0] imem84_io_bus_request_bits_address; // @[top.scala 602:22]
  wire [31:0] imem84_io_bus_response_bits_data; // @[top.scala 602:22]
  wire  dmem84_clock; // @[top.scala 603:22]
  wire  dmem84_reset; // @[top.scala 603:22]
  wire [31:0] dmem84_io_pipeline_address; // @[top.scala 603:22]
  wire  dmem84_io_pipeline_valid; // @[top.scala 603:22]
  wire [31:0] dmem84_io_pipeline_writedata; // @[top.scala 603:22]
  wire  dmem84_io_pipeline_memread; // @[top.scala 603:22]
  wire  dmem84_io_pipeline_memwrite; // @[top.scala 603:22]
  wire [1:0] dmem84_io_pipeline_maskmode; // @[top.scala 603:22]
  wire  dmem84_io_pipeline_sext; // @[top.scala 603:22]
  wire [31:0] dmem84_io_pipeline_readdata; // @[top.scala 603:22]
  wire  dmem84_io_bus_request_valid; // @[top.scala 603:22]
  wire [31:0] dmem84_io_bus_request_bits_address; // @[top.scala 603:22]
  wire [31:0] dmem84_io_bus_request_bits_writedata; // @[top.scala 603:22]
  wire [1:0] dmem84_io_bus_request_bits_operation; // @[top.scala 603:22]
  wire  dmem84_io_bus_response_valid; // @[top.scala 603:22]
  wire [31:0] dmem84_io_bus_response_bits_data; // @[top.scala 603:22]
  wire  cpu85_clock; // @[top.scala 607:21]
  wire  cpu85_reset; // @[top.scala 607:21]
  wire [31:0] cpu85_io_imem_address; // @[top.scala 607:21]
  wire [31:0] cpu85_io_imem_instruction; // @[top.scala 607:21]
  wire [31:0] cpu85_io_dmem_address; // @[top.scala 607:21]
  wire  cpu85_io_dmem_valid; // @[top.scala 607:21]
  wire [31:0] cpu85_io_dmem_writedata; // @[top.scala 607:21]
  wire  cpu85_io_dmem_memread; // @[top.scala 607:21]
  wire  cpu85_io_dmem_memwrite; // @[top.scala 607:21]
  wire [1:0] cpu85_io_dmem_maskmode; // @[top.scala 607:21]
  wire  cpu85_io_dmem_sext; // @[top.scala 607:21]
  wire [31:0] cpu85_io_dmem_readdata; // @[top.scala 607:21]
  wire  mem85_clock; // @[top.scala 608:21]
  wire  mem85_reset; // @[top.scala 608:21]
  wire [31:0] mem85_io_imem_request_bits_address; // @[top.scala 608:21]
  wire [31:0] mem85_io_imem_response_bits_data; // @[top.scala 608:21]
  wire  mem85_io_dmem_request_valid; // @[top.scala 608:21]
  wire [31:0] mem85_io_dmem_request_bits_address; // @[top.scala 608:21]
  wire [31:0] mem85_io_dmem_request_bits_writedata; // @[top.scala 608:21]
  wire [1:0] mem85_io_dmem_request_bits_operation; // @[top.scala 608:21]
  wire  mem85_io_dmem_response_valid; // @[top.scala 608:21]
  wire [31:0] mem85_io_dmem_response_bits_data; // @[top.scala 608:21]
  wire [31:0] imem85_io_pipeline_address; // @[top.scala 609:22]
  wire [31:0] imem85_io_pipeline_instruction; // @[top.scala 609:22]
  wire [31:0] imem85_io_bus_request_bits_address; // @[top.scala 609:22]
  wire [31:0] imem85_io_bus_response_bits_data; // @[top.scala 609:22]
  wire  dmem85_clock; // @[top.scala 610:22]
  wire  dmem85_reset; // @[top.scala 610:22]
  wire [31:0] dmem85_io_pipeline_address; // @[top.scala 610:22]
  wire  dmem85_io_pipeline_valid; // @[top.scala 610:22]
  wire [31:0] dmem85_io_pipeline_writedata; // @[top.scala 610:22]
  wire  dmem85_io_pipeline_memread; // @[top.scala 610:22]
  wire  dmem85_io_pipeline_memwrite; // @[top.scala 610:22]
  wire [1:0] dmem85_io_pipeline_maskmode; // @[top.scala 610:22]
  wire  dmem85_io_pipeline_sext; // @[top.scala 610:22]
  wire [31:0] dmem85_io_pipeline_readdata; // @[top.scala 610:22]
  wire  dmem85_io_bus_request_valid; // @[top.scala 610:22]
  wire [31:0] dmem85_io_bus_request_bits_address; // @[top.scala 610:22]
  wire [31:0] dmem85_io_bus_request_bits_writedata; // @[top.scala 610:22]
  wire [1:0] dmem85_io_bus_request_bits_operation; // @[top.scala 610:22]
  wire  dmem85_io_bus_response_valid; // @[top.scala 610:22]
  wire [31:0] dmem85_io_bus_response_bits_data; // @[top.scala 610:22]
  wire  cpu86_clock; // @[top.scala 614:21]
  wire  cpu86_reset; // @[top.scala 614:21]
  wire [31:0] cpu86_io_imem_address; // @[top.scala 614:21]
  wire [31:0] cpu86_io_imem_instruction; // @[top.scala 614:21]
  wire [31:0] cpu86_io_dmem_address; // @[top.scala 614:21]
  wire  cpu86_io_dmem_valid; // @[top.scala 614:21]
  wire [31:0] cpu86_io_dmem_writedata; // @[top.scala 614:21]
  wire  cpu86_io_dmem_memread; // @[top.scala 614:21]
  wire  cpu86_io_dmem_memwrite; // @[top.scala 614:21]
  wire [1:0] cpu86_io_dmem_maskmode; // @[top.scala 614:21]
  wire  cpu86_io_dmem_sext; // @[top.scala 614:21]
  wire [31:0] cpu86_io_dmem_readdata; // @[top.scala 614:21]
  wire  mem86_clock; // @[top.scala 615:21]
  wire  mem86_reset; // @[top.scala 615:21]
  wire [31:0] mem86_io_imem_request_bits_address; // @[top.scala 615:21]
  wire [31:0] mem86_io_imem_response_bits_data; // @[top.scala 615:21]
  wire  mem86_io_dmem_request_valid; // @[top.scala 615:21]
  wire [31:0] mem86_io_dmem_request_bits_address; // @[top.scala 615:21]
  wire [31:0] mem86_io_dmem_request_bits_writedata; // @[top.scala 615:21]
  wire [1:0] mem86_io_dmem_request_bits_operation; // @[top.scala 615:21]
  wire  mem86_io_dmem_response_valid; // @[top.scala 615:21]
  wire [31:0] mem86_io_dmem_response_bits_data; // @[top.scala 615:21]
  wire [31:0] imem86_io_pipeline_address; // @[top.scala 616:22]
  wire [31:0] imem86_io_pipeline_instruction; // @[top.scala 616:22]
  wire [31:0] imem86_io_bus_request_bits_address; // @[top.scala 616:22]
  wire [31:0] imem86_io_bus_response_bits_data; // @[top.scala 616:22]
  wire  dmem86_clock; // @[top.scala 617:22]
  wire  dmem86_reset; // @[top.scala 617:22]
  wire [31:0] dmem86_io_pipeline_address; // @[top.scala 617:22]
  wire  dmem86_io_pipeline_valid; // @[top.scala 617:22]
  wire [31:0] dmem86_io_pipeline_writedata; // @[top.scala 617:22]
  wire  dmem86_io_pipeline_memread; // @[top.scala 617:22]
  wire  dmem86_io_pipeline_memwrite; // @[top.scala 617:22]
  wire [1:0] dmem86_io_pipeline_maskmode; // @[top.scala 617:22]
  wire  dmem86_io_pipeline_sext; // @[top.scala 617:22]
  wire [31:0] dmem86_io_pipeline_readdata; // @[top.scala 617:22]
  wire  dmem86_io_bus_request_valid; // @[top.scala 617:22]
  wire [31:0] dmem86_io_bus_request_bits_address; // @[top.scala 617:22]
  wire [31:0] dmem86_io_bus_request_bits_writedata; // @[top.scala 617:22]
  wire [1:0] dmem86_io_bus_request_bits_operation; // @[top.scala 617:22]
  wire  dmem86_io_bus_response_valid; // @[top.scala 617:22]
  wire [31:0] dmem86_io_bus_response_bits_data; // @[top.scala 617:22]
  wire  cpu87_clock; // @[top.scala 621:21]
  wire  cpu87_reset; // @[top.scala 621:21]
  wire [31:0] cpu87_io_imem_address; // @[top.scala 621:21]
  wire [31:0] cpu87_io_imem_instruction; // @[top.scala 621:21]
  wire [31:0] cpu87_io_dmem_address; // @[top.scala 621:21]
  wire  cpu87_io_dmem_valid; // @[top.scala 621:21]
  wire [31:0] cpu87_io_dmem_writedata; // @[top.scala 621:21]
  wire  cpu87_io_dmem_memread; // @[top.scala 621:21]
  wire  cpu87_io_dmem_memwrite; // @[top.scala 621:21]
  wire [1:0] cpu87_io_dmem_maskmode; // @[top.scala 621:21]
  wire  cpu87_io_dmem_sext; // @[top.scala 621:21]
  wire [31:0] cpu87_io_dmem_readdata; // @[top.scala 621:21]
  wire  mem87_clock; // @[top.scala 622:21]
  wire  mem87_reset; // @[top.scala 622:21]
  wire [31:0] mem87_io_imem_request_bits_address; // @[top.scala 622:21]
  wire [31:0] mem87_io_imem_response_bits_data; // @[top.scala 622:21]
  wire  mem87_io_dmem_request_valid; // @[top.scala 622:21]
  wire [31:0] mem87_io_dmem_request_bits_address; // @[top.scala 622:21]
  wire [31:0] mem87_io_dmem_request_bits_writedata; // @[top.scala 622:21]
  wire [1:0] mem87_io_dmem_request_bits_operation; // @[top.scala 622:21]
  wire  mem87_io_dmem_response_valid; // @[top.scala 622:21]
  wire [31:0] mem87_io_dmem_response_bits_data; // @[top.scala 622:21]
  wire [31:0] imem87_io_pipeline_address; // @[top.scala 623:22]
  wire [31:0] imem87_io_pipeline_instruction; // @[top.scala 623:22]
  wire [31:0] imem87_io_bus_request_bits_address; // @[top.scala 623:22]
  wire [31:0] imem87_io_bus_response_bits_data; // @[top.scala 623:22]
  wire  dmem87_clock; // @[top.scala 624:22]
  wire  dmem87_reset; // @[top.scala 624:22]
  wire [31:0] dmem87_io_pipeline_address; // @[top.scala 624:22]
  wire  dmem87_io_pipeline_valid; // @[top.scala 624:22]
  wire [31:0] dmem87_io_pipeline_writedata; // @[top.scala 624:22]
  wire  dmem87_io_pipeline_memread; // @[top.scala 624:22]
  wire  dmem87_io_pipeline_memwrite; // @[top.scala 624:22]
  wire [1:0] dmem87_io_pipeline_maskmode; // @[top.scala 624:22]
  wire  dmem87_io_pipeline_sext; // @[top.scala 624:22]
  wire [31:0] dmem87_io_pipeline_readdata; // @[top.scala 624:22]
  wire  dmem87_io_bus_request_valid; // @[top.scala 624:22]
  wire [31:0] dmem87_io_bus_request_bits_address; // @[top.scala 624:22]
  wire [31:0] dmem87_io_bus_request_bits_writedata; // @[top.scala 624:22]
  wire [1:0] dmem87_io_bus_request_bits_operation; // @[top.scala 624:22]
  wire  dmem87_io_bus_response_valid; // @[top.scala 624:22]
  wire [31:0] dmem87_io_bus_response_bits_data; // @[top.scala 624:22]
  wire  cpu88_clock; // @[top.scala 628:21]
  wire  cpu88_reset; // @[top.scala 628:21]
  wire [31:0] cpu88_io_imem_address; // @[top.scala 628:21]
  wire [31:0] cpu88_io_imem_instruction; // @[top.scala 628:21]
  wire [31:0] cpu88_io_dmem_address; // @[top.scala 628:21]
  wire  cpu88_io_dmem_valid; // @[top.scala 628:21]
  wire [31:0] cpu88_io_dmem_writedata; // @[top.scala 628:21]
  wire  cpu88_io_dmem_memread; // @[top.scala 628:21]
  wire  cpu88_io_dmem_memwrite; // @[top.scala 628:21]
  wire [1:0] cpu88_io_dmem_maskmode; // @[top.scala 628:21]
  wire  cpu88_io_dmem_sext; // @[top.scala 628:21]
  wire [31:0] cpu88_io_dmem_readdata; // @[top.scala 628:21]
  wire  mem88_clock; // @[top.scala 629:21]
  wire  mem88_reset; // @[top.scala 629:21]
  wire [31:0] mem88_io_imem_request_bits_address; // @[top.scala 629:21]
  wire [31:0] mem88_io_imem_response_bits_data; // @[top.scala 629:21]
  wire  mem88_io_dmem_request_valid; // @[top.scala 629:21]
  wire [31:0] mem88_io_dmem_request_bits_address; // @[top.scala 629:21]
  wire [31:0] mem88_io_dmem_request_bits_writedata; // @[top.scala 629:21]
  wire [1:0] mem88_io_dmem_request_bits_operation; // @[top.scala 629:21]
  wire  mem88_io_dmem_response_valid; // @[top.scala 629:21]
  wire [31:0] mem88_io_dmem_response_bits_data; // @[top.scala 629:21]
  wire [31:0] imem88_io_pipeline_address; // @[top.scala 630:22]
  wire [31:0] imem88_io_pipeline_instruction; // @[top.scala 630:22]
  wire [31:0] imem88_io_bus_request_bits_address; // @[top.scala 630:22]
  wire [31:0] imem88_io_bus_response_bits_data; // @[top.scala 630:22]
  wire  dmem88_clock; // @[top.scala 631:22]
  wire  dmem88_reset; // @[top.scala 631:22]
  wire [31:0] dmem88_io_pipeline_address; // @[top.scala 631:22]
  wire  dmem88_io_pipeline_valid; // @[top.scala 631:22]
  wire [31:0] dmem88_io_pipeline_writedata; // @[top.scala 631:22]
  wire  dmem88_io_pipeline_memread; // @[top.scala 631:22]
  wire  dmem88_io_pipeline_memwrite; // @[top.scala 631:22]
  wire [1:0] dmem88_io_pipeline_maskmode; // @[top.scala 631:22]
  wire  dmem88_io_pipeline_sext; // @[top.scala 631:22]
  wire [31:0] dmem88_io_pipeline_readdata; // @[top.scala 631:22]
  wire  dmem88_io_bus_request_valid; // @[top.scala 631:22]
  wire [31:0] dmem88_io_bus_request_bits_address; // @[top.scala 631:22]
  wire [31:0] dmem88_io_bus_request_bits_writedata; // @[top.scala 631:22]
  wire [1:0] dmem88_io_bus_request_bits_operation; // @[top.scala 631:22]
  wire  dmem88_io_bus_response_valid; // @[top.scala 631:22]
  wire [31:0] dmem88_io_bus_response_bits_data; // @[top.scala 631:22]
  wire  cpu89_clock; // @[top.scala 635:21]
  wire  cpu89_reset; // @[top.scala 635:21]
  wire [31:0] cpu89_io_imem_address; // @[top.scala 635:21]
  wire [31:0] cpu89_io_imem_instruction; // @[top.scala 635:21]
  wire [31:0] cpu89_io_dmem_address; // @[top.scala 635:21]
  wire  cpu89_io_dmem_valid; // @[top.scala 635:21]
  wire [31:0] cpu89_io_dmem_writedata; // @[top.scala 635:21]
  wire  cpu89_io_dmem_memread; // @[top.scala 635:21]
  wire  cpu89_io_dmem_memwrite; // @[top.scala 635:21]
  wire [1:0] cpu89_io_dmem_maskmode; // @[top.scala 635:21]
  wire  cpu89_io_dmem_sext; // @[top.scala 635:21]
  wire [31:0] cpu89_io_dmem_readdata; // @[top.scala 635:21]
  wire  mem89_clock; // @[top.scala 636:21]
  wire  mem89_reset; // @[top.scala 636:21]
  wire [31:0] mem89_io_imem_request_bits_address; // @[top.scala 636:21]
  wire [31:0] mem89_io_imem_response_bits_data; // @[top.scala 636:21]
  wire  mem89_io_dmem_request_valid; // @[top.scala 636:21]
  wire [31:0] mem89_io_dmem_request_bits_address; // @[top.scala 636:21]
  wire [31:0] mem89_io_dmem_request_bits_writedata; // @[top.scala 636:21]
  wire [1:0] mem89_io_dmem_request_bits_operation; // @[top.scala 636:21]
  wire  mem89_io_dmem_response_valid; // @[top.scala 636:21]
  wire [31:0] mem89_io_dmem_response_bits_data; // @[top.scala 636:21]
  wire [31:0] imem89_io_pipeline_address; // @[top.scala 637:22]
  wire [31:0] imem89_io_pipeline_instruction; // @[top.scala 637:22]
  wire [31:0] imem89_io_bus_request_bits_address; // @[top.scala 637:22]
  wire [31:0] imem89_io_bus_response_bits_data; // @[top.scala 637:22]
  wire  dmem89_clock; // @[top.scala 638:22]
  wire  dmem89_reset; // @[top.scala 638:22]
  wire [31:0] dmem89_io_pipeline_address; // @[top.scala 638:22]
  wire  dmem89_io_pipeline_valid; // @[top.scala 638:22]
  wire [31:0] dmem89_io_pipeline_writedata; // @[top.scala 638:22]
  wire  dmem89_io_pipeline_memread; // @[top.scala 638:22]
  wire  dmem89_io_pipeline_memwrite; // @[top.scala 638:22]
  wire [1:0] dmem89_io_pipeline_maskmode; // @[top.scala 638:22]
  wire  dmem89_io_pipeline_sext; // @[top.scala 638:22]
  wire [31:0] dmem89_io_pipeline_readdata; // @[top.scala 638:22]
  wire  dmem89_io_bus_request_valid; // @[top.scala 638:22]
  wire [31:0] dmem89_io_bus_request_bits_address; // @[top.scala 638:22]
  wire [31:0] dmem89_io_bus_request_bits_writedata; // @[top.scala 638:22]
  wire [1:0] dmem89_io_bus_request_bits_operation; // @[top.scala 638:22]
  wire  dmem89_io_bus_response_valid; // @[top.scala 638:22]
  wire [31:0] dmem89_io_bus_response_bits_data; // @[top.scala 638:22]
  wire  cpu90_clock; // @[top.scala 642:21]
  wire  cpu90_reset; // @[top.scala 642:21]
  wire [31:0] cpu90_io_imem_address; // @[top.scala 642:21]
  wire [31:0] cpu90_io_imem_instruction; // @[top.scala 642:21]
  wire [31:0] cpu90_io_dmem_address; // @[top.scala 642:21]
  wire  cpu90_io_dmem_valid; // @[top.scala 642:21]
  wire [31:0] cpu90_io_dmem_writedata; // @[top.scala 642:21]
  wire  cpu90_io_dmem_memread; // @[top.scala 642:21]
  wire  cpu90_io_dmem_memwrite; // @[top.scala 642:21]
  wire [1:0] cpu90_io_dmem_maskmode; // @[top.scala 642:21]
  wire  cpu90_io_dmem_sext; // @[top.scala 642:21]
  wire [31:0] cpu90_io_dmem_readdata; // @[top.scala 642:21]
  wire  mem90_clock; // @[top.scala 643:21]
  wire  mem90_reset; // @[top.scala 643:21]
  wire [31:0] mem90_io_imem_request_bits_address; // @[top.scala 643:21]
  wire [31:0] mem90_io_imem_response_bits_data; // @[top.scala 643:21]
  wire  mem90_io_dmem_request_valid; // @[top.scala 643:21]
  wire [31:0] mem90_io_dmem_request_bits_address; // @[top.scala 643:21]
  wire [31:0] mem90_io_dmem_request_bits_writedata; // @[top.scala 643:21]
  wire [1:0] mem90_io_dmem_request_bits_operation; // @[top.scala 643:21]
  wire  mem90_io_dmem_response_valid; // @[top.scala 643:21]
  wire [31:0] mem90_io_dmem_response_bits_data; // @[top.scala 643:21]
  wire [31:0] imem90_io_pipeline_address; // @[top.scala 644:22]
  wire [31:0] imem90_io_pipeline_instruction; // @[top.scala 644:22]
  wire [31:0] imem90_io_bus_request_bits_address; // @[top.scala 644:22]
  wire [31:0] imem90_io_bus_response_bits_data; // @[top.scala 644:22]
  wire  dmem90_clock; // @[top.scala 645:22]
  wire  dmem90_reset; // @[top.scala 645:22]
  wire [31:0] dmem90_io_pipeline_address; // @[top.scala 645:22]
  wire  dmem90_io_pipeline_valid; // @[top.scala 645:22]
  wire [31:0] dmem90_io_pipeline_writedata; // @[top.scala 645:22]
  wire  dmem90_io_pipeline_memread; // @[top.scala 645:22]
  wire  dmem90_io_pipeline_memwrite; // @[top.scala 645:22]
  wire [1:0] dmem90_io_pipeline_maskmode; // @[top.scala 645:22]
  wire  dmem90_io_pipeline_sext; // @[top.scala 645:22]
  wire [31:0] dmem90_io_pipeline_readdata; // @[top.scala 645:22]
  wire  dmem90_io_bus_request_valid; // @[top.scala 645:22]
  wire [31:0] dmem90_io_bus_request_bits_address; // @[top.scala 645:22]
  wire [31:0] dmem90_io_bus_request_bits_writedata; // @[top.scala 645:22]
  wire [1:0] dmem90_io_bus_request_bits_operation; // @[top.scala 645:22]
  wire  dmem90_io_bus_response_valid; // @[top.scala 645:22]
  wire [31:0] dmem90_io_bus_response_bits_data; // @[top.scala 645:22]
  wire  cpu91_clock; // @[top.scala 649:21]
  wire  cpu91_reset; // @[top.scala 649:21]
  wire [31:0] cpu91_io_imem_address; // @[top.scala 649:21]
  wire [31:0] cpu91_io_imem_instruction; // @[top.scala 649:21]
  wire [31:0] cpu91_io_dmem_address; // @[top.scala 649:21]
  wire  cpu91_io_dmem_valid; // @[top.scala 649:21]
  wire [31:0] cpu91_io_dmem_writedata; // @[top.scala 649:21]
  wire  cpu91_io_dmem_memread; // @[top.scala 649:21]
  wire  cpu91_io_dmem_memwrite; // @[top.scala 649:21]
  wire [1:0] cpu91_io_dmem_maskmode; // @[top.scala 649:21]
  wire  cpu91_io_dmem_sext; // @[top.scala 649:21]
  wire [31:0] cpu91_io_dmem_readdata; // @[top.scala 649:21]
  wire  mem91_clock; // @[top.scala 650:21]
  wire  mem91_reset; // @[top.scala 650:21]
  wire [31:0] mem91_io_imem_request_bits_address; // @[top.scala 650:21]
  wire [31:0] mem91_io_imem_response_bits_data; // @[top.scala 650:21]
  wire  mem91_io_dmem_request_valid; // @[top.scala 650:21]
  wire [31:0] mem91_io_dmem_request_bits_address; // @[top.scala 650:21]
  wire [31:0] mem91_io_dmem_request_bits_writedata; // @[top.scala 650:21]
  wire [1:0] mem91_io_dmem_request_bits_operation; // @[top.scala 650:21]
  wire  mem91_io_dmem_response_valid; // @[top.scala 650:21]
  wire [31:0] mem91_io_dmem_response_bits_data; // @[top.scala 650:21]
  wire [31:0] imem91_io_pipeline_address; // @[top.scala 651:22]
  wire [31:0] imem91_io_pipeline_instruction; // @[top.scala 651:22]
  wire [31:0] imem91_io_bus_request_bits_address; // @[top.scala 651:22]
  wire [31:0] imem91_io_bus_response_bits_data; // @[top.scala 651:22]
  wire  dmem91_clock; // @[top.scala 652:22]
  wire  dmem91_reset; // @[top.scala 652:22]
  wire [31:0] dmem91_io_pipeline_address; // @[top.scala 652:22]
  wire  dmem91_io_pipeline_valid; // @[top.scala 652:22]
  wire [31:0] dmem91_io_pipeline_writedata; // @[top.scala 652:22]
  wire  dmem91_io_pipeline_memread; // @[top.scala 652:22]
  wire  dmem91_io_pipeline_memwrite; // @[top.scala 652:22]
  wire [1:0] dmem91_io_pipeline_maskmode; // @[top.scala 652:22]
  wire  dmem91_io_pipeline_sext; // @[top.scala 652:22]
  wire [31:0] dmem91_io_pipeline_readdata; // @[top.scala 652:22]
  wire  dmem91_io_bus_request_valid; // @[top.scala 652:22]
  wire [31:0] dmem91_io_bus_request_bits_address; // @[top.scala 652:22]
  wire [31:0] dmem91_io_bus_request_bits_writedata; // @[top.scala 652:22]
  wire [1:0] dmem91_io_bus_request_bits_operation; // @[top.scala 652:22]
  wire  dmem91_io_bus_response_valid; // @[top.scala 652:22]
  wire [31:0] dmem91_io_bus_response_bits_data; // @[top.scala 652:22]
  wire  cpu92_clock; // @[top.scala 656:21]
  wire  cpu92_reset; // @[top.scala 656:21]
  wire [31:0] cpu92_io_imem_address; // @[top.scala 656:21]
  wire [31:0] cpu92_io_imem_instruction; // @[top.scala 656:21]
  wire [31:0] cpu92_io_dmem_address; // @[top.scala 656:21]
  wire  cpu92_io_dmem_valid; // @[top.scala 656:21]
  wire [31:0] cpu92_io_dmem_writedata; // @[top.scala 656:21]
  wire  cpu92_io_dmem_memread; // @[top.scala 656:21]
  wire  cpu92_io_dmem_memwrite; // @[top.scala 656:21]
  wire [1:0] cpu92_io_dmem_maskmode; // @[top.scala 656:21]
  wire  cpu92_io_dmem_sext; // @[top.scala 656:21]
  wire [31:0] cpu92_io_dmem_readdata; // @[top.scala 656:21]
  wire  mem92_clock; // @[top.scala 657:21]
  wire  mem92_reset; // @[top.scala 657:21]
  wire [31:0] mem92_io_imem_request_bits_address; // @[top.scala 657:21]
  wire [31:0] mem92_io_imem_response_bits_data; // @[top.scala 657:21]
  wire  mem92_io_dmem_request_valid; // @[top.scala 657:21]
  wire [31:0] mem92_io_dmem_request_bits_address; // @[top.scala 657:21]
  wire [31:0] mem92_io_dmem_request_bits_writedata; // @[top.scala 657:21]
  wire [1:0] mem92_io_dmem_request_bits_operation; // @[top.scala 657:21]
  wire  mem92_io_dmem_response_valid; // @[top.scala 657:21]
  wire [31:0] mem92_io_dmem_response_bits_data; // @[top.scala 657:21]
  wire [31:0] imem92_io_pipeline_address; // @[top.scala 658:22]
  wire [31:0] imem92_io_pipeline_instruction; // @[top.scala 658:22]
  wire [31:0] imem92_io_bus_request_bits_address; // @[top.scala 658:22]
  wire [31:0] imem92_io_bus_response_bits_data; // @[top.scala 658:22]
  wire  dmem92_clock; // @[top.scala 659:22]
  wire  dmem92_reset; // @[top.scala 659:22]
  wire [31:0] dmem92_io_pipeline_address; // @[top.scala 659:22]
  wire  dmem92_io_pipeline_valid; // @[top.scala 659:22]
  wire [31:0] dmem92_io_pipeline_writedata; // @[top.scala 659:22]
  wire  dmem92_io_pipeline_memread; // @[top.scala 659:22]
  wire  dmem92_io_pipeline_memwrite; // @[top.scala 659:22]
  wire [1:0] dmem92_io_pipeline_maskmode; // @[top.scala 659:22]
  wire  dmem92_io_pipeline_sext; // @[top.scala 659:22]
  wire [31:0] dmem92_io_pipeline_readdata; // @[top.scala 659:22]
  wire  dmem92_io_bus_request_valid; // @[top.scala 659:22]
  wire [31:0] dmem92_io_bus_request_bits_address; // @[top.scala 659:22]
  wire [31:0] dmem92_io_bus_request_bits_writedata; // @[top.scala 659:22]
  wire [1:0] dmem92_io_bus_request_bits_operation; // @[top.scala 659:22]
  wire  dmem92_io_bus_response_valid; // @[top.scala 659:22]
  wire [31:0] dmem92_io_bus_response_bits_data; // @[top.scala 659:22]
  wire  cpu93_clock; // @[top.scala 663:21]
  wire  cpu93_reset; // @[top.scala 663:21]
  wire [31:0] cpu93_io_imem_address; // @[top.scala 663:21]
  wire [31:0] cpu93_io_imem_instruction; // @[top.scala 663:21]
  wire [31:0] cpu93_io_dmem_address; // @[top.scala 663:21]
  wire  cpu93_io_dmem_valid; // @[top.scala 663:21]
  wire [31:0] cpu93_io_dmem_writedata; // @[top.scala 663:21]
  wire  cpu93_io_dmem_memread; // @[top.scala 663:21]
  wire  cpu93_io_dmem_memwrite; // @[top.scala 663:21]
  wire [1:0] cpu93_io_dmem_maskmode; // @[top.scala 663:21]
  wire  cpu93_io_dmem_sext; // @[top.scala 663:21]
  wire [31:0] cpu93_io_dmem_readdata; // @[top.scala 663:21]
  wire  mem93_clock; // @[top.scala 664:21]
  wire  mem93_reset; // @[top.scala 664:21]
  wire [31:0] mem93_io_imem_request_bits_address; // @[top.scala 664:21]
  wire [31:0] mem93_io_imem_response_bits_data; // @[top.scala 664:21]
  wire  mem93_io_dmem_request_valid; // @[top.scala 664:21]
  wire [31:0] mem93_io_dmem_request_bits_address; // @[top.scala 664:21]
  wire [31:0] mem93_io_dmem_request_bits_writedata; // @[top.scala 664:21]
  wire [1:0] mem93_io_dmem_request_bits_operation; // @[top.scala 664:21]
  wire  mem93_io_dmem_response_valid; // @[top.scala 664:21]
  wire [31:0] mem93_io_dmem_response_bits_data; // @[top.scala 664:21]
  wire [31:0] imem93_io_pipeline_address; // @[top.scala 665:22]
  wire [31:0] imem93_io_pipeline_instruction; // @[top.scala 665:22]
  wire [31:0] imem93_io_bus_request_bits_address; // @[top.scala 665:22]
  wire [31:0] imem93_io_bus_response_bits_data; // @[top.scala 665:22]
  wire  dmem93_clock; // @[top.scala 666:22]
  wire  dmem93_reset; // @[top.scala 666:22]
  wire [31:0] dmem93_io_pipeline_address; // @[top.scala 666:22]
  wire  dmem93_io_pipeline_valid; // @[top.scala 666:22]
  wire [31:0] dmem93_io_pipeline_writedata; // @[top.scala 666:22]
  wire  dmem93_io_pipeline_memread; // @[top.scala 666:22]
  wire  dmem93_io_pipeline_memwrite; // @[top.scala 666:22]
  wire [1:0] dmem93_io_pipeline_maskmode; // @[top.scala 666:22]
  wire  dmem93_io_pipeline_sext; // @[top.scala 666:22]
  wire [31:0] dmem93_io_pipeline_readdata; // @[top.scala 666:22]
  wire  dmem93_io_bus_request_valid; // @[top.scala 666:22]
  wire [31:0] dmem93_io_bus_request_bits_address; // @[top.scala 666:22]
  wire [31:0] dmem93_io_bus_request_bits_writedata; // @[top.scala 666:22]
  wire [1:0] dmem93_io_bus_request_bits_operation; // @[top.scala 666:22]
  wire  dmem93_io_bus_response_valid; // @[top.scala 666:22]
  wire [31:0] dmem93_io_bus_response_bits_data; // @[top.scala 666:22]
  wire  cpu94_clock; // @[top.scala 670:21]
  wire  cpu94_reset; // @[top.scala 670:21]
  wire [31:0] cpu94_io_imem_address; // @[top.scala 670:21]
  wire [31:0] cpu94_io_imem_instruction; // @[top.scala 670:21]
  wire [31:0] cpu94_io_dmem_address; // @[top.scala 670:21]
  wire  cpu94_io_dmem_valid; // @[top.scala 670:21]
  wire [31:0] cpu94_io_dmem_writedata; // @[top.scala 670:21]
  wire  cpu94_io_dmem_memread; // @[top.scala 670:21]
  wire  cpu94_io_dmem_memwrite; // @[top.scala 670:21]
  wire [1:0] cpu94_io_dmem_maskmode; // @[top.scala 670:21]
  wire  cpu94_io_dmem_sext; // @[top.scala 670:21]
  wire [31:0] cpu94_io_dmem_readdata; // @[top.scala 670:21]
  wire  mem94_clock; // @[top.scala 671:21]
  wire  mem94_reset; // @[top.scala 671:21]
  wire [31:0] mem94_io_imem_request_bits_address; // @[top.scala 671:21]
  wire [31:0] mem94_io_imem_response_bits_data; // @[top.scala 671:21]
  wire  mem94_io_dmem_request_valid; // @[top.scala 671:21]
  wire [31:0] mem94_io_dmem_request_bits_address; // @[top.scala 671:21]
  wire [31:0] mem94_io_dmem_request_bits_writedata; // @[top.scala 671:21]
  wire [1:0] mem94_io_dmem_request_bits_operation; // @[top.scala 671:21]
  wire  mem94_io_dmem_response_valid; // @[top.scala 671:21]
  wire [31:0] mem94_io_dmem_response_bits_data; // @[top.scala 671:21]
  wire [31:0] imem94_io_pipeline_address; // @[top.scala 672:22]
  wire [31:0] imem94_io_pipeline_instruction; // @[top.scala 672:22]
  wire [31:0] imem94_io_bus_request_bits_address; // @[top.scala 672:22]
  wire [31:0] imem94_io_bus_response_bits_data; // @[top.scala 672:22]
  wire  dmem94_clock; // @[top.scala 673:22]
  wire  dmem94_reset; // @[top.scala 673:22]
  wire [31:0] dmem94_io_pipeline_address; // @[top.scala 673:22]
  wire  dmem94_io_pipeline_valid; // @[top.scala 673:22]
  wire [31:0] dmem94_io_pipeline_writedata; // @[top.scala 673:22]
  wire  dmem94_io_pipeline_memread; // @[top.scala 673:22]
  wire  dmem94_io_pipeline_memwrite; // @[top.scala 673:22]
  wire [1:0] dmem94_io_pipeline_maskmode; // @[top.scala 673:22]
  wire  dmem94_io_pipeline_sext; // @[top.scala 673:22]
  wire [31:0] dmem94_io_pipeline_readdata; // @[top.scala 673:22]
  wire  dmem94_io_bus_request_valid; // @[top.scala 673:22]
  wire [31:0] dmem94_io_bus_request_bits_address; // @[top.scala 673:22]
  wire [31:0] dmem94_io_bus_request_bits_writedata; // @[top.scala 673:22]
  wire [1:0] dmem94_io_bus_request_bits_operation; // @[top.scala 673:22]
  wire  dmem94_io_bus_response_valid; // @[top.scala 673:22]
  wire [31:0] dmem94_io_bus_response_bits_data; // @[top.scala 673:22]
  wire  cpu95_clock; // @[top.scala 677:21]
  wire  cpu95_reset; // @[top.scala 677:21]
  wire [31:0] cpu95_io_imem_address; // @[top.scala 677:21]
  wire [31:0] cpu95_io_imem_instruction; // @[top.scala 677:21]
  wire [31:0] cpu95_io_dmem_address; // @[top.scala 677:21]
  wire  cpu95_io_dmem_valid; // @[top.scala 677:21]
  wire [31:0] cpu95_io_dmem_writedata; // @[top.scala 677:21]
  wire  cpu95_io_dmem_memread; // @[top.scala 677:21]
  wire  cpu95_io_dmem_memwrite; // @[top.scala 677:21]
  wire [1:0] cpu95_io_dmem_maskmode; // @[top.scala 677:21]
  wire  cpu95_io_dmem_sext; // @[top.scala 677:21]
  wire [31:0] cpu95_io_dmem_readdata; // @[top.scala 677:21]
  wire  mem95_clock; // @[top.scala 678:21]
  wire  mem95_reset; // @[top.scala 678:21]
  wire [31:0] mem95_io_imem_request_bits_address; // @[top.scala 678:21]
  wire [31:0] mem95_io_imem_response_bits_data; // @[top.scala 678:21]
  wire  mem95_io_dmem_request_valid; // @[top.scala 678:21]
  wire [31:0] mem95_io_dmem_request_bits_address; // @[top.scala 678:21]
  wire [31:0] mem95_io_dmem_request_bits_writedata; // @[top.scala 678:21]
  wire [1:0] mem95_io_dmem_request_bits_operation; // @[top.scala 678:21]
  wire  mem95_io_dmem_response_valid; // @[top.scala 678:21]
  wire [31:0] mem95_io_dmem_response_bits_data; // @[top.scala 678:21]
  wire [31:0] imem95_io_pipeline_address; // @[top.scala 679:22]
  wire [31:0] imem95_io_pipeline_instruction; // @[top.scala 679:22]
  wire [31:0] imem95_io_bus_request_bits_address; // @[top.scala 679:22]
  wire [31:0] imem95_io_bus_response_bits_data; // @[top.scala 679:22]
  wire  dmem95_clock; // @[top.scala 680:22]
  wire  dmem95_reset; // @[top.scala 680:22]
  wire [31:0] dmem95_io_pipeline_address; // @[top.scala 680:22]
  wire  dmem95_io_pipeline_valid; // @[top.scala 680:22]
  wire [31:0] dmem95_io_pipeline_writedata; // @[top.scala 680:22]
  wire  dmem95_io_pipeline_memread; // @[top.scala 680:22]
  wire  dmem95_io_pipeline_memwrite; // @[top.scala 680:22]
  wire [1:0] dmem95_io_pipeline_maskmode; // @[top.scala 680:22]
  wire  dmem95_io_pipeline_sext; // @[top.scala 680:22]
  wire [31:0] dmem95_io_pipeline_readdata; // @[top.scala 680:22]
  wire  dmem95_io_bus_request_valid; // @[top.scala 680:22]
  wire [31:0] dmem95_io_bus_request_bits_address; // @[top.scala 680:22]
  wire [31:0] dmem95_io_bus_request_bits_writedata; // @[top.scala 680:22]
  wire [1:0] dmem95_io_bus_request_bits_operation; // @[top.scala 680:22]
  wire  dmem95_io_bus_response_valid; // @[top.scala 680:22]
  wire [31:0] dmem95_io_bus_response_bits_data; // @[top.scala 680:22]
  wire  cpu96_clock; // @[top.scala 684:21]
  wire  cpu96_reset; // @[top.scala 684:21]
  wire [31:0] cpu96_io_imem_address; // @[top.scala 684:21]
  wire [31:0] cpu96_io_imem_instruction; // @[top.scala 684:21]
  wire [31:0] cpu96_io_dmem_address; // @[top.scala 684:21]
  wire  cpu96_io_dmem_valid; // @[top.scala 684:21]
  wire [31:0] cpu96_io_dmem_writedata; // @[top.scala 684:21]
  wire  cpu96_io_dmem_memread; // @[top.scala 684:21]
  wire  cpu96_io_dmem_memwrite; // @[top.scala 684:21]
  wire [1:0] cpu96_io_dmem_maskmode; // @[top.scala 684:21]
  wire  cpu96_io_dmem_sext; // @[top.scala 684:21]
  wire [31:0] cpu96_io_dmem_readdata; // @[top.scala 684:21]
  wire  mem96_clock; // @[top.scala 685:21]
  wire  mem96_reset; // @[top.scala 685:21]
  wire [31:0] mem96_io_imem_request_bits_address; // @[top.scala 685:21]
  wire [31:0] mem96_io_imem_response_bits_data; // @[top.scala 685:21]
  wire  mem96_io_dmem_request_valid; // @[top.scala 685:21]
  wire [31:0] mem96_io_dmem_request_bits_address; // @[top.scala 685:21]
  wire [31:0] mem96_io_dmem_request_bits_writedata; // @[top.scala 685:21]
  wire [1:0] mem96_io_dmem_request_bits_operation; // @[top.scala 685:21]
  wire  mem96_io_dmem_response_valid; // @[top.scala 685:21]
  wire [31:0] mem96_io_dmem_response_bits_data; // @[top.scala 685:21]
  wire [31:0] imem96_io_pipeline_address; // @[top.scala 686:22]
  wire [31:0] imem96_io_pipeline_instruction; // @[top.scala 686:22]
  wire [31:0] imem96_io_bus_request_bits_address; // @[top.scala 686:22]
  wire [31:0] imem96_io_bus_response_bits_data; // @[top.scala 686:22]
  wire  dmem96_clock; // @[top.scala 687:22]
  wire  dmem96_reset; // @[top.scala 687:22]
  wire [31:0] dmem96_io_pipeline_address; // @[top.scala 687:22]
  wire  dmem96_io_pipeline_valid; // @[top.scala 687:22]
  wire [31:0] dmem96_io_pipeline_writedata; // @[top.scala 687:22]
  wire  dmem96_io_pipeline_memread; // @[top.scala 687:22]
  wire  dmem96_io_pipeline_memwrite; // @[top.scala 687:22]
  wire [1:0] dmem96_io_pipeline_maskmode; // @[top.scala 687:22]
  wire  dmem96_io_pipeline_sext; // @[top.scala 687:22]
  wire [31:0] dmem96_io_pipeline_readdata; // @[top.scala 687:22]
  wire  dmem96_io_bus_request_valid; // @[top.scala 687:22]
  wire [31:0] dmem96_io_bus_request_bits_address; // @[top.scala 687:22]
  wire [31:0] dmem96_io_bus_request_bits_writedata; // @[top.scala 687:22]
  wire [1:0] dmem96_io_bus_request_bits_operation; // @[top.scala 687:22]
  wire  dmem96_io_bus_response_valid; // @[top.scala 687:22]
  wire [31:0] dmem96_io_bus_response_bits_data; // @[top.scala 687:22]
  wire  cpu97_clock; // @[top.scala 691:21]
  wire  cpu97_reset; // @[top.scala 691:21]
  wire [31:0] cpu97_io_imem_address; // @[top.scala 691:21]
  wire [31:0] cpu97_io_imem_instruction; // @[top.scala 691:21]
  wire [31:0] cpu97_io_dmem_address; // @[top.scala 691:21]
  wire  cpu97_io_dmem_valid; // @[top.scala 691:21]
  wire [31:0] cpu97_io_dmem_writedata; // @[top.scala 691:21]
  wire  cpu97_io_dmem_memread; // @[top.scala 691:21]
  wire  cpu97_io_dmem_memwrite; // @[top.scala 691:21]
  wire [1:0] cpu97_io_dmem_maskmode; // @[top.scala 691:21]
  wire  cpu97_io_dmem_sext; // @[top.scala 691:21]
  wire [31:0] cpu97_io_dmem_readdata; // @[top.scala 691:21]
  wire  mem97_clock; // @[top.scala 692:21]
  wire  mem97_reset; // @[top.scala 692:21]
  wire [31:0] mem97_io_imem_request_bits_address; // @[top.scala 692:21]
  wire [31:0] mem97_io_imem_response_bits_data; // @[top.scala 692:21]
  wire  mem97_io_dmem_request_valid; // @[top.scala 692:21]
  wire [31:0] mem97_io_dmem_request_bits_address; // @[top.scala 692:21]
  wire [31:0] mem97_io_dmem_request_bits_writedata; // @[top.scala 692:21]
  wire [1:0] mem97_io_dmem_request_bits_operation; // @[top.scala 692:21]
  wire  mem97_io_dmem_response_valid; // @[top.scala 692:21]
  wire [31:0] mem97_io_dmem_response_bits_data; // @[top.scala 692:21]
  wire [31:0] imem97_io_pipeline_address; // @[top.scala 693:22]
  wire [31:0] imem97_io_pipeline_instruction; // @[top.scala 693:22]
  wire [31:0] imem97_io_bus_request_bits_address; // @[top.scala 693:22]
  wire [31:0] imem97_io_bus_response_bits_data; // @[top.scala 693:22]
  wire  dmem97_clock; // @[top.scala 694:22]
  wire  dmem97_reset; // @[top.scala 694:22]
  wire [31:0] dmem97_io_pipeline_address; // @[top.scala 694:22]
  wire  dmem97_io_pipeline_valid; // @[top.scala 694:22]
  wire [31:0] dmem97_io_pipeline_writedata; // @[top.scala 694:22]
  wire  dmem97_io_pipeline_memread; // @[top.scala 694:22]
  wire  dmem97_io_pipeline_memwrite; // @[top.scala 694:22]
  wire [1:0] dmem97_io_pipeline_maskmode; // @[top.scala 694:22]
  wire  dmem97_io_pipeline_sext; // @[top.scala 694:22]
  wire [31:0] dmem97_io_pipeline_readdata; // @[top.scala 694:22]
  wire  dmem97_io_bus_request_valid; // @[top.scala 694:22]
  wire [31:0] dmem97_io_bus_request_bits_address; // @[top.scala 694:22]
  wire [31:0] dmem97_io_bus_request_bits_writedata; // @[top.scala 694:22]
  wire [1:0] dmem97_io_bus_request_bits_operation; // @[top.scala 694:22]
  wire  dmem97_io_bus_response_valid; // @[top.scala 694:22]
  wire [31:0] dmem97_io_bus_response_bits_data; // @[top.scala 694:22]
  wire  cpu98_clock; // @[top.scala 698:21]
  wire  cpu98_reset; // @[top.scala 698:21]
  wire [31:0] cpu98_io_imem_address; // @[top.scala 698:21]
  wire [31:0] cpu98_io_imem_instruction; // @[top.scala 698:21]
  wire [31:0] cpu98_io_dmem_address; // @[top.scala 698:21]
  wire  cpu98_io_dmem_valid; // @[top.scala 698:21]
  wire [31:0] cpu98_io_dmem_writedata; // @[top.scala 698:21]
  wire  cpu98_io_dmem_memread; // @[top.scala 698:21]
  wire  cpu98_io_dmem_memwrite; // @[top.scala 698:21]
  wire [1:0] cpu98_io_dmem_maskmode; // @[top.scala 698:21]
  wire  cpu98_io_dmem_sext; // @[top.scala 698:21]
  wire [31:0] cpu98_io_dmem_readdata; // @[top.scala 698:21]
  wire  mem98_clock; // @[top.scala 699:21]
  wire  mem98_reset; // @[top.scala 699:21]
  wire [31:0] mem98_io_imem_request_bits_address; // @[top.scala 699:21]
  wire [31:0] mem98_io_imem_response_bits_data; // @[top.scala 699:21]
  wire  mem98_io_dmem_request_valid; // @[top.scala 699:21]
  wire [31:0] mem98_io_dmem_request_bits_address; // @[top.scala 699:21]
  wire [31:0] mem98_io_dmem_request_bits_writedata; // @[top.scala 699:21]
  wire [1:0] mem98_io_dmem_request_bits_operation; // @[top.scala 699:21]
  wire  mem98_io_dmem_response_valid; // @[top.scala 699:21]
  wire [31:0] mem98_io_dmem_response_bits_data; // @[top.scala 699:21]
  wire [31:0] imem98_io_pipeline_address; // @[top.scala 700:22]
  wire [31:0] imem98_io_pipeline_instruction; // @[top.scala 700:22]
  wire [31:0] imem98_io_bus_request_bits_address; // @[top.scala 700:22]
  wire [31:0] imem98_io_bus_response_bits_data; // @[top.scala 700:22]
  wire  dmem98_clock; // @[top.scala 701:22]
  wire  dmem98_reset; // @[top.scala 701:22]
  wire [31:0] dmem98_io_pipeline_address; // @[top.scala 701:22]
  wire  dmem98_io_pipeline_valid; // @[top.scala 701:22]
  wire [31:0] dmem98_io_pipeline_writedata; // @[top.scala 701:22]
  wire  dmem98_io_pipeline_memread; // @[top.scala 701:22]
  wire  dmem98_io_pipeline_memwrite; // @[top.scala 701:22]
  wire [1:0] dmem98_io_pipeline_maskmode; // @[top.scala 701:22]
  wire  dmem98_io_pipeline_sext; // @[top.scala 701:22]
  wire [31:0] dmem98_io_pipeline_readdata; // @[top.scala 701:22]
  wire  dmem98_io_bus_request_valid; // @[top.scala 701:22]
  wire [31:0] dmem98_io_bus_request_bits_address; // @[top.scala 701:22]
  wire [31:0] dmem98_io_bus_request_bits_writedata; // @[top.scala 701:22]
  wire [1:0] dmem98_io_bus_request_bits_operation; // @[top.scala 701:22]
  wire  dmem98_io_bus_response_valid; // @[top.scala 701:22]
  wire [31:0] dmem98_io_bus_response_bits_data; // @[top.scala 701:22]
  wire  cpu99_clock; // @[top.scala 705:21]
  wire  cpu99_reset; // @[top.scala 705:21]
  wire [31:0] cpu99_io_imem_address; // @[top.scala 705:21]
  wire [31:0] cpu99_io_imem_instruction; // @[top.scala 705:21]
  wire [31:0] cpu99_io_dmem_address; // @[top.scala 705:21]
  wire  cpu99_io_dmem_valid; // @[top.scala 705:21]
  wire [31:0] cpu99_io_dmem_writedata; // @[top.scala 705:21]
  wire  cpu99_io_dmem_memread; // @[top.scala 705:21]
  wire  cpu99_io_dmem_memwrite; // @[top.scala 705:21]
  wire [1:0] cpu99_io_dmem_maskmode; // @[top.scala 705:21]
  wire  cpu99_io_dmem_sext; // @[top.scala 705:21]
  wire [31:0] cpu99_io_dmem_readdata; // @[top.scala 705:21]
  wire  mem99_clock; // @[top.scala 706:21]
  wire  mem99_reset; // @[top.scala 706:21]
  wire [31:0] mem99_io_imem_request_bits_address; // @[top.scala 706:21]
  wire [31:0] mem99_io_imem_response_bits_data; // @[top.scala 706:21]
  wire  mem99_io_dmem_request_valid; // @[top.scala 706:21]
  wire [31:0] mem99_io_dmem_request_bits_address; // @[top.scala 706:21]
  wire [31:0] mem99_io_dmem_request_bits_writedata; // @[top.scala 706:21]
  wire [1:0] mem99_io_dmem_request_bits_operation; // @[top.scala 706:21]
  wire  mem99_io_dmem_response_valid; // @[top.scala 706:21]
  wire [31:0] mem99_io_dmem_response_bits_data; // @[top.scala 706:21]
  wire [31:0] imem99_io_pipeline_address; // @[top.scala 707:22]
  wire [31:0] imem99_io_pipeline_instruction; // @[top.scala 707:22]
  wire [31:0] imem99_io_bus_request_bits_address; // @[top.scala 707:22]
  wire [31:0] imem99_io_bus_response_bits_data; // @[top.scala 707:22]
  wire  dmem99_clock; // @[top.scala 708:22]
  wire  dmem99_reset; // @[top.scala 708:22]
  wire [31:0] dmem99_io_pipeline_address; // @[top.scala 708:22]
  wire  dmem99_io_pipeline_valid; // @[top.scala 708:22]
  wire [31:0] dmem99_io_pipeline_writedata; // @[top.scala 708:22]
  wire  dmem99_io_pipeline_memread; // @[top.scala 708:22]
  wire  dmem99_io_pipeline_memwrite; // @[top.scala 708:22]
  wire [1:0] dmem99_io_pipeline_maskmode; // @[top.scala 708:22]
  wire  dmem99_io_pipeline_sext; // @[top.scala 708:22]
  wire [31:0] dmem99_io_pipeline_readdata; // @[top.scala 708:22]
  wire  dmem99_io_bus_request_valid; // @[top.scala 708:22]
  wire [31:0] dmem99_io_bus_request_bits_address; // @[top.scala 708:22]
  wire [31:0] dmem99_io_bus_request_bits_writedata; // @[top.scala 708:22]
  wire [1:0] dmem99_io_bus_request_bits_operation; // @[top.scala 708:22]
  wire  dmem99_io_bus_response_valid; // @[top.scala 708:22]
  wire [31:0] dmem99_io_bus_response_bits_data; // @[top.scala 708:22]
  wire  cpu100_clock; // @[top.scala 712:22]
  wire  cpu100_reset; // @[top.scala 712:22]
  wire [31:0] cpu100_io_imem_address; // @[top.scala 712:22]
  wire [31:0] cpu100_io_imem_instruction; // @[top.scala 712:22]
  wire [31:0] cpu100_io_dmem_address; // @[top.scala 712:22]
  wire  cpu100_io_dmem_valid; // @[top.scala 712:22]
  wire [31:0] cpu100_io_dmem_writedata; // @[top.scala 712:22]
  wire  cpu100_io_dmem_memread; // @[top.scala 712:22]
  wire  cpu100_io_dmem_memwrite; // @[top.scala 712:22]
  wire [1:0] cpu100_io_dmem_maskmode; // @[top.scala 712:22]
  wire  cpu100_io_dmem_sext; // @[top.scala 712:22]
  wire [31:0] cpu100_io_dmem_readdata; // @[top.scala 712:22]
  wire  mem100_clock; // @[top.scala 713:22]
  wire  mem100_reset; // @[top.scala 713:22]
  wire [31:0] mem100_io_imem_request_bits_address; // @[top.scala 713:22]
  wire [31:0] mem100_io_imem_response_bits_data; // @[top.scala 713:22]
  wire  mem100_io_dmem_request_valid; // @[top.scala 713:22]
  wire [31:0] mem100_io_dmem_request_bits_address; // @[top.scala 713:22]
  wire [31:0] mem100_io_dmem_request_bits_writedata; // @[top.scala 713:22]
  wire [1:0] mem100_io_dmem_request_bits_operation; // @[top.scala 713:22]
  wire  mem100_io_dmem_response_valid; // @[top.scala 713:22]
  wire [31:0] mem100_io_dmem_response_bits_data; // @[top.scala 713:22]
  wire [31:0] imem100_io_pipeline_address; // @[top.scala 714:23]
  wire [31:0] imem100_io_pipeline_instruction; // @[top.scala 714:23]
  wire [31:0] imem100_io_bus_request_bits_address; // @[top.scala 714:23]
  wire [31:0] imem100_io_bus_response_bits_data; // @[top.scala 714:23]
  wire  dmem100_clock; // @[top.scala 715:23]
  wire  dmem100_reset; // @[top.scala 715:23]
  wire [31:0] dmem100_io_pipeline_address; // @[top.scala 715:23]
  wire  dmem100_io_pipeline_valid; // @[top.scala 715:23]
  wire [31:0] dmem100_io_pipeline_writedata; // @[top.scala 715:23]
  wire  dmem100_io_pipeline_memread; // @[top.scala 715:23]
  wire  dmem100_io_pipeline_memwrite; // @[top.scala 715:23]
  wire [1:0] dmem100_io_pipeline_maskmode; // @[top.scala 715:23]
  wire  dmem100_io_pipeline_sext; // @[top.scala 715:23]
  wire [31:0] dmem100_io_pipeline_readdata; // @[top.scala 715:23]
  wire  dmem100_io_bus_request_valid; // @[top.scala 715:23]
  wire [31:0] dmem100_io_bus_request_bits_address; // @[top.scala 715:23]
  wire [31:0] dmem100_io_bus_request_bits_writedata; // @[top.scala 715:23]
  wire [1:0] dmem100_io_bus_request_bits_operation; // @[top.scala 715:23]
  wire  dmem100_io_bus_response_valid; // @[top.scala 715:23]
  wire [31:0] dmem100_io_bus_response_bits_data; // @[top.scala 715:23]
  wire  cpu101_clock; // @[top.scala 719:22]
  wire  cpu101_reset; // @[top.scala 719:22]
  wire [31:0] cpu101_io_imem_address; // @[top.scala 719:22]
  wire [31:0] cpu101_io_imem_instruction; // @[top.scala 719:22]
  wire [31:0] cpu101_io_dmem_address; // @[top.scala 719:22]
  wire  cpu101_io_dmem_valid; // @[top.scala 719:22]
  wire [31:0] cpu101_io_dmem_writedata; // @[top.scala 719:22]
  wire  cpu101_io_dmem_memread; // @[top.scala 719:22]
  wire  cpu101_io_dmem_memwrite; // @[top.scala 719:22]
  wire [1:0] cpu101_io_dmem_maskmode; // @[top.scala 719:22]
  wire  cpu101_io_dmem_sext; // @[top.scala 719:22]
  wire [31:0] cpu101_io_dmem_readdata; // @[top.scala 719:22]
  wire  mem101_clock; // @[top.scala 720:22]
  wire  mem101_reset; // @[top.scala 720:22]
  wire [31:0] mem101_io_imem_request_bits_address; // @[top.scala 720:22]
  wire [31:0] mem101_io_imem_response_bits_data; // @[top.scala 720:22]
  wire  mem101_io_dmem_request_valid; // @[top.scala 720:22]
  wire [31:0] mem101_io_dmem_request_bits_address; // @[top.scala 720:22]
  wire [31:0] mem101_io_dmem_request_bits_writedata; // @[top.scala 720:22]
  wire [1:0] mem101_io_dmem_request_bits_operation; // @[top.scala 720:22]
  wire  mem101_io_dmem_response_valid; // @[top.scala 720:22]
  wire [31:0] mem101_io_dmem_response_bits_data; // @[top.scala 720:22]
  wire [31:0] imem101_io_pipeline_address; // @[top.scala 721:23]
  wire [31:0] imem101_io_pipeline_instruction; // @[top.scala 721:23]
  wire [31:0] imem101_io_bus_request_bits_address; // @[top.scala 721:23]
  wire [31:0] imem101_io_bus_response_bits_data; // @[top.scala 721:23]
  wire  dmem101_clock; // @[top.scala 722:23]
  wire  dmem101_reset; // @[top.scala 722:23]
  wire [31:0] dmem101_io_pipeline_address; // @[top.scala 722:23]
  wire  dmem101_io_pipeline_valid; // @[top.scala 722:23]
  wire [31:0] dmem101_io_pipeline_writedata; // @[top.scala 722:23]
  wire  dmem101_io_pipeline_memread; // @[top.scala 722:23]
  wire  dmem101_io_pipeline_memwrite; // @[top.scala 722:23]
  wire [1:0] dmem101_io_pipeline_maskmode; // @[top.scala 722:23]
  wire  dmem101_io_pipeline_sext; // @[top.scala 722:23]
  wire [31:0] dmem101_io_pipeline_readdata; // @[top.scala 722:23]
  wire  dmem101_io_bus_request_valid; // @[top.scala 722:23]
  wire [31:0] dmem101_io_bus_request_bits_address; // @[top.scala 722:23]
  wire [31:0] dmem101_io_bus_request_bits_writedata; // @[top.scala 722:23]
  wire [1:0] dmem101_io_bus_request_bits_operation; // @[top.scala 722:23]
  wire  dmem101_io_bus_response_valid; // @[top.scala 722:23]
  wire [31:0] dmem101_io_bus_response_bits_data; // @[top.scala 722:23]
  wire  cpu102_clock; // @[top.scala 726:22]
  wire  cpu102_reset; // @[top.scala 726:22]
  wire [31:0] cpu102_io_imem_address; // @[top.scala 726:22]
  wire [31:0] cpu102_io_imem_instruction; // @[top.scala 726:22]
  wire [31:0] cpu102_io_dmem_address; // @[top.scala 726:22]
  wire  cpu102_io_dmem_valid; // @[top.scala 726:22]
  wire [31:0] cpu102_io_dmem_writedata; // @[top.scala 726:22]
  wire  cpu102_io_dmem_memread; // @[top.scala 726:22]
  wire  cpu102_io_dmem_memwrite; // @[top.scala 726:22]
  wire [1:0] cpu102_io_dmem_maskmode; // @[top.scala 726:22]
  wire  cpu102_io_dmem_sext; // @[top.scala 726:22]
  wire [31:0] cpu102_io_dmem_readdata; // @[top.scala 726:22]
  wire  mem102_clock; // @[top.scala 727:22]
  wire  mem102_reset; // @[top.scala 727:22]
  wire [31:0] mem102_io_imem_request_bits_address; // @[top.scala 727:22]
  wire [31:0] mem102_io_imem_response_bits_data; // @[top.scala 727:22]
  wire  mem102_io_dmem_request_valid; // @[top.scala 727:22]
  wire [31:0] mem102_io_dmem_request_bits_address; // @[top.scala 727:22]
  wire [31:0] mem102_io_dmem_request_bits_writedata; // @[top.scala 727:22]
  wire [1:0] mem102_io_dmem_request_bits_operation; // @[top.scala 727:22]
  wire  mem102_io_dmem_response_valid; // @[top.scala 727:22]
  wire [31:0] mem102_io_dmem_response_bits_data; // @[top.scala 727:22]
  wire [31:0] imem102_io_pipeline_address; // @[top.scala 728:23]
  wire [31:0] imem102_io_pipeline_instruction; // @[top.scala 728:23]
  wire [31:0] imem102_io_bus_request_bits_address; // @[top.scala 728:23]
  wire [31:0] imem102_io_bus_response_bits_data; // @[top.scala 728:23]
  wire  dmem102_clock; // @[top.scala 729:23]
  wire  dmem102_reset; // @[top.scala 729:23]
  wire [31:0] dmem102_io_pipeline_address; // @[top.scala 729:23]
  wire  dmem102_io_pipeline_valid; // @[top.scala 729:23]
  wire [31:0] dmem102_io_pipeline_writedata; // @[top.scala 729:23]
  wire  dmem102_io_pipeline_memread; // @[top.scala 729:23]
  wire  dmem102_io_pipeline_memwrite; // @[top.scala 729:23]
  wire [1:0] dmem102_io_pipeline_maskmode; // @[top.scala 729:23]
  wire  dmem102_io_pipeline_sext; // @[top.scala 729:23]
  wire [31:0] dmem102_io_pipeline_readdata; // @[top.scala 729:23]
  wire  dmem102_io_bus_request_valid; // @[top.scala 729:23]
  wire [31:0] dmem102_io_bus_request_bits_address; // @[top.scala 729:23]
  wire [31:0] dmem102_io_bus_request_bits_writedata; // @[top.scala 729:23]
  wire [1:0] dmem102_io_bus_request_bits_operation; // @[top.scala 729:23]
  wire  dmem102_io_bus_response_valid; // @[top.scala 729:23]
  wire [31:0] dmem102_io_bus_response_bits_data; // @[top.scala 729:23]
  wire  cpu103_clock; // @[top.scala 733:22]
  wire  cpu103_reset; // @[top.scala 733:22]
  wire [31:0] cpu103_io_imem_address; // @[top.scala 733:22]
  wire [31:0] cpu103_io_imem_instruction; // @[top.scala 733:22]
  wire [31:0] cpu103_io_dmem_address; // @[top.scala 733:22]
  wire  cpu103_io_dmem_valid; // @[top.scala 733:22]
  wire [31:0] cpu103_io_dmem_writedata; // @[top.scala 733:22]
  wire  cpu103_io_dmem_memread; // @[top.scala 733:22]
  wire  cpu103_io_dmem_memwrite; // @[top.scala 733:22]
  wire [1:0] cpu103_io_dmem_maskmode; // @[top.scala 733:22]
  wire  cpu103_io_dmem_sext; // @[top.scala 733:22]
  wire [31:0] cpu103_io_dmem_readdata; // @[top.scala 733:22]
  wire  mem103_clock; // @[top.scala 734:22]
  wire  mem103_reset; // @[top.scala 734:22]
  wire [31:0] mem103_io_imem_request_bits_address; // @[top.scala 734:22]
  wire [31:0] mem103_io_imem_response_bits_data; // @[top.scala 734:22]
  wire  mem103_io_dmem_request_valid; // @[top.scala 734:22]
  wire [31:0] mem103_io_dmem_request_bits_address; // @[top.scala 734:22]
  wire [31:0] mem103_io_dmem_request_bits_writedata; // @[top.scala 734:22]
  wire [1:0] mem103_io_dmem_request_bits_operation; // @[top.scala 734:22]
  wire  mem103_io_dmem_response_valid; // @[top.scala 734:22]
  wire [31:0] mem103_io_dmem_response_bits_data; // @[top.scala 734:22]
  wire [31:0] imem103_io_pipeline_address; // @[top.scala 735:23]
  wire [31:0] imem103_io_pipeline_instruction; // @[top.scala 735:23]
  wire [31:0] imem103_io_bus_request_bits_address; // @[top.scala 735:23]
  wire [31:0] imem103_io_bus_response_bits_data; // @[top.scala 735:23]
  wire  dmem103_clock; // @[top.scala 736:23]
  wire  dmem103_reset; // @[top.scala 736:23]
  wire [31:0] dmem103_io_pipeline_address; // @[top.scala 736:23]
  wire  dmem103_io_pipeline_valid; // @[top.scala 736:23]
  wire [31:0] dmem103_io_pipeline_writedata; // @[top.scala 736:23]
  wire  dmem103_io_pipeline_memread; // @[top.scala 736:23]
  wire  dmem103_io_pipeline_memwrite; // @[top.scala 736:23]
  wire [1:0] dmem103_io_pipeline_maskmode; // @[top.scala 736:23]
  wire  dmem103_io_pipeline_sext; // @[top.scala 736:23]
  wire [31:0] dmem103_io_pipeline_readdata; // @[top.scala 736:23]
  wire  dmem103_io_bus_request_valid; // @[top.scala 736:23]
  wire [31:0] dmem103_io_bus_request_bits_address; // @[top.scala 736:23]
  wire [31:0] dmem103_io_bus_request_bits_writedata; // @[top.scala 736:23]
  wire [1:0] dmem103_io_bus_request_bits_operation; // @[top.scala 736:23]
  wire  dmem103_io_bus_response_valid; // @[top.scala 736:23]
  wire [31:0] dmem103_io_bus_response_bits_data; // @[top.scala 736:23]
  wire  cpu104_clock; // @[top.scala 740:22]
  wire  cpu104_reset; // @[top.scala 740:22]
  wire [31:0] cpu104_io_imem_address; // @[top.scala 740:22]
  wire [31:0] cpu104_io_imem_instruction; // @[top.scala 740:22]
  wire [31:0] cpu104_io_dmem_address; // @[top.scala 740:22]
  wire  cpu104_io_dmem_valid; // @[top.scala 740:22]
  wire [31:0] cpu104_io_dmem_writedata; // @[top.scala 740:22]
  wire  cpu104_io_dmem_memread; // @[top.scala 740:22]
  wire  cpu104_io_dmem_memwrite; // @[top.scala 740:22]
  wire [1:0] cpu104_io_dmem_maskmode; // @[top.scala 740:22]
  wire  cpu104_io_dmem_sext; // @[top.scala 740:22]
  wire [31:0] cpu104_io_dmem_readdata; // @[top.scala 740:22]
  wire  mem104_clock; // @[top.scala 741:22]
  wire  mem104_reset; // @[top.scala 741:22]
  wire [31:0] mem104_io_imem_request_bits_address; // @[top.scala 741:22]
  wire [31:0] mem104_io_imem_response_bits_data; // @[top.scala 741:22]
  wire  mem104_io_dmem_request_valid; // @[top.scala 741:22]
  wire [31:0] mem104_io_dmem_request_bits_address; // @[top.scala 741:22]
  wire [31:0] mem104_io_dmem_request_bits_writedata; // @[top.scala 741:22]
  wire [1:0] mem104_io_dmem_request_bits_operation; // @[top.scala 741:22]
  wire  mem104_io_dmem_response_valid; // @[top.scala 741:22]
  wire [31:0] mem104_io_dmem_response_bits_data; // @[top.scala 741:22]
  wire [31:0] imem104_io_pipeline_address; // @[top.scala 742:23]
  wire [31:0] imem104_io_pipeline_instruction; // @[top.scala 742:23]
  wire [31:0] imem104_io_bus_request_bits_address; // @[top.scala 742:23]
  wire [31:0] imem104_io_bus_response_bits_data; // @[top.scala 742:23]
  wire  dmem104_clock; // @[top.scala 743:23]
  wire  dmem104_reset; // @[top.scala 743:23]
  wire [31:0] dmem104_io_pipeline_address; // @[top.scala 743:23]
  wire  dmem104_io_pipeline_valid; // @[top.scala 743:23]
  wire [31:0] dmem104_io_pipeline_writedata; // @[top.scala 743:23]
  wire  dmem104_io_pipeline_memread; // @[top.scala 743:23]
  wire  dmem104_io_pipeline_memwrite; // @[top.scala 743:23]
  wire [1:0] dmem104_io_pipeline_maskmode; // @[top.scala 743:23]
  wire  dmem104_io_pipeline_sext; // @[top.scala 743:23]
  wire [31:0] dmem104_io_pipeline_readdata; // @[top.scala 743:23]
  wire  dmem104_io_bus_request_valid; // @[top.scala 743:23]
  wire [31:0] dmem104_io_bus_request_bits_address; // @[top.scala 743:23]
  wire [31:0] dmem104_io_bus_request_bits_writedata; // @[top.scala 743:23]
  wire [1:0] dmem104_io_bus_request_bits_operation; // @[top.scala 743:23]
  wire  dmem104_io_bus_response_valid; // @[top.scala 743:23]
  wire [31:0] dmem104_io_bus_response_bits_data; // @[top.scala 743:23]
  wire  cpu105_clock; // @[top.scala 747:22]
  wire  cpu105_reset; // @[top.scala 747:22]
  wire [31:0] cpu105_io_imem_address; // @[top.scala 747:22]
  wire [31:0] cpu105_io_imem_instruction; // @[top.scala 747:22]
  wire [31:0] cpu105_io_dmem_address; // @[top.scala 747:22]
  wire  cpu105_io_dmem_valid; // @[top.scala 747:22]
  wire [31:0] cpu105_io_dmem_writedata; // @[top.scala 747:22]
  wire  cpu105_io_dmem_memread; // @[top.scala 747:22]
  wire  cpu105_io_dmem_memwrite; // @[top.scala 747:22]
  wire [1:0] cpu105_io_dmem_maskmode; // @[top.scala 747:22]
  wire  cpu105_io_dmem_sext; // @[top.scala 747:22]
  wire [31:0] cpu105_io_dmem_readdata; // @[top.scala 747:22]
  wire  mem105_clock; // @[top.scala 748:22]
  wire  mem105_reset; // @[top.scala 748:22]
  wire [31:0] mem105_io_imem_request_bits_address; // @[top.scala 748:22]
  wire [31:0] mem105_io_imem_response_bits_data; // @[top.scala 748:22]
  wire  mem105_io_dmem_request_valid; // @[top.scala 748:22]
  wire [31:0] mem105_io_dmem_request_bits_address; // @[top.scala 748:22]
  wire [31:0] mem105_io_dmem_request_bits_writedata; // @[top.scala 748:22]
  wire [1:0] mem105_io_dmem_request_bits_operation; // @[top.scala 748:22]
  wire  mem105_io_dmem_response_valid; // @[top.scala 748:22]
  wire [31:0] mem105_io_dmem_response_bits_data; // @[top.scala 748:22]
  wire [31:0] imem105_io_pipeline_address; // @[top.scala 749:23]
  wire [31:0] imem105_io_pipeline_instruction; // @[top.scala 749:23]
  wire [31:0] imem105_io_bus_request_bits_address; // @[top.scala 749:23]
  wire [31:0] imem105_io_bus_response_bits_data; // @[top.scala 749:23]
  wire  dmem105_clock; // @[top.scala 750:23]
  wire  dmem105_reset; // @[top.scala 750:23]
  wire [31:0] dmem105_io_pipeline_address; // @[top.scala 750:23]
  wire  dmem105_io_pipeline_valid; // @[top.scala 750:23]
  wire [31:0] dmem105_io_pipeline_writedata; // @[top.scala 750:23]
  wire  dmem105_io_pipeline_memread; // @[top.scala 750:23]
  wire  dmem105_io_pipeline_memwrite; // @[top.scala 750:23]
  wire [1:0] dmem105_io_pipeline_maskmode; // @[top.scala 750:23]
  wire  dmem105_io_pipeline_sext; // @[top.scala 750:23]
  wire [31:0] dmem105_io_pipeline_readdata; // @[top.scala 750:23]
  wire  dmem105_io_bus_request_valid; // @[top.scala 750:23]
  wire [31:0] dmem105_io_bus_request_bits_address; // @[top.scala 750:23]
  wire [31:0] dmem105_io_bus_request_bits_writedata; // @[top.scala 750:23]
  wire [1:0] dmem105_io_bus_request_bits_operation; // @[top.scala 750:23]
  wire  dmem105_io_bus_response_valid; // @[top.scala 750:23]
  wire [31:0] dmem105_io_bus_response_bits_data; // @[top.scala 750:23]
  wire  cpu106_clock; // @[top.scala 754:22]
  wire  cpu106_reset; // @[top.scala 754:22]
  wire [31:0] cpu106_io_imem_address; // @[top.scala 754:22]
  wire [31:0] cpu106_io_imem_instruction; // @[top.scala 754:22]
  wire [31:0] cpu106_io_dmem_address; // @[top.scala 754:22]
  wire  cpu106_io_dmem_valid; // @[top.scala 754:22]
  wire [31:0] cpu106_io_dmem_writedata; // @[top.scala 754:22]
  wire  cpu106_io_dmem_memread; // @[top.scala 754:22]
  wire  cpu106_io_dmem_memwrite; // @[top.scala 754:22]
  wire [1:0] cpu106_io_dmem_maskmode; // @[top.scala 754:22]
  wire  cpu106_io_dmem_sext; // @[top.scala 754:22]
  wire [31:0] cpu106_io_dmem_readdata; // @[top.scala 754:22]
  wire  mem106_clock; // @[top.scala 755:22]
  wire  mem106_reset; // @[top.scala 755:22]
  wire [31:0] mem106_io_imem_request_bits_address; // @[top.scala 755:22]
  wire [31:0] mem106_io_imem_response_bits_data; // @[top.scala 755:22]
  wire  mem106_io_dmem_request_valid; // @[top.scala 755:22]
  wire [31:0] mem106_io_dmem_request_bits_address; // @[top.scala 755:22]
  wire [31:0] mem106_io_dmem_request_bits_writedata; // @[top.scala 755:22]
  wire [1:0] mem106_io_dmem_request_bits_operation; // @[top.scala 755:22]
  wire  mem106_io_dmem_response_valid; // @[top.scala 755:22]
  wire [31:0] mem106_io_dmem_response_bits_data; // @[top.scala 755:22]
  wire [31:0] imem106_io_pipeline_address; // @[top.scala 756:23]
  wire [31:0] imem106_io_pipeline_instruction; // @[top.scala 756:23]
  wire [31:0] imem106_io_bus_request_bits_address; // @[top.scala 756:23]
  wire [31:0] imem106_io_bus_response_bits_data; // @[top.scala 756:23]
  wire  dmem106_clock; // @[top.scala 757:23]
  wire  dmem106_reset; // @[top.scala 757:23]
  wire [31:0] dmem106_io_pipeline_address; // @[top.scala 757:23]
  wire  dmem106_io_pipeline_valid; // @[top.scala 757:23]
  wire [31:0] dmem106_io_pipeline_writedata; // @[top.scala 757:23]
  wire  dmem106_io_pipeline_memread; // @[top.scala 757:23]
  wire  dmem106_io_pipeline_memwrite; // @[top.scala 757:23]
  wire [1:0] dmem106_io_pipeline_maskmode; // @[top.scala 757:23]
  wire  dmem106_io_pipeline_sext; // @[top.scala 757:23]
  wire [31:0] dmem106_io_pipeline_readdata; // @[top.scala 757:23]
  wire  dmem106_io_bus_request_valid; // @[top.scala 757:23]
  wire [31:0] dmem106_io_bus_request_bits_address; // @[top.scala 757:23]
  wire [31:0] dmem106_io_bus_request_bits_writedata; // @[top.scala 757:23]
  wire [1:0] dmem106_io_bus_request_bits_operation; // @[top.scala 757:23]
  wire  dmem106_io_bus_response_valid; // @[top.scala 757:23]
  wire [31:0] dmem106_io_bus_response_bits_data; // @[top.scala 757:23]
  wire  cpu107_clock; // @[top.scala 761:22]
  wire  cpu107_reset; // @[top.scala 761:22]
  wire [31:0] cpu107_io_imem_address; // @[top.scala 761:22]
  wire [31:0] cpu107_io_imem_instruction; // @[top.scala 761:22]
  wire [31:0] cpu107_io_dmem_address; // @[top.scala 761:22]
  wire  cpu107_io_dmem_valid; // @[top.scala 761:22]
  wire [31:0] cpu107_io_dmem_writedata; // @[top.scala 761:22]
  wire  cpu107_io_dmem_memread; // @[top.scala 761:22]
  wire  cpu107_io_dmem_memwrite; // @[top.scala 761:22]
  wire [1:0] cpu107_io_dmem_maskmode; // @[top.scala 761:22]
  wire  cpu107_io_dmem_sext; // @[top.scala 761:22]
  wire [31:0] cpu107_io_dmem_readdata; // @[top.scala 761:22]
  wire  mem107_clock; // @[top.scala 762:22]
  wire  mem107_reset; // @[top.scala 762:22]
  wire [31:0] mem107_io_imem_request_bits_address; // @[top.scala 762:22]
  wire [31:0] mem107_io_imem_response_bits_data; // @[top.scala 762:22]
  wire  mem107_io_dmem_request_valid; // @[top.scala 762:22]
  wire [31:0] mem107_io_dmem_request_bits_address; // @[top.scala 762:22]
  wire [31:0] mem107_io_dmem_request_bits_writedata; // @[top.scala 762:22]
  wire [1:0] mem107_io_dmem_request_bits_operation; // @[top.scala 762:22]
  wire  mem107_io_dmem_response_valid; // @[top.scala 762:22]
  wire [31:0] mem107_io_dmem_response_bits_data; // @[top.scala 762:22]
  wire [31:0] imem107_io_pipeline_address; // @[top.scala 763:23]
  wire [31:0] imem107_io_pipeline_instruction; // @[top.scala 763:23]
  wire [31:0] imem107_io_bus_request_bits_address; // @[top.scala 763:23]
  wire [31:0] imem107_io_bus_response_bits_data; // @[top.scala 763:23]
  wire  dmem107_clock; // @[top.scala 764:23]
  wire  dmem107_reset; // @[top.scala 764:23]
  wire [31:0] dmem107_io_pipeline_address; // @[top.scala 764:23]
  wire  dmem107_io_pipeline_valid; // @[top.scala 764:23]
  wire [31:0] dmem107_io_pipeline_writedata; // @[top.scala 764:23]
  wire  dmem107_io_pipeline_memread; // @[top.scala 764:23]
  wire  dmem107_io_pipeline_memwrite; // @[top.scala 764:23]
  wire [1:0] dmem107_io_pipeline_maskmode; // @[top.scala 764:23]
  wire  dmem107_io_pipeline_sext; // @[top.scala 764:23]
  wire [31:0] dmem107_io_pipeline_readdata; // @[top.scala 764:23]
  wire  dmem107_io_bus_request_valid; // @[top.scala 764:23]
  wire [31:0] dmem107_io_bus_request_bits_address; // @[top.scala 764:23]
  wire [31:0] dmem107_io_bus_request_bits_writedata; // @[top.scala 764:23]
  wire [1:0] dmem107_io_bus_request_bits_operation; // @[top.scala 764:23]
  wire  dmem107_io_bus_response_valid; // @[top.scala 764:23]
  wire [31:0] dmem107_io_bus_response_bits_data; // @[top.scala 764:23]
  wire  cpu108_clock; // @[top.scala 768:22]
  wire  cpu108_reset; // @[top.scala 768:22]
  wire [31:0] cpu108_io_imem_address; // @[top.scala 768:22]
  wire [31:0] cpu108_io_imem_instruction; // @[top.scala 768:22]
  wire [31:0] cpu108_io_dmem_address; // @[top.scala 768:22]
  wire  cpu108_io_dmem_valid; // @[top.scala 768:22]
  wire [31:0] cpu108_io_dmem_writedata; // @[top.scala 768:22]
  wire  cpu108_io_dmem_memread; // @[top.scala 768:22]
  wire  cpu108_io_dmem_memwrite; // @[top.scala 768:22]
  wire [1:0] cpu108_io_dmem_maskmode; // @[top.scala 768:22]
  wire  cpu108_io_dmem_sext; // @[top.scala 768:22]
  wire [31:0] cpu108_io_dmem_readdata; // @[top.scala 768:22]
  wire  mem108_clock; // @[top.scala 769:22]
  wire  mem108_reset; // @[top.scala 769:22]
  wire [31:0] mem108_io_imem_request_bits_address; // @[top.scala 769:22]
  wire [31:0] mem108_io_imem_response_bits_data; // @[top.scala 769:22]
  wire  mem108_io_dmem_request_valid; // @[top.scala 769:22]
  wire [31:0] mem108_io_dmem_request_bits_address; // @[top.scala 769:22]
  wire [31:0] mem108_io_dmem_request_bits_writedata; // @[top.scala 769:22]
  wire [1:0] mem108_io_dmem_request_bits_operation; // @[top.scala 769:22]
  wire  mem108_io_dmem_response_valid; // @[top.scala 769:22]
  wire [31:0] mem108_io_dmem_response_bits_data; // @[top.scala 769:22]
  wire [31:0] imem108_io_pipeline_address; // @[top.scala 770:23]
  wire [31:0] imem108_io_pipeline_instruction; // @[top.scala 770:23]
  wire [31:0] imem108_io_bus_request_bits_address; // @[top.scala 770:23]
  wire [31:0] imem108_io_bus_response_bits_data; // @[top.scala 770:23]
  wire  dmem108_clock; // @[top.scala 771:23]
  wire  dmem108_reset; // @[top.scala 771:23]
  wire [31:0] dmem108_io_pipeline_address; // @[top.scala 771:23]
  wire  dmem108_io_pipeline_valid; // @[top.scala 771:23]
  wire [31:0] dmem108_io_pipeline_writedata; // @[top.scala 771:23]
  wire  dmem108_io_pipeline_memread; // @[top.scala 771:23]
  wire  dmem108_io_pipeline_memwrite; // @[top.scala 771:23]
  wire [1:0] dmem108_io_pipeline_maskmode; // @[top.scala 771:23]
  wire  dmem108_io_pipeline_sext; // @[top.scala 771:23]
  wire [31:0] dmem108_io_pipeline_readdata; // @[top.scala 771:23]
  wire  dmem108_io_bus_request_valid; // @[top.scala 771:23]
  wire [31:0] dmem108_io_bus_request_bits_address; // @[top.scala 771:23]
  wire [31:0] dmem108_io_bus_request_bits_writedata; // @[top.scala 771:23]
  wire [1:0] dmem108_io_bus_request_bits_operation; // @[top.scala 771:23]
  wire  dmem108_io_bus_response_valid; // @[top.scala 771:23]
  wire [31:0] dmem108_io_bus_response_bits_data; // @[top.scala 771:23]
  wire  cpu109_clock; // @[top.scala 775:22]
  wire  cpu109_reset; // @[top.scala 775:22]
  wire [31:0] cpu109_io_imem_address; // @[top.scala 775:22]
  wire [31:0] cpu109_io_imem_instruction; // @[top.scala 775:22]
  wire [31:0] cpu109_io_dmem_address; // @[top.scala 775:22]
  wire  cpu109_io_dmem_valid; // @[top.scala 775:22]
  wire [31:0] cpu109_io_dmem_writedata; // @[top.scala 775:22]
  wire  cpu109_io_dmem_memread; // @[top.scala 775:22]
  wire  cpu109_io_dmem_memwrite; // @[top.scala 775:22]
  wire [1:0] cpu109_io_dmem_maskmode; // @[top.scala 775:22]
  wire  cpu109_io_dmem_sext; // @[top.scala 775:22]
  wire [31:0] cpu109_io_dmem_readdata; // @[top.scala 775:22]
  wire  mem109_clock; // @[top.scala 776:22]
  wire  mem109_reset; // @[top.scala 776:22]
  wire [31:0] mem109_io_imem_request_bits_address; // @[top.scala 776:22]
  wire [31:0] mem109_io_imem_response_bits_data; // @[top.scala 776:22]
  wire  mem109_io_dmem_request_valid; // @[top.scala 776:22]
  wire [31:0] mem109_io_dmem_request_bits_address; // @[top.scala 776:22]
  wire [31:0] mem109_io_dmem_request_bits_writedata; // @[top.scala 776:22]
  wire [1:0] mem109_io_dmem_request_bits_operation; // @[top.scala 776:22]
  wire  mem109_io_dmem_response_valid; // @[top.scala 776:22]
  wire [31:0] mem109_io_dmem_response_bits_data; // @[top.scala 776:22]
  wire [31:0] imem109_io_pipeline_address; // @[top.scala 777:23]
  wire [31:0] imem109_io_pipeline_instruction; // @[top.scala 777:23]
  wire [31:0] imem109_io_bus_request_bits_address; // @[top.scala 777:23]
  wire [31:0] imem109_io_bus_response_bits_data; // @[top.scala 777:23]
  wire  dmem109_clock; // @[top.scala 778:23]
  wire  dmem109_reset; // @[top.scala 778:23]
  wire [31:0] dmem109_io_pipeline_address; // @[top.scala 778:23]
  wire  dmem109_io_pipeline_valid; // @[top.scala 778:23]
  wire [31:0] dmem109_io_pipeline_writedata; // @[top.scala 778:23]
  wire  dmem109_io_pipeline_memread; // @[top.scala 778:23]
  wire  dmem109_io_pipeline_memwrite; // @[top.scala 778:23]
  wire [1:0] dmem109_io_pipeline_maskmode; // @[top.scala 778:23]
  wire  dmem109_io_pipeline_sext; // @[top.scala 778:23]
  wire [31:0] dmem109_io_pipeline_readdata; // @[top.scala 778:23]
  wire  dmem109_io_bus_request_valid; // @[top.scala 778:23]
  wire [31:0] dmem109_io_bus_request_bits_address; // @[top.scala 778:23]
  wire [31:0] dmem109_io_bus_request_bits_writedata; // @[top.scala 778:23]
  wire [1:0] dmem109_io_bus_request_bits_operation; // @[top.scala 778:23]
  wire  dmem109_io_bus_response_valid; // @[top.scala 778:23]
  wire [31:0] dmem109_io_bus_response_bits_data; // @[top.scala 778:23]
  wire  cpu110_clock; // @[top.scala 782:22]
  wire  cpu110_reset; // @[top.scala 782:22]
  wire [31:0] cpu110_io_imem_address; // @[top.scala 782:22]
  wire [31:0] cpu110_io_imem_instruction; // @[top.scala 782:22]
  wire [31:0] cpu110_io_dmem_address; // @[top.scala 782:22]
  wire  cpu110_io_dmem_valid; // @[top.scala 782:22]
  wire [31:0] cpu110_io_dmem_writedata; // @[top.scala 782:22]
  wire  cpu110_io_dmem_memread; // @[top.scala 782:22]
  wire  cpu110_io_dmem_memwrite; // @[top.scala 782:22]
  wire [1:0] cpu110_io_dmem_maskmode; // @[top.scala 782:22]
  wire  cpu110_io_dmem_sext; // @[top.scala 782:22]
  wire [31:0] cpu110_io_dmem_readdata; // @[top.scala 782:22]
  wire  mem110_clock; // @[top.scala 783:22]
  wire  mem110_reset; // @[top.scala 783:22]
  wire [31:0] mem110_io_imem_request_bits_address; // @[top.scala 783:22]
  wire [31:0] mem110_io_imem_response_bits_data; // @[top.scala 783:22]
  wire  mem110_io_dmem_request_valid; // @[top.scala 783:22]
  wire [31:0] mem110_io_dmem_request_bits_address; // @[top.scala 783:22]
  wire [31:0] mem110_io_dmem_request_bits_writedata; // @[top.scala 783:22]
  wire [1:0] mem110_io_dmem_request_bits_operation; // @[top.scala 783:22]
  wire  mem110_io_dmem_response_valid; // @[top.scala 783:22]
  wire [31:0] mem110_io_dmem_response_bits_data; // @[top.scala 783:22]
  wire [31:0] imem110_io_pipeline_address; // @[top.scala 784:23]
  wire [31:0] imem110_io_pipeline_instruction; // @[top.scala 784:23]
  wire [31:0] imem110_io_bus_request_bits_address; // @[top.scala 784:23]
  wire [31:0] imem110_io_bus_response_bits_data; // @[top.scala 784:23]
  wire  dmem110_clock; // @[top.scala 785:23]
  wire  dmem110_reset; // @[top.scala 785:23]
  wire [31:0] dmem110_io_pipeline_address; // @[top.scala 785:23]
  wire  dmem110_io_pipeline_valid; // @[top.scala 785:23]
  wire [31:0] dmem110_io_pipeline_writedata; // @[top.scala 785:23]
  wire  dmem110_io_pipeline_memread; // @[top.scala 785:23]
  wire  dmem110_io_pipeline_memwrite; // @[top.scala 785:23]
  wire [1:0] dmem110_io_pipeline_maskmode; // @[top.scala 785:23]
  wire  dmem110_io_pipeline_sext; // @[top.scala 785:23]
  wire [31:0] dmem110_io_pipeline_readdata; // @[top.scala 785:23]
  wire  dmem110_io_bus_request_valid; // @[top.scala 785:23]
  wire [31:0] dmem110_io_bus_request_bits_address; // @[top.scala 785:23]
  wire [31:0] dmem110_io_bus_request_bits_writedata; // @[top.scala 785:23]
  wire [1:0] dmem110_io_bus_request_bits_operation; // @[top.scala 785:23]
  wire  dmem110_io_bus_response_valid; // @[top.scala 785:23]
  wire [31:0] dmem110_io_bus_response_bits_data; // @[top.scala 785:23]
  wire  cpu111_clock; // @[top.scala 789:22]
  wire  cpu111_reset; // @[top.scala 789:22]
  wire [31:0] cpu111_io_imem_address; // @[top.scala 789:22]
  wire [31:0] cpu111_io_imem_instruction; // @[top.scala 789:22]
  wire [31:0] cpu111_io_dmem_address; // @[top.scala 789:22]
  wire  cpu111_io_dmem_valid; // @[top.scala 789:22]
  wire [31:0] cpu111_io_dmem_writedata; // @[top.scala 789:22]
  wire  cpu111_io_dmem_memread; // @[top.scala 789:22]
  wire  cpu111_io_dmem_memwrite; // @[top.scala 789:22]
  wire [1:0] cpu111_io_dmem_maskmode; // @[top.scala 789:22]
  wire  cpu111_io_dmem_sext; // @[top.scala 789:22]
  wire [31:0] cpu111_io_dmem_readdata; // @[top.scala 789:22]
  wire  mem111_clock; // @[top.scala 790:22]
  wire  mem111_reset; // @[top.scala 790:22]
  wire [31:0] mem111_io_imem_request_bits_address; // @[top.scala 790:22]
  wire [31:0] mem111_io_imem_response_bits_data; // @[top.scala 790:22]
  wire  mem111_io_dmem_request_valid; // @[top.scala 790:22]
  wire [31:0] mem111_io_dmem_request_bits_address; // @[top.scala 790:22]
  wire [31:0] mem111_io_dmem_request_bits_writedata; // @[top.scala 790:22]
  wire [1:0] mem111_io_dmem_request_bits_operation; // @[top.scala 790:22]
  wire  mem111_io_dmem_response_valid; // @[top.scala 790:22]
  wire [31:0] mem111_io_dmem_response_bits_data; // @[top.scala 790:22]
  wire [31:0] imem111_io_pipeline_address; // @[top.scala 791:23]
  wire [31:0] imem111_io_pipeline_instruction; // @[top.scala 791:23]
  wire [31:0] imem111_io_bus_request_bits_address; // @[top.scala 791:23]
  wire [31:0] imem111_io_bus_response_bits_data; // @[top.scala 791:23]
  wire  dmem111_clock; // @[top.scala 792:23]
  wire  dmem111_reset; // @[top.scala 792:23]
  wire [31:0] dmem111_io_pipeline_address; // @[top.scala 792:23]
  wire  dmem111_io_pipeline_valid; // @[top.scala 792:23]
  wire [31:0] dmem111_io_pipeline_writedata; // @[top.scala 792:23]
  wire  dmem111_io_pipeline_memread; // @[top.scala 792:23]
  wire  dmem111_io_pipeline_memwrite; // @[top.scala 792:23]
  wire [1:0] dmem111_io_pipeline_maskmode; // @[top.scala 792:23]
  wire  dmem111_io_pipeline_sext; // @[top.scala 792:23]
  wire [31:0] dmem111_io_pipeline_readdata; // @[top.scala 792:23]
  wire  dmem111_io_bus_request_valid; // @[top.scala 792:23]
  wire [31:0] dmem111_io_bus_request_bits_address; // @[top.scala 792:23]
  wire [31:0] dmem111_io_bus_request_bits_writedata; // @[top.scala 792:23]
  wire [1:0] dmem111_io_bus_request_bits_operation; // @[top.scala 792:23]
  wire  dmem111_io_bus_response_valid; // @[top.scala 792:23]
  wire [31:0] dmem111_io_bus_response_bits_data; // @[top.scala 792:23]
  wire  cpu112_clock; // @[top.scala 796:22]
  wire  cpu112_reset; // @[top.scala 796:22]
  wire [31:0] cpu112_io_imem_address; // @[top.scala 796:22]
  wire [31:0] cpu112_io_imem_instruction; // @[top.scala 796:22]
  wire [31:0] cpu112_io_dmem_address; // @[top.scala 796:22]
  wire  cpu112_io_dmem_valid; // @[top.scala 796:22]
  wire [31:0] cpu112_io_dmem_writedata; // @[top.scala 796:22]
  wire  cpu112_io_dmem_memread; // @[top.scala 796:22]
  wire  cpu112_io_dmem_memwrite; // @[top.scala 796:22]
  wire [1:0] cpu112_io_dmem_maskmode; // @[top.scala 796:22]
  wire  cpu112_io_dmem_sext; // @[top.scala 796:22]
  wire [31:0] cpu112_io_dmem_readdata; // @[top.scala 796:22]
  wire  mem112_clock; // @[top.scala 797:22]
  wire  mem112_reset; // @[top.scala 797:22]
  wire [31:0] mem112_io_imem_request_bits_address; // @[top.scala 797:22]
  wire [31:0] mem112_io_imem_response_bits_data; // @[top.scala 797:22]
  wire  mem112_io_dmem_request_valid; // @[top.scala 797:22]
  wire [31:0] mem112_io_dmem_request_bits_address; // @[top.scala 797:22]
  wire [31:0] mem112_io_dmem_request_bits_writedata; // @[top.scala 797:22]
  wire [1:0] mem112_io_dmem_request_bits_operation; // @[top.scala 797:22]
  wire  mem112_io_dmem_response_valid; // @[top.scala 797:22]
  wire [31:0] mem112_io_dmem_response_bits_data; // @[top.scala 797:22]
  wire [31:0] imem112_io_pipeline_address; // @[top.scala 798:23]
  wire [31:0] imem112_io_pipeline_instruction; // @[top.scala 798:23]
  wire [31:0] imem112_io_bus_request_bits_address; // @[top.scala 798:23]
  wire [31:0] imem112_io_bus_response_bits_data; // @[top.scala 798:23]
  wire  dmem112_clock; // @[top.scala 799:23]
  wire  dmem112_reset; // @[top.scala 799:23]
  wire [31:0] dmem112_io_pipeline_address; // @[top.scala 799:23]
  wire  dmem112_io_pipeline_valid; // @[top.scala 799:23]
  wire [31:0] dmem112_io_pipeline_writedata; // @[top.scala 799:23]
  wire  dmem112_io_pipeline_memread; // @[top.scala 799:23]
  wire  dmem112_io_pipeline_memwrite; // @[top.scala 799:23]
  wire [1:0] dmem112_io_pipeline_maskmode; // @[top.scala 799:23]
  wire  dmem112_io_pipeline_sext; // @[top.scala 799:23]
  wire [31:0] dmem112_io_pipeline_readdata; // @[top.scala 799:23]
  wire  dmem112_io_bus_request_valid; // @[top.scala 799:23]
  wire [31:0] dmem112_io_bus_request_bits_address; // @[top.scala 799:23]
  wire [31:0] dmem112_io_bus_request_bits_writedata; // @[top.scala 799:23]
  wire [1:0] dmem112_io_bus_request_bits_operation; // @[top.scala 799:23]
  wire  dmem112_io_bus_response_valid; // @[top.scala 799:23]
  wire [31:0] dmem112_io_bus_response_bits_data; // @[top.scala 799:23]
  wire  cpu113_clock; // @[top.scala 803:22]
  wire  cpu113_reset; // @[top.scala 803:22]
  wire [31:0] cpu113_io_imem_address; // @[top.scala 803:22]
  wire [31:0] cpu113_io_imem_instruction; // @[top.scala 803:22]
  wire [31:0] cpu113_io_dmem_address; // @[top.scala 803:22]
  wire  cpu113_io_dmem_valid; // @[top.scala 803:22]
  wire [31:0] cpu113_io_dmem_writedata; // @[top.scala 803:22]
  wire  cpu113_io_dmem_memread; // @[top.scala 803:22]
  wire  cpu113_io_dmem_memwrite; // @[top.scala 803:22]
  wire [1:0] cpu113_io_dmem_maskmode; // @[top.scala 803:22]
  wire  cpu113_io_dmem_sext; // @[top.scala 803:22]
  wire [31:0] cpu113_io_dmem_readdata; // @[top.scala 803:22]
  wire  mem113_clock; // @[top.scala 804:22]
  wire  mem113_reset; // @[top.scala 804:22]
  wire [31:0] mem113_io_imem_request_bits_address; // @[top.scala 804:22]
  wire [31:0] mem113_io_imem_response_bits_data; // @[top.scala 804:22]
  wire  mem113_io_dmem_request_valid; // @[top.scala 804:22]
  wire [31:0] mem113_io_dmem_request_bits_address; // @[top.scala 804:22]
  wire [31:0] mem113_io_dmem_request_bits_writedata; // @[top.scala 804:22]
  wire [1:0] mem113_io_dmem_request_bits_operation; // @[top.scala 804:22]
  wire  mem113_io_dmem_response_valid; // @[top.scala 804:22]
  wire [31:0] mem113_io_dmem_response_bits_data; // @[top.scala 804:22]
  wire [31:0] imem113_io_pipeline_address; // @[top.scala 805:23]
  wire [31:0] imem113_io_pipeline_instruction; // @[top.scala 805:23]
  wire [31:0] imem113_io_bus_request_bits_address; // @[top.scala 805:23]
  wire [31:0] imem113_io_bus_response_bits_data; // @[top.scala 805:23]
  wire  dmem113_clock; // @[top.scala 806:23]
  wire  dmem113_reset; // @[top.scala 806:23]
  wire [31:0] dmem113_io_pipeline_address; // @[top.scala 806:23]
  wire  dmem113_io_pipeline_valid; // @[top.scala 806:23]
  wire [31:0] dmem113_io_pipeline_writedata; // @[top.scala 806:23]
  wire  dmem113_io_pipeline_memread; // @[top.scala 806:23]
  wire  dmem113_io_pipeline_memwrite; // @[top.scala 806:23]
  wire [1:0] dmem113_io_pipeline_maskmode; // @[top.scala 806:23]
  wire  dmem113_io_pipeline_sext; // @[top.scala 806:23]
  wire [31:0] dmem113_io_pipeline_readdata; // @[top.scala 806:23]
  wire  dmem113_io_bus_request_valid; // @[top.scala 806:23]
  wire [31:0] dmem113_io_bus_request_bits_address; // @[top.scala 806:23]
  wire [31:0] dmem113_io_bus_request_bits_writedata; // @[top.scala 806:23]
  wire [1:0] dmem113_io_bus_request_bits_operation; // @[top.scala 806:23]
  wire  dmem113_io_bus_response_valid; // @[top.scala 806:23]
  wire [31:0] dmem113_io_bus_response_bits_data; // @[top.scala 806:23]
  wire  cpu114_clock; // @[top.scala 810:22]
  wire  cpu114_reset; // @[top.scala 810:22]
  wire [31:0] cpu114_io_imem_address; // @[top.scala 810:22]
  wire [31:0] cpu114_io_imem_instruction; // @[top.scala 810:22]
  wire [31:0] cpu114_io_dmem_address; // @[top.scala 810:22]
  wire  cpu114_io_dmem_valid; // @[top.scala 810:22]
  wire [31:0] cpu114_io_dmem_writedata; // @[top.scala 810:22]
  wire  cpu114_io_dmem_memread; // @[top.scala 810:22]
  wire  cpu114_io_dmem_memwrite; // @[top.scala 810:22]
  wire [1:0] cpu114_io_dmem_maskmode; // @[top.scala 810:22]
  wire  cpu114_io_dmem_sext; // @[top.scala 810:22]
  wire [31:0] cpu114_io_dmem_readdata; // @[top.scala 810:22]
  wire  mem114_clock; // @[top.scala 811:22]
  wire  mem114_reset; // @[top.scala 811:22]
  wire [31:0] mem114_io_imem_request_bits_address; // @[top.scala 811:22]
  wire [31:0] mem114_io_imem_response_bits_data; // @[top.scala 811:22]
  wire  mem114_io_dmem_request_valid; // @[top.scala 811:22]
  wire [31:0] mem114_io_dmem_request_bits_address; // @[top.scala 811:22]
  wire [31:0] mem114_io_dmem_request_bits_writedata; // @[top.scala 811:22]
  wire [1:0] mem114_io_dmem_request_bits_operation; // @[top.scala 811:22]
  wire  mem114_io_dmem_response_valid; // @[top.scala 811:22]
  wire [31:0] mem114_io_dmem_response_bits_data; // @[top.scala 811:22]
  wire [31:0] imem114_io_pipeline_address; // @[top.scala 812:23]
  wire [31:0] imem114_io_pipeline_instruction; // @[top.scala 812:23]
  wire [31:0] imem114_io_bus_request_bits_address; // @[top.scala 812:23]
  wire [31:0] imem114_io_bus_response_bits_data; // @[top.scala 812:23]
  wire  dmem114_clock; // @[top.scala 813:23]
  wire  dmem114_reset; // @[top.scala 813:23]
  wire [31:0] dmem114_io_pipeline_address; // @[top.scala 813:23]
  wire  dmem114_io_pipeline_valid; // @[top.scala 813:23]
  wire [31:0] dmem114_io_pipeline_writedata; // @[top.scala 813:23]
  wire  dmem114_io_pipeline_memread; // @[top.scala 813:23]
  wire  dmem114_io_pipeline_memwrite; // @[top.scala 813:23]
  wire [1:0] dmem114_io_pipeline_maskmode; // @[top.scala 813:23]
  wire  dmem114_io_pipeline_sext; // @[top.scala 813:23]
  wire [31:0] dmem114_io_pipeline_readdata; // @[top.scala 813:23]
  wire  dmem114_io_bus_request_valid; // @[top.scala 813:23]
  wire [31:0] dmem114_io_bus_request_bits_address; // @[top.scala 813:23]
  wire [31:0] dmem114_io_bus_request_bits_writedata; // @[top.scala 813:23]
  wire [1:0] dmem114_io_bus_request_bits_operation; // @[top.scala 813:23]
  wire  dmem114_io_bus_response_valid; // @[top.scala 813:23]
  wire [31:0] dmem114_io_bus_response_bits_data; // @[top.scala 813:23]
  wire  cpu115_clock; // @[top.scala 817:22]
  wire  cpu115_reset; // @[top.scala 817:22]
  wire [31:0] cpu115_io_imem_address; // @[top.scala 817:22]
  wire [31:0] cpu115_io_imem_instruction; // @[top.scala 817:22]
  wire [31:0] cpu115_io_dmem_address; // @[top.scala 817:22]
  wire  cpu115_io_dmem_valid; // @[top.scala 817:22]
  wire [31:0] cpu115_io_dmem_writedata; // @[top.scala 817:22]
  wire  cpu115_io_dmem_memread; // @[top.scala 817:22]
  wire  cpu115_io_dmem_memwrite; // @[top.scala 817:22]
  wire [1:0] cpu115_io_dmem_maskmode; // @[top.scala 817:22]
  wire  cpu115_io_dmem_sext; // @[top.scala 817:22]
  wire [31:0] cpu115_io_dmem_readdata; // @[top.scala 817:22]
  wire  mem115_clock; // @[top.scala 818:22]
  wire  mem115_reset; // @[top.scala 818:22]
  wire [31:0] mem115_io_imem_request_bits_address; // @[top.scala 818:22]
  wire [31:0] mem115_io_imem_response_bits_data; // @[top.scala 818:22]
  wire  mem115_io_dmem_request_valid; // @[top.scala 818:22]
  wire [31:0] mem115_io_dmem_request_bits_address; // @[top.scala 818:22]
  wire [31:0] mem115_io_dmem_request_bits_writedata; // @[top.scala 818:22]
  wire [1:0] mem115_io_dmem_request_bits_operation; // @[top.scala 818:22]
  wire  mem115_io_dmem_response_valid; // @[top.scala 818:22]
  wire [31:0] mem115_io_dmem_response_bits_data; // @[top.scala 818:22]
  wire [31:0] imem115_io_pipeline_address; // @[top.scala 819:23]
  wire [31:0] imem115_io_pipeline_instruction; // @[top.scala 819:23]
  wire [31:0] imem115_io_bus_request_bits_address; // @[top.scala 819:23]
  wire [31:0] imem115_io_bus_response_bits_data; // @[top.scala 819:23]
  wire  dmem115_clock; // @[top.scala 820:23]
  wire  dmem115_reset; // @[top.scala 820:23]
  wire [31:0] dmem115_io_pipeline_address; // @[top.scala 820:23]
  wire  dmem115_io_pipeline_valid; // @[top.scala 820:23]
  wire [31:0] dmem115_io_pipeline_writedata; // @[top.scala 820:23]
  wire  dmem115_io_pipeline_memread; // @[top.scala 820:23]
  wire  dmem115_io_pipeline_memwrite; // @[top.scala 820:23]
  wire [1:0] dmem115_io_pipeline_maskmode; // @[top.scala 820:23]
  wire  dmem115_io_pipeline_sext; // @[top.scala 820:23]
  wire [31:0] dmem115_io_pipeline_readdata; // @[top.scala 820:23]
  wire  dmem115_io_bus_request_valid; // @[top.scala 820:23]
  wire [31:0] dmem115_io_bus_request_bits_address; // @[top.scala 820:23]
  wire [31:0] dmem115_io_bus_request_bits_writedata; // @[top.scala 820:23]
  wire [1:0] dmem115_io_bus_request_bits_operation; // @[top.scala 820:23]
  wire  dmem115_io_bus_response_valid; // @[top.scala 820:23]
  wire [31:0] dmem115_io_bus_response_bits_data; // @[top.scala 820:23]
  wire  cpu116_clock; // @[top.scala 824:22]
  wire  cpu116_reset; // @[top.scala 824:22]
  wire [31:0] cpu116_io_imem_address; // @[top.scala 824:22]
  wire [31:0] cpu116_io_imem_instruction; // @[top.scala 824:22]
  wire [31:0] cpu116_io_dmem_address; // @[top.scala 824:22]
  wire  cpu116_io_dmem_valid; // @[top.scala 824:22]
  wire [31:0] cpu116_io_dmem_writedata; // @[top.scala 824:22]
  wire  cpu116_io_dmem_memread; // @[top.scala 824:22]
  wire  cpu116_io_dmem_memwrite; // @[top.scala 824:22]
  wire [1:0] cpu116_io_dmem_maskmode; // @[top.scala 824:22]
  wire  cpu116_io_dmem_sext; // @[top.scala 824:22]
  wire [31:0] cpu116_io_dmem_readdata; // @[top.scala 824:22]
  wire  mem116_clock; // @[top.scala 825:22]
  wire  mem116_reset; // @[top.scala 825:22]
  wire [31:0] mem116_io_imem_request_bits_address; // @[top.scala 825:22]
  wire [31:0] mem116_io_imem_response_bits_data; // @[top.scala 825:22]
  wire  mem116_io_dmem_request_valid; // @[top.scala 825:22]
  wire [31:0] mem116_io_dmem_request_bits_address; // @[top.scala 825:22]
  wire [31:0] mem116_io_dmem_request_bits_writedata; // @[top.scala 825:22]
  wire [1:0] mem116_io_dmem_request_bits_operation; // @[top.scala 825:22]
  wire  mem116_io_dmem_response_valid; // @[top.scala 825:22]
  wire [31:0] mem116_io_dmem_response_bits_data; // @[top.scala 825:22]
  wire [31:0] imem116_io_pipeline_address; // @[top.scala 826:23]
  wire [31:0] imem116_io_pipeline_instruction; // @[top.scala 826:23]
  wire [31:0] imem116_io_bus_request_bits_address; // @[top.scala 826:23]
  wire [31:0] imem116_io_bus_response_bits_data; // @[top.scala 826:23]
  wire  dmem116_clock; // @[top.scala 827:23]
  wire  dmem116_reset; // @[top.scala 827:23]
  wire [31:0] dmem116_io_pipeline_address; // @[top.scala 827:23]
  wire  dmem116_io_pipeline_valid; // @[top.scala 827:23]
  wire [31:0] dmem116_io_pipeline_writedata; // @[top.scala 827:23]
  wire  dmem116_io_pipeline_memread; // @[top.scala 827:23]
  wire  dmem116_io_pipeline_memwrite; // @[top.scala 827:23]
  wire [1:0] dmem116_io_pipeline_maskmode; // @[top.scala 827:23]
  wire  dmem116_io_pipeline_sext; // @[top.scala 827:23]
  wire [31:0] dmem116_io_pipeline_readdata; // @[top.scala 827:23]
  wire  dmem116_io_bus_request_valid; // @[top.scala 827:23]
  wire [31:0] dmem116_io_bus_request_bits_address; // @[top.scala 827:23]
  wire [31:0] dmem116_io_bus_request_bits_writedata; // @[top.scala 827:23]
  wire [1:0] dmem116_io_bus_request_bits_operation; // @[top.scala 827:23]
  wire  dmem116_io_bus_response_valid; // @[top.scala 827:23]
  wire [31:0] dmem116_io_bus_response_bits_data; // @[top.scala 827:23]
  wire  cpu117_clock; // @[top.scala 831:22]
  wire  cpu117_reset; // @[top.scala 831:22]
  wire [31:0] cpu117_io_imem_address; // @[top.scala 831:22]
  wire [31:0] cpu117_io_imem_instruction; // @[top.scala 831:22]
  wire [31:0] cpu117_io_dmem_address; // @[top.scala 831:22]
  wire  cpu117_io_dmem_valid; // @[top.scala 831:22]
  wire [31:0] cpu117_io_dmem_writedata; // @[top.scala 831:22]
  wire  cpu117_io_dmem_memread; // @[top.scala 831:22]
  wire  cpu117_io_dmem_memwrite; // @[top.scala 831:22]
  wire [1:0] cpu117_io_dmem_maskmode; // @[top.scala 831:22]
  wire  cpu117_io_dmem_sext; // @[top.scala 831:22]
  wire [31:0] cpu117_io_dmem_readdata; // @[top.scala 831:22]
  wire  mem117_clock; // @[top.scala 832:22]
  wire  mem117_reset; // @[top.scala 832:22]
  wire [31:0] mem117_io_imem_request_bits_address; // @[top.scala 832:22]
  wire [31:0] mem117_io_imem_response_bits_data; // @[top.scala 832:22]
  wire  mem117_io_dmem_request_valid; // @[top.scala 832:22]
  wire [31:0] mem117_io_dmem_request_bits_address; // @[top.scala 832:22]
  wire [31:0] mem117_io_dmem_request_bits_writedata; // @[top.scala 832:22]
  wire [1:0] mem117_io_dmem_request_bits_operation; // @[top.scala 832:22]
  wire  mem117_io_dmem_response_valid; // @[top.scala 832:22]
  wire [31:0] mem117_io_dmem_response_bits_data; // @[top.scala 832:22]
  wire [31:0] imem117_io_pipeline_address; // @[top.scala 833:23]
  wire [31:0] imem117_io_pipeline_instruction; // @[top.scala 833:23]
  wire [31:0] imem117_io_bus_request_bits_address; // @[top.scala 833:23]
  wire [31:0] imem117_io_bus_response_bits_data; // @[top.scala 833:23]
  wire  dmem117_clock; // @[top.scala 834:23]
  wire  dmem117_reset; // @[top.scala 834:23]
  wire [31:0] dmem117_io_pipeline_address; // @[top.scala 834:23]
  wire  dmem117_io_pipeline_valid; // @[top.scala 834:23]
  wire [31:0] dmem117_io_pipeline_writedata; // @[top.scala 834:23]
  wire  dmem117_io_pipeline_memread; // @[top.scala 834:23]
  wire  dmem117_io_pipeline_memwrite; // @[top.scala 834:23]
  wire [1:0] dmem117_io_pipeline_maskmode; // @[top.scala 834:23]
  wire  dmem117_io_pipeline_sext; // @[top.scala 834:23]
  wire [31:0] dmem117_io_pipeline_readdata; // @[top.scala 834:23]
  wire  dmem117_io_bus_request_valid; // @[top.scala 834:23]
  wire [31:0] dmem117_io_bus_request_bits_address; // @[top.scala 834:23]
  wire [31:0] dmem117_io_bus_request_bits_writedata; // @[top.scala 834:23]
  wire [1:0] dmem117_io_bus_request_bits_operation; // @[top.scala 834:23]
  wire  dmem117_io_bus_response_valid; // @[top.scala 834:23]
  wire [31:0] dmem117_io_bus_response_bits_data; // @[top.scala 834:23]
  wire  cpu118_clock; // @[top.scala 838:22]
  wire  cpu118_reset; // @[top.scala 838:22]
  wire [31:0] cpu118_io_imem_address; // @[top.scala 838:22]
  wire [31:0] cpu118_io_imem_instruction; // @[top.scala 838:22]
  wire [31:0] cpu118_io_dmem_address; // @[top.scala 838:22]
  wire  cpu118_io_dmem_valid; // @[top.scala 838:22]
  wire [31:0] cpu118_io_dmem_writedata; // @[top.scala 838:22]
  wire  cpu118_io_dmem_memread; // @[top.scala 838:22]
  wire  cpu118_io_dmem_memwrite; // @[top.scala 838:22]
  wire [1:0] cpu118_io_dmem_maskmode; // @[top.scala 838:22]
  wire  cpu118_io_dmem_sext; // @[top.scala 838:22]
  wire [31:0] cpu118_io_dmem_readdata; // @[top.scala 838:22]
  wire  mem118_clock; // @[top.scala 839:22]
  wire  mem118_reset; // @[top.scala 839:22]
  wire [31:0] mem118_io_imem_request_bits_address; // @[top.scala 839:22]
  wire [31:0] mem118_io_imem_response_bits_data; // @[top.scala 839:22]
  wire  mem118_io_dmem_request_valid; // @[top.scala 839:22]
  wire [31:0] mem118_io_dmem_request_bits_address; // @[top.scala 839:22]
  wire [31:0] mem118_io_dmem_request_bits_writedata; // @[top.scala 839:22]
  wire [1:0] mem118_io_dmem_request_bits_operation; // @[top.scala 839:22]
  wire  mem118_io_dmem_response_valid; // @[top.scala 839:22]
  wire [31:0] mem118_io_dmem_response_bits_data; // @[top.scala 839:22]
  wire [31:0] imem118_io_pipeline_address; // @[top.scala 840:23]
  wire [31:0] imem118_io_pipeline_instruction; // @[top.scala 840:23]
  wire [31:0] imem118_io_bus_request_bits_address; // @[top.scala 840:23]
  wire [31:0] imem118_io_bus_response_bits_data; // @[top.scala 840:23]
  wire  dmem118_clock; // @[top.scala 841:23]
  wire  dmem118_reset; // @[top.scala 841:23]
  wire [31:0] dmem118_io_pipeline_address; // @[top.scala 841:23]
  wire  dmem118_io_pipeline_valid; // @[top.scala 841:23]
  wire [31:0] dmem118_io_pipeline_writedata; // @[top.scala 841:23]
  wire  dmem118_io_pipeline_memread; // @[top.scala 841:23]
  wire  dmem118_io_pipeline_memwrite; // @[top.scala 841:23]
  wire [1:0] dmem118_io_pipeline_maskmode; // @[top.scala 841:23]
  wire  dmem118_io_pipeline_sext; // @[top.scala 841:23]
  wire [31:0] dmem118_io_pipeline_readdata; // @[top.scala 841:23]
  wire  dmem118_io_bus_request_valid; // @[top.scala 841:23]
  wire [31:0] dmem118_io_bus_request_bits_address; // @[top.scala 841:23]
  wire [31:0] dmem118_io_bus_request_bits_writedata; // @[top.scala 841:23]
  wire [1:0] dmem118_io_bus_request_bits_operation; // @[top.scala 841:23]
  wire  dmem118_io_bus_response_valid; // @[top.scala 841:23]
  wire [31:0] dmem118_io_bus_response_bits_data; // @[top.scala 841:23]
  wire  cpu119_clock; // @[top.scala 845:22]
  wire  cpu119_reset; // @[top.scala 845:22]
  wire [31:0] cpu119_io_imem_address; // @[top.scala 845:22]
  wire [31:0] cpu119_io_imem_instruction; // @[top.scala 845:22]
  wire [31:0] cpu119_io_dmem_address; // @[top.scala 845:22]
  wire  cpu119_io_dmem_valid; // @[top.scala 845:22]
  wire [31:0] cpu119_io_dmem_writedata; // @[top.scala 845:22]
  wire  cpu119_io_dmem_memread; // @[top.scala 845:22]
  wire  cpu119_io_dmem_memwrite; // @[top.scala 845:22]
  wire [1:0] cpu119_io_dmem_maskmode; // @[top.scala 845:22]
  wire  cpu119_io_dmem_sext; // @[top.scala 845:22]
  wire [31:0] cpu119_io_dmem_readdata; // @[top.scala 845:22]
  wire  mem119_clock; // @[top.scala 846:22]
  wire  mem119_reset; // @[top.scala 846:22]
  wire [31:0] mem119_io_imem_request_bits_address; // @[top.scala 846:22]
  wire [31:0] mem119_io_imem_response_bits_data; // @[top.scala 846:22]
  wire  mem119_io_dmem_request_valid; // @[top.scala 846:22]
  wire [31:0] mem119_io_dmem_request_bits_address; // @[top.scala 846:22]
  wire [31:0] mem119_io_dmem_request_bits_writedata; // @[top.scala 846:22]
  wire [1:0] mem119_io_dmem_request_bits_operation; // @[top.scala 846:22]
  wire  mem119_io_dmem_response_valid; // @[top.scala 846:22]
  wire [31:0] mem119_io_dmem_response_bits_data; // @[top.scala 846:22]
  wire [31:0] imem119_io_pipeline_address; // @[top.scala 847:23]
  wire [31:0] imem119_io_pipeline_instruction; // @[top.scala 847:23]
  wire [31:0] imem119_io_bus_request_bits_address; // @[top.scala 847:23]
  wire [31:0] imem119_io_bus_response_bits_data; // @[top.scala 847:23]
  wire  dmem119_clock; // @[top.scala 848:23]
  wire  dmem119_reset; // @[top.scala 848:23]
  wire [31:0] dmem119_io_pipeline_address; // @[top.scala 848:23]
  wire  dmem119_io_pipeline_valid; // @[top.scala 848:23]
  wire [31:0] dmem119_io_pipeline_writedata; // @[top.scala 848:23]
  wire  dmem119_io_pipeline_memread; // @[top.scala 848:23]
  wire  dmem119_io_pipeline_memwrite; // @[top.scala 848:23]
  wire [1:0] dmem119_io_pipeline_maskmode; // @[top.scala 848:23]
  wire  dmem119_io_pipeline_sext; // @[top.scala 848:23]
  wire [31:0] dmem119_io_pipeline_readdata; // @[top.scala 848:23]
  wire  dmem119_io_bus_request_valid; // @[top.scala 848:23]
  wire [31:0] dmem119_io_bus_request_bits_address; // @[top.scala 848:23]
  wire [31:0] dmem119_io_bus_request_bits_writedata; // @[top.scala 848:23]
  wire [1:0] dmem119_io_bus_request_bits_operation; // @[top.scala 848:23]
  wire  dmem119_io_bus_response_valid; // @[top.scala 848:23]
  wire [31:0] dmem119_io_bus_response_bits_data; // @[top.scala 848:23]
  wire  cpu120_clock; // @[top.scala 852:22]
  wire  cpu120_reset; // @[top.scala 852:22]
  wire [31:0] cpu120_io_imem_address; // @[top.scala 852:22]
  wire [31:0] cpu120_io_imem_instruction; // @[top.scala 852:22]
  wire [31:0] cpu120_io_dmem_address; // @[top.scala 852:22]
  wire  cpu120_io_dmem_valid; // @[top.scala 852:22]
  wire [31:0] cpu120_io_dmem_writedata; // @[top.scala 852:22]
  wire  cpu120_io_dmem_memread; // @[top.scala 852:22]
  wire  cpu120_io_dmem_memwrite; // @[top.scala 852:22]
  wire [1:0] cpu120_io_dmem_maskmode; // @[top.scala 852:22]
  wire  cpu120_io_dmem_sext; // @[top.scala 852:22]
  wire [31:0] cpu120_io_dmem_readdata; // @[top.scala 852:22]
  wire  mem120_clock; // @[top.scala 853:22]
  wire  mem120_reset; // @[top.scala 853:22]
  wire [31:0] mem120_io_imem_request_bits_address; // @[top.scala 853:22]
  wire [31:0] mem120_io_imem_response_bits_data; // @[top.scala 853:22]
  wire  mem120_io_dmem_request_valid; // @[top.scala 853:22]
  wire [31:0] mem120_io_dmem_request_bits_address; // @[top.scala 853:22]
  wire [31:0] mem120_io_dmem_request_bits_writedata; // @[top.scala 853:22]
  wire [1:0] mem120_io_dmem_request_bits_operation; // @[top.scala 853:22]
  wire  mem120_io_dmem_response_valid; // @[top.scala 853:22]
  wire [31:0] mem120_io_dmem_response_bits_data; // @[top.scala 853:22]
  wire [31:0] imem120_io_pipeline_address; // @[top.scala 854:23]
  wire [31:0] imem120_io_pipeline_instruction; // @[top.scala 854:23]
  wire [31:0] imem120_io_bus_request_bits_address; // @[top.scala 854:23]
  wire [31:0] imem120_io_bus_response_bits_data; // @[top.scala 854:23]
  wire  dmem120_clock; // @[top.scala 855:23]
  wire  dmem120_reset; // @[top.scala 855:23]
  wire [31:0] dmem120_io_pipeline_address; // @[top.scala 855:23]
  wire  dmem120_io_pipeline_valid; // @[top.scala 855:23]
  wire [31:0] dmem120_io_pipeline_writedata; // @[top.scala 855:23]
  wire  dmem120_io_pipeline_memread; // @[top.scala 855:23]
  wire  dmem120_io_pipeline_memwrite; // @[top.scala 855:23]
  wire [1:0] dmem120_io_pipeline_maskmode; // @[top.scala 855:23]
  wire  dmem120_io_pipeline_sext; // @[top.scala 855:23]
  wire [31:0] dmem120_io_pipeline_readdata; // @[top.scala 855:23]
  wire  dmem120_io_bus_request_valid; // @[top.scala 855:23]
  wire [31:0] dmem120_io_bus_request_bits_address; // @[top.scala 855:23]
  wire [31:0] dmem120_io_bus_request_bits_writedata; // @[top.scala 855:23]
  wire [1:0] dmem120_io_bus_request_bits_operation; // @[top.scala 855:23]
  wire  dmem120_io_bus_response_valid; // @[top.scala 855:23]
  wire [31:0] dmem120_io_bus_response_bits_data; // @[top.scala 855:23]
  wire  cpu121_clock; // @[top.scala 859:22]
  wire  cpu121_reset; // @[top.scala 859:22]
  wire [31:0] cpu121_io_imem_address; // @[top.scala 859:22]
  wire [31:0] cpu121_io_imem_instruction; // @[top.scala 859:22]
  wire [31:0] cpu121_io_dmem_address; // @[top.scala 859:22]
  wire  cpu121_io_dmem_valid; // @[top.scala 859:22]
  wire [31:0] cpu121_io_dmem_writedata; // @[top.scala 859:22]
  wire  cpu121_io_dmem_memread; // @[top.scala 859:22]
  wire  cpu121_io_dmem_memwrite; // @[top.scala 859:22]
  wire [1:0] cpu121_io_dmem_maskmode; // @[top.scala 859:22]
  wire  cpu121_io_dmem_sext; // @[top.scala 859:22]
  wire [31:0] cpu121_io_dmem_readdata; // @[top.scala 859:22]
  wire  mem121_clock; // @[top.scala 860:22]
  wire  mem121_reset; // @[top.scala 860:22]
  wire [31:0] mem121_io_imem_request_bits_address; // @[top.scala 860:22]
  wire [31:0] mem121_io_imem_response_bits_data; // @[top.scala 860:22]
  wire  mem121_io_dmem_request_valid; // @[top.scala 860:22]
  wire [31:0] mem121_io_dmem_request_bits_address; // @[top.scala 860:22]
  wire [31:0] mem121_io_dmem_request_bits_writedata; // @[top.scala 860:22]
  wire [1:0] mem121_io_dmem_request_bits_operation; // @[top.scala 860:22]
  wire  mem121_io_dmem_response_valid; // @[top.scala 860:22]
  wire [31:0] mem121_io_dmem_response_bits_data; // @[top.scala 860:22]
  wire [31:0] imem121_io_pipeline_address; // @[top.scala 861:23]
  wire [31:0] imem121_io_pipeline_instruction; // @[top.scala 861:23]
  wire [31:0] imem121_io_bus_request_bits_address; // @[top.scala 861:23]
  wire [31:0] imem121_io_bus_response_bits_data; // @[top.scala 861:23]
  wire  dmem121_clock; // @[top.scala 862:23]
  wire  dmem121_reset; // @[top.scala 862:23]
  wire [31:0] dmem121_io_pipeline_address; // @[top.scala 862:23]
  wire  dmem121_io_pipeline_valid; // @[top.scala 862:23]
  wire [31:0] dmem121_io_pipeline_writedata; // @[top.scala 862:23]
  wire  dmem121_io_pipeline_memread; // @[top.scala 862:23]
  wire  dmem121_io_pipeline_memwrite; // @[top.scala 862:23]
  wire [1:0] dmem121_io_pipeline_maskmode; // @[top.scala 862:23]
  wire  dmem121_io_pipeline_sext; // @[top.scala 862:23]
  wire [31:0] dmem121_io_pipeline_readdata; // @[top.scala 862:23]
  wire  dmem121_io_bus_request_valid; // @[top.scala 862:23]
  wire [31:0] dmem121_io_bus_request_bits_address; // @[top.scala 862:23]
  wire [31:0] dmem121_io_bus_request_bits_writedata; // @[top.scala 862:23]
  wire [1:0] dmem121_io_bus_request_bits_operation; // @[top.scala 862:23]
  wire  dmem121_io_bus_response_valid; // @[top.scala 862:23]
  wire [31:0] dmem121_io_bus_response_bits_data; // @[top.scala 862:23]
  wire  cpu122_clock; // @[top.scala 866:22]
  wire  cpu122_reset; // @[top.scala 866:22]
  wire [31:0] cpu122_io_imem_address; // @[top.scala 866:22]
  wire [31:0] cpu122_io_imem_instruction; // @[top.scala 866:22]
  wire [31:0] cpu122_io_dmem_address; // @[top.scala 866:22]
  wire  cpu122_io_dmem_valid; // @[top.scala 866:22]
  wire [31:0] cpu122_io_dmem_writedata; // @[top.scala 866:22]
  wire  cpu122_io_dmem_memread; // @[top.scala 866:22]
  wire  cpu122_io_dmem_memwrite; // @[top.scala 866:22]
  wire [1:0] cpu122_io_dmem_maskmode; // @[top.scala 866:22]
  wire  cpu122_io_dmem_sext; // @[top.scala 866:22]
  wire [31:0] cpu122_io_dmem_readdata; // @[top.scala 866:22]
  wire  mem122_clock; // @[top.scala 867:22]
  wire  mem122_reset; // @[top.scala 867:22]
  wire [31:0] mem122_io_imem_request_bits_address; // @[top.scala 867:22]
  wire [31:0] mem122_io_imem_response_bits_data; // @[top.scala 867:22]
  wire  mem122_io_dmem_request_valid; // @[top.scala 867:22]
  wire [31:0] mem122_io_dmem_request_bits_address; // @[top.scala 867:22]
  wire [31:0] mem122_io_dmem_request_bits_writedata; // @[top.scala 867:22]
  wire [1:0] mem122_io_dmem_request_bits_operation; // @[top.scala 867:22]
  wire  mem122_io_dmem_response_valid; // @[top.scala 867:22]
  wire [31:0] mem122_io_dmem_response_bits_data; // @[top.scala 867:22]
  wire [31:0] imem122_io_pipeline_address; // @[top.scala 868:23]
  wire [31:0] imem122_io_pipeline_instruction; // @[top.scala 868:23]
  wire [31:0] imem122_io_bus_request_bits_address; // @[top.scala 868:23]
  wire [31:0] imem122_io_bus_response_bits_data; // @[top.scala 868:23]
  wire  dmem122_clock; // @[top.scala 869:23]
  wire  dmem122_reset; // @[top.scala 869:23]
  wire [31:0] dmem122_io_pipeline_address; // @[top.scala 869:23]
  wire  dmem122_io_pipeline_valid; // @[top.scala 869:23]
  wire [31:0] dmem122_io_pipeline_writedata; // @[top.scala 869:23]
  wire  dmem122_io_pipeline_memread; // @[top.scala 869:23]
  wire  dmem122_io_pipeline_memwrite; // @[top.scala 869:23]
  wire [1:0] dmem122_io_pipeline_maskmode; // @[top.scala 869:23]
  wire  dmem122_io_pipeline_sext; // @[top.scala 869:23]
  wire [31:0] dmem122_io_pipeline_readdata; // @[top.scala 869:23]
  wire  dmem122_io_bus_request_valid; // @[top.scala 869:23]
  wire [31:0] dmem122_io_bus_request_bits_address; // @[top.scala 869:23]
  wire [31:0] dmem122_io_bus_request_bits_writedata; // @[top.scala 869:23]
  wire [1:0] dmem122_io_bus_request_bits_operation; // @[top.scala 869:23]
  wire  dmem122_io_bus_response_valid; // @[top.scala 869:23]
  wire [31:0] dmem122_io_bus_response_bits_data; // @[top.scala 869:23]
  wire  cpu123_clock; // @[top.scala 873:22]
  wire  cpu123_reset; // @[top.scala 873:22]
  wire [31:0] cpu123_io_imem_address; // @[top.scala 873:22]
  wire [31:0] cpu123_io_imem_instruction; // @[top.scala 873:22]
  wire [31:0] cpu123_io_dmem_address; // @[top.scala 873:22]
  wire  cpu123_io_dmem_valid; // @[top.scala 873:22]
  wire [31:0] cpu123_io_dmem_writedata; // @[top.scala 873:22]
  wire  cpu123_io_dmem_memread; // @[top.scala 873:22]
  wire  cpu123_io_dmem_memwrite; // @[top.scala 873:22]
  wire [1:0] cpu123_io_dmem_maskmode; // @[top.scala 873:22]
  wire  cpu123_io_dmem_sext; // @[top.scala 873:22]
  wire [31:0] cpu123_io_dmem_readdata; // @[top.scala 873:22]
  wire  mem123_clock; // @[top.scala 874:22]
  wire  mem123_reset; // @[top.scala 874:22]
  wire [31:0] mem123_io_imem_request_bits_address; // @[top.scala 874:22]
  wire [31:0] mem123_io_imem_response_bits_data; // @[top.scala 874:22]
  wire  mem123_io_dmem_request_valid; // @[top.scala 874:22]
  wire [31:0] mem123_io_dmem_request_bits_address; // @[top.scala 874:22]
  wire [31:0] mem123_io_dmem_request_bits_writedata; // @[top.scala 874:22]
  wire [1:0] mem123_io_dmem_request_bits_operation; // @[top.scala 874:22]
  wire  mem123_io_dmem_response_valid; // @[top.scala 874:22]
  wire [31:0] mem123_io_dmem_response_bits_data; // @[top.scala 874:22]
  wire [31:0] imem123_io_pipeline_address; // @[top.scala 875:23]
  wire [31:0] imem123_io_pipeline_instruction; // @[top.scala 875:23]
  wire [31:0] imem123_io_bus_request_bits_address; // @[top.scala 875:23]
  wire [31:0] imem123_io_bus_response_bits_data; // @[top.scala 875:23]
  wire  dmem123_clock; // @[top.scala 876:23]
  wire  dmem123_reset; // @[top.scala 876:23]
  wire [31:0] dmem123_io_pipeline_address; // @[top.scala 876:23]
  wire  dmem123_io_pipeline_valid; // @[top.scala 876:23]
  wire [31:0] dmem123_io_pipeline_writedata; // @[top.scala 876:23]
  wire  dmem123_io_pipeline_memread; // @[top.scala 876:23]
  wire  dmem123_io_pipeline_memwrite; // @[top.scala 876:23]
  wire [1:0] dmem123_io_pipeline_maskmode; // @[top.scala 876:23]
  wire  dmem123_io_pipeline_sext; // @[top.scala 876:23]
  wire [31:0] dmem123_io_pipeline_readdata; // @[top.scala 876:23]
  wire  dmem123_io_bus_request_valid; // @[top.scala 876:23]
  wire [31:0] dmem123_io_bus_request_bits_address; // @[top.scala 876:23]
  wire [31:0] dmem123_io_bus_request_bits_writedata; // @[top.scala 876:23]
  wire [1:0] dmem123_io_bus_request_bits_operation; // @[top.scala 876:23]
  wire  dmem123_io_bus_response_valid; // @[top.scala 876:23]
  wire [31:0] dmem123_io_bus_response_bits_data; // @[top.scala 876:23]
  wire  cpu124_clock; // @[top.scala 880:22]
  wire  cpu124_reset; // @[top.scala 880:22]
  wire [31:0] cpu124_io_imem_address; // @[top.scala 880:22]
  wire [31:0] cpu124_io_imem_instruction; // @[top.scala 880:22]
  wire [31:0] cpu124_io_dmem_address; // @[top.scala 880:22]
  wire  cpu124_io_dmem_valid; // @[top.scala 880:22]
  wire [31:0] cpu124_io_dmem_writedata; // @[top.scala 880:22]
  wire  cpu124_io_dmem_memread; // @[top.scala 880:22]
  wire  cpu124_io_dmem_memwrite; // @[top.scala 880:22]
  wire [1:0] cpu124_io_dmem_maskmode; // @[top.scala 880:22]
  wire  cpu124_io_dmem_sext; // @[top.scala 880:22]
  wire [31:0] cpu124_io_dmem_readdata; // @[top.scala 880:22]
  wire  mem124_clock; // @[top.scala 881:22]
  wire  mem124_reset; // @[top.scala 881:22]
  wire [31:0] mem124_io_imem_request_bits_address; // @[top.scala 881:22]
  wire [31:0] mem124_io_imem_response_bits_data; // @[top.scala 881:22]
  wire  mem124_io_dmem_request_valid; // @[top.scala 881:22]
  wire [31:0] mem124_io_dmem_request_bits_address; // @[top.scala 881:22]
  wire [31:0] mem124_io_dmem_request_bits_writedata; // @[top.scala 881:22]
  wire [1:0] mem124_io_dmem_request_bits_operation; // @[top.scala 881:22]
  wire  mem124_io_dmem_response_valid; // @[top.scala 881:22]
  wire [31:0] mem124_io_dmem_response_bits_data; // @[top.scala 881:22]
  wire [31:0] imem124_io_pipeline_address; // @[top.scala 882:23]
  wire [31:0] imem124_io_pipeline_instruction; // @[top.scala 882:23]
  wire [31:0] imem124_io_bus_request_bits_address; // @[top.scala 882:23]
  wire [31:0] imem124_io_bus_response_bits_data; // @[top.scala 882:23]
  wire  dmem124_clock; // @[top.scala 883:23]
  wire  dmem124_reset; // @[top.scala 883:23]
  wire [31:0] dmem124_io_pipeline_address; // @[top.scala 883:23]
  wire  dmem124_io_pipeline_valid; // @[top.scala 883:23]
  wire [31:0] dmem124_io_pipeline_writedata; // @[top.scala 883:23]
  wire  dmem124_io_pipeline_memread; // @[top.scala 883:23]
  wire  dmem124_io_pipeline_memwrite; // @[top.scala 883:23]
  wire [1:0] dmem124_io_pipeline_maskmode; // @[top.scala 883:23]
  wire  dmem124_io_pipeline_sext; // @[top.scala 883:23]
  wire [31:0] dmem124_io_pipeline_readdata; // @[top.scala 883:23]
  wire  dmem124_io_bus_request_valid; // @[top.scala 883:23]
  wire [31:0] dmem124_io_bus_request_bits_address; // @[top.scala 883:23]
  wire [31:0] dmem124_io_bus_request_bits_writedata; // @[top.scala 883:23]
  wire [1:0] dmem124_io_bus_request_bits_operation; // @[top.scala 883:23]
  wire  dmem124_io_bus_response_valid; // @[top.scala 883:23]
  wire [31:0] dmem124_io_bus_response_bits_data; // @[top.scala 883:23]
  wire  cpu125_clock; // @[top.scala 887:22]
  wire  cpu125_reset; // @[top.scala 887:22]
  wire [31:0] cpu125_io_imem_address; // @[top.scala 887:22]
  wire [31:0] cpu125_io_imem_instruction; // @[top.scala 887:22]
  wire [31:0] cpu125_io_dmem_address; // @[top.scala 887:22]
  wire  cpu125_io_dmem_valid; // @[top.scala 887:22]
  wire [31:0] cpu125_io_dmem_writedata; // @[top.scala 887:22]
  wire  cpu125_io_dmem_memread; // @[top.scala 887:22]
  wire  cpu125_io_dmem_memwrite; // @[top.scala 887:22]
  wire [1:0] cpu125_io_dmem_maskmode; // @[top.scala 887:22]
  wire  cpu125_io_dmem_sext; // @[top.scala 887:22]
  wire [31:0] cpu125_io_dmem_readdata; // @[top.scala 887:22]
  wire  mem125_clock; // @[top.scala 888:22]
  wire  mem125_reset; // @[top.scala 888:22]
  wire [31:0] mem125_io_imem_request_bits_address; // @[top.scala 888:22]
  wire [31:0] mem125_io_imem_response_bits_data; // @[top.scala 888:22]
  wire  mem125_io_dmem_request_valid; // @[top.scala 888:22]
  wire [31:0] mem125_io_dmem_request_bits_address; // @[top.scala 888:22]
  wire [31:0] mem125_io_dmem_request_bits_writedata; // @[top.scala 888:22]
  wire [1:0] mem125_io_dmem_request_bits_operation; // @[top.scala 888:22]
  wire  mem125_io_dmem_response_valid; // @[top.scala 888:22]
  wire [31:0] mem125_io_dmem_response_bits_data; // @[top.scala 888:22]
  wire [31:0] imem125_io_pipeline_address; // @[top.scala 889:23]
  wire [31:0] imem125_io_pipeline_instruction; // @[top.scala 889:23]
  wire [31:0] imem125_io_bus_request_bits_address; // @[top.scala 889:23]
  wire [31:0] imem125_io_bus_response_bits_data; // @[top.scala 889:23]
  wire  dmem125_clock; // @[top.scala 890:23]
  wire  dmem125_reset; // @[top.scala 890:23]
  wire [31:0] dmem125_io_pipeline_address; // @[top.scala 890:23]
  wire  dmem125_io_pipeline_valid; // @[top.scala 890:23]
  wire [31:0] dmem125_io_pipeline_writedata; // @[top.scala 890:23]
  wire  dmem125_io_pipeline_memread; // @[top.scala 890:23]
  wire  dmem125_io_pipeline_memwrite; // @[top.scala 890:23]
  wire [1:0] dmem125_io_pipeline_maskmode; // @[top.scala 890:23]
  wire  dmem125_io_pipeline_sext; // @[top.scala 890:23]
  wire [31:0] dmem125_io_pipeline_readdata; // @[top.scala 890:23]
  wire  dmem125_io_bus_request_valid; // @[top.scala 890:23]
  wire [31:0] dmem125_io_bus_request_bits_address; // @[top.scala 890:23]
  wire [31:0] dmem125_io_bus_request_bits_writedata; // @[top.scala 890:23]
  wire [1:0] dmem125_io_bus_request_bits_operation; // @[top.scala 890:23]
  wire  dmem125_io_bus_response_valid; // @[top.scala 890:23]
  wire [31:0] dmem125_io_bus_response_bits_data; // @[top.scala 890:23]
  wire  cpu126_clock; // @[top.scala 894:22]
  wire  cpu126_reset; // @[top.scala 894:22]
  wire [31:0] cpu126_io_imem_address; // @[top.scala 894:22]
  wire [31:0] cpu126_io_imem_instruction; // @[top.scala 894:22]
  wire [31:0] cpu126_io_dmem_address; // @[top.scala 894:22]
  wire  cpu126_io_dmem_valid; // @[top.scala 894:22]
  wire [31:0] cpu126_io_dmem_writedata; // @[top.scala 894:22]
  wire  cpu126_io_dmem_memread; // @[top.scala 894:22]
  wire  cpu126_io_dmem_memwrite; // @[top.scala 894:22]
  wire [1:0] cpu126_io_dmem_maskmode; // @[top.scala 894:22]
  wire  cpu126_io_dmem_sext; // @[top.scala 894:22]
  wire [31:0] cpu126_io_dmem_readdata; // @[top.scala 894:22]
  wire  mem126_clock; // @[top.scala 895:22]
  wire  mem126_reset; // @[top.scala 895:22]
  wire [31:0] mem126_io_imem_request_bits_address; // @[top.scala 895:22]
  wire [31:0] mem126_io_imem_response_bits_data; // @[top.scala 895:22]
  wire  mem126_io_dmem_request_valid; // @[top.scala 895:22]
  wire [31:0] mem126_io_dmem_request_bits_address; // @[top.scala 895:22]
  wire [31:0] mem126_io_dmem_request_bits_writedata; // @[top.scala 895:22]
  wire [1:0] mem126_io_dmem_request_bits_operation; // @[top.scala 895:22]
  wire  mem126_io_dmem_response_valid; // @[top.scala 895:22]
  wire [31:0] mem126_io_dmem_response_bits_data; // @[top.scala 895:22]
  wire [31:0] imem126_io_pipeline_address; // @[top.scala 896:23]
  wire [31:0] imem126_io_pipeline_instruction; // @[top.scala 896:23]
  wire [31:0] imem126_io_bus_request_bits_address; // @[top.scala 896:23]
  wire [31:0] imem126_io_bus_response_bits_data; // @[top.scala 896:23]
  wire  dmem126_clock; // @[top.scala 897:23]
  wire  dmem126_reset; // @[top.scala 897:23]
  wire [31:0] dmem126_io_pipeline_address; // @[top.scala 897:23]
  wire  dmem126_io_pipeline_valid; // @[top.scala 897:23]
  wire [31:0] dmem126_io_pipeline_writedata; // @[top.scala 897:23]
  wire  dmem126_io_pipeline_memread; // @[top.scala 897:23]
  wire  dmem126_io_pipeline_memwrite; // @[top.scala 897:23]
  wire [1:0] dmem126_io_pipeline_maskmode; // @[top.scala 897:23]
  wire  dmem126_io_pipeline_sext; // @[top.scala 897:23]
  wire [31:0] dmem126_io_pipeline_readdata; // @[top.scala 897:23]
  wire  dmem126_io_bus_request_valid; // @[top.scala 897:23]
  wire [31:0] dmem126_io_bus_request_bits_address; // @[top.scala 897:23]
  wire [31:0] dmem126_io_bus_request_bits_writedata; // @[top.scala 897:23]
  wire [1:0] dmem126_io_bus_request_bits_operation; // @[top.scala 897:23]
  wire  dmem126_io_bus_response_valid; // @[top.scala 897:23]
  wire [31:0] dmem126_io_bus_response_bits_data; // @[top.scala 897:23]
  wire  cpu127_clock; // @[top.scala 901:22]
  wire  cpu127_reset; // @[top.scala 901:22]
  wire [31:0] cpu127_io_imem_address; // @[top.scala 901:22]
  wire [31:0] cpu127_io_imem_instruction; // @[top.scala 901:22]
  wire [31:0] cpu127_io_dmem_address; // @[top.scala 901:22]
  wire  cpu127_io_dmem_valid; // @[top.scala 901:22]
  wire [31:0] cpu127_io_dmem_writedata; // @[top.scala 901:22]
  wire  cpu127_io_dmem_memread; // @[top.scala 901:22]
  wire  cpu127_io_dmem_memwrite; // @[top.scala 901:22]
  wire [1:0] cpu127_io_dmem_maskmode; // @[top.scala 901:22]
  wire  cpu127_io_dmem_sext; // @[top.scala 901:22]
  wire [31:0] cpu127_io_dmem_readdata; // @[top.scala 901:22]
  wire  mem127_clock; // @[top.scala 902:22]
  wire  mem127_reset; // @[top.scala 902:22]
  wire [31:0] mem127_io_imem_request_bits_address; // @[top.scala 902:22]
  wire [31:0] mem127_io_imem_response_bits_data; // @[top.scala 902:22]
  wire  mem127_io_dmem_request_valid; // @[top.scala 902:22]
  wire [31:0] mem127_io_dmem_request_bits_address; // @[top.scala 902:22]
  wire [31:0] mem127_io_dmem_request_bits_writedata; // @[top.scala 902:22]
  wire [1:0] mem127_io_dmem_request_bits_operation; // @[top.scala 902:22]
  wire  mem127_io_dmem_response_valid; // @[top.scala 902:22]
  wire [31:0] mem127_io_dmem_response_bits_data; // @[top.scala 902:22]
  wire [31:0] imem127_io_pipeline_address; // @[top.scala 903:23]
  wire [31:0] imem127_io_pipeline_instruction; // @[top.scala 903:23]
  wire [31:0] imem127_io_bus_request_bits_address; // @[top.scala 903:23]
  wire [31:0] imem127_io_bus_response_bits_data; // @[top.scala 903:23]
  wire  dmem127_clock; // @[top.scala 904:23]
  wire  dmem127_reset; // @[top.scala 904:23]
  wire [31:0] dmem127_io_pipeline_address; // @[top.scala 904:23]
  wire  dmem127_io_pipeline_valid; // @[top.scala 904:23]
  wire [31:0] dmem127_io_pipeline_writedata; // @[top.scala 904:23]
  wire  dmem127_io_pipeline_memread; // @[top.scala 904:23]
  wire  dmem127_io_pipeline_memwrite; // @[top.scala 904:23]
  wire [1:0] dmem127_io_pipeline_maskmode; // @[top.scala 904:23]
  wire  dmem127_io_pipeline_sext; // @[top.scala 904:23]
  wire [31:0] dmem127_io_pipeline_readdata; // @[top.scala 904:23]
  wire  dmem127_io_bus_request_valid; // @[top.scala 904:23]
  wire [31:0] dmem127_io_bus_request_bits_address; // @[top.scala 904:23]
  wire [31:0] dmem127_io_bus_request_bits_writedata; // @[top.scala 904:23]
  wire [1:0] dmem127_io_bus_request_bits_operation; // @[top.scala 904:23]
  wire  dmem127_io_bus_response_valid; // @[top.scala 904:23]
  wire [31:0] dmem127_io_bus_response_bits_data; // @[top.scala 904:23]
  PipelinedCPUBP cpu0 ( // @[top.scala 12:20]
    .clock(cpu0_clock),
    .reset(cpu0_reset),
    .io_imem_address(cpu0_io_imem_address),
    .io_imem_instruction(cpu0_io_imem_instruction),
    .io_dmem_address(cpu0_io_dmem_address),
    .io_dmem_valid(cpu0_io_dmem_valid),
    .io_dmem_writedata(cpu0_io_dmem_writedata),
    .io_dmem_memread(cpu0_io_dmem_memread),
    .io_dmem_memwrite(cpu0_io_dmem_memwrite),
    .io_dmem_maskmode(cpu0_io_dmem_maskmode),
    .io_dmem_sext(cpu0_io_dmem_sext),
    .io_dmem_readdata(cpu0_io_dmem_readdata)
  );
  DualPortedCombinMemory mem0 ( // @[top.scala 13:20]
    .clock(mem0_clock),
    .reset(mem0_reset),
    .io_imem_request_bits_address(mem0_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem0_io_imem_response_bits_data),
    .io_dmem_request_valid(mem0_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem0_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem0_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem0_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem0_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem0_io_dmem_response_bits_data)
  );
  ICombinMemPort imem0 ( // @[top.scala 14:21]
    .io_pipeline_address(imem0_io_pipeline_address),
    .io_pipeline_instruction(imem0_io_pipeline_instruction),
    .io_bus_request_bits_address(imem0_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem0_io_bus_response_bits_data)
  );
  DCombinMemPort dmem0 ( // @[top.scala 15:21]
    .clock(dmem0_clock),
    .reset(dmem0_reset),
    .io_pipeline_address(dmem0_io_pipeline_address),
    .io_pipeline_valid(dmem0_io_pipeline_valid),
    .io_pipeline_writedata(dmem0_io_pipeline_writedata),
    .io_pipeline_memread(dmem0_io_pipeline_memread),
    .io_pipeline_memwrite(dmem0_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem0_io_pipeline_maskmode),
    .io_pipeline_sext(dmem0_io_pipeline_sext),
    .io_pipeline_readdata(dmem0_io_pipeline_readdata),
    .io_bus_request_valid(dmem0_io_bus_request_valid),
    .io_bus_request_bits_address(dmem0_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem0_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem0_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem0_io_bus_response_valid),
    .io_bus_response_bits_data(dmem0_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu1 ( // @[top.scala 19:20]
    .clock(cpu1_clock),
    .reset(cpu1_reset),
    .io_imem_address(cpu1_io_imem_address),
    .io_imem_instruction(cpu1_io_imem_instruction),
    .io_dmem_address(cpu1_io_dmem_address),
    .io_dmem_valid(cpu1_io_dmem_valid),
    .io_dmem_writedata(cpu1_io_dmem_writedata),
    .io_dmem_memread(cpu1_io_dmem_memread),
    .io_dmem_memwrite(cpu1_io_dmem_memwrite),
    .io_dmem_maskmode(cpu1_io_dmem_maskmode),
    .io_dmem_sext(cpu1_io_dmem_sext),
    .io_dmem_readdata(cpu1_io_dmem_readdata)
  );
  DualPortedCombinMemory mem1 ( // @[top.scala 20:20]
    .clock(mem1_clock),
    .reset(mem1_reset),
    .io_imem_request_bits_address(mem1_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem1_io_imem_response_bits_data),
    .io_dmem_request_valid(mem1_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem1_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem1_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem1_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem1_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem1_io_dmem_response_bits_data)
  );
  ICombinMemPort imem1 ( // @[top.scala 21:21]
    .io_pipeline_address(imem1_io_pipeline_address),
    .io_pipeline_instruction(imem1_io_pipeline_instruction),
    .io_bus_request_bits_address(imem1_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem1_io_bus_response_bits_data)
  );
  DCombinMemPort dmem1 ( // @[top.scala 22:21]
    .clock(dmem1_clock),
    .reset(dmem1_reset),
    .io_pipeline_address(dmem1_io_pipeline_address),
    .io_pipeline_valid(dmem1_io_pipeline_valid),
    .io_pipeline_writedata(dmem1_io_pipeline_writedata),
    .io_pipeline_memread(dmem1_io_pipeline_memread),
    .io_pipeline_memwrite(dmem1_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem1_io_pipeline_maskmode),
    .io_pipeline_sext(dmem1_io_pipeline_sext),
    .io_pipeline_readdata(dmem1_io_pipeline_readdata),
    .io_bus_request_valid(dmem1_io_bus_request_valid),
    .io_bus_request_bits_address(dmem1_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem1_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem1_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem1_io_bus_response_valid),
    .io_bus_response_bits_data(dmem1_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu2 ( // @[top.scala 26:20]
    .clock(cpu2_clock),
    .reset(cpu2_reset),
    .io_imem_address(cpu2_io_imem_address),
    .io_imem_instruction(cpu2_io_imem_instruction),
    .io_dmem_address(cpu2_io_dmem_address),
    .io_dmem_valid(cpu2_io_dmem_valid),
    .io_dmem_writedata(cpu2_io_dmem_writedata),
    .io_dmem_memread(cpu2_io_dmem_memread),
    .io_dmem_memwrite(cpu2_io_dmem_memwrite),
    .io_dmem_maskmode(cpu2_io_dmem_maskmode),
    .io_dmem_sext(cpu2_io_dmem_sext),
    .io_dmem_readdata(cpu2_io_dmem_readdata)
  );
  DualPortedCombinMemory mem2 ( // @[top.scala 27:20]
    .clock(mem2_clock),
    .reset(mem2_reset),
    .io_imem_request_bits_address(mem2_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem2_io_imem_response_bits_data),
    .io_dmem_request_valid(mem2_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem2_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem2_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem2_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem2_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem2_io_dmem_response_bits_data)
  );
  ICombinMemPort imem2 ( // @[top.scala 28:21]
    .io_pipeline_address(imem2_io_pipeline_address),
    .io_pipeline_instruction(imem2_io_pipeline_instruction),
    .io_bus_request_bits_address(imem2_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem2_io_bus_response_bits_data)
  );
  DCombinMemPort dmem2 ( // @[top.scala 29:21]
    .clock(dmem2_clock),
    .reset(dmem2_reset),
    .io_pipeline_address(dmem2_io_pipeline_address),
    .io_pipeline_valid(dmem2_io_pipeline_valid),
    .io_pipeline_writedata(dmem2_io_pipeline_writedata),
    .io_pipeline_memread(dmem2_io_pipeline_memread),
    .io_pipeline_memwrite(dmem2_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem2_io_pipeline_maskmode),
    .io_pipeline_sext(dmem2_io_pipeline_sext),
    .io_pipeline_readdata(dmem2_io_pipeline_readdata),
    .io_bus_request_valid(dmem2_io_bus_request_valid),
    .io_bus_request_bits_address(dmem2_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem2_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem2_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem2_io_bus_response_valid),
    .io_bus_response_bits_data(dmem2_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu3 ( // @[top.scala 33:20]
    .clock(cpu3_clock),
    .reset(cpu3_reset),
    .io_imem_address(cpu3_io_imem_address),
    .io_imem_instruction(cpu3_io_imem_instruction),
    .io_dmem_address(cpu3_io_dmem_address),
    .io_dmem_valid(cpu3_io_dmem_valid),
    .io_dmem_writedata(cpu3_io_dmem_writedata),
    .io_dmem_memread(cpu3_io_dmem_memread),
    .io_dmem_memwrite(cpu3_io_dmem_memwrite),
    .io_dmem_maskmode(cpu3_io_dmem_maskmode),
    .io_dmem_sext(cpu3_io_dmem_sext),
    .io_dmem_readdata(cpu3_io_dmem_readdata)
  );
  DualPortedCombinMemory mem3 ( // @[top.scala 34:20]
    .clock(mem3_clock),
    .reset(mem3_reset),
    .io_imem_request_bits_address(mem3_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem3_io_imem_response_bits_data),
    .io_dmem_request_valid(mem3_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem3_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem3_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem3_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem3_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem3_io_dmem_response_bits_data)
  );
  ICombinMemPort imem3 ( // @[top.scala 35:21]
    .io_pipeline_address(imem3_io_pipeline_address),
    .io_pipeline_instruction(imem3_io_pipeline_instruction),
    .io_bus_request_bits_address(imem3_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem3_io_bus_response_bits_data)
  );
  DCombinMemPort dmem3 ( // @[top.scala 36:21]
    .clock(dmem3_clock),
    .reset(dmem3_reset),
    .io_pipeline_address(dmem3_io_pipeline_address),
    .io_pipeline_valid(dmem3_io_pipeline_valid),
    .io_pipeline_writedata(dmem3_io_pipeline_writedata),
    .io_pipeline_memread(dmem3_io_pipeline_memread),
    .io_pipeline_memwrite(dmem3_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem3_io_pipeline_maskmode),
    .io_pipeline_sext(dmem3_io_pipeline_sext),
    .io_pipeline_readdata(dmem3_io_pipeline_readdata),
    .io_bus_request_valid(dmem3_io_bus_request_valid),
    .io_bus_request_bits_address(dmem3_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem3_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem3_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem3_io_bus_response_valid),
    .io_bus_response_bits_data(dmem3_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu4 ( // @[top.scala 40:20]
    .clock(cpu4_clock),
    .reset(cpu4_reset),
    .io_imem_address(cpu4_io_imem_address),
    .io_imem_instruction(cpu4_io_imem_instruction),
    .io_dmem_address(cpu4_io_dmem_address),
    .io_dmem_valid(cpu4_io_dmem_valid),
    .io_dmem_writedata(cpu4_io_dmem_writedata),
    .io_dmem_memread(cpu4_io_dmem_memread),
    .io_dmem_memwrite(cpu4_io_dmem_memwrite),
    .io_dmem_maskmode(cpu4_io_dmem_maskmode),
    .io_dmem_sext(cpu4_io_dmem_sext),
    .io_dmem_readdata(cpu4_io_dmem_readdata)
  );
  DualPortedCombinMemory mem4 ( // @[top.scala 41:20]
    .clock(mem4_clock),
    .reset(mem4_reset),
    .io_imem_request_bits_address(mem4_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem4_io_imem_response_bits_data),
    .io_dmem_request_valid(mem4_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem4_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem4_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem4_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem4_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem4_io_dmem_response_bits_data)
  );
  ICombinMemPort imem4 ( // @[top.scala 42:21]
    .io_pipeline_address(imem4_io_pipeline_address),
    .io_pipeline_instruction(imem4_io_pipeline_instruction),
    .io_bus_request_bits_address(imem4_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem4_io_bus_response_bits_data)
  );
  DCombinMemPort dmem4 ( // @[top.scala 43:21]
    .clock(dmem4_clock),
    .reset(dmem4_reset),
    .io_pipeline_address(dmem4_io_pipeline_address),
    .io_pipeline_valid(dmem4_io_pipeline_valid),
    .io_pipeline_writedata(dmem4_io_pipeline_writedata),
    .io_pipeline_memread(dmem4_io_pipeline_memread),
    .io_pipeline_memwrite(dmem4_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem4_io_pipeline_maskmode),
    .io_pipeline_sext(dmem4_io_pipeline_sext),
    .io_pipeline_readdata(dmem4_io_pipeline_readdata),
    .io_bus_request_valid(dmem4_io_bus_request_valid),
    .io_bus_request_bits_address(dmem4_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem4_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem4_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem4_io_bus_response_valid),
    .io_bus_response_bits_data(dmem4_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu5 ( // @[top.scala 47:20]
    .clock(cpu5_clock),
    .reset(cpu5_reset),
    .io_imem_address(cpu5_io_imem_address),
    .io_imem_instruction(cpu5_io_imem_instruction),
    .io_dmem_address(cpu5_io_dmem_address),
    .io_dmem_valid(cpu5_io_dmem_valid),
    .io_dmem_writedata(cpu5_io_dmem_writedata),
    .io_dmem_memread(cpu5_io_dmem_memread),
    .io_dmem_memwrite(cpu5_io_dmem_memwrite),
    .io_dmem_maskmode(cpu5_io_dmem_maskmode),
    .io_dmem_sext(cpu5_io_dmem_sext),
    .io_dmem_readdata(cpu5_io_dmem_readdata)
  );
  DualPortedCombinMemory mem5 ( // @[top.scala 48:20]
    .clock(mem5_clock),
    .reset(mem5_reset),
    .io_imem_request_bits_address(mem5_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem5_io_imem_response_bits_data),
    .io_dmem_request_valid(mem5_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem5_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem5_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem5_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem5_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem5_io_dmem_response_bits_data)
  );
  ICombinMemPort imem5 ( // @[top.scala 49:21]
    .io_pipeline_address(imem5_io_pipeline_address),
    .io_pipeline_instruction(imem5_io_pipeline_instruction),
    .io_bus_request_bits_address(imem5_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem5_io_bus_response_bits_data)
  );
  DCombinMemPort dmem5 ( // @[top.scala 50:21]
    .clock(dmem5_clock),
    .reset(dmem5_reset),
    .io_pipeline_address(dmem5_io_pipeline_address),
    .io_pipeline_valid(dmem5_io_pipeline_valid),
    .io_pipeline_writedata(dmem5_io_pipeline_writedata),
    .io_pipeline_memread(dmem5_io_pipeline_memread),
    .io_pipeline_memwrite(dmem5_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem5_io_pipeline_maskmode),
    .io_pipeline_sext(dmem5_io_pipeline_sext),
    .io_pipeline_readdata(dmem5_io_pipeline_readdata),
    .io_bus_request_valid(dmem5_io_bus_request_valid),
    .io_bus_request_bits_address(dmem5_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem5_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem5_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem5_io_bus_response_valid),
    .io_bus_response_bits_data(dmem5_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu6 ( // @[top.scala 54:20]
    .clock(cpu6_clock),
    .reset(cpu6_reset),
    .io_imem_address(cpu6_io_imem_address),
    .io_imem_instruction(cpu6_io_imem_instruction),
    .io_dmem_address(cpu6_io_dmem_address),
    .io_dmem_valid(cpu6_io_dmem_valid),
    .io_dmem_writedata(cpu6_io_dmem_writedata),
    .io_dmem_memread(cpu6_io_dmem_memread),
    .io_dmem_memwrite(cpu6_io_dmem_memwrite),
    .io_dmem_maskmode(cpu6_io_dmem_maskmode),
    .io_dmem_sext(cpu6_io_dmem_sext),
    .io_dmem_readdata(cpu6_io_dmem_readdata)
  );
  DualPortedCombinMemory mem6 ( // @[top.scala 55:20]
    .clock(mem6_clock),
    .reset(mem6_reset),
    .io_imem_request_bits_address(mem6_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem6_io_imem_response_bits_data),
    .io_dmem_request_valid(mem6_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem6_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem6_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem6_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem6_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem6_io_dmem_response_bits_data)
  );
  ICombinMemPort imem6 ( // @[top.scala 56:21]
    .io_pipeline_address(imem6_io_pipeline_address),
    .io_pipeline_instruction(imem6_io_pipeline_instruction),
    .io_bus_request_bits_address(imem6_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem6_io_bus_response_bits_data)
  );
  DCombinMemPort dmem6 ( // @[top.scala 57:21]
    .clock(dmem6_clock),
    .reset(dmem6_reset),
    .io_pipeline_address(dmem6_io_pipeline_address),
    .io_pipeline_valid(dmem6_io_pipeline_valid),
    .io_pipeline_writedata(dmem6_io_pipeline_writedata),
    .io_pipeline_memread(dmem6_io_pipeline_memread),
    .io_pipeline_memwrite(dmem6_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem6_io_pipeline_maskmode),
    .io_pipeline_sext(dmem6_io_pipeline_sext),
    .io_pipeline_readdata(dmem6_io_pipeline_readdata),
    .io_bus_request_valid(dmem6_io_bus_request_valid),
    .io_bus_request_bits_address(dmem6_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem6_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem6_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem6_io_bus_response_valid),
    .io_bus_response_bits_data(dmem6_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu7 ( // @[top.scala 61:20]
    .clock(cpu7_clock),
    .reset(cpu7_reset),
    .io_imem_address(cpu7_io_imem_address),
    .io_imem_instruction(cpu7_io_imem_instruction),
    .io_dmem_address(cpu7_io_dmem_address),
    .io_dmem_valid(cpu7_io_dmem_valid),
    .io_dmem_writedata(cpu7_io_dmem_writedata),
    .io_dmem_memread(cpu7_io_dmem_memread),
    .io_dmem_memwrite(cpu7_io_dmem_memwrite),
    .io_dmem_maskmode(cpu7_io_dmem_maskmode),
    .io_dmem_sext(cpu7_io_dmem_sext),
    .io_dmem_readdata(cpu7_io_dmem_readdata)
  );
  DualPortedCombinMemory mem7 ( // @[top.scala 62:20]
    .clock(mem7_clock),
    .reset(mem7_reset),
    .io_imem_request_bits_address(mem7_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem7_io_imem_response_bits_data),
    .io_dmem_request_valid(mem7_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem7_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem7_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem7_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem7_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem7_io_dmem_response_bits_data)
  );
  ICombinMemPort imem7 ( // @[top.scala 63:21]
    .io_pipeline_address(imem7_io_pipeline_address),
    .io_pipeline_instruction(imem7_io_pipeline_instruction),
    .io_bus_request_bits_address(imem7_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem7_io_bus_response_bits_data)
  );
  DCombinMemPort dmem7 ( // @[top.scala 64:21]
    .clock(dmem7_clock),
    .reset(dmem7_reset),
    .io_pipeline_address(dmem7_io_pipeline_address),
    .io_pipeline_valid(dmem7_io_pipeline_valid),
    .io_pipeline_writedata(dmem7_io_pipeline_writedata),
    .io_pipeline_memread(dmem7_io_pipeline_memread),
    .io_pipeline_memwrite(dmem7_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem7_io_pipeline_maskmode),
    .io_pipeline_sext(dmem7_io_pipeline_sext),
    .io_pipeline_readdata(dmem7_io_pipeline_readdata),
    .io_bus_request_valid(dmem7_io_bus_request_valid),
    .io_bus_request_bits_address(dmem7_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem7_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem7_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem7_io_bus_response_valid),
    .io_bus_response_bits_data(dmem7_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu8 ( // @[top.scala 68:20]
    .clock(cpu8_clock),
    .reset(cpu8_reset),
    .io_imem_address(cpu8_io_imem_address),
    .io_imem_instruction(cpu8_io_imem_instruction),
    .io_dmem_address(cpu8_io_dmem_address),
    .io_dmem_valid(cpu8_io_dmem_valid),
    .io_dmem_writedata(cpu8_io_dmem_writedata),
    .io_dmem_memread(cpu8_io_dmem_memread),
    .io_dmem_memwrite(cpu8_io_dmem_memwrite),
    .io_dmem_maskmode(cpu8_io_dmem_maskmode),
    .io_dmem_sext(cpu8_io_dmem_sext),
    .io_dmem_readdata(cpu8_io_dmem_readdata)
  );
  DualPortedCombinMemory mem8 ( // @[top.scala 69:20]
    .clock(mem8_clock),
    .reset(mem8_reset),
    .io_imem_request_bits_address(mem8_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem8_io_imem_response_bits_data),
    .io_dmem_request_valid(mem8_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem8_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem8_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem8_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem8_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem8_io_dmem_response_bits_data)
  );
  ICombinMemPort imem8 ( // @[top.scala 70:21]
    .io_pipeline_address(imem8_io_pipeline_address),
    .io_pipeline_instruction(imem8_io_pipeline_instruction),
    .io_bus_request_bits_address(imem8_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem8_io_bus_response_bits_data)
  );
  DCombinMemPort dmem8 ( // @[top.scala 71:21]
    .clock(dmem8_clock),
    .reset(dmem8_reset),
    .io_pipeline_address(dmem8_io_pipeline_address),
    .io_pipeline_valid(dmem8_io_pipeline_valid),
    .io_pipeline_writedata(dmem8_io_pipeline_writedata),
    .io_pipeline_memread(dmem8_io_pipeline_memread),
    .io_pipeline_memwrite(dmem8_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem8_io_pipeline_maskmode),
    .io_pipeline_sext(dmem8_io_pipeline_sext),
    .io_pipeline_readdata(dmem8_io_pipeline_readdata),
    .io_bus_request_valid(dmem8_io_bus_request_valid),
    .io_bus_request_bits_address(dmem8_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem8_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem8_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem8_io_bus_response_valid),
    .io_bus_response_bits_data(dmem8_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu9 ( // @[top.scala 75:20]
    .clock(cpu9_clock),
    .reset(cpu9_reset),
    .io_imem_address(cpu9_io_imem_address),
    .io_imem_instruction(cpu9_io_imem_instruction),
    .io_dmem_address(cpu9_io_dmem_address),
    .io_dmem_valid(cpu9_io_dmem_valid),
    .io_dmem_writedata(cpu9_io_dmem_writedata),
    .io_dmem_memread(cpu9_io_dmem_memread),
    .io_dmem_memwrite(cpu9_io_dmem_memwrite),
    .io_dmem_maskmode(cpu9_io_dmem_maskmode),
    .io_dmem_sext(cpu9_io_dmem_sext),
    .io_dmem_readdata(cpu9_io_dmem_readdata)
  );
  DualPortedCombinMemory mem9 ( // @[top.scala 76:20]
    .clock(mem9_clock),
    .reset(mem9_reset),
    .io_imem_request_bits_address(mem9_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem9_io_imem_response_bits_data),
    .io_dmem_request_valid(mem9_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem9_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem9_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem9_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem9_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem9_io_dmem_response_bits_data)
  );
  ICombinMemPort imem9 ( // @[top.scala 77:21]
    .io_pipeline_address(imem9_io_pipeline_address),
    .io_pipeline_instruction(imem9_io_pipeline_instruction),
    .io_bus_request_bits_address(imem9_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem9_io_bus_response_bits_data)
  );
  DCombinMemPort dmem9 ( // @[top.scala 78:21]
    .clock(dmem9_clock),
    .reset(dmem9_reset),
    .io_pipeline_address(dmem9_io_pipeline_address),
    .io_pipeline_valid(dmem9_io_pipeline_valid),
    .io_pipeline_writedata(dmem9_io_pipeline_writedata),
    .io_pipeline_memread(dmem9_io_pipeline_memread),
    .io_pipeline_memwrite(dmem9_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem9_io_pipeline_maskmode),
    .io_pipeline_sext(dmem9_io_pipeline_sext),
    .io_pipeline_readdata(dmem9_io_pipeline_readdata),
    .io_bus_request_valid(dmem9_io_bus_request_valid),
    .io_bus_request_bits_address(dmem9_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem9_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem9_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem9_io_bus_response_valid),
    .io_bus_response_bits_data(dmem9_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu10 ( // @[top.scala 82:21]
    .clock(cpu10_clock),
    .reset(cpu10_reset),
    .io_imem_address(cpu10_io_imem_address),
    .io_imem_instruction(cpu10_io_imem_instruction),
    .io_dmem_address(cpu10_io_dmem_address),
    .io_dmem_valid(cpu10_io_dmem_valid),
    .io_dmem_writedata(cpu10_io_dmem_writedata),
    .io_dmem_memread(cpu10_io_dmem_memread),
    .io_dmem_memwrite(cpu10_io_dmem_memwrite),
    .io_dmem_maskmode(cpu10_io_dmem_maskmode),
    .io_dmem_sext(cpu10_io_dmem_sext),
    .io_dmem_readdata(cpu10_io_dmem_readdata)
  );
  DualPortedCombinMemory mem10 ( // @[top.scala 83:21]
    .clock(mem10_clock),
    .reset(mem10_reset),
    .io_imem_request_bits_address(mem10_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem10_io_imem_response_bits_data),
    .io_dmem_request_valid(mem10_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem10_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem10_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem10_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem10_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem10_io_dmem_response_bits_data)
  );
  ICombinMemPort imem10 ( // @[top.scala 84:22]
    .io_pipeline_address(imem10_io_pipeline_address),
    .io_pipeline_instruction(imem10_io_pipeline_instruction),
    .io_bus_request_bits_address(imem10_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem10_io_bus_response_bits_data)
  );
  DCombinMemPort dmem10 ( // @[top.scala 85:22]
    .clock(dmem10_clock),
    .reset(dmem10_reset),
    .io_pipeline_address(dmem10_io_pipeline_address),
    .io_pipeline_valid(dmem10_io_pipeline_valid),
    .io_pipeline_writedata(dmem10_io_pipeline_writedata),
    .io_pipeline_memread(dmem10_io_pipeline_memread),
    .io_pipeline_memwrite(dmem10_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem10_io_pipeline_maskmode),
    .io_pipeline_sext(dmem10_io_pipeline_sext),
    .io_pipeline_readdata(dmem10_io_pipeline_readdata),
    .io_bus_request_valid(dmem10_io_bus_request_valid),
    .io_bus_request_bits_address(dmem10_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem10_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem10_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem10_io_bus_response_valid),
    .io_bus_response_bits_data(dmem10_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu11 ( // @[top.scala 89:21]
    .clock(cpu11_clock),
    .reset(cpu11_reset),
    .io_imem_address(cpu11_io_imem_address),
    .io_imem_instruction(cpu11_io_imem_instruction),
    .io_dmem_address(cpu11_io_dmem_address),
    .io_dmem_valid(cpu11_io_dmem_valid),
    .io_dmem_writedata(cpu11_io_dmem_writedata),
    .io_dmem_memread(cpu11_io_dmem_memread),
    .io_dmem_memwrite(cpu11_io_dmem_memwrite),
    .io_dmem_maskmode(cpu11_io_dmem_maskmode),
    .io_dmem_sext(cpu11_io_dmem_sext),
    .io_dmem_readdata(cpu11_io_dmem_readdata)
  );
  DualPortedCombinMemory mem11 ( // @[top.scala 90:21]
    .clock(mem11_clock),
    .reset(mem11_reset),
    .io_imem_request_bits_address(mem11_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem11_io_imem_response_bits_data),
    .io_dmem_request_valid(mem11_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem11_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem11_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem11_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem11_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem11_io_dmem_response_bits_data)
  );
  ICombinMemPort imem11 ( // @[top.scala 91:22]
    .io_pipeline_address(imem11_io_pipeline_address),
    .io_pipeline_instruction(imem11_io_pipeline_instruction),
    .io_bus_request_bits_address(imem11_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem11_io_bus_response_bits_data)
  );
  DCombinMemPort dmem11 ( // @[top.scala 92:22]
    .clock(dmem11_clock),
    .reset(dmem11_reset),
    .io_pipeline_address(dmem11_io_pipeline_address),
    .io_pipeline_valid(dmem11_io_pipeline_valid),
    .io_pipeline_writedata(dmem11_io_pipeline_writedata),
    .io_pipeline_memread(dmem11_io_pipeline_memread),
    .io_pipeline_memwrite(dmem11_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem11_io_pipeline_maskmode),
    .io_pipeline_sext(dmem11_io_pipeline_sext),
    .io_pipeline_readdata(dmem11_io_pipeline_readdata),
    .io_bus_request_valid(dmem11_io_bus_request_valid),
    .io_bus_request_bits_address(dmem11_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem11_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem11_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem11_io_bus_response_valid),
    .io_bus_response_bits_data(dmem11_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu12 ( // @[top.scala 96:21]
    .clock(cpu12_clock),
    .reset(cpu12_reset),
    .io_imem_address(cpu12_io_imem_address),
    .io_imem_instruction(cpu12_io_imem_instruction),
    .io_dmem_address(cpu12_io_dmem_address),
    .io_dmem_valid(cpu12_io_dmem_valid),
    .io_dmem_writedata(cpu12_io_dmem_writedata),
    .io_dmem_memread(cpu12_io_dmem_memread),
    .io_dmem_memwrite(cpu12_io_dmem_memwrite),
    .io_dmem_maskmode(cpu12_io_dmem_maskmode),
    .io_dmem_sext(cpu12_io_dmem_sext),
    .io_dmem_readdata(cpu12_io_dmem_readdata)
  );
  DualPortedCombinMemory mem12 ( // @[top.scala 97:21]
    .clock(mem12_clock),
    .reset(mem12_reset),
    .io_imem_request_bits_address(mem12_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem12_io_imem_response_bits_data),
    .io_dmem_request_valid(mem12_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem12_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem12_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem12_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem12_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem12_io_dmem_response_bits_data)
  );
  ICombinMemPort imem12 ( // @[top.scala 98:22]
    .io_pipeline_address(imem12_io_pipeline_address),
    .io_pipeline_instruction(imem12_io_pipeline_instruction),
    .io_bus_request_bits_address(imem12_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem12_io_bus_response_bits_data)
  );
  DCombinMemPort dmem12 ( // @[top.scala 99:22]
    .clock(dmem12_clock),
    .reset(dmem12_reset),
    .io_pipeline_address(dmem12_io_pipeline_address),
    .io_pipeline_valid(dmem12_io_pipeline_valid),
    .io_pipeline_writedata(dmem12_io_pipeline_writedata),
    .io_pipeline_memread(dmem12_io_pipeline_memread),
    .io_pipeline_memwrite(dmem12_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem12_io_pipeline_maskmode),
    .io_pipeline_sext(dmem12_io_pipeline_sext),
    .io_pipeline_readdata(dmem12_io_pipeline_readdata),
    .io_bus_request_valid(dmem12_io_bus_request_valid),
    .io_bus_request_bits_address(dmem12_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem12_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem12_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem12_io_bus_response_valid),
    .io_bus_response_bits_data(dmem12_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu13 ( // @[top.scala 103:21]
    .clock(cpu13_clock),
    .reset(cpu13_reset),
    .io_imem_address(cpu13_io_imem_address),
    .io_imem_instruction(cpu13_io_imem_instruction),
    .io_dmem_address(cpu13_io_dmem_address),
    .io_dmem_valid(cpu13_io_dmem_valid),
    .io_dmem_writedata(cpu13_io_dmem_writedata),
    .io_dmem_memread(cpu13_io_dmem_memread),
    .io_dmem_memwrite(cpu13_io_dmem_memwrite),
    .io_dmem_maskmode(cpu13_io_dmem_maskmode),
    .io_dmem_sext(cpu13_io_dmem_sext),
    .io_dmem_readdata(cpu13_io_dmem_readdata)
  );
  DualPortedCombinMemory mem13 ( // @[top.scala 104:21]
    .clock(mem13_clock),
    .reset(mem13_reset),
    .io_imem_request_bits_address(mem13_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem13_io_imem_response_bits_data),
    .io_dmem_request_valid(mem13_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem13_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem13_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem13_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem13_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem13_io_dmem_response_bits_data)
  );
  ICombinMemPort imem13 ( // @[top.scala 105:22]
    .io_pipeline_address(imem13_io_pipeline_address),
    .io_pipeline_instruction(imem13_io_pipeline_instruction),
    .io_bus_request_bits_address(imem13_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem13_io_bus_response_bits_data)
  );
  DCombinMemPort dmem13 ( // @[top.scala 106:22]
    .clock(dmem13_clock),
    .reset(dmem13_reset),
    .io_pipeline_address(dmem13_io_pipeline_address),
    .io_pipeline_valid(dmem13_io_pipeline_valid),
    .io_pipeline_writedata(dmem13_io_pipeline_writedata),
    .io_pipeline_memread(dmem13_io_pipeline_memread),
    .io_pipeline_memwrite(dmem13_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem13_io_pipeline_maskmode),
    .io_pipeline_sext(dmem13_io_pipeline_sext),
    .io_pipeline_readdata(dmem13_io_pipeline_readdata),
    .io_bus_request_valid(dmem13_io_bus_request_valid),
    .io_bus_request_bits_address(dmem13_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem13_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem13_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem13_io_bus_response_valid),
    .io_bus_response_bits_data(dmem13_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu14 ( // @[top.scala 110:21]
    .clock(cpu14_clock),
    .reset(cpu14_reset),
    .io_imem_address(cpu14_io_imem_address),
    .io_imem_instruction(cpu14_io_imem_instruction),
    .io_dmem_address(cpu14_io_dmem_address),
    .io_dmem_valid(cpu14_io_dmem_valid),
    .io_dmem_writedata(cpu14_io_dmem_writedata),
    .io_dmem_memread(cpu14_io_dmem_memread),
    .io_dmem_memwrite(cpu14_io_dmem_memwrite),
    .io_dmem_maskmode(cpu14_io_dmem_maskmode),
    .io_dmem_sext(cpu14_io_dmem_sext),
    .io_dmem_readdata(cpu14_io_dmem_readdata)
  );
  DualPortedCombinMemory mem14 ( // @[top.scala 111:21]
    .clock(mem14_clock),
    .reset(mem14_reset),
    .io_imem_request_bits_address(mem14_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem14_io_imem_response_bits_data),
    .io_dmem_request_valid(mem14_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem14_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem14_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem14_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem14_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem14_io_dmem_response_bits_data)
  );
  ICombinMemPort imem14 ( // @[top.scala 112:22]
    .io_pipeline_address(imem14_io_pipeline_address),
    .io_pipeline_instruction(imem14_io_pipeline_instruction),
    .io_bus_request_bits_address(imem14_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem14_io_bus_response_bits_data)
  );
  DCombinMemPort dmem14 ( // @[top.scala 113:22]
    .clock(dmem14_clock),
    .reset(dmem14_reset),
    .io_pipeline_address(dmem14_io_pipeline_address),
    .io_pipeline_valid(dmem14_io_pipeline_valid),
    .io_pipeline_writedata(dmem14_io_pipeline_writedata),
    .io_pipeline_memread(dmem14_io_pipeline_memread),
    .io_pipeline_memwrite(dmem14_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem14_io_pipeline_maskmode),
    .io_pipeline_sext(dmem14_io_pipeline_sext),
    .io_pipeline_readdata(dmem14_io_pipeline_readdata),
    .io_bus_request_valid(dmem14_io_bus_request_valid),
    .io_bus_request_bits_address(dmem14_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem14_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem14_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem14_io_bus_response_valid),
    .io_bus_response_bits_data(dmem14_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu15 ( // @[top.scala 117:21]
    .clock(cpu15_clock),
    .reset(cpu15_reset),
    .io_imem_address(cpu15_io_imem_address),
    .io_imem_instruction(cpu15_io_imem_instruction),
    .io_dmem_address(cpu15_io_dmem_address),
    .io_dmem_valid(cpu15_io_dmem_valid),
    .io_dmem_writedata(cpu15_io_dmem_writedata),
    .io_dmem_memread(cpu15_io_dmem_memread),
    .io_dmem_memwrite(cpu15_io_dmem_memwrite),
    .io_dmem_maskmode(cpu15_io_dmem_maskmode),
    .io_dmem_sext(cpu15_io_dmem_sext),
    .io_dmem_readdata(cpu15_io_dmem_readdata)
  );
  DualPortedCombinMemory mem15 ( // @[top.scala 118:21]
    .clock(mem15_clock),
    .reset(mem15_reset),
    .io_imem_request_bits_address(mem15_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem15_io_imem_response_bits_data),
    .io_dmem_request_valid(mem15_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem15_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem15_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem15_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem15_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem15_io_dmem_response_bits_data)
  );
  ICombinMemPort imem15 ( // @[top.scala 119:22]
    .io_pipeline_address(imem15_io_pipeline_address),
    .io_pipeline_instruction(imem15_io_pipeline_instruction),
    .io_bus_request_bits_address(imem15_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem15_io_bus_response_bits_data)
  );
  DCombinMemPort dmem15 ( // @[top.scala 120:22]
    .clock(dmem15_clock),
    .reset(dmem15_reset),
    .io_pipeline_address(dmem15_io_pipeline_address),
    .io_pipeline_valid(dmem15_io_pipeline_valid),
    .io_pipeline_writedata(dmem15_io_pipeline_writedata),
    .io_pipeline_memread(dmem15_io_pipeline_memread),
    .io_pipeline_memwrite(dmem15_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem15_io_pipeline_maskmode),
    .io_pipeline_sext(dmem15_io_pipeline_sext),
    .io_pipeline_readdata(dmem15_io_pipeline_readdata),
    .io_bus_request_valid(dmem15_io_bus_request_valid),
    .io_bus_request_bits_address(dmem15_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem15_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem15_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem15_io_bus_response_valid),
    .io_bus_response_bits_data(dmem15_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu16 ( // @[top.scala 124:21]
    .clock(cpu16_clock),
    .reset(cpu16_reset),
    .io_imem_address(cpu16_io_imem_address),
    .io_imem_instruction(cpu16_io_imem_instruction),
    .io_dmem_address(cpu16_io_dmem_address),
    .io_dmem_valid(cpu16_io_dmem_valid),
    .io_dmem_writedata(cpu16_io_dmem_writedata),
    .io_dmem_memread(cpu16_io_dmem_memread),
    .io_dmem_memwrite(cpu16_io_dmem_memwrite),
    .io_dmem_maskmode(cpu16_io_dmem_maskmode),
    .io_dmem_sext(cpu16_io_dmem_sext),
    .io_dmem_readdata(cpu16_io_dmem_readdata)
  );
  DualPortedCombinMemory mem16 ( // @[top.scala 125:21]
    .clock(mem16_clock),
    .reset(mem16_reset),
    .io_imem_request_bits_address(mem16_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem16_io_imem_response_bits_data),
    .io_dmem_request_valid(mem16_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem16_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem16_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem16_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem16_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem16_io_dmem_response_bits_data)
  );
  ICombinMemPort imem16 ( // @[top.scala 126:22]
    .io_pipeline_address(imem16_io_pipeline_address),
    .io_pipeline_instruction(imem16_io_pipeline_instruction),
    .io_bus_request_bits_address(imem16_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem16_io_bus_response_bits_data)
  );
  DCombinMemPort dmem16 ( // @[top.scala 127:22]
    .clock(dmem16_clock),
    .reset(dmem16_reset),
    .io_pipeline_address(dmem16_io_pipeline_address),
    .io_pipeline_valid(dmem16_io_pipeline_valid),
    .io_pipeline_writedata(dmem16_io_pipeline_writedata),
    .io_pipeline_memread(dmem16_io_pipeline_memread),
    .io_pipeline_memwrite(dmem16_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem16_io_pipeline_maskmode),
    .io_pipeline_sext(dmem16_io_pipeline_sext),
    .io_pipeline_readdata(dmem16_io_pipeline_readdata),
    .io_bus_request_valid(dmem16_io_bus_request_valid),
    .io_bus_request_bits_address(dmem16_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem16_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem16_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem16_io_bus_response_valid),
    .io_bus_response_bits_data(dmem16_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu17 ( // @[top.scala 131:21]
    .clock(cpu17_clock),
    .reset(cpu17_reset),
    .io_imem_address(cpu17_io_imem_address),
    .io_imem_instruction(cpu17_io_imem_instruction),
    .io_dmem_address(cpu17_io_dmem_address),
    .io_dmem_valid(cpu17_io_dmem_valid),
    .io_dmem_writedata(cpu17_io_dmem_writedata),
    .io_dmem_memread(cpu17_io_dmem_memread),
    .io_dmem_memwrite(cpu17_io_dmem_memwrite),
    .io_dmem_maskmode(cpu17_io_dmem_maskmode),
    .io_dmem_sext(cpu17_io_dmem_sext),
    .io_dmem_readdata(cpu17_io_dmem_readdata)
  );
  DualPortedCombinMemory mem17 ( // @[top.scala 132:21]
    .clock(mem17_clock),
    .reset(mem17_reset),
    .io_imem_request_bits_address(mem17_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem17_io_imem_response_bits_data),
    .io_dmem_request_valid(mem17_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem17_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem17_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem17_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem17_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem17_io_dmem_response_bits_data)
  );
  ICombinMemPort imem17 ( // @[top.scala 133:22]
    .io_pipeline_address(imem17_io_pipeline_address),
    .io_pipeline_instruction(imem17_io_pipeline_instruction),
    .io_bus_request_bits_address(imem17_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem17_io_bus_response_bits_data)
  );
  DCombinMemPort dmem17 ( // @[top.scala 134:22]
    .clock(dmem17_clock),
    .reset(dmem17_reset),
    .io_pipeline_address(dmem17_io_pipeline_address),
    .io_pipeline_valid(dmem17_io_pipeline_valid),
    .io_pipeline_writedata(dmem17_io_pipeline_writedata),
    .io_pipeline_memread(dmem17_io_pipeline_memread),
    .io_pipeline_memwrite(dmem17_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem17_io_pipeline_maskmode),
    .io_pipeline_sext(dmem17_io_pipeline_sext),
    .io_pipeline_readdata(dmem17_io_pipeline_readdata),
    .io_bus_request_valid(dmem17_io_bus_request_valid),
    .io_bus_request_bits_address(dmem17_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem17_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem17_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem17_io_bus_response_valid),
    .io_bus_response_bits_data(dmem17_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu18 ( // @[top.scala 138:21]
    .clock(cpu18_clock),
    .reset(cpu18_reset),
    .io_imem_address(cpu18_io_imem_address),
    .io_imem_instruction(cpu18_io_imem_instruction),
    .io_dmem_address(cpu18_io_dmem_address),
    .io_dmem_valid(cpu18_io_dmem_valid),
    .io_dmem_writedata(cpu18_io_dmem_writedata),
    .io_dmem_memread(cpu18_io_dmem_memread),
    .io_dmem_memwrite(cpu18_io_dmem_memwrite),
    .io_dmem_maskmode(cpu18_io_dmem_maskmode),
    .io_dmem_sext(cpu18_io_dmem_sext),
    .io_dmem_readdata(cpu18_io_dmem_readdata)
  );
  DualPortedCombinMemory mem18 ( // @[top.scala 139:21]
    .clock(mem18_clock),
    .reset(mem18_reset),
    .io_imem_request_bits_address(mem18_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem18_io_imem_response_bits_data),
    .io_dmem_request_valid(mem18_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem18_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem18_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem18_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem18_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem18_io_dmem_response_bits_data)
  );
  ICombinMemPort imem18 ( // @[top.scala 140:22]
    .io_pipeline_address(imem18_io_pipeline_address),
    .io_pipeline_instruction(imem18_io_pipeline_instruction),
    .io_bus_request_bits_address(imem18_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem18_io_bus_response_bits_data)
  );
  DCombinMemPort dmem18 ( // @[top.scala 141:22]
    .clock(dmem18_clock),
    .reset(dmem18_reset),
    .io_pipeline_address(dmem18_io_pipeline_address),
    .io_pipeline_valid(dmem18_io_pipeline_valid),
    .io_pipeline_writedata(dmem18_io_pipeline_writedata),
    .io_pipeline_memread(dmem18_io_pipeline_memread),
    .io_pipeline_memwrite(dmem18_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem18_io_pipeline_maskmode),
    .io_pipeline_sext(dmem18_io_pipeline_sext),
    .io_pipeline_readdata(dmem18_io_pipeline_readdata),
    .io_bus_request_valid(dmem18_io_bus_request_valid),
    .io_bus_request_bits_address(dmem18_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem18_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem18_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem18_io_bus_response_valid),
    .io_bus_response_bits_data(dmem18_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu19 ( // @[top.scala 145:21]
    .clock(cpu19_clock),
    .reset(cpu19_reset),
    .io_imem_address(cpu19_io_imem_address),
    .io_imem_instruction(cpu19_io_imem_instruction),
    .io_dmem_address(cpu19_io_dmem_address),
    .io_dmem_valid(cpu19_io_dmem_valid),
    .io_dmem_writedata(cpu19_io_dmem_writedata),
    .io_dmem_memread(cpu19_io_dmem_memread),
    .io_dmem_memwrite(cpu19_io_dmem_memwrite),
    .io_dmem_maskmode(cpu19_io_dmem_maskmode),
    .io_dmem_sext(cpu19_io_dmem_sext),
    .io_dmem_readdata(cpu19_io_dmem_readdata)
  );
  DualPortedCombinMemory mem19 ( // @[top.scala 146:21]
    .clock(mem19_clock),
    .reset(mem19_reset),
    .io_imem_request_bits_address(mem19_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem19_io_imem_response_bits_data),
    .io_dmem_request_valid(mem19_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem19_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem19_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem19_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem19_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem19_io_dmem_response_bits_data)
  );
  ICombinMemPort imem19 ( // @[top.scala 147:22]
    .io_pipeline_address(imem19_io_pipeline_address),
    .io_pipeline_instruction(imem19_io_pipeline_instruction),
    .io_bus_request_bits_address(imem19_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem19_io_bus_response_bits_data)
  );
  DCombinMemPort dmem19 ( // @[top.scala 148:22]
    .clock(dmem19_clock),
    .reset(dmem19_reset),
    .io_pipeline_address(dmem19_io_pipeline_address),
    .io_pipeline_valid(dmem19_io_pipeline_valid),
    .io_pipeline_writedata(dmem19_io_pipeline_writedata),
    .io_pipeline_memread(dmem19_io_pipeline_memread),
    .io_pipeline_memwrite(dmem19_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem19_io_pipeline_maskmode),
    .io_pipeline_sext(dmem19_io_pipeline_sext),
    .io_pipeline_readdata(dmem19_io_pipeline_readdata),
    .io_bus_request_valid(dmem19_io_bus_request_valid),
    .io_bus_request_bits_address(dmem19_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem19_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem19_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem19_io_bus_response_valid),
    .io_bus_response_bits_data(dmem19_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu20 ( // @[top.scala 152:21]
    .clock(cpu20_clock),
    .reset(cpu20_reset),
    .io_imem_address(cpu20_io_imem_address),
    .io_imem_instruction(cpu20_io_imem_instruction),
    .io_dmem_address(cpu20_io_dmem_address),
    .io_dmem_valid(cpu20_io_dmem_valid),
    .io_dmem_writedata(cpu20_io_dmem_writedata),
    .io_dmem_memread(cpu20_io_dmem_memread),
    .io_dmem_memwrite(cpu20_io_dmem_memwrite),
    .io_dmem_maskmode(cpu20_io_dmem_maskmode),
    .io_dmem_sext(cpu20_io_dmem_sext),
    .io_dmem_readdata(cpu20_io_dmem_readdata)
  );
  DualPortedCombinMemory mem20 ( // @[top.scala 153:21]
    .clock(mem20_clock),
    .reset(mem20_reset),
    .io_imem_request_bits_address(mem20_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem20_io_imem_response_bits_data),
    .io_dmem_request_valid(mem20_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem20_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem20_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem20_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem20_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem20_io_dmem_response_bits_data)
  );
  ICombinMemPort imem20 ( // @[top.scala 154:22]
    .io_pipeline_address(imem20_io_pipeline_address),
    .io_pipeline_instruction(imem20_io_pipeline_instruction),
    .io_bus_request_bits_address(imem20_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem20_io_bus_response_bits_data)
  );
  DCombinMemPort dmem20 ( // @[top.scala 155:22]
    .clock(dmem20_clock),
    .reset(dmem20_reset),
    .io_pipeline_address(dmem20_io_pipeline_address),
    .io_pipeline_valid(dmem20_io_pipeline_valid),
    .io_pipeline_writedata(dmem20_io_pipeline_writedata),
    .io_pipeline_memread(dmem20_io_pipeline_memread),
    .io_pipeline_memwrite(dmem20_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem20_io_pipeline_maskmode),
    .io_pipeline_sext(dmem20_io_pipeline_sext),
    .io_pipeline_readdata(dmem20_io_pipeline_readdata),
    .io_bus_request_valid(dmem20_io_bus_request_valid),
    .io_bus_request_bits_address(dmem20_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem20_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem20_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem20_io_bus_response_valid),
    .io_bus_response_bits_data(dmem20_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu21 ( // @[top.scala 159:21]
    .clock(cpu21_clock),
    .reset(cpu21_reset),
    .io_imem_address(cpu21_io_imem_address),
    .io_imem_instruction(cpu21_io_imem_instruction),
    .io_dmem_address(cpu21_io_dmem_address),
    .io_dmem_valid(cpu21_io_dmem_valid),
    .io_dmem_writedata(cpu21_io_dmem_writedata),
    .io_dmem_memread(cpu21_io_dmem_memread),
    .io_dmem_memwrite(cpu21_io_dmem_memwrite),
    .io_dmem_maskmode(cpu21_io_dmem_maskmode),
    .io_dmem_sext(cpu21_io_dmem_sext),
    .io_dmem_readdata(cpu21_io_dmem_readdata)
  );
  DualPortedCombinMemory mem21 ( // @[top.scala 160:21]
    .clock(mem21_clock),
    .reset(mem21_reset),
    .io_imem_request_bits_address(mem21_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem21_io_imem_response_bits_data),
    .io_dmem_request_valid(mem21_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem21_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem21_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem21_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem21_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem21_io_dmem_response_bits_data)
  );
  ICombinMemPort imem21 ( // @[top.scala 161:22]
    .io_pipeline_address(imem21_io_pipeline_address),
    .io_pipeline_instruction(imem21_io_pipeline_instruction),
    .io_bus_request_bits_address(imem21_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem21_io_bus_response_bits_data)
  );
  DCombinMemPort dmem21 ( // @[top.scala 162:22]
    .clock(dmem21_clock),
    .reset(dmem21_reset),
    .io_pipeline_address(dmem21_io_pipeline_address),
    .io_pipeline_valid(dmem21_io_pipeline_valid),
    .io_pipeline_writedata(dmem21_io_pipeline_writedata),
    .io_pipeline_memread(dmem21_io_pipeline_memread),
    .io_pipeline_memwrite(dmem21_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem21_io_pipeline_maskmode),
    .io_pipeline_sext(dmem21_io_pipeline_sext),
    .io_pipeline_readdata(dmem21_io_pipeline_readdata),
    .io_bus_request_valid(dmem21_io_bus_request_valid),
    .io_bus_request_bits_address(dmem21_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem21_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem21_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem21_io_bus_response_valid),
    .io_bus_response_bits_data(dmem21_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu22 ( // @[top.scala 166:21]
    .clock(cpu22_clock),
    .reset(cpu22_reset),
    .io_imem_address(cpu22_io_imem_address),
    .io_imem_instruction(cpu22_io_imem_instruction),
    .io_dmem_address(cpu22_io_dmem_address),
    .io_dmem_valid(cpu22_io_dmem_valid),
    .io_dmem_writedata(cpu22_io_dmem_writedata),
    .io_dmem_memread(cpu22_io_dmem_memread),
    .io_dmem_memwrite(cpu22_io_dmem_memwrite),
    .io_dmem_maskmode(cpu22_io_dmem_maskmode),
    .io_dmem_sext(cpu22_io_dmem_sext),
    .io_dmem_readdata(cpu22_io_dmem_readdata)
  );
  DualPortedCombinMemory mem22 ( // @[top.scala 167:21]
    .clock(mem22_clock),
    .reset(mem22_reset),
    .io_imem_request_bits_address(mem22_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem22_io_imem_response_bits_data),
    .io_dmem_request_valid(mem22_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem22_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem22_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem22_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem22_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem22_io_dmem_response_bits_data)
  );
  ICombinMemPort imem22 ( // @[top.scala 168:22]
    .io_pipeline_address(imem22_io_pipeline_address),
    .io_pipeline_instruction(imem22_io_pipeline_instruction),
    .io_bus_request_bits_address(imem22_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem22_io_bus_response_bits_data)
  );
  DCombinMemPort dmem22 ( // @[top.scala 169:22]
    .clock(dmem22_clock),
    .reset(dmem22_reset),
    .io_pipeline_address(dmem22_io_pipeline_address),
    .io_pipeline_valid(dmem22_io_pipeline_valid),
    .io_pipeline_writedata(dmem22_io_pipeline_writedata),
    .io_pipeline_memread(dmem22_io_pipeline_memread),
    .io_pipeline_memwrite(dmem22_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem22_io_pipeline_maskmode),
    .io_pipeline_sext(dmem22_io_pipeline_sext),
    .io_pipeline_readdata(dmem22_io_pipeline_readdata),
    .io_bus_request_valid(dmem22_io_bus_request_valid),
    .io_bus_request_bits_address(dmem22_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem22_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem22_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem22_io_bus_response_valid),
    .io_bus_response_bits_data(dmem22_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu23 ( // @[top.scala 173:21]
    .clock(cpu23_clock),
    .reset(cpu23_reset),
    .io_imem_address(cpu23_io_imem_address),
    .io_imem_instruction(cpu23_io_imem_instruction),
    .io_dmem_address(cpu23_io_dmem_address),
    .io_dmem_valid(cpu23_io_dmem_valid),
    .io_dmem_writedata(cpu23_io_dmem_writedata),
    .io_dmem_memread(cpu23_io_dmem_memread),
    .io_dmem_memwrite(cpu23_io_dmem_memwrite),
    .io_dmem_maskmode(cpu23_io_dmem_maskmode),
    .io_dmem_sext(cpu23_io_dmem_sext),
    .io_dmem_readdata(cpu23_io_dmem_readdata)
  );
  DualPortedCombinMemory mem23 ( // @[top.scala 174:21]
    .clock(mem23_clock),
    .reset(mem23_reset),
    .io_imem_request_bits_address(mem23_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem23_io_imem_response_bits_data),
    .io_dmem_request_valid(mem23_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem23_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem23_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem23_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem23_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem23_io_dmem_response_bits_data)
  );
  ICombinMemPort imem23 ( // @[top.scala 175:22]
    .io_pipeline_address(imem23_io_pipeline_address),
    .io_pipeline_instruction(imem23_io_pipeline_instruction),
    .io_bus_request_bits_address(imem23_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem23_io_bus_response_bits_data)
  );
  DCombinMemPort dmem23 ( // @[top.scala 176:22]
    .clock(dmem23_clock),
    .reset(dmem23_reset),
    .io_pipeline_address(dmem23_io_pipeline_address),
    .io_pipeline_valid(dmem23_io_pipeline_valid),
    .io_pipeline_writedata(dmem23_io_pipeline_writedata),
    .io_pipeline_memread(dmem23_io_pipeline_memread),
    .io_pipeline_memwrite(dmem23_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem23_io_pipeline_maskmode),
    .io_pipeline_sext(dmem23_io_pipeline_sext),
    .io_pipeline_readdata(dmem23_io_pipeline_readdata),
    .io_bus_request_valid(dmem23_io_bus_request_valid),
    .io_bus_request_bits_address(dmem23_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem23_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem23_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem23_io_bus_response_valid),
    .io_bus_response_bits_data(dmem23_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu24 ( // @[top.scala 180:21]
    .clock(cpu24_clock),
    .reset(cpu24_reset),
    .io_imem_address(cpu24_io_imem_address),
    .io_imem_instruction(cpu24_io_imem_instruction),
    .io_dmem_address(cpu24_io_dmem_address),
    .io_dmem_valid(cpu24_io_dmem_valid),
    .io_dmem_writedata(cpu24_io_dmem_writedata),
    .io_dmem_memread(cpu24_io_dmem_memread),
    .io_dmem_memwrite(cpu24_io_dmem_memwrite),
    .io_dmem_maskmode(cpu24_io_dmem_maskmode),
    .io_dmem_sext(cpu24_io_dmem_sext),
    .io_dmem_readdata(cpu24_io_dmem_readdata)
  );
  DualPortedCombinMemory mem24 ( // @[top.scala 181:21]
    .clock(mem24_clock),
    .reset(mem24_reset),
    .io_imem_request_bits_address(mem24_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem24_io_imem_response_bits_data),
    .io_dmem_request_valid(mem24_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem24_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem24_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem24_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem24_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem24_io_dmem_response_bits_data)
  );
  ICombinMemPort imem24 ( // @[top.scala 182:22]
    .io_pipeline_address(imem24_io_pipeline_address),
    .io_pipeline_instruction(imem24_io_pipeline_instruction),
    .io_bus_request_bits_address(imem24_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem24_io_bus_response_bits_data)
  );
  DCombinMemPort dmem24 ( // @[top.scala 183:22]
    .clock(dmem24_clock),
    .reset(dmem24_reset),
    .io_pipeline_address(dmem24_io_pipeline_address),
    .io_pipeline_valid(dmem24_io_pipeline_valid),
    .io_pipeline_writedata(dmem24_io_pipeline_writedata),
    .io_pipeline_memread(dmem24_io_pipeline_memread),
    .io_pipeline_memwrite(dmem24_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem24_io_pipeline_maskmode),
    .io_pipeline_sext(dmem24_io_pipeline_sext),
    .io_pipeline_readdata(dmem24_io_pipeline_readdata),
    .io_bus_request_valid(dmem24_io_bus_request_valid),
    .io_bus_request_bits_address(dmem24_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem24_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem24_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem24_io_bus_response_valid),
    .io_bus_response_bits_data(dmem24_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu25 ( // @[top.scala 187:21]
    .clock(cpu25_clock),
    .reset(cpu25_reset),
    .io_imem_address(cpu25_io_imem_address),
    .io_imem_instruction(cpu25_io_imem_instruction),
    .io_dmem_address(cpu25_io_dmem_address),
    .io_dmem_valid(cpu25_io_dmem_valid),
    .io_dmem_writedata(cpu25_io_dmem_writedata),
    .io_dmem_memread(cpu25_io_dmem_memread),
    .io_dmem_memwrite(cpu25_io_dmem_memwrite),
    .io_dmem_maskmode(cpu25_io_dmem_maskmode),
    .io_dmem_sext(cpu25_io_dmem_sext),
    .io_dmem_readdata(cpu25_io_dmem_readdata)
  );
  DualPortedCombinMemory mem25 ( // @[top.scala 188:21]
    .clock(mem25_clock),
    .reset(mem25_reset),
    .io_imem_request_bits_address(mem25_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem25_io_imem_response_bits_data),
    .io_dmem_request_valid(mem25_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem25_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem25_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem25_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem25_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem25_io_dmem_response_bits_data)
  );
  ICombinMemPort imem25 ( // @[top.scala 189:22]
    .io_pipeline_address(imem25_io_pipeline_address),
    .io_pipeline_instruction(imem25_io_pipeline_instruction),
    .io_bus_request_bits_address(imem25_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem25_io_bus_response_bits_data)
  );
  DCombinMemPort dmem25 ( // @[top.scala 190:22]
    .clock(dmem25_clock),
    .reset(dmem25_reset),
    .io_pipeline_address(dmem25_io_pipeline_address),
    .io_pipeline_valid(dmem25_io_pipeline_valid),
    .io_pipeline_writedata(dmem25_io_pipeline_writedata),
    .io_pipeline_memread(dmem25_io_pipeline_memread),
    .io_pipeline_memwrite(dmem25_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem25_io_pipeline_maskmode),
    .io_pipeline_sext(dmem25_io_pipeline_sext),
    .io_pipeline_readdata(dmem25_io_pipeline_readdata),
    .io_bus_request_valid(dmem25_io_bus_request_valid),
    .io_bus_request_bits_address(dmem25_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem25_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem25_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem25_io_bus_response_valid),
    .io_bus_response_bits_data(dmem25_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu26 ( // @[top.scala 194:21]
    .clock(cpu26_clock),
    .reset(cpu26_reset),
    .io_imem_address(cpu26_io_imem_address),
    .io_imem_instruction(cpu26_io_imem_instruction),
    .io_dmem_address(cpu26_io_dmem_address),
    .io_dmem_valid(cpu26_io_dmem_valid),
    .io_dmem_writedata(cpu26_io_dmem_writedata),
    .io_dmem_memread(cpu26_io_dmem_memread),
    .io_dmem_memwrite(cpu26_io_dmem_memwrite),
    .io_dmem_maskmode(cpu26_io_dmem_maskmode),
    .io_dmem_sext(cpu26_io_dmem_sext),
    .io_dmem_readdata(cpu26_io_dmem_readdata)
  );
  DualPortedCombinMemory mem26 ( // @[top.scala 195:21]
    .clock(mem26_clock),
    .reset(mem26_reset),
    .io_imem_request_bits_address(mem26_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem26_io_imem_response_bits_data),
    .io_dmem_request_valid(mem26_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem26_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem26_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem26_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem26_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem26_io_dmem_response_bits_data)
  );
  ICombinMemPort imem26 ( // @[top.scala 196:22]
    .io_pipeline_address(imem26_io_pipeline_address),
    .io_pipeline_instruction(imem26_io_pipeline_instruction),
    .io_bus_request_bits_address(imem26_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem26_io_bus_response_bits_data)
  );
  DCombinMemPort dmem26 ( // @[top.scala 197:22]
    .clock(dmem26_clock),
    .reset(dmem26_reset),
    .io_pipeline_address(dmem26_io_pipeline_address),
    .io_pipeline_valid(dmem26_io_pipeline_valid),
    .io_pipeline_writedata(dmem26_io_pipeline_writedata),
    .io_pipeline_memread(dmem26_io_pipeline_memread),
    .io_pipeline_memwrite(dmem26_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem26_io_pipeline_maskmode),
    .io_pipeline_sext(dmem26_io_pipeline_sext),
    .io_pipeline_readdata(dmem26_io_pipeline_readdata),
    .io_bus_request_valid(dmem26_io_bus_request_valid),
    .io_bus_request_bits_address(dmem26_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem26_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem26_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem26_io_bus_response_valid),
    .io_bus_response_bits_data(dmem26_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu27 ( // @[top.scala 201:21]
    .clock(cpu27_clock),
    .reset(cpu27_reset),
    .io_imem_address(cpu27_io_imem_address),
    .io_imem_instruction(cpu27_io_imem_instruction),
    .io_dmem_address(cpu27_io_dmem_address),
    .io_dmem_valid(cpu27_io_dmem_valid),
    .io_dmem_writedata(cpu27_io_dmem_writedata),
    .io_dmem_memread(cpu27_io_dmem_memread),
    .io_dmem_memwrite(cpu27_io_dmem_memwrite),
    .io_dmem_maskmode(cpu27_io_dmem_maskmode),
    .io_dmem_sext(cpu27_io_dmem_sext),
    .io_dmem_readdata(cpu27_io_dmem_readdata)
  );
  DualPortedCombinMemory mem27 ( // @[top.scala 202:21]
    .clock(mem27_clock),
    .reset(mem27_reset),
    .io_imem_request_bits_address(mem27_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem27_io_imem_response_bits_data),
    .io_dmem_request_valid(mem27_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem27_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem27_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem27_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem27_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem27_io_dmem_response_bits_data)
  );
  ICombinMemPort imem27 ( // @[top.scala 203:22]
    .io_pipeline_address(imem27_io_pipeline_address),
    .io_pipeline_instruction(imem27_io_pipeline_instruction),
    .io_bus_request_bits_address(imem27_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem27_io_bus_response_bits_data)
  );
  DCombinMemPort dmem27 ( // @[top.scala 204:22]
    .clock(dmem27_clock),
    .reset(dmem27_reset),
    .io_pipeline_address(dmem27_io_pipeline_address),
    .io_pipeline_valid(dmem27_io_pipeline_valid),
    .io_pipeline_writedata(dmem27_io_pipeline_writedata),
    .io_pipeline_memread(dmem27_io_pipeline_memread),
    .io_pipeline_memwrite(dmem27_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem27_io_pipeline_maskmode),
    .io_pipeline_sext(dmem27_io_pipeline_sext),
    .io_pipeline_readdata(dmem27_io_pipeline_readdata),
    .io_bus_request_valid(dmem27_io_bus_request_valid),
    .io_bus_request_bits_address(dmem27_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem27_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem27_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem27_io_bus_response_valid),
    .io_bus_response_bits_data(dmem27_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu28 ( // @[top.scala 208:21]
    .clock(cpu28_clock),
    .reset(cpu28_reset),
    .io_imem_address(cpu28_io_imem_address),
    .io_imem_instruction(cpu28_io_imem_instruction),
    .io_dmem_address(cpu28_io_dmem_address),
    .io_dmem_valid(cpu28_io_dmem_valid),
    .io_dmem_writedata(cpu28_io_dmem_writedata),
    .io_dmem_memread(cpu28_io_dmem_memread),
    .io_dmem_memwrite(cpu28_io_dmem_memwrite),
    .io_dmem_maskmode(cpu28_io_dmem_maskmode),
    .io_dmem_sext(cpu28_io_dmem_sext),
    .io_dmem_readdata(cpu28_io_dmem_readdata)
  );
  DualPortedCombinMemory mem28 ( // @[top.scala 209:21]
    .clock(mem28_clock),
    .reset(mem28_reset),
    .io_imem_request_bits_address(mem28_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem28_io_imem_response_bits_data),
    .io_dmem_request_valid(mem28_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem28_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem28_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem28_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem28_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem28_io_dmem_response_bits_data)
  );
  ICombinMemPort imem28 ( // @[top.scala 210:22]
    .io_pipeline_address(imem28_io_pipeline_address),
    .io_pipeline_instruction(imem28_io_pipeline_instruction),
    .io_bus_request_bits_address(imem28_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem28_io_bus_response_bits_data)
  );
  DCombinMemPort dmem28 ( // @[top.scala 211:22]
    .clock(dmem28_clock),
    .reset(dmem28_reset),
    .io_pipeline_address(dmem28_io_pipeline_address),
    .io_pipeline_valid(dmem28_io_pipeline_valid),
    .io_pipeline_writedata(dmem28_io_pipeline_writedata),
    .io_pipeline_memread(dmem28_io_pipeline_memread),
    .io_pipeline_memwrite(dmem28_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem28_io_pipeline_maskmode),
    .io_pipeline_sext(dmem28_io_pipeline_sext),
    .io_pipeline_readdata(dmem28_io_pipeline_readdata),
    .io_bus_request_valid(dmem28_io_bus_request_valid),
    .io_bus_request_bits_address(dmem28_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem28_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem28_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem28_io_bus_response_valid),
    .io_bus_response_bits_data(dmem28_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu29 ( // @[top.scala 215:21]
    .clock(cpu29_clock),
    .reset(cpu29_reset),
    .io_imem_address(cpu29_io_imem_address),
    .io_imem_instruction(cpu29_io_imem_instruction),
    .io_dmem_address(cpu29_io_dmem_address),
    .io_dmem_valid(cpu29_io_dmem_valid),
    .io_dmem_writedata(cpu29_io_dmem_writedata),
    .io_dmem_memread(cpu29_io_dmem_memread),
    .io_dmem_memwrite(cpu29_io_dmem_memwrite),
    .io_dmem_maskmode(cpu29_io_dmem_maskmode),
    .io_dmem_sext(cpu29_io_dmem_sext),
    .io_dmem_readdata(cpu29_io_dmem_readdata)
  );
  DualPortedCombinMemory mem29 ( // @[top.scala 216:21]
    .clock(mem29_clock),
    .reset(mem29_reset),
    .io_imem_request_bits_address(mem29_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem29_io_imem_response_bits_data),
    .io_dmem_request_valid(mem29_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem29_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem29_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem29_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem29_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem29_io_dmem_response_bits_data)
  );
  ICombinMemPort imem29 ( // @[top.scala 217:22]
    .io_pipeline_address(imem29_io_pipeline_address),
    .io_pipeline_instruction(imem29_io_pipeline_instruction),
    .io_bus_request_bits_address(imem29_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem29_io_bus_response_bits_data)
  );
  DCombinMemPort dmem29 ( // @[top.scala 218:22]
    .clock(dmem29_clock),
    .reset(dmem29_reset),
    .io_pipeline_address(dmem29_io_pipeline_address),
    .io_pipeline_valid(dmem29_io_pipeline_valid),
    .io_pipeline_writedata(dmem29_io_pipeline_writedata),
    .io_pipeline_memread(dmem29_io_pipeline_memread),
    .io_pipeline_memwrite(dmem29_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem29_io_pipeline_maskmode),
    .io_pipeline_sext(dmem29_io_pipeline_sext),
    .io_pipeline_readdata(dmem29_io_pipeline_readdata),
    .io_bus_request_valid(dmem29_io_bus_request_valid),
    .io_bus_request_bits_address(dmem29_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem29_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem29_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem29_io_bus_response_valid),
    .io_bus_response_bits_data(dmem29_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu30 ( // @[top.scala 222:21]
    .clock(cpu30_clock),
    .reset(cpu30_reset),
    .io_imem_address(cpu30_io_imem_address),
    .io_imem_instruction(cpu30_io_imem_instruction),
    .io_dmem_address(cpu30_io_dmem_address),
    .io_dmem_valid(cpu30_io_dmem_valid),
    .io_dmem_writedata(cpu30_io_dmem_writedata),
    .io_dmem_memread(cpu30_io_dmem_memread),
    .io_dmem_memwrite(cpu30_io_dmem_memwrite),
    .io_dmem_maskmode(cpu30_io_dmem_maskmode),
    .io_dmem_sext(cpu30_io_dmem_sext),
    .io_dmem_readdata(cpu30_io_dmem_readdata)
  );
  DualPortedCombinMemory mem30 ( // @[top.scala 223:21]
    .clock(mem30_clock),
    .reset(mem30_reset),
    .io_imem_request_bits_address(mem30_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem30_io_imem_response_bits_data),
    .io_dmem_request_valid(mem30_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem30_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem30_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem30_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem30_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem30_io_dmem_response_bits_data)
  );
  ICombinMemPort imem30 ( // @[top.scala 224:22]
    .io_pipeline_address(imem30_io_pipeline_address),
    .io_pipeline_instruction(imem30_io_pipeline_instruction),
    .io_bus_request_bits_address(imem30_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem30_io_bus_response_bits_data)
  );
  DCombinMemPort dmem30 ( // @[top.scala 225:22]
    .clock(dmem30_clock),
    .reset(dmem30_reset),
    .io_pipeline_address(dmem30_io_pipeline_address),
    .io_pipeline_valid(dmem30_io_pipeline_valid),
    .io_pipeline_writedata(dmem30_io_pipeline_writedata),
    .io_pipeline_memread(dmem30_io_pipeline_memread),
    .io_pipeline_memwrite(dmem30_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem30_io_pipeline_maskmode),
    .io_pipeline_sext(dmem30_io_pipeline_sext),
    .io_pipeline_readdata(dmem30_io_pipeline_readdata),
    .io_bus_request_valid(dmem30_io_bus_request_valid),
    .io_bus_request_bits_address(dmem30_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem30_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem30_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem30_io_bus_response_valid),
    .io_bus_response_bits_data(dmem30_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu31 ( // @[top.scala 229:21]
    .clock(cpu31_clock),
    .reset(cpu31_reset),
    .io_imem_address(cpu31_io_imem_address),
    .io_imem_instruction(cpu31_io_imem_instruction),
    .io_dmem_address(cpu31_io_dmem_address),
    .io_dmem_valid(cpu31_io_dmem_valid),
    .io_dmem_writedata(cpu31_io_dmem_writedata),
    .io_dmem_memread(cpu31_io_dmem_memread),
    .io_dmem_memwrite(cpu31_io_dmem_memwrite),
    .io_dmem_maskmode(cpu31_io_dmem_maskmode),
    .io_dmem_sext(cpu31_io_dmem_sext),
    .io_dmem_readdata(cpu31_io_dmem_readdata)
  );
  DualPortedCombinMemory mem31 ( // @[top.scala 230:21]
    .clock(mem31_clock),
    .reset(mem31_reset),
    .io_imem_request_bits_address(mem31_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem31_io_imem_response_bits_data),
    .io_dmem_request_valid(mem31_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem31_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem31_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem31_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem31_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem31_io_dmem_response_bits_data)
  );
  ICombinMemPort imem31 ( // @[top.scala 231:22]
    .io_pipeline_address(imem31_io_pipeline_address),
    .io_pipeline_instruction(imem31_io_pipeline_instruction),
    .io_bus_request_bits_address(imem31_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem31_io_bus_response_bits_data)
  );
  DCombinMemPort dmem31 ( // @[top.scala 232:22]
    .clock(dmem31_clock),
    .reset(dmem31_reset),
    .io_pipeline_address(dmem31_io_pipeline_address),
    .io_pipeline_valid(dmem31_io_pipeline_valid),
    .io_pipeline_writedata(dmem31_io_pipeline_writedata),
    .io_pipeline_memread(dmem31_io_pipeline_memread),
    .io_pipeline_memwrite(dmem31_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem31_io_pipeline_maskmode),
    .io_pipeline_sext(dmem31_io_pipeline_sext),
    .io_pipeline_readdata(dmem31_io_pipeline_readdata),
    .io_bus_request_valid(dmem31_io_bus_request_valid),
    .io_bus_request_bits_address(dmem31_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem31_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem31_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem31_io_bus_response_valid),
    .io_bus_response_bits_data(dmem31_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu32 ( // @[top.scala 236:21]
    .clock(cpu32_clock),
    .reset(cpu32_reset),
    .io_imem_address(cpu32_io_imem_address),
    .io_imem_instruction(cpu32_io_imem_instruction),
    .io_dmem_address(cpu32_io_dmem_address),
    .io_dmem_valid(cpu32_io_dmem_valid),
    .io_dmem_writedata(cpu32_io_dmem_writedata),
    .io_dmem_memread(cpu32_io_dmem_memread),
    .io_dmem_memwrite(cpu32_io_dmem_memwrite),
    .io_dmem_maskmode(cpu32_io_dmem_maskmode),
    .io_dmem_sext(cpu32_io_dmem_sext),
    .io_dmem_readdata(cpu32_io_dmem_readdata)
  );
  DualPortedCombinMemory mem32 ( // @[top.scala 237:21]
    .clock(mem32_clock),
    .reset(mem32_reset),
    .io_imem_request_bits_address(mem32_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem32_io_imem_response_bits_data),
    .io_dmem_request_valid(mem32_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem32_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem32_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem32_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem32_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem32_io_dmem_response_bits_data)
  );
  ICombinMemPort imem32 ( // @[top.scala 238:22]
    .io_pipeline_address(imem32_io_pipeline_address),
    .io_pipeline_instruction(imem32_io_pipeline_instruction),
    .io_bus_request_bits_address(imem32_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem32_io_bus_response_bits_data)
  );
  DCombinMemPort dmem32 ( // @[top.scala 239:22]
    .clock(dmem32_clock),
    .reset(dmem32_reset),
    .io_pipeline_address(dmem32_io_pipeline_address),
    .io_pipeline_valid(dmem32_io_pipeline_valid),
    .io_pipeline_writedata(dmem32_io_pipeline_writedata),
    .io_pipeline_memread(dmem32_io_pipeline_memread),
    .io_pipeline_memwrite(dmem32_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem32_io_pipeline_maskmode),
    .io_pipeline_sext(dmem32_io_pipeline_sext),
    .io_pipeline_readdata(dmem32_io_pipeline_readdata),
    .io_bus_request_valid(dmem32_io_bus_request_valid),
    .io_bus_request_bits_address(dmem32_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem32_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem32_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem32_io_bus_response_valid),
    .io_bus_response_bits_data(dmem32_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu33 ( // @[top.scala 243:21]
    .clock(cpu33_clock),
    .reset(cpu33_reset),
    .io_imem_address(cpu33_io_imem_address),
    .io_imem_instruction(cpu33_io_imem_instruction),
    .io_dmem_address(cpu33_io_dmem_address),
    .io_dmem_valid(cpu33_io_dmem_valid),
    .io_dmem_writedata(cpu33_io_dmem_writedata),
    .io_dmem_memread(cpu33_io_dmem_memread),
    .io_dmem_memwrite(cpu33_io_dmem_memwrite),
    .io_dmem_maskmode(cpu33_io_dmem_maskmode),
    .io_dmem_sext(cpu33_io_dmem_sext),
    .io_dmem_readdata(cpu33_io_dmem_readdata)
  );
  DualPortedCombinMemory mem33 ( // @[top.scala 244:21]
    .clock(mem33_clock),
    .reset(mem33_reset),
    .io_imem_request_bits_address(mem33_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem33_io_imem_response_bits_data),
    .io_dmem_request_valid(mem33_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem33_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem33_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem33_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem33_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem33_io_dmem_response_bits_data)
  );
  ICombinMemPort imem33 ( // @[top.scala 245:22]
    .io_pipeline_address(imem33_io_pipeline_address),
    .io_pipeline_instruction(imem33_io_pipeline_instruction),
    .io_bus_request_bits_address(imem33_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem33_io_bus_response_bits_data)
  );
  DCombinMemPort dmem33 ( // @[top.scala 246:22]
    .clock(dmem33_clock),
    .reset(dmem33_reset),
    .io_pipeline_address(dmem33_io_pipeline_address),
    .io_pipeline_valid(dmem33_io_pipeline_valid),
    .io_pipeline_writedata(dmem33_io_pipeline_writedata),
    .io_pipeline_memread(dmem33_io_pipeline_memread),
    .io_pipeline_memwrite(dmem33_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem33_io_pipeline_maskmode),
    .io_pipeline_sext(dmem33_io_pipeline_sext),
    .io_pipeline_readdata(dmem33_io_pipeline_readdata),
    .io_bus_request_valid(dmem33_io_bus_request_valid),
    .io_bus_request_bits_address(dmem33_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem33_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem33_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem33_io_bus_response_valid),
    .io_bus_response_bits_data(dmem33_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu34 ( // @[top.scala 250:21]
    .clock(cpu34_clock),
    .reset(cpu34_reset),
    .io_imem_address(cpu34_io_imem_address),
    .io_imem_instruction(cpu34_io_imem_instruction),
    .io_dmem_address(cpu34_io_dmem_address),
    .io_dmem_valid(cpu34_io_dmem_valid),
    .io_dmem_writedata(cpu34_io_dmem_writedata),
    .io_dmem_memread(cpu34_io_dmem_memread),
    .io_dmem_memwrite(cpu34_io_dmem_memwrite),
    .io_dmem_maskmode(cpu34_io_dmem_maskmode),
    .io_dmem_sext(cpu34_io_dmem_sext),
    .io_dmem_readdata(cpu34_io_dmem_readdata)
  );
  DualPortedCombinMemory mem34 ( // @[top.scala 251:21]
    .clock(mem34_clock),
    .reset(mem34_reset),
    .io_imem_request_bits_address(mem34_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem34_io_imem_response_bits_data),
    .io_dmem_request_valid(mem34_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem34_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem34_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem34_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem34_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem34_io_dmem_response_bits_data)
  );
  ICombinMemPort imem34 ( // @[top.scala 252:22]
    .io_pipeline_address(imem34_io_pipeline_address),
    .io_pipeline_instruction(imem34_io_pipeline_instruction),
    .io_bus_request_bits_address(imem34_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem34_io_bus_response_bits_data)
  );
  DCombinMemPort dmem34 ( // @[top.scala 253:22]
    .clock(dmem34_clock),
    .reset(dmem34_reset),
    .io_pipeline_address(dmem34_io_pipeline_address),
    .io_pipeline_valid(dmem34_io_pipeline_valid),
    .io_pipeline_writedata(dmem34_io_pipeline_writedata),
    .io_pipeline_memread(dmem34_io_pipeline_memread),
    .io_pipeline_memwrite(dmem34_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem34_io_pipeline_maskmode),
    .io_pipeline_sext(dmem34_io_pipeline_sext),
    .io_pipeline_readdata(dmem34_io_pipeline_readdata),
    .io_bus_request_valid(dmem34_io_bus_request_valid),
    .io_bus_request_bits_address(dmem34_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem34_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem34_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem34_io_bus_response_valid),
    .io_bus_response_bits_data(dmem34_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu35 ( // @[top.scala 257:21]
    .clock(cpu35_clock),
    .reset(cpu35_reset),
    .io_imem_address(cpu35_io_imem_address),
    .io_imem_instruction(cpu35_io_imem_instruction),
    .io_dmem_address(cpu35_io_dmem_address),
    .io_dmem_valid(cpu35_io_dmem_valid),
    .io_dmem_writedata(cpu35_io_dmem_writedata),
    .io_dmem_memread(cpu35_io_dmem_memread),
    .io_dmem_memwrite(cpu35_io_dmem_memwrite),
    .io_dmem_maskmode(cpu35_io_dmem_maskmode),
    .io_dmem_sext(cpu35_io_dmem_sext),
    .io_dmem_readdata(cpu35_io_dmem_readdata)
  );
  DualPortedCombinMemory mem35 ( // @[top.scala 258:21]
    .clock(mem35_clock),
    .reset(mem35_reset),
    .io_imem_request_bits_address(mem35_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem35_io_imem_response_bits_data),
    .io_dmem_request_valid(mem35_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem35_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem35_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem35_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem35_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem35_io_dmem_response_bits_data)
  );
  ICombinMemPort imem35 ( // @[top.scala 259:22]
    .io_pipeline_address(imem35_io_pipeline_address),
    .io_pipeline_instruction(imem35_io_pipeline_instruction),
    .io_bus_request_bits_address(imem35_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem35_io_bus_response_bits_data)
  );
  DCombinMemPort dmem35 ( // @[top.scala 260:22]
    .clock(dmem35_clock),
    .reset(dmem35_reset),
    .io_pipeline_address(dmem35_io_pipeline_address),
    .io_pipeline_valid(dmem35_io_pipeline_valid),
    .io_pipeline_writedata(dmem35_io_pipeline_writedata),
    .io_pipeline_memread(dmem35_io_pipeline_memread),
    .io_pipeline_memwrite(dmem35_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem35_io_pipeline_maskmode),
    .io_pipeline_sext(dmem35_io_pipeline_sext),
    .io_pipeline_readdata(dmem35_io_pipeline_readdata),
    .io_bus_request_valid(dmem35_io_bus_request_valid),
    .io_bus_request_bits_address(dmem35_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem35_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem35_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem35_io_bus_response_valid),
    .io_bus_response_bits_data(dmem35_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu36 ( // @[top.scala 264:21]
    .clock(cpu36_clock),
    .reset(cpu36_reset),
    .io_imem_address(cpu36_io_imem_address),
    .io_imem_instruction(cpu36_io_imem_instruction),
    .io_dmem_address(cpu36_io_dmem_address),
    .io_dmem_valid(cpu36_io_dmem_valid),
    .io_dmem_writedata(cpu36_io_dmem_writedata),
    .io_dmem_memread(cpu36_io_dmem_memread),
    .io_dmem_memwrite(cpu36_io_dmem_memwrite),
    .io_dmem_maskmode(cpu36_io_dmem_maskmode),
    .io_dmem_sext(cpu36_io_dmem_sext),
    .io_dmem_readdata(cpu36_io_dmem_readdata)
  );
  DualPortedCombinMemory mem36 ( // @[top.scala 265:21]
    .clock(mem36_clock),
    .reset(mem36_reset),
    .io_imem_request_bits_address(mem36_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem36_io_imem_response_bits_data),
    .io_dmem_request_valid(mem36_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem36_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem36_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem36_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem36_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem36_io_dmem_response_bits_data)
  );
  ICombinMemPort imem36 ( // @[top.scala 266:22]
    .io_pipeline_address(imem36_io_pipeline_address),
    .io_pipeline_instruction(imem36_io_pipeline_instruction),
    .io_bus_request_bits_address(imem36_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem36_io_bus_response_bits_data)
  );
  DCombinMemPort dmem36 ( // @[top.scala 267:22]
    .clock(dmem36_clock),
    .reset(dmem36_reset),
    .io_pipeline_address(dmem36_io_pipeline_address),
    .io_pipeline_valid(dmem36_io_pipeline_valid),
    .io_pipeline_writedata(dmem36_io_pipeline_writedata),
    .io_pipeline_memread(dmem36_io_pipeline_memread),
    .io_pipeline_memwrite(dmem36_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem36_io_pipeline_maskmode),
    .io_pipeline_sext(dmem36_io_pipeline_sext),
    .io_pipeline_readdata(dmem36_io_pipeline_readdata),
    .io_bus_request_valid(dmem36_io_bus_request_valid),
    .io_bus_request_bits_address(dmem36_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem36_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem36_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem36_io_bus_response_valid),
    .io_bus_response_bits_data(dmem36_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu37 ( // @[top.scala 271:21]
    .clock(cpu37_clock),
    .reset(cpu37_reset),
    .io_imem_address(cpu37_io_imem_address),
    .io_imem_instruction(cpu37_io_imem_instruction),
    .io_dmem_address(cpu37_io_dmem_address),
    .io_dmem_valid(cpu37_io_dmem_valid),
    .io_dmem_writedata(cpu37_io_dmem_writedata),
    .io_dmem_memread(cpu37_io_dmem_memread),
    .io_dmem_memwrite(cpu37_io_dmem_memwrite),
    .io_dmem_maskmode(cpu37_io_dmem_maskmode),
    .io_dmem_sext(cpu37_io_dmem_sext),
    .io_dmem_readdata(cpu37_io_dmem_readdata)
  );
  DualPortedCombinMemory mem37 ( // @[top.scala 272:21]
    .clock(mem37_clock),
    .reset(mem37_reset),
    .io_imem_request_bits_address(mem37_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem37_io_imem_response_bits_data),
    .io_dmem_request_valid(mem37_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem37_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem37_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem37_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem37_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem37_io_dmem_response_bits_data)
  );
  ICombinMemPort imem37 ( // @[top.scala 273:22]
    .io_pipeline_address(imem37_io_pipeline_address),
    .io_pipeline_instruction(imem37_io_pipeline_instruction),
    .io_bus_request_bits_address(imem37_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem37_io_bus_response_bits_data)
  );
  DCombinMemPort dmem37 ( // @[top.scala 274:22]
    .clock(dmem37_clock),
    .reset(dmem37_reset),
    .io_pipeline_address(dmem37_io_pipeline_address),
    .io_pipeline_valid(dmem37_io_pipeline_valid),
    .io_pipeline_writedata(dmem37_io_pipeline_writedata),
    .io_pipeline_memread(dmem37_io_pipeline_memread),
    .io_pipeline_memwrite(dmem37_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem37_io_pipeline_maskmode),
    .io_pipeline_sext(dmem37_io_pipeline_sext),
    .io_pipeline_readdata(dmem37_io_pipeline_readdata),
    .io_bus_request_valid(dmem37_io_bus_request_valid),
    .io_bus_request_bits_address(dmem37_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem37_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem37_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem37_io_bus_response_valid),
    .io_bus_response_bits_data(dmem37_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu38 ( // @[top.scala 278:21]
    .clock(cpu38_clock),
    .reset(cpu38_reset),
    .io_imem_address(cpu38_io_imem_address),
    .io_imem_instruction(cpu38_io_imem_instruction),
    .io_dmem_address(cpu38_io_dmem_address),
    .io_dmem_valid(cpu38_io_dmem_valid),
    .io_dmem_writedata(cpu38_io_dmem_writedata),
    .io_dmem_memread(cpu38_io_dmem_memread),
    .io_dmem_memwrite(cpu38_io_dmem_memwrite),
    .io_dmem_maskmode(cpu38_io_dmem_maskmode),
    .io_dmem_sext(cpu38_io_dmem_sext),
    .io_dmem_readdata(cpu38_io_dmem_readdata)
  );
  DualPortedCombinMemory mem38 ( // @[top.scala 279:21]
    .clock(mem38_clock),
    .reset(mem38_reset),
    .io_imem_request_bits_address(mem38_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem38_io_imem_response_bits_data),
    .io_dmem_request_valid(mem38_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem38_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem38_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem38_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem38_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem38_io_dmem_response_bits_data)
  );
  ICombinMemPort imem38 ( // @[top.scala 280:22]
    .io_pipeline_address(imem38_io_pipeline_address),
    .io_pipeline_instruction(imem38_io_pipeline_instruction),
    .io_bus_request_bits_address(imem38_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem38_io_bus_response_bits_data)
  );
  DCombinMemPort dmem38 ( // @[top.scala 281:22]
    .clock(dmem38_clock),
    .reset(dmem38_reset),
    .io_pipeline_address(dmem38_io_pipeline_address),
    .io_pipeline_valid(dmem38_io_pipeline_valid),
    .io_pipeline_writedata(dmem38_io_pipeline_writedata),
    .io_pipeline_memread(dmem38_io_pipeline_memread),
    .io_pipeline_memwrite(dmem38_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem38_io_pipeline_maskmode),
    .io_pipeline_sext(dmem38_io_pipeline_sext),
    .io_pipeline_readdata(dmem38_io_pipeline_readdata),
    .io_bus_request_valid(dmem38_io_bus_request_valid),
    .io_bus_request_bits_address(dmem38_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem38_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem38_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem38_io_bus_response_valid),
    .io_bus_response_bits_data(dmem38_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu39 ( // @[top.scala 285:21]
    .clock(cpu39_clock),
    .reset(cpu39_reset),
    .io_imem_address(cpu39_io_imem_address),
    .io_imem_instruction(cpu39_io_imem_instruction),
    .io_dmem_address(cpu39_io_dmem_address),
    .io_dmem_valid(cpu39_io_dmem_valid),
    .io_dmem_writedata(cpu39_io_dmem_writedata),
    .io_dmem_memread(cpu39_io_dmem_memread),
    .io_dmem_memwrite(cpu39_io_dmem_memwrite),
    .io_dmem_maskmode(cpu39_io_dmem_maskmode),
    .io_dmem_sext(cpu39_io_dmem_sext),
    .io_dmem_readdata(cpu39_io_dmem_readdata)
  );
  DualPortedCombinMemory mem39 ( // @[top.scala 286:21]
    .clock(mem39_clock),
    .reset(mem39_reset),
    .io_imem_request_bits_address(mem39_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem39_io_imem_response_bits_data),
    .io_dmem_request_valid(mem39_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem39_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem39_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem39_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem39_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem39_io_dmem_response_bits_data)
  );
  ICombinMemPort imem39 ( // @[top.scala 287:22]
    .io_pipeline_address(imem39_io_pipeline_address),
    .io_pipeline_instruction(imem39_io_pipeline_instruction),
    .io_bus_request_bits_address(imem39_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem39_io_bus_response_bits_data)
  );
  DCombinMemPort dmem39 ( // @[top.scala 288:22]
    .clock(dmem39_clock),
    .reset(dmem39_reset),
    .io_pipeline_address(dmem39_io_pipeline_address),
    .io_pipeline_valid(dmem39_io_pipeline_valid),
    .io_pipeline_writedata(dmem39_io_pipeline_writedata),
    .io_pipeline_memread(dmem39_io_pipeline_memread),
    .io_pipeline_memwrite(dmem39_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem39_io_pipeline_maskmode),
    .io_pipeline_sext(dmem39_io_pipeline_sext),
    .io_pipeline_readdata(dmem39_io_pipeline_readdata),
    .io_bus_request_valid(dmem39_io_bus_request_valid),
    .io_bus_request_bits_address(dmem39_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem39_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem39_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem39_io_bus_response_valid),
    .io_bus_response_bits_data(dmem39_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu40 ( // @[top.scala 292:21]
    .clock(cpu40_clock),
    .reset(cpu40_reset),
    .io_imem_address(cpu40_io_imem_address),
    .io_imem_instruction(cpu40_io_imem_instruction),
    .io_dmem_address(cpu40_io_dmem_address),
    .io_dmem_valid(cpu40_io_dmem_valid),
    .io_dmem_writedata(cpu40_io_dmem_writedata),
    .io_dmem_memread(cpu40_io_dmem_memread),
    .io_dmem_memwrite(cpu40_io_dmem_memwrite),
    .io_dmem_maskmode(cpu40_io_dmem_maskmode),
    .io_dmem_sext(cpu40_io_dmem_sext),
    .io_dmem_readdata(cpu40_io_dmem_readdata)
  );
  DualPortedCombinMemory mem40 ( // @[top.scala 293:21]
    .clock(mem40_clock),
    .reset(mem40_reset),
    .io_imem_request_bits_address(mem40_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem40_io_imem_response_bits_data),
    .io_dmem_request_valid(mem40_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem40_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem40_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem40_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem40_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem40_io_dmem_response_bits_data)
  );
  ICombinMemPort imem40 ( // @[top.scala 294:22]
    .io_pipeline_address(imem40_io_pipeline_address),
    .io_pipeline_instruction(imem40_io_pipeline_instruction),
    .io_bus_request_bits_address(imem40_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem40_io_bus_response_bits_data)
  );
  DCombinMemPort dmem40 ( // @[top.scala 295:22]
    .clock(dmem40_clock),
    .reset(dmem40_reset),
    .io_pipeline_address(dmem40_io_pipeline_address),
    .io_pipeline_valid(dmem40_io_pipeline_valid),
    .io_pipeline_writedata(dmem40_io_pipeline_writedata),
    .io_pipeline_memread(dmem40_io_pipeline_memread),
    .io_pipeline_memwrite(dmem40_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem40_io_pipeline_maskmode),
    .io_pipeline_sext(dmem40_io_pipeline_sext),
    .io_pipeline_readdata(dmem40_io_pipeline_readdata),
    .io_bus_request_valid(dmem40_io_bus_request_valid),
    .io_bus_request_bits_address(dmem40_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem40_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem40_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem40_io_bus_response_valid),
    .io_bus_response_bits_data(dmem40_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu41 ( // @[top.scala 299:21]
    .clock(cpu41_clock),
    .reset(cpu41_reset),
    .io_imem_address(cpu41_io_imem_address),
    .io_imem_instruction(cpu41_io_imem_instruction),
    .io_dmem_address(cpu41_io_dmem_address),
    .io_dmem_valid(cpu41_io_dmem_valid),
    .io_dmem_writedata(cpu41_io_dmem_writedata),
    .io_dmem_memread(cpu41_io_dmem_memread),
    .io_dmem_memwrite(cpu41_io_dmem_memwrite),
    .io_dmem_maskmode(cpu41_io_dmem_maskmode),
    .io_dmem_sext(cpu41_io_dmem_sext),
    .io_dmem_readdata(cpu41_io_dmem_readdata)
  );
  DualPortedCombinMemory mem41 ( // @[top.scala 300:21]
    .clock(mem41_clock),
    .reset(mem41_reset),
    .io_imem_request_bits_address(mem41_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem41_io_imem_response_bits_data),
    .io_dmem_request_valid(mem41_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem41_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem41_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem41_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem41_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem41_io_dmem_response_bits_data)
  );
  ICombinMemPort imem41 ( // @[top.scala 301:22]
    .io_pipeline_address(imem41_io_pipeline_address),
    .io_pipeline_instruction(imem41_io_pipeline_instruction),
    .io_bus_request_bits_address(imem41_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem41_io_bus_response_bits_data)
  );
  DCombinMemPort dmem41 ( // @[top.scala 302:22]
    .clock(dmem41_clock),
    .reset(dmem41_reset),
    .io_pipeline_address(dmem41_io_pipeline_address),
    .io_pipeline_valid(dmem41_io_pipeline_valid),
    .io_pipeline_writedata(dmem41_io_pipeline_writedata),
    .io_pipeline_memread(dmem41_io_pipeline_memread),
    .io_pipeline_memwrite(dmem41_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem41_io_pipeline_maskmode),
    .io_pipeline_sext(dmem41_io_pipeline_sext),
    .io_pipeline_readdata(dmem41_io_pipeline_readdata),
    .io_bus_request_valid(dmem41_io_bus_request_valid),
    .io_bus_request_bits_address(dmem41_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem41_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem41_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem41_io_bus_response_valid),
    .io_bus_response_bits_data(dmem41_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu42 ( // @[top.scala 306:21]
    .clock(cpu42_clock),
    .reset(cpu42_reset),
    .io_imem_address(cpu42_io_imem_address),
    .io_imem_instruction(cpu42_io_imem_instruction),
    .io_dmem_address(cpu42_io_dmem_address),
    .io_dmem_valid(cpu42_io_dmem_valid),
    .io_dmem_writedata(cpu42_io_dmem_writedata),
    .io_dmem_memread(cpu42_io_dmem_memread),
    .io_dmem_memwrite(cpu42_io_dmem_memwrite),
    .io_dmem_maskmode(cpu42_io_dmem_maskmode),
    .io_dmem_sext(cpu42_io_dmem_sext),
    .io_dmem_readdata(cpu42_io_dmem_readdata)
  );
  DualPortedCombinMemory mem42 ( // @[top.scala 307:21]
    .clock(mem42_clock),
    .reset(mem42_reset),
    .io_imem_request_bits_address(mem42_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem42_io_imem_response_bits_data),
    .io_dmem_request_valid(mem42_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem42_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem42_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem42_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem42_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem42_io_dmem_response_bits_data)
  );
  ICombinMemPort imem42 ( // @[top.scala 308:22]
    .io_pipeline_address(imem42_io_pipeline_address),
    .io_pipeline_instruction(imem42_io_pipeline_instruction),
    .io_bus_request_bits_address(imem42_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem42_io_bus_response_bits_data)
  );
  DCombinMemPort dmem42 ( // @[top.scala 309:22]
    .clock(dmem42_clock),
    .reset(dmem42_reset),
    .io_pipeline_address(dmem42_io_pipeline_address),
    .io_pipeline_valid(dmem42_io_pipeline_valid),
    .io_pipeline_writedata(dmem42_io_pipeline_writedata),
    .io_pipeline_memread(dmem42_io_pipeline_memread),
    .io_pipeline_memwrite(dmem42_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem42_io_pipeline_maskmode),
    .io_pipeline_sext(dmem42_io_pipeline_sext),
    .io_pipeline_readdata(dmem42_io_pipeline_readdata),
    .io_bus_request_valid(dmem42_io_bus_request_valid),
    .io_bus_request_bits_address(dmem42_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem42_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem42_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem42_io_bus_response_valid),
    .io_bus_response_bits_data(dmem42_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu43 ( // @[top.scala 313:21]
    .clock(cpu43_clock),
    .reset(cpu43_reset),
    .io_imem_address(cpu43_io_imem_address),
    .io_imem_instruction(cpu43_io_imem_instruction),
    .io_dmem_address(cpu43_io_dmem_address),
    .io_dmem_valid(cpu43_io_dmem_valid),
    .io_dmem_writedata(cpu43_io_dmem_writedata),
    .io_dmem_memread(cpu43_io_dmem_memread),
    .io_dmem_memwrite(cpu43_io_dmem_memwrite),
    .io_dmem_maskmode(cpu43_io_dmem_maskmode),
    .io_dmem_sext(cpu43_io_dmem_sext),
    .io_dmem_readdata(cpu43_io_dmem_readdata)
  );
  DualPortedCombinMemory mem43 ( // @[top.scala 314:21]
    .clock(mem43_clock),
    .reset(mem43_reset),
    .io_imem_request_bits_address(mem43_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem43_io_imem_response_bits_data),
    .io_dmem_request_valid(mem43_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem43_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem43_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem43_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem43_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem43_io_dmem_response_bits_data)
  );
  ICombinMemPort imem43 ( // @[top.scala 315:22]
    .io_pipeline_address(imem43_io_pipeline_address),
    .io_pipeline_instruction(imem43_io_pipeline_instruction),
    .io_bus_request_bits_address(imem43_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem43_io_bus_response_bits_data)
  );
  DCombinMemPort dmem43 ( // @[top.scala 316:22]
    .clock(dmem43_clock),
    .reset(dmem43_reset),
    .io_pipeline_address(dmem43_io_pipeline_address),
    .io_pipeline_valid(dmem43_io_pipeline_valid),
    .io_pipeline_writedata(dmem43_io_pipeline_writedata),
    .io_pipeline_memread(dmem43_io_pipeline_memread),
    .io_pipeline_memwrite(dmem43_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem43_io_pipeline_maskmode),
    .io_pipeline_sext(dmem43_io_pipeline_sext),
    .io_pipeline_readdata(dmem43_io_pipeline_readdata),
    .io_bus_request_valid(dmem43_io_bus_request_valid),
    .io_bus_request_bits_address(dmem43_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem43_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem43_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem43_io_bus_response_valid),
    .io_bus_response_bits_data(dmem43_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu44 ( // @[top.scala 320:21]
    .clock(cpu44_clock),
    .reset(cpu44_reset),
    .io_imem_address(cpu44_io_imem_address),
    .io_imem_instruction(cpu44_io_imem_instruction),
    .io_dmem_address(cpu44_io_dmem_address),
    .io_dmem_valid(cpu44_io_dmem_valid),
    .io_dmem_writedata(cpu44_io_dmem_writedata),
    .io_dmem_memread(cpu44_io_dmem_memread),
    .io_dmem_memwrite(cpu44_io_dmem_memwrite),
    .io_dmem_maskmode(cpu44_io_dmem_maskmode),
    .io_dmem_sext(cpu44_io_dmem_sext),
    .io_dmem_readdata(cpu44_io_dmem_readdata)
  );
  DualPortedCombinMemory mem44 ( // @[top.scala 321:21]
    .clock(mem44_clock),
    .reset(mem44_reset),
    .io_imem_request_bits_address(mem44_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem44_io_imem_response_bits_data),
    .io_dmem_request_valid(mem44_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem44_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem44_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem44_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem44_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem44_io_dmem_response_bits_data)
  );
  ICombinMemPort imem44 ( // @[top.scala 322:22]
    .io_pipeline_address(imem44_io_pipeline_address),
    .io_pipeline_instruction(imem44_io_pipeline_instruction),
    .io_bus_request_bits_address(imem44_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem44_io_bus_response_bits_data)
  );
  DCombinMemPort dmem44 ( // @[top.scala 323:22]
    .clock(dmem44_clock),
    .reset(dmem44_reset),
    .io_pipeline_address(dmem44_io_pipeline_address),
    .io_pipeline_valid(dmem44_io_pipeline_valid),
    .io_pipeline_writedata(dmem44_io_pipeline_writedata),
    .io_pipeline_memread(dmem44_io_pipeline_memread),
    .io_pipeline_memwrite(dmem44_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem44_io_pipeline_maskmode),
    .io_pipeline_sext(dmem44_io_pipeline_sext),
    .io_pipeline_readdata(dmem44_io_pipeline_readdata),
    .io_bus_request_valid(dmem44_io_bus_request_valid),
    .io_bus_request_bits_address(dmem44_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem44_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem44_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem44_io_bus_response_valid),
    .io_bus_response_bits_data(dmem44_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu45 ( // @[top.scala 327:21]
    .clock(cpu45_clock),
    .reset(cpu45_reset),
    .io_imem_address(cpu45_io_imem_address),
    .io_imem_instruction(cpu45_io_imem_instruction),
    .io_dmem_address(cpu45_io_dmem_address),
    .io_dmem_valid(cpu45_io_dmem_valid),
    .io_dmem_writedata(cpu45_io_dmem_writedata),
    .io_dmem_memread(cpu45_io_dmem_memread),
    .io_dmem_memwrite(cpu45_io_dmem_memwrite),
    .io_dmem_maskmode(cpu45_io_dmem_maskmode),
    .io_dmem_sext(cpu45_io_dmem_sext),
    .io_dmem_readdata(cpu45_io_dmem_readdata)
  );
  DualPortedCombinMemory mem45 ( // @[top.scala 328:21]
    .clock(mem45_clock),
    .reset(mem45_reset),
    .io_imem_request_bits_address(mem45_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem45_io_imem_response_bits_data),
    .io_dmem_request_valid(mem45_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem45_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem45_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem45_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem45_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem45_io_dmem_response_bits_data)
  );
  ICombinMemPort imem45 ( // @[top.scala 329:22]
    .io_pipeline_address(imem45_io_pipeline_address),
    .io_pipeline_instruction(imem45_io_pipeline_instruction),
    .io_bus_request_bits_address(imem45_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem45_io_bus_response_bits_data)
  );
  DCombinMemPort dmem45 ( // @[top.scala 330:22]
    .clock(dmem45_clock),
    .reset(dmem45_reset),
    .io_pipeline_address(dmem45_io_pipeline_address),
    .io_pipeline_valid(dmem45_io_pipeline_valid),
    .io_pipeline_writedata(dmem45_io_pipeline_writedata),
    .io_pipeline_memread(dmem45_io_pipeline_memread),
    .io_pipeline_memwrite(dmem45_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem45_io_pipeline_maskmode),
    .io_pipeline_sext(dmem45_io_pipeline_sext),
    .io_pipeline_readdata(dmem45_io_pipeline_readdata),
    .io_bus_request_valid(dmem45_io_bus_request_valid),
    .io_bus_request_bits_address(dmem45_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem45_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem45_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem45_io_bus_response_valid),
    .io_bus_response_bits_data(dmem45_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu46 ( // @[top.scala 334:21]
    .clock(cpu46_clock),
    .reset(cpu46_reset),
    .io_imem_address(cpu46_io_imem_address),
    .io_imem_instruction(cpu46_io_imem_instruction),
    .io_dmem_address(cpu46_io_dmem_address),
    .io_dmem_valid(cpu46_io_dmem_valid),
    .io_dmem_writedata(cpu46_io_dmem_writedata),
    .io_dmem_memread(cpu46_io_dmem_memread),
    .io_dmem_memwrite(cpu46_io_dmem_memwrite),
    .io_dmem_maskmode(cpu46_io_dmem_maskmode),
    .io_dmem_sext(cpu46_io_dmem_sext),
    .io_dmem_readdata(cpu46_io_dmem_readdata)
  );
  DualPortedCombinMemory mem46 ( // @[top.scala 335:21]
    .clock(mem46_clock),
    .reset(mem46_reset),
    .io_imem_request_bits_address(mem46_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem46_io_imem_response_bits_data),
    .io_dmem_request_valid(mem46_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem46_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem46_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem46_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem46_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem46_io_dmem_response_bits_data)
  );
  ICombinMemPort imem46 ( // @[top.scala 336:22]
    .io_pipeline_address(imem46_io_pipeline_address),
    .io_pipeline_instruction(imem46_io_pipeline_instruction),
    .io_bus_request_bits_address(imem46_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem46_io_bus_response_bits_data)
  );
  DCombinMemPort dmem46 ( // @[top.scala 337:22]
    .clock(dmem46_clock),
    .reset(dmem46_reset),
    .io_pipeline_address(dmem46_io_pipeline_address),
    .io_pipeline_valid(dmem46_io_pipeline_valid),
    .io_pipeline_writedata(dmem46_io_pipeline_writedata),
    .io_pipeline_memread(dmem46_io_pipeline_memread),
    .io_pipeline_memwrite(dmem46_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem46_io_pipeline_maskmode),
    .io_pipeline_sext(dmem46_io_pipeline_sext),
    .io_pipeline_readdata(dmem46_io_pipeline_readdata),
    .io_bus_request_valid(dmem46_io_bus_request_valid),
    .io_bus_request_bits_address(dmem46_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem46_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem46_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem46_io_bus_response_valid),
    .io_bus_response_bits_data(dmem46_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu47 ( // @[top.scala 341:21]
    .clock(cpu47_clock),
    .reset(cpu47_reset),
    .io_imem_address(cpu47_io_imem_address),
    .io_imem_instruction(cpu47_io_imem_instruction),
    .io_dmem_address(cpu47_io_dmem_address),
    .io_dmem_valid(cpu47_io_dmem_valid),
    .io_dmem_writedata(cpu47_io_dmem_writedata),
    .io_dmem_memread(cpu47_io_dmem_memread),
    .io_dmem_memwrite(cpu47_io_dmem_memwrite),
    .io_dmem_maskmode(cpu47_io_dmem_maskmode),
    .io_dmem_sext(cpu47_io_dmem_sext),
    .io_dmem_readdata(cpu47_io_dmem_readdata)
  );
  DualPortedCombinMemory mem47 ( // @[top.scala 342:21]
    .clock(mem47_clock),
    .reset(mem47_reset),
    .io_imem_request_bits_address(mem47_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem47_io_imem_response_bits_data),
    .io_dmem_request_valid(mem47_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem47_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem47_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem47_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem47_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem47_io_dmem_response_bits_data)
  );
  ICombinMemPort imem47 ( // @[top.scala 343:22]
    .io_pipeline_address(imem47_io_pipeline_address),
    .io_pipeline_instruction(imem47_io_pipeline_instruction),
    .io_bus_request_bits_address(imem47_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem47_io_bus_response_bits_data)
  );
  DCombinMemPort dmem47 ( // @[top.scala 344:22]
    .clock(dmem47_clock),
    .reset(dmem47_reset),
    .io_pipeline_address(dmem47_io_pipeline_address),
    .io_pipeline_valid(dmem47_io_pipeline_valid),
    .io_pipeline_writedata(dmem47_io_pipeline_writedata),
    .io_pipeline_memread(dmem47_io_pipeline_memread),
    .io_pipeline_memwrite(dmem47_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem47_io_pipeline_maskmode),
    .io_pipeline_sext(dmem47_io_pipeline_sext),
    .io_pipeline_readdata(dmem47_io_pipeline_readdata),
    .io_bus_request_valid(dmem47_io_bus_request_valid),
    .io_bus_request_bits_address(dmem47_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem47_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem47_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem47_io_bus_response_valid),
    .io_bus_response_bits_data(dmem47_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu48 ( // @[top.scala 348:21]
    .clock(cpu48_clock),
    .reset(cpu48_reset),
    .io_imem_address(cpu48_io_imem_address),
    .io_imem_instruction(cpu48_io_imem_instruction),
    .io_dmem_address(cpu48_io_dmem_address),
    .io_dmem_valid(cpu48_io_dmem_valid),
    .io_dmem_writedata(cpu48_io_dmem_writedata),
    .io_dmem_memread(cpu48_io_dmem_memread),
    .io_dmem_memwrite(cpu48_io_dmem_memwrite),
    .io_dmem_maskmode(cpu48_io_dmem_maskmode),
    .io_dmem_sext(cpu48_io_dmem_sext),
    .io_dmem_readdata(cpu48_io_dmem_readdata)
  );
  DualPortedCombinMemory mem48 ( // @[top.scala 349:21]
    .clock(mem48_clock),
    .reset(mem48_reset),
    .io_imem_request_bits_address(mem48_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem48_io_imem_response_bits_data),
    .io_dmem_request_valid(mem48_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem48_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem48_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem48_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem48_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem48_io_dmem_response_bits_data)
  );
  ICombinMemPort imem48 ( // @[top.scala 350:22]
    .io_pipeline_address(imem48_io_pipeline_address),
    .io_pipeline_instruction(imem48_io_pipeline_instruction),
    .io_bus_request_bits_address(imem48_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem48_io_bus_response_bits_data)
  );
  DCombinMemPort dmem48 ( // @[top.scala 351:22]
    .clock(dmem48_clock),
    .reset(dmem48_reset),
    .io_pipeline_address(dmem48_io_pipeline_address),
    .io_pipeline_valid(dmem48_io_pipeline_valid),
    .io_pipeline_writedata(dmem48_io_pipeline_writedata),
    .io_pipeline_memread(dmem48_io_pipeline_memread),
    .io_pipeline_memwrite(dmem48_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem48_io_pipeline_maskmode),
    .io_pipeline_sext(dmem48_io_pipeline_sext),
    .io_pipeline_readdata(dmem48_io_pipeline_readdata),
    .io_bus_request_valid(dmem48_io_bus_request_valid),
    .io_bus_request_bits_address(dmem48_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem48_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem48_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem48_io_bus_response_valid),
    .io_bus_response_bits_data(dmem48_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu49 ( // @[top.scala 355:21]
    .clock(cpu49_clock),
    .reset(cpu49_reset),
    .io_imem_address(cpu49_io_imem_address),
    .io_imem_instruction(cpu49_io_imem_instruction),
    .io_dmem_address(cpu49_io_dmem_address),
    .io_dmem_valid(cpu49_io_dmem_valid),
    .io_dmem_writedata(cpu49_io_dmem_writedata),
    .io_dmem_memread(cpu49_io_dmem_memread),
    .io_dmem_memwrite(cpu49_io_dmem_memwrite),
    .io_dmem_maskmode(cpu49_io_dmem_maskmode),
    .io_dmem_sext(cpu49_io_dmem_sext),
    .io_dmem_readdata(cpu49_io_dmem_readdata)
  );
  DualPortedCombinMemory mem49 ( // @[top.scala 356:21]
    .clock(mem49_clock),
    .reset(mem49_reset),
    .io_imem_request_bits_address(mem49_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem49_io_imem_response_bits_data),
    .io_dmem_request_valid(mem49_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem49_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem49_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem49_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem49_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem49_io_dmem_response_bits_data)
  );
  ICombinMemPort imem49 ( // @[top.scala 357:22]
    .io_pipeline_address(imem49_io_pipeline_address),
    .io_pipeline_instruction(imem49_io_pipeline_instruction),
    .io_bus_request_bits_address(imem49_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem49_io_bus_response_bits_data)
  );
  DCombinMemPort dmem49 ( // @[top.scala 358:22]
    .clock(dmem49_clock),
    .reset(dmem49_reset),
    .io_pipeline_address(dmem49_io_pipeline_address),
    .io_pipeline_valid(dmem49_io_pipeline_valid),
    .io_pipeline_writedata(dmem49_io_pipeline_writedata),
    .io_pipeline_memread(dmem49_io_pipeline_memread),
    .io_pipeline_memwrite(dmem49_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem49_io_pipeline_maskmode),
    .io_pipeline_sext(dmem49_io_pipeline_sext),
    .io_pipeline_readdata(dmem49_io_pipeline_readdata),
    .io_bus_request_valid(dmem49_io_bus_request_valid),
    .io_bus_request_bits_address(dmem49_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem49_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem49_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem49_io_bus_response_valid),
    .io_bus_response_bits_data(dmem49_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu50 ( // @[top.scala 362:21]
    .clock(cpu50_clock),
    .reset(cpu50_reset),
    .io_imem_address(cpu50_io_imem_address),
    .io_imem_instruction(cpu50_io_imem_instruction),
    .io_dmem_address(cpu50_io_dmem_address),
    .io_dmem_valid(cpu50_io_dmem_valid),
    .io_dmem_writedata(cpu50_io_dmem_writedata),
    .io_dmem_memread(cpu50_io_dmem_memread),
    .io_dmem_memwrite(cpu50_io_dmem_memwrite),
    .io_dmem_maskmode(cpu50_io_dmem_maskmode),
    .io_dmem_sext(cpu50_io_dmem_sext),
    .io_dmem_readdata(cpu50_io_dmem_readdata)
  );
  DualPortedCombinMemory mem50 ( // @[top.scala 363:21]
    .clock(mem50_clock),
    .reset(mem50_reset),
    .io_imem_request_bits_address(mem50_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem50_io_imem_response_bits_data),
    .io_dmem_request_valid(mem50_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem50_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem50_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem50_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem50_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem50_io_dmem_response_bits_data)
  );
  ICombinMemPort imem50 ( // @[top.scala 364:22]
    .io_pipeline_address(imem50_io_pipeline_address),
    .io_pipeline_instruction(imem50_io_pipeline_instruction),
    .io_bus_request_bits_address(imem50_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem50_io_bus_response_bits_data)
  );
  DCombinMemPort dmem50 ( // @[top.scala 365:22]
    .clock(dmem50_clock),
    .reset(dmem50_reset),
    .io_pipeline_address(dmem50_io_pipeline_address),
    .io_pipeline_valid(dmem50_io_pipeline_valid),
    .io_pipeline_writedata(dmem50_io_pipeline_writedata),
    .io_pipeline_memread(dmem50_io_pipeline_memread),
    .io_pipeline_memwrite(dmem50_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem50_io_pipeline_maskmode),
    .io_pipeline_sext(dmem50_io_pipeline_sext),
    .io_pipeline_readdata(dmem50_io_pipeline_readdata),
    .io_bus_request_valid(dmem50_io_bus_request_valid),
    .io_bus_request_bits_address(dmem50_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem50_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem50_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem50_io_bus_response_valid),
    .io_bus_response_bits_data(dmem50_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu51 ( // @[top.scala 369:21]
    .clock(cpu51_clock),
    .reset(cpu51_reset),
    .io_imem_address(cpu51_io_imem_address),
    .io_imem_instruction(cpu51_io_imem_instruction),
    .io_dmem_address(cpu51_io_dmem_address),
    .io_dmem_valid(cpu51_io_dmem_valid),
    .io_dmem_writedata(cpu51_io_dmem_writedata),
    .io_dmem_memread(cpu51_io_dmem_memread),
    .io_dmem_memwrite(cpu51_io_dmem_memwrite),
    .io_dmem_maskmode(cpu51_io_dmem_maskmode),
    .io_dmem_sext(cpu51_io_dmem_sext),
    .io_dmem_readdata(cpu51_io_dmem_readdata)
  );
  DualPortedCombinMemory mem51 ( // @[top.scala 370:21]
    .clock(mem51_clock),
    .reset(mem51_reset),
    .io_imem_request_bits_address(mem51_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem51_io_imem_response_bits_data),
    .io_dmem_request_valid(mem51_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem51_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem51_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem51_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem51_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem51_io_dmem_response_bits_data)
  );
  ICombinMemPort imem51 ( // @[top.scala 371:22]
    .io_pipeline_address(imem51_io_pipeline_address),
    .io_pipeline_instruction(imem51_io_pipeline_instruction),
    .io_bus_request_bits_address(imem51_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem51_io_bus_response_bits_data)
  );
  DCombinMemPort dmem51 ( // @[top.scala 372:22]
    .clock(dmem51_clock),
    .reset(dmem51_reset),
    .io_pipeline_address(dmem51_io_pipeline_address),
    .io_pipeline_valid(dmem51_io_pipeline_valid),
    .io_pipeline_writedata(dmem51_io_pipeline_writedata),
    .io_pipeline_memread(dmem51_io_pipeline_memread),
    .io_pipeline_memwrite(dmem51_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem51_io_pipeline_maskmode),
    .io_pipeline_sext(dmem51_io_pipeline_sext),
    .io_pipeline_readdata(dmem51_io_pipeline_readdata),
    .io_bus_request_valid(dmem51_io_bus_request_valid),
    .io_bus_request_bits_address(dmem51_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem51_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem51_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem51_io_bus_response_valid),
    .io_bus_response_bits_data(dmem51_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu52 ( // @[top.scala 376:21]
    .clock(cpu52_clock),
    .reset(cpu52_reset),
    .io_imem_address(cpu52_io_imem_address),
    .io_imem_instruction(cpu52_io_imem_instruction),
    .io_dmem_address(cpu52_io_dmem_address),
    .io_dmem_valid(cpu52_io_dmem_valid),
    .io_dmem_writedata(cpu52_io_dmem_writedata),
    .io_dmem_memread(cpu52_io_dmem_memread),
    .io_dmem_memwrite(cpu52_io_dmem_memwrite),
    .io_dmem_maskmode(cpu52_io_dmem_maskmode),
    .io_dmem_sext(cpu52_io_dmem_sext),
    .io_dmem_readdata(cpu52_io_dmem_readdata)
  );
  DualPortedCombinMemory mem52 ( // @[top.scala 377:21]
    .clock(mem52_clock),
    .reset(mem52_reset),
    .io_imem_request_bits_address(mem52_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem52_io_imem_response_bits_data),
    .io_dmem_request_valid(mem52_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem52_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem52_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem52_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem52_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem52_io_dmem_response_bits_data)
  );
  ICombinMemPort imem52 ( // @[top.scala 378:22]
    .io_pipeline_address(imem52_io_pipeline_address),
    .io_pipeline_instruction(imem52_io_pipeline_instruction),
    .io_bus_request_bits_address(imem52_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem52_io_bus_response_bits_data)
  );
  DCombinMemPort dmem52 ( // @[top.scala 379:22]
    .clock(dmem52_clock),
    .reset(dmem52_reset),
    .io_pipeline_address(dmem52_io_pipeline_address),
    .io_pipeline_valid(dmem52_io_pipeline_valid),
    .io_pipeline_writedata(dmem52_io_pipeline_writedata),
    .io_pipeline_memread(dmem52_io_pipeline_memread),
    .io_pipeline_memwrite(dmem52_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem52_io_pipeline_maskmode),
    .io_pipeline_sext(dmem52_io_pipeline_sext),
    .io_pipeline_readdata(dmem52_io_pipeline_readdata),
    .io_bus_request_valid(dmem52_io_bus_request_valid),
    .io_bus_request_bits_address(dmem52_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem52_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem52_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem52_io_bus_response_valid),
    .io_bus_response_bits_data(dmem52_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu53 ( // @[top.scala 383:21]
    .clock(cpu53_clock),
    .reset(cpu53_reset),
    .io_imem_address(cpu53_io_imem_address),
    .io_imem_instruction(cpu53_io_imem_instruction),
    .io_dmem_address(cpu53_io_dmem_address),
    .io_dmem_valid(cpu53_io_dmem_valid),
    .io_dmem_writedata(cpu53_io_dmem_writedata),
    .io_dmem_memread(cpu53_io_dmem_memread),
    .io_dmem_memwrite(cpu53_io_dmem_memwrite),
    .io_dmem_maskmode(cpu53_io_dmem_maskmode),
    .io_dmem_sext(cpu53_io_dmem_sext),
    .io_dmem_readdata(cpu53_io_dmem_readdata)
  );
  DualPortedCombinMemory mem53 ( // @[top.scala 384:21]
    .clock(mem53_clock),
    .reset(mem53_reset),
    .io_imem_request_bits_address(mem53_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem53_io_imem_response_bits_data),
    .io_dmem_request_valid(mem53_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem53_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem53_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem53_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem53_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem53_io_dmem_response_bits_data)
  );
  ICombinMemPort imem53 ( // @[top.scala 385:22]
    .io_pipeline_address(imem53_io_pipeline_address),
    .io_pipeline_instruction(imem53_io_pipeline_instruction),
    .io_bus_request_bits_address(imem53_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem53_io_bus_response_bits_data)
  );
  DCombinMemPort dmem53 ( // @[top.scala 386:22]
    .clock(dmem53_clock),
    .reset(dmem53_reset),
    .io_pipeline_address(dmem53_io_pipeline_address),
    .io_pipeline_valid(dmem53_io_pipeline_valid),
    .io_pipeline_writedata(dmem53_io_pipeline_writedata),
    .io_pipeline_memread(dmem53_io_pipeline_memread),
    .io_pipeline_memwrite(dmem53_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem53_io_pipeline_maskmode),
    .io_pipeline_sext(dmem53_io_pipeline_sext),
    .io_pipeline_readdata(dmem53_io_pipeline_readdata),
    .io_bus_request_valid(dmem53_io_bus_request_valid),
    .io_bus_request_bits_address(dmem53_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem53_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem53_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem53_io_bus_response_valid),
    .io_bus_response_bits_data(dmem53_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu54 ( // @[top.scala 390:21]
    .clock(cpu54_clock),
    .reset(cpu54_reset),
    .io_imem_address(cpu54_io_imem_address),
    .io_imem_instruction(cpu54_io_imem_instruction),
    .io_dmem_address(cpu54_io_dmem_address),
    .io_dmem_valid(cpu54_io_dmem_valid),
    .io_dmem_writedata(cpu54_io_dmem_writedata),
    .io_dmem_memread(cpu54_io_dmem_memread),
    .io_dmem_memwrite(cpu54_io_dmem_memwrite),
    .io_dmem_maskmode(cpu54_io_dmem_maskmode),
    .io_dmem_sext(cpu54_io_dmem_sext),
    .io_dmem_readdata(cpu54_io_dmem_readdata)
  );
  DualPortedCombinMemory mem54 ( // @[top.scala 391:21]
    .clock(mem54_clock),
    .reset(mem54_reset),
    .io_imem_request_bits_address(mem54_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem54_io_imem_response_bits_data),
    .io_dmem_request_valid(mem54_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem54_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem54_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem54_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem54_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem54_io_dmem_response_bits_data)
  );
  ICombinMemPort imem54 ( // @[top.scala 392:22]
    .io_pipeline_address(imem54_io_pipeline_address),
    .io_pipeline_instruction(imem54_io_pipeline_instruction),
    .io_bus_request_bits_address(imem54_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem54_io_bus_response_bits_data)
  );
  DCombinMemPort dmem54 ( // @[top.scala 393:22]
    .clock(dmem54_clock),
    .reset(dmem54_reset),
    .io_pipeline_address(dmem54_io_pipeline_address),
    .io_pipeline_valid(dmem54_io_pipeline_valid),
    .io_pipeline_writedata(dmem54_io_pipeline_writedata),
    .io_pipeline_memread(dmem54_io_pipeline_memread),
    .io_pipeline_memwrite(dmem54_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem54_io_pipeline_maskmode),
    .io_pipeline_sext(dmem54_io_pipeline_sext),
    .io_pipeline_readdata(dmem54_io_pipeline_readdata),
    .io_bus_request_valid(dmem54_io_bus_request_valid),
    .io_bus_request_bits_address(dmem54_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem54_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem54_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem54_io_bus_response_valid),
    .io_bus_response_bits_data(dmem54_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu55 ( // @[top.scala 397:21]
    .clock(cpu55_clock),
    .reset(cpu55_reset),
    .io_imem_address(cpu55_io_imem_address),
    .io_imem_instruction(cpu55_io_imem_instruction),
    .io_dmem_address(cpu55_io_dmem_address),
    .io_dmem_valid(cpu55_io_dmem_valid),
    .io_dmem_writedata(cpu55_io_dmem_writedata),
    .io_dmem_memread(cpu55_io_dmem_memread),
    .io_dmem_memwrite(cpu55_io_dmem_memwrite),
    .io_dmem_maskmode(cpu55_io_dmem_maskmode),
    .io_dmem_sext(cpu55_io_dmem_sext),
    .io_dmem_readdata(cpu55_io_dmem_readdata)
  );
  DualPortedCombinMemory mem55 ( // @[top.scala 398:21]
    .clock(mem55_clock),
    .reset(mem55_reset),
    .io_imem_request_bits_address(mem55_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem55_io_imem_response_bits_data),
    .io_dmem_request_valid(mem55_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem55_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem55_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem55_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem55_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem55_io_dmem_response_bits_data)
  );
  ICombinMemPort imem55 ( // @[top.scala 399:22]
    .io_pipeline_address(imem55_io_pipeline_address),
    .io_pipeline_instruction(imem55_io_pipeline_instruction),
    .io_bus_request_bits_address(imem55_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem55_io_bus_response_bits_data)
  );
  DCombinMemPort dmem55 ( // @[top.scala 400:22]
    .clock(dmem55_clock),
    .reset(dmem55_reset),
    .io_pipeline_address(dmem55_io_pipeline_address),
    .io_pipeline_valid(dmem55_io_pipeline_valid),
    .io_pipeline_writedata(dmem55_io_pipeline_writedata),
    .io_pipeline_memread(dmem55_io_pipeline_memread),
    .io_pipeline_memwrite(dmem55_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem55_io_pipeline_maskmode),
    .io_pipeline_sext(dmem55_io_pipeline_sext),
    .io_pipeline_readdata(dmem55_io_pipeline_readdata),
    .io_bus_request_valid(dmem55_io_bus_request_valid),
    .io_bus_request_bits_address(dmem55_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem55_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem55_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem55_io_bus_response_valid),
    .io_bus_response_bits_data(dmem55_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu56 ( // @[top.scala 404:21]
    .clock(cpu56_clock),
    .reset(cpu56_reset),
    .io_imem_address(cpu56_io_imem_address),
    .io_imem_instruction(cpu56_io_imem_instruction),
    .io_dmem_address(cpu56_io_dmem_address),
    .io_dmem_valid(cpu56_io_dmem_valid),
    .io_dmem_writedata(cpu56_io_dmem_writedata),
    .io_dmem_memread(cpu56_io_dmem_memread),
    .io_dmem_memwrite(cpu56_io_dmem_memwrite),
    .io_dmem_maskmode(cpu56_io_dmem_maskmode),
    .io_dmem_sext(cpu56_io_dmem_sext),
    .io_dmem_readdata(cpu56_io_dmem_readdata)
  );
  DualPortedCombinMemory mem56 ( // @[top.scala 405:21]
    .clock(mem56_clock),
    .reset(mem56_reset),
    .io_imem_request_bits_address(mem56_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem56_io_imem_response_bits_data),
    .io_dmem_request_valid(mem56_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem56_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem56_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem56_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem56_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem56_io_dmem_response_bits_data)
  );
  ICombinMemPort imem56 ( // @[top.scala 406:22]
    .io_pipeline_address(imem56_io_pipeline_address),
    .io_pipeline_instruction(imem56_io_pipeline_instruction),
    .io_bus_request_bits_address(imem56_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem56_io_bus_response_bits_data)
  );
  DCombinMemPort dmem56 ( // @[top.scala 407:22]
    .clock(dmem56_clock),
    .reset(dmem56_reset),
    .io_pipeline_address(dmem56_io_pipeline_address),
    .io_pipeline_valid(dmem56_io_pipeline_valid),
    .io_pipeline_writedata(dmem56_io_pipeline_writedata),
    .io_pipeline_memread(dmem56_io_pipeline_memread),
    .io_pipeline_memwrite(dmem56_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem56_io_pipeline_maskmode),
    .io_pipeline_sext(dmem56_io_pipeline_sext),
    .io_pipeline_readdata(dmem56_io_pipeline_readdata),
    .io_bus_request_valid(dmem56_io_bus_request_valid),
    .io_bus_request_bits_address(dmem56_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem56_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem56_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem56_io_bus_response_valid),
    .io_bus_response_bits_data(dmem56_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu57 ( // @[top.scala 411:21]
    .clock(cpu57_clock),
    .reset(cpu57_reset),
    .io_imem_address(cpu57_io_imem_address),
    .io_imem_instruction(cpu57_io_imem_instruction),
    .io_dmem_address(cpu57_io_dmem_address),
    .io_dmem_valid(cpu57_io_dmem_valid),
    .io_dmem_writedata(cpu57_io_dmem_writedata),
    .io_dmem_memread(cpu57_io_dmem_memread),
    .io_dmem_memwrite(cpu57_io_dmem_memwrite),
    .io_dmem_maskmode(cpu57_io_dmem_maskmode),
    .io_dmem_sext(cpu57_io_dmem_sext),
    .io_dmem_readdata(cpu57_io_dmem_readdata)
  );
  DualPortedCombinMemory mem57 ( // @[top.scala 412:21]
    .clock(mem57_clock),
    .reset(mem57_reset),
    .io_imem_request_bits_address(mem57_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem57_io_imem_response_bits_data),
    .io_dmem_request_valid(mem57_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem57_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem57_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem57_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem57_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem57_io_dmem_response_bits_data)
  );
  ICombinMemPort imem57 ( // @[top.scala 413:22]
    .io_pipeline_address(imem57_io_pipeline_address),
    .io_pipeline_instruction(imem57_io_pipeline_instruction),
    .io_bus_request_bits_address(imem57_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem57_io_bus_response_bits_data)
  );
  DCombinMemPort dmem57 ( // @[top.scala 414:22]
    .clock(dmem57_clock),
    .reset(dmem57_reset),
    .io_pipeline_address(dmem57_io_pipeline_address),
    .io_pipeline_valid(dmem57_io_pipeline_valid),
    .io_pipeline_writedata(dmem57_io_pipeline_writedata),
    .io_pipeline_memread(dmem57_io_pipeline_memread),
    .io_pipeline_memwrite(dmem57_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem57_io_pipeline_maskmode),
    .io_pipeline_sext(dmem57_io_pipeline_sext),
    .io_pipeline_readdata(dmem57_io_pipeline_readdata),
    .io_bus_request_valid(dmem57_io_bus_request_valid),
    .io_bus_request_bits_address(dmem57_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem57_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem57_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem57_io_bus_response_valid),
    .io_bus_response_bits_data(dmem57_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu58 ( // @[top.scala 418:21]
    .clock(cpu58_clock),
    .reset(cpu58_reset),
    .io_imem_address(cpu58_io_imem_address),
    .io_imem_instruction(cpu58_io_imem_instruction),
    .io_dmem_address(cpu58_io_dmem_address),
    .io_dmem_valid(cpu58_io_dmem_valid),
    .io_dmem_writedata(cpu58_io_dmem_writedata),
    .io_dmem_memread(cpu58_io_dmem_memread),
    .io_dmem_memwrite(cpu58_io_dmem_memwrite),
    .io_dmem_maskmode(cpu58_io_dmem_maskmode),
    .io_dmem_sext(cpu58_io_dmem_sext),
    .io_dmem_readdata(cpu58_io_dmem_readdata)
  );
  DualPortedCombinMemory mem58 ( // @[top.scala 419:21]
    .clock(mem58_clock),
    .reset(mem58_reset),
    .io_imem_request_bits_address(mem58_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem58_io_imem_response_bits_data),
    .io_dmem_request_valid(mem58_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem58_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem58_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem58_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem58_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem58_io_dmem_response_bits_data)
  );
  ICombinMemPort imem58 ( // @[top.scala 420:22]
    .io_pipeline_address(imem58_io_pipeline_address),
    .io_pipeline_instruction(imem58_io_pipeline_instruction),
    .io_bus_request_bits_address(imem58_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem58_io_bus_response_bits_data)
  );
  DCombinMemPort dmem58 ( // @[top.scala 421:22]
    .clock(dmem58_clock),
    .reset(dmem58_reset),
    .io_pipeline_address(dmem58_io_pipeline_address),
    .io_pipeline_valid(dmem58_io_pipeline_valid),
    .io_pipeline_writedata(dmem58_io_pipeline_writedata),
    .io_pipeline_memread(dmem58_io_pipeline_memread),
    .io_pipeline_memwrite(dmem58_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem58_io_pipeline_maskmode),
    .io_pipeline_sext(dmem58_io_pipeline_sext),
    .io_pipeline_readdata(dmem58_io_pipeline_readdata),
    .io_bus_request_valid(dmem58_io_bus_request_valid),
    .io_bus_request_bits_address(dmem58_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem58_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem58_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem58_io_bus_response_valid),
    .io_bus_response_bits_data(dmem58_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu59 ( // @[top.scala 425:21]
    .clock(cpu59_clock),
    .reset(cpu59_reset),
    .io_imem_address(cpu59_io_imem_address),
    .io_imem_instruction(cpu59_io_imem_instruction),
    .io_dmem_address(cpu59_io_dmem_address),
    .io_dmem_valid(cpu59_io_dmem_valid),
    .io_dmem_writedata(cpu59_io_dmem_writedata),
    .io_dmem_memread(cpu59_io_dmem_memread),
    .io_dmem_memwrite(cpu59_io_dmem_memwrite),
    .io_dmem_maskmode(cpu59_io_dmem_maskmode),
    .io_dmem_sext(cpu59_io_dmem_sext),
    .io_dmem_readdata(cpu59_io_dmem_readdata)
  );
  DualPortedCombinMemory mem59 ( // @[top.scala 426:21]
    .clock(mem59_clock),
    .reset(mem59_reset),
    .io_imem_request_bits_address(mem59_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem59_io_imem_response_bits_data),
    .io_dmem_request_valid(mem59_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem59_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem59_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem59_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem59_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem59_io_dmem_response_bits_data)
  );
  ICombinMemPort imem59 ( // @[top.scala 427:22]
    .io_pipeline_address(imem59_io_pipeline_address),
    .io_pipeline_instruction(imem59_io_pipeline_instruction),
    .io_bus_request_bits_address(imem59_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem59_io_bus_response_bits_data)
  );
  DCombinMemPort dmem59 ( // @[top.scala 428:22]
    .clock(dmem59_clock),
    .reset(dmem59_reset),
    .io_pipeline_address(dmem59_io_pipeline_address),
    .io_pipeline_valid(dmem59_io_pipeline_valid),
    .io_pipeline_writedata(dmem59_io_pipeline_writedata),
    .io_pipeline_memread(dmem59_io_pipeline_memread),
    .io_pipeline_memwrite(dmem59_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem59_io_pipeline_maskmode),
    .io_pipeline_sext(dmem59_io_pipeline_sext),
    .io_pipeline_readdata(dmem59_io_pipeline_readdata),
    .io_bus_request_valid(dmem59_io_bus_request_valid),
    .io_bus_request_bits_address(dmem59_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem59_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem59_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem59_io_bus_response_valid),
    .io_bus_response_bits_data(dmem59_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu60 ( // @[top.scala 432:21]
    .clock(cpu60_clock),
    .reset(cpu60_reset),
    .io_imem_address(cpu60_io_imem_address),
    .io_imem_instruction(cpu60_io_imem_instruction),
    .io_dmem_address(cpu60_io_dmem_address),
    .io_dmem_valid(cpu60_io_dmem_valid),
    .io_dmem_writedata(cpu60_io_dmem_writedata),
    .io_dmem_memread(cpu60_io_dmem_memread),
    .io_dmem_memwrite(cpu60_io_dmem_memwrite),
    .io_dmem_maskmode(cpu60_io_dmem_maskmode),
    .io_dmem_sext(cpu60_io_dmem_sext),
    .io_dmem_readdata(cpu60_io_dmem_readdata)
  );
  DualPortedCombinMemory mem60 ( // @[top.scala 433:21]
    .clock(mem60_clock),
    .reset(mem60_reset),
    .io_imem_request_bits_address(mem60_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem60_io_imem_response_bits_data),
    .io_dmem_request_valid(mem60_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem60_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem60_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem60_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem60_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem60_io_dmem_response_bits_data)
  );
  ICombinMemPort imem60 ( // @[top.scala 434:22]
    .io_pipeline_address(imem60_io_pipeline_address),
    .io_pipeline_instruction(imem60_io_pipeline_instruction),
    .io_bus_request_bits_address(imem60_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem60_io_bus_response_bits_data)
  );
  DCombinMemPort dmem60 ( // @[top.scala 435:22]
    .clock(dmem60_clock),
    .reset(dmem60_reset),
    .io_pipeline_address(dmem60_io_pipeline_address),
    .io_pipeline_valid(dmem60_io_pipeline_valid),
    .io_pipeline_writedata(dmem60_io_pipeline_writedata),
    .io_pipeline_memread(dmem60_io_pipeline_memread),
    .io_pipeline_memwrite(dmem60_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem60_io_pipeline_maskmode),
    .io_pipeline_sext(dmem60_io_pipeline_sext),
    .io_pipeline_readdata(dmem60_io_pipeline_readdata),
    .io_bus_request_valid(dmem60_io_bus_request_valid),
    .io_bus_request_bits_address(dmem60_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem60_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem60_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem60_io_bus_response_valid),
    .io_bus_response_bits_data(dmem60_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu61 ( // @[top.scala 439:21]
    .clock(cpu61_clock),
    .reset(cpu61_reset),
    .io_imem_address(cpu61_io_imem_address),
    .io_imem_instruction(cpu61_io_imem_instruction),
    .io_dmem_address(cpu61_io_dmem_address),
    .io_dmem_valid(cpu61_io_dmem_valid),
    .io_dmem_writedata(cpu61_io_dmem_writedata),
    .io_dmem_memread(cpu61_io_dmem_memread),
    .io_dmem_memwrite(cpu61_io_dmem_memwrite),
    .io_dmem_maskmode(cpu61_io_dmem_maskmode),
    .io_dmem_sext(cpu61_io_dmem_sext),
    .io_dmem_readdata(cpu61_io_dmem_readdata)
  );
  DualPortedCombinMemory mem61 ( // @[top.scala 440:21]
    .clock(mem61_clock),
    .reset(mem61_reset),
    .io_imem_request_bits_address(mem61_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem61_io_imem_response_bits_data),
    .io_dmem_request_valid(mem61_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem61_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem61_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem61_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem61_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem61_io_dmem_response_bits_data)
  );
  ICombinMemPort imem61 ( // @[top.scala 441:22]
    .io_pipeline_address(imem61_io_pipeline_address),
    .io_pipeline_instruction(imem61_io_pipeline_instruction),
    .io_bus_request_bits_address(imem61_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem61_io_bus_response_bits_data)
  );
  DCombinMemPort dmem61 ( // @[top.scala 442:22]
    .clock(dmem61_clock),
    .reset(dmem61_reset),
    .io_pipeline_address(dmem61_io_pipeline_address),
    .io_pipeline_valid(dmem61_io_pipeline_valid),
    .io_pipeline_writedata(dmem61_io_pipeline_writedata),
    .io_pipeline_memread(dmem61_io_pipeline_memread),
    .io_pipeline_memwrite(dmem61_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem61_io_pipeline_maskmode),
    .io_pipeline_sext(dmem61_io_pipeline_sext),
    .io_pipeline_readdata(dmem61_io_pipeline_readdata),
    .io_bus_request_valid(dmem61_io_bus_request_valid),
    .io_bus_request_bits_address(dmem61_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem61_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem61_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem61_io_bus_response_valid),
    .io_bus_response_bits_data(dmem61_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu62 ( // @[top.scala 446:21]
    .clock(cpu62_clock),
    .reset(cpu62_reset),
    .io_imem_address(cpu62_io_imem_address),
    .io_imem_instruction(cpu62_io_imem_instruction),
    .io_dmem_address(cpu62_io_dmem_address),
    .io_dmem_valid(cpu62_io_dmem_valid),
    .io_dmem_writedata(cpu62_io_dmem_writedata),
    .io_dmem_memread(cpu62_io_dmem_memread),
    .io_dmem_memwrite(cpu62_io_dmem_memwrite),
    .io_dmem_maskmode(cpu62_io_dmem_maskmode),
    .io_dmem_sext(cpu62_io_dmem_sext),
    .io_dmem_readdata(cpu62_io_dmem_readdata)
  );
  DualPortedCombinMemory mem62 ( // @[top.scala 447:21]
    .clock(mem62_clock),
    .reset(mem62_reset),
    .io_imem_request_bits_address(mem62_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem62_io_imem_response_bits_data),
    .io_dmem_request_valid(mem62_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem62_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem62_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem62_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem62_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem62_io_dmem_response_bits_data)
  );
  ICombinMemPort imem62 ( // @[top.scala 448:22]
    .io_pipeline_address(imem62_io_pipeline_address),
    .io_pipeline_instruction(imem62_io_pipeline_instruction),
    .io_bus_request_bits_address(imem62_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem62_io_bus_response_bits_data)
  );
  DCombinMemPort dmem62 ( // @[top.scala 449:22]
    .clock(dmem62_clock),
    .reset(dmem62_reset),
    .io_pipeline_address(dmem62_io_pipeline_address),
    .io_pipeline_valid(dmem62_io_pipeline_valid),
    .io_pipeline_writedata(dmem62_io_pipeline_writedata),
    .io_pipeline_memread(dmem62_io_pipeline_memread),
    .io_pipeline_memwrite(dmem62_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem62_io_pipeline_maskmode),
    .io_pipeline_sext(dmem62_io_pipeline_sext),
    .io_pipeline_readdata(dmem62_io_pipeline_readdata),
    .io_bus_request_valid(dmem62_io_bus_request_valid),
    .io_bus_request_bits_address(dmem62_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem62_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem62_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem62_io_bus_response_valid),
    .io_bus_response_bits_data(dmem62_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu63 ( // @[top.scala 453:21]
    .clock(cpu63_clock),
    .reset(cpu63_reset),
    .io_imem_address(cpu63_io_imem_address),
    .io_imem_instruction(cpu63_io_imem_instruction),
    .io_dmem_address(cpu63_io_dmem_address),
    .io_dmem_valid(cpu63_io_dmem_valid),
    .io_dmem_writedata(cpu63_io_dmem_writedata),
    .io_dmem_memread(cpu63_io_dmem_memread),
    .io_dmem_memwrite(cpu63_io_dmem_memwrite),
    .io_dmem_maskmode(cpu63_io_dmem_maskmode),
    .io_dmem_sext(cpu63_io_dmem_sext),
    .io_dmem_readdata(cpu63_io_dmem_readdata)
  );
  DualPortedCombinMemory mem63 ( // @[top.scala 454:21]
    .clock(mem63_clock),
    .reset(mem63_reset),
    .io_imem_request_bits_address(mem63_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem63_io_imem_response_bits_data),
    .io_dmem_request_valid(mem63_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem63_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem63_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem63_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem63_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem63_io_dmem_response_bits_data)
  );
  ICombinMemPort imem63 ( // @[top.scala 455:22]
    .io_pipeline_address(imem63_io_pipeline_address),
    .io_pipeline_instruction(imem63_io_pipeline_instruction),
    .io_bus_request_bits_address(imem63_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem63_io_bus_response_bits_data)
  );
  DCombinMemPort dmem63 ( // @[top.scala 456:22]
    .clock(dmem63_clock),
    .reset(dmem63_reset),
    .io_pipeline_address(dmem63_io_pipeline_address),
    .io_pipeline_valid(dmem63_io_pipeline_valid),
    .io_pipeline_writedata(dmem63_io_pipeline_writedata),
    .io_pipeline_memread(dmem63_io_pipeline_memread),
    .io_pipeline_memwrite(dmem63_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem63_io_pipeline_maskmode),
    .io_pipeline_sext(dmem63_io_pipeline_sext),
    .io_pipeline_readdata(dmem63_io_pipeline_readdata),
    .io_bus_request_valid(dmem63_io_bus_request_valid),
    .io_bus_request_bits_address(dmem63_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem63_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem63_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem63_io_bus_response_valid),
    .io_bus_response_bits_data(dmem63_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu64 ( // @[top.scala 460:21]
    .clock(cpu64_clock),
    .reset(cpu64_reset),
    .io_imem_address(cpu64_io_imem_address),
    .io_imem_instruction(cpu64_io_imem_instruction),
    .io_dmem_address(cpu64_io_dmem_address),
    .io_dmem_valid(cpu64_io_dmem_valid),
    .io_dmem_writedata(cpu64_io_dmem_writedata),
    .io_dmem_memread(cpu64_io_dmem_memread),
    .io_dmem_memwrite(cpu64_io_dmem_memwrite),
    .io_dmem_maskmode(cpu64_io_dmem_maskmode),
    .io_dmem_sext(cpu64_io_dmem_sext),
    .io_dmem_readdata(cpu64_io_dmem_readdata)
  );
  DualPortedCombinMemory mem64 ( // @[top.scala 461:21]
    .clock(mem64_clock),
    .reset(mem64_reset),
    .io_imem_request_bits_address(mem64_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem64_io_imem_response_bits_data),
    .io_dmem_request_valid(mem64_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem64_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem64_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem64_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem64_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem64_io_dmem_response_bits_data)
  );
  ICombinMemPort imem64 ( // @[top.scala 462:22]
    .io_pipeline_address(imem64_io_pipeline_address),
    .io_pipeline_instruction(imem64_io_pipeline_instruction),
    .io_bus_request_bits_address(imem64_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem64_io_bus_response_bits_data)
  );
  DCombinMemPort dmem64 ( // @[top.scala 463:22]
    .clock(dmem64_clock),
    .reset(dmem64_reset),
    .io_pipeline_address(dmem64_io_pipeline_address),
    .io_pipeline_valid(dmem64_io_pipeline_valid),
    .io_pipeline_writedata(dmem64_io_pipeline_writedata),
    .io_pipeline_memread(dmem64_io_pipeline_memread),
    .io_pipeline_memwrite(dmem64_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem64_io_pipeline_maskmode),
    .io_pipeline_sext(dmem64_io_pipeline_sext),
    .io_pipeline_readdata(dmem64_io_pipeline_readdata),
    .io_bus_request_valid(dmem64_io_bus_request_valid),
    .io_bus_request_bits_address(dmem64_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem64_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem64_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem64_io_bus_response_valid),
    .io_bus_response_bits_data(dmem64_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu65 ( // @[top.scala 467:21]
    .clock(cpu65_clock),
    .reset(cpu65_reset),
    .io_imem_address(cpu65_io_imem_address),
    .io_imem_instruction(cpu65_io_imem_instruction),
    .io_dmem_address(cpu65_io_dmem_address),
    .io_dmem_valid(cpu65_io_dmem_valid),
    .io_dmem_writedata(cpu65_io_dmem_writedata),
    .io_dmem_memread(cpu65_io_dmem_memread),
    .io_dmem_memwrite(cpu65_io_dmem_memwrite),
    .io_dmem_maskmode(cpu65_io_dmem_maskmode),
    .io_dmem_sext(cpu65_io_dmem_sext),
    .io_dmem_readdata(cpu65_io_dmem_readdata)
  );
  DualPortedCombinMemory mem65 ( // @[top.scala 468:21]
    .clock(mem65_clock),
    .reset(mem65_reset),
    .io_imem_request_bits_address(mem65_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem65_io_imem_response_bits_data),
    .io_dmem_request_valid(mem65_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem65_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem65_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem65_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem65_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem65_io_dmem_response_bits_data)
  );
  ICombinMemPort imem65 ( // @[top.scala 469:22]
    .io_pipeline_address(imem65_io_pipeline_address),
    .io_pipeline_instruction(imem65_io_pipeline_instruction),
    .io_bus_request_bits_address(imem65_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem65_io_bus_response_bits_data)
  );
  DCombinMemPort dmem65 ( // @[top.scala 470:22]
    .clock(dmem65_clock),
    .reset(dmem65_reset),
    .io_pipeline_address(dmem65_io_pipeline_address),
    .io_pipeline_valid(dmem65_io_pipeline_valid),
    .io_pipeline_writedata(dmem65_io_pipeline_writedata),
    .io_pipeline_memread(dmem65_io_pipeline_memread),
    .io_pipeline_memwrite(dmem65_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem65_io_pipeline_maskmode),
    .io_pipeline_sext(dmem65_io_pipeline_sext),
    .io_pipeline_readdata(dmem65_io_pipeline_readdata),
    .io_bus_request_valid(dmem65_io_bus_request_valid),
    .io_bus_request_bits_address(dmem65_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem65_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem65_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem65_io_bus_response_valid),
    .io_bus_response_bits_data(dmem65_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu66 ( // @[top.scala 474:21]
    .clock(cpu66_clock),
    .reset(cpu66_reset),
    .io_imem_address(cpu66_io_imem_address),
    .io_imem_instruction(cpu66_io_imem_instruction),
    .io_dmem_address(cpu66_io_dmem_address),
    .io_dmem_valid(cpu66_io_dmem_valid),
    .io_dmem_writedata(cpu66_io_dmem_writedata),
    .io_dmem_memread(cpu66_io_dmem_memread),
    .io_dmem_memwrite(cpu66_io_dmem_memwrite),
    .io_dmem_maskmode(cpu66_io_dmem_maskmode),
    .io_dmem_sext(cpu66_io_dmem_sext),
    .io_dmem_readdata(cpu66_io_dmem_readdata)
  );
  DualPortedCombinMemory mem66 ( // @[top.scala 475:21]
    .clock(mem66_clock),
    .reset(mem66_reset),
    .io_imem_request_bits_address(mem66_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem66_io_imem_response_bits_data),
    .io_dmem_request_valid(mem66_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem66_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem66_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem66_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem66_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem66_io_dmem_response_bits_data)
  );
  ICombinMemPort imem66 ( // @[top.scala 476:22]
    .io_pipeline_address(imem66_io_pipeline_address),
    .io_pipeline_instruction(imem66_io_pipeline_instruction),
    .io_bus_request_bits_address(imem66_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem66_io_bus_response_bits_data)
  );
  DCombinMemPort dmem66 ( // @[top.scala 477:22]
    .clock(dmem66_clock),
    .reset(dmem66_reset),
    .io_pipeline_address(dmem66_io_pipeline_address),
    .io_pipeline_valid(dmem66_io_pipeline_valid),
    .io_pipeline_writedata(dmem66_io_pipeline_writedata),
    .io_pipeline_memread(dmem66_io_pipeline_memread),
    .io_pipeline_memwrite(dmem66_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem66_io_pipeline_maskmode),
    .io_pipeline_sext(dmem66_io_pipeline_sext),
    .io_pipeline_readdata(dmem66_io_pipeline_readdata),
    .io_bus_request_valid(dmem66_io_bus_request_valid),
    .io_bus_request_bits_address(dmem66_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem66_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem66_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem66_io_bus_response_valid),
    .io_bus_response_bits_data(dmem66_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu67 ( // @[top.scala 481:21]
    .clock(cpu67_clock),
    .reset(cpu67_reset),
    .io_imem_address(cpu67_io_imem_address),
    .io_imem_instruction(cpu67_io_imem_instruction),
    .io_dmem_address(cpu67_io_dmem_address),
    .io_dmem_valid(cpu67_io_dmem_valid),
    .io_dmem_writedata(cpu67_io_dmem_writedata),
    .io_dmem_memread(cpu67_io_dmem_memread),
    .io_dmem_memwrite(cpu67_io_dmem_memwrite),
    .io_dmem_maskmode(cpu67_io_dmem_maskmode),
    .io_dmem_sext(cpu67_io_dmem_sext),
    .io_dmem_readdata(cpu67_io_dmem_readdata)
  );
  DualPortedCombinMemory mem67 ( // @[top.scala 482:21]
    .clock(mem67_clock),
    .reset(mem67_reset),
    .io_imem_request_bits_address(mem67_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem67_io_imem_response_bits_data),
    .io_dmem_request_valid(mem67_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem67_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem67_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem67_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem67_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem67_io_dmem_response_bits_data)
  );
  ICombinMemPort imem67 ( // @[top.scala 483:22]
    .io_pipeline_address(imem67_io_pipeline_address),
    .io_pipeline_instruction(imem67_io_pipeline_instruction),
    .io_bus_request_bits_address(imem67_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem67_io_bus_response_bits_data)
  );
  DCombinMemPort dmem67 ( // @[top.scala 484:22]
    .clock(dmem67_clock),
    .reset(dmem67_reset),
    .io_pipeline_address(dmem67_io_pipeline_address),
    .io_pipeline_valid(dmem67_io_pipeline_valid),
    .io_pipeline_writedata(dmem67_io_pipeline_writedata),
    .io_pipeline_memread(dmem67_io_pipeline_memread),
    .io_pipeline_memwrite(dmem67_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem67_io_pipeline_maskmode),
    .io_pipeline_sext(dmem67_io_pipeline_sext),
    .io_pipeline_readdata(dmem67_io_pipeline_readdata),
    .io_bus_request_valid(dmem67_io_bus_request_valid),
    .io_bus_request_bits_address(dmem67_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem67_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem67_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem67_io_bus_response_valid),
    .io_bus_response_bits_data(dmem67_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu68 ( // @[top.scala 488:21]
    .clock(cpu68_clock),
    .reset(cpu68_reset),
    .io_imem_address(cpu68_io_imem_address),
    .io_imem_instruction(cpu68_io_imem_instruction),
    .io_dmem_address(cpu68_io_dmem_address),
    .io_dmem_valid(cpu68_io_dmem_valid),
    .io_dmem_writedata(cpu68_io_dmem_writedata),
    .io_dmem_memread(cpu68_io_dmem_memread),
    .io_dmem_memwrite(cpu68_io_dmem_memwrite),
    .io_dmem_maskmode(cpu68_io_dmem_maskmode),
    .io_dmem_sext(cpu68_io_dmem_sext),
    .io_dmem_readdata(cpu68_io_dmem_readdata)
  );
  DualPortedCombinMemory mem68 ( // @[top.scala 489:21]
    .clock(mem68_clock),
    .reset(mem68_reset),
    .io_imem_request_bits_address(mem68_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem68_io_imem_response_bits_data),
    .io_dmem_request_valid(mem68_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem68_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem68_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem68_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem68_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem68_io_dmem_response_bits_data)
  );
  ICombinMemPort imem68 ( // @[top.scala 490:22]
    .io_pipeline_address(imem68_io_pipeline_address),
    .io_pipeline_instruction(imem68_io_pipeline_instruction),
    .io_bus_request_bits_address(imem68_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem68_io_bus_response_bits_data)
  );
  DCombinMemPort dmem68 ( // @[top.scala 491:22]
    .clock(dmem68_clock),
    .reset(dmem68_reset),
    .io_pipeline_address(dmem68_io_pipeline_address),
    .io_pipeline_valid(dmem68_io_pipeline_valid),
    .io_pipeline_writedata(dmem68_io_pipeline_writedata),
    .io_pipeline_memread(dmem68_io_pipeline_memread),
    .io_pipeline_memwrite(dmem68_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem68_io_pipeline_maskmode),
    .io_pipeline_sext(dmem68_io_pipeline_sext),
    .io_pipeline_readdata(dmem68_io_pipeline_readdata),
    .io_bus_request_valid(dmem68_io_bus_request_valid),
    .io_bus_request_bits_address(dmem68_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem68_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem68_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem68_io_bus_response_valid),
    .io_bus_response_bits_data(dmem68_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu69 ( // @[top.scala 495:21]
    .clock(cpu69_clock),
    .reset(cpu69_reset),
    .io_imem_address(cpu69_io_imem_address),
    .io_imem_instruction(cpu69_io_imem_instruction),
    .io_dmem_address(cpu69_io_dmem_address),
    .io_dmem_valid(cpu69_io_dmem_valid),
    .io_dmem_writedata(cpu69_io_dmem_writedata),
    .io_dmem_memread(cpu69_io_dmem_memread),
    .io_dmem_memwrite(cpu69_io_dmem_memwrite),
    .io_dmem_maskmode(cpu69_io_dmem_maskmode),
    .io_dmem_sext(cpu69_io_dmem_sext),
    .io_dmem_readdata(cpu69_io_dmem_readdata)
  );
  DualPortedCombinMemory mem69 ( // @[top.scala 496:21]
    .clock(mem69_clock),
    .reset(mem69_reset),
    .io_imem_request_bits_address(mem69_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem69_io_imem_response_bits_data),
    .io_dmem_request_valid(mem69_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem69_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem69_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem69_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem69_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem69_io_dmem_response_bits_data)
  );
  ICombinMemPort imem69 ( // @[top.scala 497:22]
    .io_pipeline_address(imem69_io_pipeline_address),
    .io_pipeline_instruction(imem69_io_pipeline_instruction),
    .io_bus_request_bits_address(imem69_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem69_io_bus_response_bits_data)
  );
  DCombinMemPort dmem69 ( // @[top.scala 498:22]
    .clock(dmem69_clock),
    .reset(dmem69_reset),
    .io_pipeline_address(dmem69_io_pipeline_address),
    .io_pipeline_valid(dmem69_io_pipeline_valid),
    .io_pipeline_writedata(dmem69_io_pipeline_writedata),
    .io_pipeline_memread(dmem69_io_pipeline_memread),
    .io_pipeline_memwrite(dmem69_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem69_io_pipeline_maskmode),
    .io_pipeline_sext(dmem69_io_pipeline_sext),
    .io_pipeline_readdata(dmem69_io_pipeline_readdata),
    .io_bus_request_valid(dmem69_io_bus_request_valid),
    .io_bus_request_bits_address(dmem69_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem69_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem69_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem69_io_bus_response_valid),
    .io_bus_response_bits_data(dmem69_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu70 ( // @[top.scala 502:21]
    .clock(cpu70_clock),
    .reset(cpu70_reset),
    .io_imem_address(cpu70_io_imem_address),
    .io_imem_instruction(cpu70_io_imem_instruction),
    .io_dmem_address(cpu70_io_dmem_address),
    .io_dmem_valid(cpu70_io_dmem_valid),
    .io_dmem_writedata(cpu70_io_dmem_writedata),
    .io_dmem_memread(cpu70_io_dmem_memread),
    .io_dmem_memwrite(cpu70_io_dmem_memwrite),
    .io_dmem_maskmode(cpu70_io_dmem_maskmode),
    .io_dmem_sext(cpu70_io_dmem_sext),
    .io_dmem_readdata(cpu70_io_dmem_readdata)
  );
  DualPortedCombinMemory mem70 ( // @[top.scala 503:21]
    .clock(mem70_clock),
    .reset(mem70_reset),
    .io_imem_request_bits_address(mem70_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem70_io_imem_response_bits_data),
    .io_dmem_request_valid(mem70_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem70_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem70_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem70_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem70_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem70_io_dmem_response_bits_data)
  );
  ICombinMemPort imem70 ( // @[top.scala 504:22]
    .io_pipeline_address(imem70_io_pipeline_address),
    .io_pipeline_instruction(imem70_io_pipeline_instruction),
    .io_bus_request_bits_address(imem70_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem70_io_bus_response_bits_data)
  );
  DCombinMemPort dmem70 ( // @[top.scala 505:22]
    .clock(dmem70_clock),
    .reset(dmem70_reset),
    .io_pipeline_address(dmem70_io_pipeline_address),
    .io_pipeline_valid(dmem70_io_pipeline_valid),
    .io_pipeline_writedata(dmem70_io_pipeline_writedata),
    .io_pipeline_memread(dmem70_io_pipeline_memread),
    .io_pipeline_memwrite(dmem70_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem70_io_pipeline_maskmode),
    .io_pipeline_sext(dmem70_io_pipeline_sext),
    .io_pipeline_readdata(dmem70_io_pipeline_readdata),
    .io_bus_request_valid(dmem70_io_bus_request_valid),
    .io_bus_request_bits_address(dmem70_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem70_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem70_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem70_io_bus_response_valid),
    .io_bus_response_bits_data(dmem70_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu71 ( // @[top.scala 509:21]
    .clock(cpu71_clock),
    .reset(cpu71_reset),
    .io_imem_address(cpu71_io_imem_address),
    .io_imem_instruction(cpu71_io_imem_instruction),
    .io_dmem_address(cpu71_io_dmem_address),
    .io_dmem_valid(cpu71_io_dmem_valid),
    .io_dmem_writedata(cpu71_io_dmem_writedata),
    .io_dmem_memread(cpu71_io_dmem_memread),
    .io_dmem_memwrite(cpu71_io_dmem_memwrite),
    .io_dmem_maskmode(cpu71_io_dmem_maskmode),
    .io_dmem_sext(cpu71_io_dmem_sext),
    .io_dmem_readdata(cpu71_io_dmem_readdata)
  );
  DualPortedCombinMemory mem71 ( // @[top.scala 510:21]
    .clock(mem71_clock),
    .reset(mem71_reset),
    .io_imem_request_bits_address(mem71_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem71_io_imem_response_bits_data),
    .io_dmem_request_valid(mem71_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem71_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem71_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem71_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem71_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem71_io_dmem_response_bits_data)
  );
  ICombinMemPort imem71 ( // @[top.scala 511:22]
    .io_pipeline_address(imem71_io_pipeline_address),
    .io_pipeline_instruction(imem71_io_pipeline_instruction),
    .io_bus_request_bits_address(imem71_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem71_io_bus_response_bits_data)
  );
  DCombinMemPort dmem71 ( // @[top.scala 512:22]
    .clock(dmem71_clock),
    .reset(dmem71_reset),
    .io_pipeline_address(dmem71_io_pipeline_address),
    .io_pipeline_valid(dmem71_io_pipeline_valid),
    .io_pipeline_writedata(dmem71_io_pipeline_writedata),
    .io_pipeline_memread(dmem71_io_pipeline_memread),
    .io_pipeline_memwrite(dmem71_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem71_io_pipeline_maskmode),
    .io_pipeline_sext(dmem71_io_pipeline_sext),
    .io_pipeline_readdata(dmem71_io_pipeline_readdata),
    .io_bus_request_valid(dmem71_io_bus_request_valid),
    .io_bus_request_bits_address(dmem71_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem71_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem71_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem71_io_bus_response_valid),
    .io_bus_response_bits_data(dmem71_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu72 ( // @[top.scala 516:21]
    .clock(cpu72_clock),
    .reset(cpu72_reset),
    .io_imem_address(cpu72_io_imem_address),
    .io_imem_instruction(cpu72_io_imem_instruction),
    .io_dmem_address(cpu72_io_dmem_address),
    .io_dmem_valid(cpu72_io_dmem_valid),
    .io_dmem_writedata(cpu72_io_dmem_writedata),
    .io_dmem_memread(cpu72_io_dmem_memread),
    .io_dmem_memwrite(cpu72_io_dmem_memwrite),
    .io_dmem_maskmode(cpu72_io_dmem_maskmode),
    .io_dmem_sext(cpu72_io_dmem_sext),
    .io_dmem_readdata(cpu72_io_dmem_readdata)
  );
  DualPortedCombinMemory mem72 ( // @[top.scala 517:21]
    .clock(mem72_clock),
    .reset(mem72_reset),
    .io_imem_request_bits_address(mem72_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem72_io_imem_response_bits_data),
    .io_dmem_request_valid(mem72_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem72_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem72_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem72_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem72_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem72_io_dmem_response_bits_data)
  );
  ICombinMemPort imem72 ( // @[top.scala 518:22]
    .io_pipeline_address(imem72_io_pipeline_address),
    .io_pipeline_instruction(imem72_io_pipeline_instruction),
    .io_bus_request_bits_address(imem72_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem72_io_bus_response_bits_data)
  );
  DCombinMemPort dmem72 ( // @[top.scala 519:22]
    .clock(dmem72_clock),
    .reset(dmem72_reset),
    .io_pipeline_address(dmem72_io_pipeline_address),
    .io_pipeline_valid(dmem72_io_pipeline_valid),
    .io_pipeline_writedata(dmem72_io_pipeline_writedata),
    .io_pipeline_memread(dmem72_io_pipeline_memread),
    .io_pipeline_memwrite(dmem72_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem72_io_pipeline_maskmode),
    .io_pipeline_sext(dmem72_io_pipeline_sext),
    .io_pipeline_readdata(dmem72_io_pipeline_readdata),
    .io_bus_request_valid(dmem72_io_bus_request_valid),
    .io_bus_request_bits_address(dmem72_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem72_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem72_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem72_io_bus_response_valid),
    .io_bus_response_bits_data(dmem72_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu73 ( // @[top.scala 523:21]
    .clock(cpu73_clock),
    .reset(cpu73_reset),
    .io_imem_address(cpu73_io_imem_address),
    .io_imem_instruction(cpu73_io_imem_instruction),
    .io_dmem_address(cpu73_io_dmem_address),
    .io_dmem_valid(cpu73_io_dmem_valid),
    .io_dmem_writedata(cpu73_io_dmem_writedata),
    .io_dmem_memread(cpu73_io_dmem_memread),
    .io_dmem_memwrite(cpu73_io_dmem_memwrite),
    .io_dmem_maskmode(cpu73_io_dmem_maskmode),
    .io_dmem_sext(cpu73_io_dmem_sext),
    .io_dmem_readdata(cpu73_io_dmem_readdata)
  );
  DualPortedCombinMemory mem73 ( // @[top.scala 524:21]
    .clock(mem73_clock),
    .reset(mem73_reset),
    .io_imem_request_bits_address(mem73_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem73_io_imem_response_bits_data),
    .io_dmem_request_valid(mem73_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem73_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem73_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem73_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem73_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem73_io_dmem_response_bits_data)
  );
  ICombinMemPort imem73 ( // @[top.scala 525:22]
    .io_pipeline_address(imem73_io_pipeline_address),
    .io_pipeline_instruction(imem73_io_pipeline_instruction),
    .io_bus_request_bits_address(imem73_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem73_io_bus_response_bits_data)
  );
  DCombinMemPort dmem73 ( // @[top.scala 526:22]
    .clock(dmem73_clock),
    .reset(dmem73_reset),
    .io_pipeline_address(dmem73_io_pipeline_address),
    .io_pipeline_valid(dmem73_io_pipeline_valid),
    .io_pipeline_writedata(dmem73_io_pipeline_writedata),
    .io_pipeline_memread(dmem73_io_pipeline_memread),
    .io_pipeline_memwrite(dmem73_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem73_io_pipeline_maskmode),
    .io_pipeline_sext(dmem73_io_pipeline_sext),
    .io_pipeline_readdata(dmem73_io_pipeline_readdata),
    .io_bus_request_valid(dmem73_io_bus_request_valid),
    .io_bus_request_bits_address(dmem73_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem73_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem73_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem73_io_bus_response_valid),
    .io_bus_response_bits_data(dmem73_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu74 ( // @[top.scala 530:21]
    .clock(cpu74_clock),
    .reset(cpu74_reset),
    .io_imem_address(cpu74_io_imem_address),
    .io_imem_instruction(cpu74_io_imem_instruction),
    .io_dmem_address(cpu74_io_dmem_address),
    .io_dmem_valid(cpu74_io_dmem_valid),
    .io_dmem_writedata(cpu74_io_dmem_writedata),
    .io_dmem_memread(cpu74_io_dmem_memread),
    .io_dmem_memwrite(cpu74_io_dmem_memwrite),
    .io_dmem_maskmode(cpu74_io_dmem_maskmode),
    .io_dmem_sext(cpu74_io_dmem_sext),
    .io_dmem_readdata(cpu74_io_dmem_readdata)
  );
  DualPortedCombinMemory mem74 ( // @[top.scala 531:21]
    .clock(mem74_clock),
    .reset(mem74_reset),
    .io_imem_request_bits_address(mem74_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem74_io_imem_response_bits_data),
    .io_dmem_request_valid(mem74_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem74_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem74_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem74_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem74_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem74_io_dmem_response_bits_data)
  );
  ICombinMemPort imem74 ( // @[top.scala 532:22]
    .io_pipeline_address(imem74_io_pipeline_address),
    .io_pipeline_instruction(imem74_io_pipeline_instruction),
    .io_bus_request_bits_address(imem74_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem74_io_bus_response_bits_data)
  );
  DCombinMemPort dmem74 ( // @[top.scala 533:22]
    .clock(dmem74_clock),
    .reset(dmem74_reset),
    .io_pipeline_address(dmem74_io_pipeline_address),
    .io_pipeline_valid(dmem74_io_pipeline_valid),
    .io_pipeline_writedata(dmem74_io_pipeline_writedata),
    .io_pipeline_memread(dmem74_io_pipeline_memread),
    .io_pipeline_memwrite(dmem74_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem74_io_pipeline_maskmode),
    .io_pipeline_sext(dmem74_io_pipeline_sext),
    .io_pipeline_readdata(dmem74_io_pipeline_readdata),
    .io_bus_request_valid(dmem74_io_bus_request_valid),
    .io_bus_request_bits_address(dmem74_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem74_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem74_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem74_io_bus_response_valid),
    .io_bus_response_bits_data(dmem74_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu75 ( // @[top.scala 537:21]
    .clock(cpu75_clock),
    .reset(cpu75_reset),
    .io_imem_address(cpu75_io_imem_address),
    .io_imem_instruction(cpu75_io_imem_instruction),
    .io_dmem_address(cpu75_io_dmem_address),
    .io_dmem_valid(cpu75_io_dmem_valid),
    .io_dmem_writedata(cpu75_io_dmem_writedata),
    .io_dmem_memread(cpu75_io_dmem_memread),
    .io_dmem_memwrite(cpu75_io_dmem_memwrite),
    .io_dmem_maskmode(cpu75_io_dmem_maskmode),
    .io_dmem_sext(cpu75_io_dmem_sext),
    .io_dmem_readdata(cpu75_io_dmem_readdata)
  );
  DualPortedCombinMemory mem75 ( // @[top.scala 538:21]
    .clock(mem75_clock),
    .reset(mem75_reset),
    .io_imem_request_bits_address(mem75_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem75_io_imem_response_bits_data),
    .io_dmem_request_valid(mem75_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem75_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem75_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem75_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem75_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem75_io_dmem_response_bits_data)
  );
  ICombinMemPort imem75 ( // @[top.scala 539:22]
    .io_pipeline_address(imem75_io_pipeline_address),
    .io_pipeline_instruction(imem75_io_pipeline_instruction),
    .io_bus_request_bits_address(imem75_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem75_io_bus_response_bits_data)
  );
  DCombinMemPort dmem75 ( // @[top.scala 540:22]
    .clock(dmem75_clock),
    .reset(dmem75_reset),
    .io_pipeline_address(dmem75_io_pipeline_address),
    .io_pipeline_valid(dmem75_io_pipeline_valid),
    .io_pipeline_writedata(dmem75_io_pipeline_writedata),
    .io_pipeline_memread(dmem75_io_pipeline_memread),
    .io_pipeline_memwrite(dmem75_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem75_io_pipeline_maskmode),
    .io_pipeline_sext(dmem75_io_pipeline_sext),
    .io_pipeline_readdata(dmem75_io_pipeline_readdata),
    .io_bus_request_valid(dmem75_io_bus_request_valid),
    .io_bus_request_bits_address(dmem75_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem75_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem75_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem75_io_bus_response_valid),
    .io_bus_response_bits_data(dmem75_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu76 ( // @[top.scala 544:21]
    .clock(cpu76_clock),
    .reset(cpu76_reset),
    .io_imem_address(cpu76_io_imem_address),
    .io_imem_instruction(cpu76_io_imem_instruction),
    .io_dmem_address(cpu76_io_dmem_address),
    .io_dmem_valid(cpu76_io_dmem_valid),
    .io_dmem_writedata(cpu76_io_dmem_writedata),
    .io_dmem_memread(cpu76_io_dmem_memread),
    .io_dmem_memwrite(cpu76_io_dmem_memwrite),
    .io_dmem_maskmode(cpu76_io_dmem_maskmode),
    .io_dmem_sext(cpu76_io_dmem_sext),
    .io_dmem_readdata(cpu76_io_dmem_readdata)
  );
  DualPortedCombinMemory mem76 ( // @[top.scala 545:21]
    .clock(mem76_clock),
    .reset(mem76_reset),
    .io_imem_request_bits_address(mem76_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem76_io_imem_response_bits_data),
    .io_dmem_request_valid(mem76_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem76_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem76_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem76_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem76_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem76_io_dmem_response_bits_data)
  );
  ICombinMemPort imem76 ( // @[top.scala 546:22]
    .io_pipeline_address(imem76_io_pipeline_address),
    .io_pipeline_instruction(imem76_io_pipeline_instruction),
    .io_bus_request_bits_address(imem76_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem76_io_bus_response_bits_data)
  );
  DCombinMemPort dmem76 ( // @[top.scala 547:22]
    .clock(dmem76_clock),
    .reset(dmem76_reset),
    .io_pipeline_address(dmem76_io_pipeline_address),
    .io_pipeline_valid(dmem76_io_pipeline_valid),
    .io_pipeline_writedata(dmem76_io_pipeline_writedata),
    .io_pipeline_memread(dmem76_io_pipeline_memread),
    .io_pipeline_memwrite(dmem76_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem76_io_pipeline_maskmode),
    .io_pipeline_sext(dmem76_io_pipeline_sext),
    .io_pipeline_readdata(dmem76_io_pipeline_readdata),
    .io_bus_request_valid(dmem76_io_bus_request_valid),
    .io_bus_request_bits_address(dmem76_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem76_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem76_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem76_io_bus_response_valid),
    .io_bus_response_bits_data(dmem76_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu77 ( // @[top.scala 551:21]
    .clock(cpu77_clock),
    .reset(cpu77_reset),
    .io_imem_address(cpu77_io_imem_address),
    .io_imem_instruction(cpu77_io_imem_instruction),
    .io_dmem_address(cpu77_io_dmem_address),
    .io_dmem_valid(cpu77_io_dmem_valid),
    .io_dmem_writedata(cpu77_io_dmem_writedata),
    .io_dmem_memread(cpu77_io_dmem_memread),
    .io_dmem_memwrite(cpu77_io_dmem_memwrite),
    .io_dmem_maskmode(cpu77_io_dmem_maskmode),
    .io_dmem_sext(cpu77_io_dmem_sext),
    .io_dmem_readdata(cpu77_io_dmem_readdata)
  );
  DualPortedCombinMemory mem77 ( // @[top.scala 552:21]
    .clock(mem77_clock),
    .reset(mem77_reset),
    .io_imem_request_bits_address(mem77_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem77_io_imem_response_bits_data),
    .io_dmem_request_valid(mem77_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem77_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem77_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem77_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem77_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem77_io_dmem_response_bits_data)
  );
  ICombinMemPort imem77 ( // @[top.scala 553:22]
    .io_pipeline_address(imem77_io_pipeline_address),
    .io_pipeline_instruction(imem77_io_pipeline_instruction),
    .io_bus_request_bits_address(imem77_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem77_io_bus_response_bits_data)
  );
  DCombinMemPort dmem77 ( // @[top.scala 554:22]
    .clock(dmem77_clock),
    .reset(dmem77_reset),
    .io_pipeline_address(dmem77_io_pipeline_address),
    .io_pipeline_valid(dmem77_io_pipeline_valid),
    .io_pipeline_writedata(dmem77_io_pipeline_writedata),
    .io_pipeline_memread(dmem77_io_pipeline_memread),
    .io_pipeline_memwrite(dmem77_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem77_io_pipeline_maskmode),
    .io_pipeline_sext(dmem77_io_pipeline_sext),
    .io_pipeline_readdata(dmem77_io_pipeline_readdata),
    .io_bus_request_valid(dmem77_io_bus_request_valid),
    .io_bus_request_bits_address(dmem77_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem77_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem77_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem77_io_bus_response_valid),
    .io_bus_response_bits_data(dmem77_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu78 ( // @[top.scala 558:21]
    .clock(cpu78_clock),
    .reset(cpu78_reset),
    .io_imem_address(cpu78_io_imem_address),
    .io_imem_instruction(cpu78_io_imem_instruction),
    .io_dmem_address(cpu78_io_dmem_address),
    .io_dmem_valid(cpu78_io_dmem_valid),
    .io_dmem_writedata(cpu78_io_dmem_writedata),
    .io_dmem_memread(cpu78_io_dmem_memread),
    .io_dmem_memwrite(cpu78_io_dmem_memwrite),
    .io_dmem_maskmode(cpu78_io_dmem_maskmode),
    .io_dmem_sext(cpu78_io_dmem_sext),
    .io_dmem_readdata(cpu78_io_dmem_readdata)
  );
  DualPortedCombinMemory mem78 ( // @[top.scala 559:21]
    .clock(mem78_clock),
    .reset(mem78_reset),
    .io_imem_request_bits_address(mem78_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem78_io_imem_response_bits_data),
    .io_dmem_request_valid(mem78_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem78_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem78_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem78_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem78_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem78_io_dmem_response_bits_data)
  );
  ICombinMemPort imem78 ( // @[top.scala 560:22]
    .io_pipeline_address(imem78_io_pipeline_address),
    .io_pipeline_instruction(imem78_io_pipeline_instruction),
    .io_bus_request_bits_address(imem78_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem78_io_bus_response_bits_data)
  );
  DCombinMemPort dmem78 ( // @[top.scala 561:22]
    .clock(dmem78_clock),
    .reset(dmem78_reset),
    .io_pipeline_address(dmem78_io_pipeline_address),
    .io_pipeline_valid(dmem78_io_pipeline_valid),
    .io_pipeline_writedata(dmem78_io_pipeline_writedata),
    .io_pipeline_memread(dmem78_io_pipeline_memread),
    .io_pipeline_memwrite(dmem78_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem78_io_pipeline_maskmode),
    .io_pipeline_sext(dmem78_io_pipeline_sext),
    .io_pipeline_readdata(dmem78_io_pipeline_readdata),
    .io_bus_request_valid(dmem78_io_bus_request_valid),
    .io_bus_request_bits_address(dmem78_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem78_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem78_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem78_io_bus_response_valid),
    .io_bus_response_bits_data(dmem78_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu79 ( // @[top.scala 565:21]
    .clock(cpu79_clock),
    .reset(cpu79_reset),
    .io_imem_address(cpu79_io_imem_address),
    .io_imem_instruction(cpu79_io_imem_instruction),
    .io_dmem_address(cpu79_io_dmem_address),
    .io_dmem_valid(cpu79_io_dmem_valid),
    .io_dmem_writedata(cpu79_io_dmem_writedata),
    .io_dmem_memread(cpu79_io_dmem_memread),
    .io_dmem_memwrite(cpu79_io_dmem_memwrite),
    .io_dmem_maskmode(cpu79_io_dmem_maskmode),
    .io_dmem_sext(cpu79_io_dmem_sext),
    .io_dmem_readdata(cpu79_io_dmem_readdata)
  );
  DualPortedCombinMemory mem79 ( // @[top.scala 566:21]
    .clock(mem79_clock),
    .reset(mem79_reset),
    .io_imem_request_bits_address(mem79_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem79_io_imem_response_bits_data),
    .io_dmem_request_valid(mem79_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem79_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem79_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem79_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem79_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem79_io_dmem_response_bits_data)
  );
  ICombinMemPort imem79 ( // @[top.scala 567:22]
    .io_pipeline_address(imem79_io_pipeline_address),
    .io_pipeline_instruction(imem79_io_pipeline_instruction),
    .io_bus_request_bits_address(imem79_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem79_io_bus_response_bits_data)
  );
  DCombinMemPort dmem79 ( // @[top.scala 568:22]
    .clock(dmem79_clock),
    .reset(dmem79_reset),
    .io_pipeline_address(dmem79_io_pipeline_address),
    .io_pipeline_valid(dmem79_io_pipeline_valid),
    .io_pipeline_writedata(dmem79_io_pipeline_writedata),
    .io_pipeline_memread(dmem79_io_pipeline_memread),
    .io_pipeline_memwrite(dmem79_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem79_io_pipeline_maskmode),
    .io_pipeline_sext(dmem79_io_pipeline_sext),
    .io_pipeline_readdata(dmem79_io_pipeline_readdata),
    .io_bus_request_valid(dmem79_io_bus_request_valid),
    .io_bus_request_bits_address(dmem79_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem79_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem79_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem79_io_bus_response_valid),
    .io_bus_response_bits_data(dmem79_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu80 ( // @[top.scala 572:21]
    .clock(cpu80_clock),
    .reset(cpu80_reset),
    .io_imem_address(cpu80_io_imem_address),
    .io_imem_instruction(cpu80_io_imem_instruction),
    .io_dmem_address(cpu80_io_dmem_address),
    .io_dmem_valid(cpu80_io_dmem_valid),
    .io_dmem_writedata(cpu80_io_dmem_writedata),
    .io_dmem_memread(cpu80_io_dmem_memread),
    .io_dmem_memwrite(cpu80_io_dmem_memwrite),
    .io_dmem_maskmode(cpu80_io_dmem_maskmode),
    .io_dmem_sext(cpu80_io_dmem_sext),
    .io_dmem_readdata(cpu80_io_dmem_readdata)
  );
  DualPortedCombinMemory mem80 ( // @[top.scala 573:21]
    .clock(mem80_clock),
    .reset(mem80_reset),
    .io_imem_request_bits_address(mem80_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem80_io_imem_response_bits_data),
    .io_dmem_request_valid(mem80_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem80_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem80_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem80_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem80_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem80_io_dmem_response_bits_data)
  );
  ICombinMemPort imem80 ( // @[top.scala 574:22]
    .io_pipeline_address(imem80_io_pipeline_address),
    .io_pipeline_instruction(imem80_io_pipeline_instruction),
    .io_bus_request_bits_address(imem80_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem80_io_bus_response_bits_data)
  );
  DCombinMemPort dmem80 ( // @[top.scala 575:22]
    .clock(dmem80_clock),
    .reset(dmem80_reset),
    .io_pipeline_address(dmem80_io_pipeline_address),
    .io_pipeline_valid(dmem80_io_pipeline_valid),
    .io_pipeline_writedata(dmem80_io_pipeline_writedata),
    .io_pipeline_memread(dmem80_io_pipeline_memread),
    .io_pipeline_memwrite(dmem80_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem80_io_pipeline_maskmode),
    .io_pipeline_sext(dmem80_io_pipeline_sext),
    .io_pipeline_readdata(dmem80_io_pipeline_readdata),
    .io_bus_request_valid(dmem80_io_bus_request_valid),
    .io_bus_request_bits_address(dmem80_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem80_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem80_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem80_io_bus_response_valid),
    .io_bus_response_bits_data(dmem80_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu81 ( // @[top.scala 579:21]
    .clock(cpu81_clock),
    .reset(cpu81_reset),
    .io_imem_address(cpu81_io_imem_address),
    .io_imem_instruction(cpu81_io_imem_instruction),
    .io_dmem_address(cpu81_io_dmem_address),
    .io_dmem_valid(cpu81_io_dmem_valid),
    .io_dmem_writedata(cpu81_io_dmem_writedata),
    .io_dmem_memread(cpu81_io_dmem_memread),
    .io_dmem_memwrite(cpu81_io_dmem_memwrite),
    .io_dmem_maskmode(cpu81_io_dmem_maskmode),
    .io_dmem_sext(cpu81_io_dmem_sext),
    .io_dmem_readdata(cpu81_io_dmem_readdata)
  );
  DualPortedCombinMemory mem81 ( // @[top.scala 580:21]
    .clock(mem81_clock),
    .reset(mem81_reset),
    .io_imem_request_bits_address(mem81_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem81_io_imem_response_bits_data),
    .io_dmem_request_valid(mem81_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem81_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem81_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem81_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem81_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem81_io_dmem_response_bits_data)
  );
  ICombinMemPort imem81 ( // @[top.scala 581:22]
    .io_pipeline_address(imem81_io_pipeline_address),
    .io_pipeline_instruction(imem81_io_pipeline_instruction),
    .io_bus_request_bits_address(imem81_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem81_io_bus_response_bits_data)
  );
  DCombinMemPort dmem81 ( // @[top.scala 582:22]
    .clock(dmem81_clock),
    .reset(dmem81_reset),
    .io_pipeline_address(dmem81_io_pipeline_address),
    .io_pipeline_valid(dmem81_io_pipeline_valid),
    .io_pipeline_writedata(dmem81_io_pipeline_writedata),
    .io_pipeline_memread(dmem81_io_pipeline_memread),
    .io_pipeline_memwrite(dmem81_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem81_io_pipeline_maskmode),
    .io_pipeline_sext(dmem81_io_pipeline_sext),
    .io_pipeline_readdata(dmem81_io_pipeline_readdata),
    .io_bus_request_valid(dmem81_io_bus_request_valid),
    .io_bus_request_bits_address(dmem81_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem81_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem81_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem81_io_bus_response_valid),
    .io_bus_response_bits_data(dmem81_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu82 ( // @[top.scala 586:21]
    .clock(cpu82_clock),
    .reset(cpu82_reset),
    .io_imem_address(cpu82_io_imem_address),
    .io_imem_instruction(cpu82_io_imem_instruction),
    .io_dmem_address(cpu82_io_dmem_address),
    .io_dmem_valid(cpu82_io_dmem_valid),
    .io_dmem_writedata(cpu82_io_dmem_writedata),
    .io_dmem_memread(cpu82_io_dmem_memread),
    .io_dmem_memwrite(cpu82_io_dmem_memwrite),
    .io_dmem_maskmode(cpu82_io_dmem_maskmode),
    .io_dmem_sext(cpu82_io_dmem_sext),
    .io_dmem_readdata(cpu82_io_dmem_readdata)
  );
  DualPortedCombinMemory mem82 ( // @[top.scala 587:21]
    .clock(mem82_clock),
    .reset(mem82_reset),
    .io_imem_request_bits_address(mem82_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem82_io_imem_response_bits_data),
    .io_dmem_request_valid(mem82_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem82_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem82_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem82_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem82_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem82_io_dmem_response_bits_data)
  );
  ICombinMemPort imem82 ( // @[top.scala 588:22]
    .io_pipeline_address(imem82_io_pipeline_address),
    .io_pipeline_instruction(imem82_io_pipeline_instruction),
    .io_bus_request_bits_address(imem82_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem82_io_bus_response_bits_data)
  );
  DCombinMemPort dmem82 ( // @[top.scala 589:22]
    .clock(dmem82_clock),
    .reset(dmem82_reset),
    .io_pipeline_address(dmem82_io_pipeline_address),
    .io_pipeline_valid(dmem82_io_pipeline_valid),
    .io_pipeline_writedata(dmem82_io_pipeline_writedata),
    .io_pipeline_memread(dmem82_io_pipeline_memread),
    .io_pipeline_memwrite(dmem82_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem82_io_pipeline_maskmode),
    .io_pipeline_sext(dmem82_io_pipeline_sext),
    .io_pipeline_readdata(dmem82_io_pipeline_readdata),
    .io_bus_request_valid(dmem82_io_bus_request_valid),
    .io_bus_request_bits_address(dmem82_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem82_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem82_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem82_io_bus_response_valid),
    .io_bus_response_bits_data(dmem82_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu83 ( // @[top.scala 593:21]
    .clock(cpu83_clock),
    .reset(cpu83_reset),
    .io_imem_address(cpu83_io_imem_address),
    .io_imem_instruction(cpu83_io_imem_instruction),
    .io_dmem_address(cpu83_io_dmem_address),
    .io_dmem_valid(cpu83_io_dmem_valid),
    .io_dmem_writedata(cpu83_io_dmem_writedata),
    .io_dmem_memread(cpu83_io_dmem_memread),
    .io_dmem_memwrite(cpu83_io_dmem_memwrite),
    .io_dmem_maskmode(cpu83_io_dmem_maskmode),
    .io_dmem_sext(cpu83_io_dmem_sext),
    .io_dmem_readdata(cpu83_io_dmem_readdata)
  );
  DualPortedCombinMemory mem83 ( // @[top.scala 594:21]
    .clock(mem83_clock),
    .reset(mem83_reset),
    .io_imem_request_bits_address(mem83_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem83_io_imem_response_bits_data),
    .io_dmem_request_valid(mem83_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem83_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem83_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem83_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem83_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem83_io_dmem_response_bits_data)
  );
  ICombinMemPort imem83 ( // @[top.scala 595:22]
    .io_pipeline_address(imem83_io_pipeline_address),
    .io_pipeline_instruction(imem83_io_pipeline_instruction),
    .io_bus_request_bits_address(imem83_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem83_io_bus_response_bits_data)
  );
  DCombinMemPort dmem83 ( // @[top.scala 596:22]
    .clock(dmem83_clock),
    .reset(dmem83_reset),
    .io_pipeline_address(dmem83_io_pipeline_address),
    .io_pipeline_valid(dmem83_io_pipeline_valid),
    .io_pipeline_writedata(dmem83_io_pipeline_writedata),
    .io_pipeline_memread(dmem83_io_pipeline_memread),
    .io_pipeline_memwrite(dmem83_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem83_io_pipeline_maskmode),
    .io_pipeline_sext(dmem83_io_pipeline_sext),
    .io_pipeline_readdata(dmem83_io_pipeline_readdata),
    .io_bus_request_valid(dmem83_io_bus_request_valid),
    .io_bus_request_bits_address(dmem83_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem83_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem83_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem83_io_bus_response_valid),
    .io_bus_response_bits_data(dmem83_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu84 ( // @[top.scala 600:21]
    .clock(cpu84_clock),
    .reset(cpu84_reset),
    .io_imem_address(cpu84_io_imem_address),
    .io_imem_instruction(cpu84_io_imem_instruction),
    .io_dmem_address(cpu84_io_dmem_address),
    .io_dmem_valid(cpu84_io_dmem_valid),
    .io_dmem_writedata(cpu84_io_dmem_writedata),
    .io_dmem_memread(cpu84_io_dmem_memread),
    .io_dmem_memwrite(cpu84_io_dmem_memwrite),
    .io_dmem_maskmode(cpu84_io_dmem_maskmode),
    .io_dmem_sext(cpu84_io_dmem_sext),
    .io_dmem_readdata(cpu84_io_dmem_readdata)
  );
  DualPortedCombinMemory mem84 ( // @[top.scala 601:21]
    .clock(mem84_clock),
    .reset(mem84_reset),
    .io_imem_request_bits_address(mem84_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem84_io_imem_response_bits_data),
    .io_dmem_request_valid(mem84_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem84_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem84_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem84_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem84_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem84_io_dmem_response_bits_data)
  );
  ICombinMemPort imem84 ( // @[top.scala 602:22]
    .io_pipeline_address(imem84_io_pipeline_address),
    .io_pipeline_instruction(imem84_io_pipeline_instruction),
    .io_bus_request_bits_address(imem84_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem84_io_bus_response_bits_data)
  );
  DCombinMemPort dmem84 ( // @[top.scala 603:22]
    .clock(dmem84_clock),
    .reset(dmem84_reset),
    .io_pipeline_address(dmem84_io_pipeline_address),
    .io_pipeline_valid(dmem84_io_pipeline_valid),
    .io_pipeline_writedata(dmem84_io_pipeline_writedata),
    .io_pipeline_memread(dmem84_io_pipeline_memread),
    .io_pipeline_memwrite(dmem84_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem84_io_pipeline_maskmode),
    .io_pipeline_sext(dmem84_io_pipeline_sext),
    .io_pipeline_readdata(dmem84_io_pipeline_readdata),
    .io_bus_request_valid(dmem84_io_bus_request_valid),
    .io_bus_request_bits_address(dmem84_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem84_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem84_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem84_io_bus_response_valid),
    .io_bus_response_bits_data(dmem84_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu85 ( // @[top.scala 607:21]
    .clock(cpu85_clock),
    .reset(cpu85_reset),
    .io_imem_address(cpu85_io_imem_address),
    .io_imem_instruction(cpu85_io_imem_instruction),
    .io_dmem_address(cpu85_io_dmem_address),
    .io_dmem_valid(cpu85_io_dmem_valid),
    .io_dmem_writedata(cpu85_io_dmem_writedata),
    .io_dmem_memread(cpu85_io_dmem_memread),
    .io_dmem_memwrite(cpu85_io_dmem_memwrite),
    .io_dmem_maskmode(cpu85_io_dmem_maskmode),
    .io_dmem_sext(cpu85_io_dmem_sext),
    .io_dmem_readdata(cpu85_io_dmem_readdata)
  );
  DualPortedCombinMemory mem85 ( // @[top.scala 608:21]
    .clock(mem85_clock),
    .reset(mem85_reset),
    .io_imem_request_bits_address(mem85_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem85_io_imem_response_bits_data),
    .io_dmem_request_valid(mem85_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem85_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem85_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem85_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem85_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem85_io_dmem_response_bits_data)
  );
  ICombinMemPort imem85 ( // @[top.scala 609:22]
    .io_pipeline_address(imem85_io_pipeline_address),
    .io_pipeline_instruction(imem85_io_pipeline_instruction),
    .io_bus_request_bits_address(imem85_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem85_io_bus_response_bits_data)
  );
  DCombinMemPort dmem85 ( // @[top.scala 610:22]
    .clock(dmem85_clock),
    .reset(dmem85_reset),
    .io_pipeline_address(dmem85_io_pipeline_address),
    .io_pipeline_valid(dmem85_io_pipeline_valid),
    .io_pipeline_writedata(dmem85_io_pipeline_writedata),
    .io_pipeline_memread(dmem85_io_pipeline_memread),
    .io_pipeline_memwrite(dmem85_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem85_io_pipeline_maskmode),
    .io_pipeline_sext(dmem85_io_pipeline_sext),
    .io_pipeline_readdata(dmem85_io_pipeline_readdata),
    .io_bus_request_valid(dmem85_io_bus_request_valid),
    .io_bus_request_bits_address(dmem85_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem85_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem85_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem85_io_bus_response_valid),
    .io_bus_response_bits_data(dmem85_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu86 ( // @[top.scala 614:21]
    .clock(cpu86_clock),
    .reset(cpu86_reset),
    .io_imem_address(cpu86_io_imem_address),
    .io_imem_instruction(cpu86_io_imem_instruction),
    .io_dmem_address(cpu86_io_dmem_address),
    .io_dmem_valid(cpu86_io_dmem_valid),
    .io_dmem_writedata(cpu86_io_dmem_writedata),
    .io_dmem_memread(cpu86_io_dmem_memread),
    .io_dmem_memwrite(cpu86_io_dmem_memwrite),
    .io_dmem_maskmode(cpu86_io_dmem_maskmode),
    .io_dmem_sext(cpu86_io_dmem_sext),
    .io_dmem_readdata(cpu86_io_dmem_readdata)
  );
  DualPortedCombinMemory mem86 ( // @[top.scala 615:21]
    .clock(mem86_clock),
    .reset(mem86_reset),
    .io_imem_request_bits_address(mem86_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem86_io_imem_response_bits_data),
    .io_dmem_request_valid(mem86_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem86_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem86_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem86_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem86_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem86_io_dmem_response_bits_data)
  );
  ICombinMemPort imem86 ( // @[top.scala 616:22]
    .io_pipeline_address(imem86_io_pipeline_address),
    .io_pipeline_instruction(imem86_io_pipeline_instruction),
    .io_bus_request_bits_address(imem86_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem86_io_bus_response_bits_data)
  );
  DCombinMemPort dmem86 ( // @[top.scala 617:22]
    .clock(dmem86_clock),
    .reset(dmem86_reset),
    .io_pipeline_address(dmem86_io_pipeline_address),
    .io_pipeline_valid(dmem86_io_pipeline_valid),
    .io_pipeline_writedata(dmem86_io_pipeline_writedata),
    .io_pipeline_memread(dmem86_io_pipeline_memread),
    .io_pipeline_memwrite(dmem86_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem86_io_pipeline_maskmode),
    .io_pipeline_sext(dmem86_io_pipeline_sext),
    .io_pipeline_readdata(dmem86_io_pipeline_readdata),
    .io_bus_request_valid(dmem86_io_bus_request_valid),
    .io_bus_request_bits_address(dmem86_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem86_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem86_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem86_io_bus_response_valid),
    .io_bus_response_bits_data(dmem86_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu87 ( // @[top.scala 621:21]
    .clock(cpu87_clock),
    .reset(cpu87_reset),
    .io_imem_address(cpu87_io_imem_address),
    .io_imem_instruction(cpu87_io_imem_instruction),
    .io_dmem_address(cpu87_io_dmem_address),
    .io_dmem_valid(cpu87_io_dmem_valid),
    .io_dmem_writedata(cpu87_io_dmem_writedata),
    .io_dmem_memread(cpu87_io_dmem_memread),
    .io_dmem_memwrite(cpu87_io_dmem_memwrite),
    .io_dmem_maskmode(cpu87_io_dmem_maskmode),
    .io_dmem_sext(cpu87_io_dmem_sext),
    .io_dmem_readdata(cpu87_io_dmem_readdata)
  );
  DualPortedCombinMemory mem87 ( // @[top.scala 622:21]
    .clock(mem87_clock),
    .reset(mem87_reset),
    .io_imem_request_bits_address(mem87_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem87_io_imem_response_bits_data),
    .io_dmem_request_valid(mem87_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem87_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem87_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem87_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem87_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem87_io_dmem_response_bits_data)
  );
  ICombinMemPort imem87 ( // @[top.scala 623:22]
    .io_pipeline_address(imem87_io_pipeline_address),
    .io_pipeline_instruction(imem87_io_pipeline_instruction),
    .io_bus_request_bits_address(imem87_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem87_io_bus_response_bits_data)
  );
  DCombinMemPort dmem87 ( // @[top.scala 624:22]
    .clock(dmem87_clock),
    .reset(dmem87_reset),
    .io_pipeline_address(dmem87_io_pipeline_address),
    .io_pipeline_valid(dmem87_io_pipeline_valid),
    .io_pipeline_writedata(dmem87_io_pipeline_writedata),
    .io_pipeline_memread(dmem87_io_pipeline_memread),
    .io_pipeline_memwrite(dmem87_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem87_io_pipeline_maskmode),
    .io_pipeline_sext(dmem87_io_pipeline_sext),
    .io_pipeline_readdata(dmem87_io_pipeline_readdata),
    .io_bus_request_valid(dmem87_io_bus_request_valid),
    .io_bus_request_bits_address(dmem87_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem87_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem87_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem87_io_bus_response_valid),
    .io_bus_response_bits_data(dmem87_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu88 ( // @[top.scala 628:21]
    .clock(cpu88_clock),
    .reset(cpu88_reset),
    .io_imem_address(cpu88_io_imem_address),
    .io_imem_instruction(cpu88_io_imem_instruction),
    .io_dmem_address(cpu88_io_dmem_address),
    .io_dmem_valid(cpu88_io_dmem_valid),
    .io_dmem_writedata(cpu88_io_dmem_writedata),
    .io_dmem_memread(cpu88_io_dmem_memread),
    .io_dmem_memwrite(cpu88_io_dmem_memwrite),
    .io_dmem_maskmode(cpu88_io_dmem_maskmode),
    .io_dmem_sext(cpu88_io_dmem_sext),
    .io_dmem_readdata(cpu88_io_dmem_readdata)
  );
  DualPortedCombinMemory mem88 ( // @[top.scala 629:21]
    .clock(mem88_clock),
    .reset(mem88_reset),
    .io_imem_request_bits_address(mem88_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem88_io_imem_response_bits_data),
    .io_dmem_request_valid(mem88_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem88_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem88_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem88_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem88_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem88_io_dmem_response_bits_data)
  );
  ICombinMemPort imem88 ( // @[top.scala 630:22]
    .io_pipeline_address(imem88_io_pipeline_address),
    .io_pipeline_instruction(imem88_io_pipeline_instruction),
    .io_bus_request_bits_address(imem88_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem88_io_bus_response_bits_data)
  );
  DCombinMemPort dmem88 ( // @[top.scala 631:22]
    .clock(dmem88_clock),
    .reset(dmem88_reset),
    .io_pipeline_address(dmem88_io_pipeline_address),
    .io_pipeline_valid(dmem88_io_pipeline_valid),
    .io_pipeline_writedata(dmem88_io_pipeline_writedata),
    .io_pipeline_memread(dmem88_io_pipeline_memread),
    .io_pipeline_memwrite(dmem88_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem88_io_pipeline_maskmode),
    .io_pipeline_sext(dmem88_io_pipeline_sext),
    .io_pipeline_readdata(dmem88_io_pipeline_readdata),
    .io_bus_request_valid(dmem88_io_bus_request_valid),
    .io_bus_request_bits_address(dmem88_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem88_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem88_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem88_io_bus_response_valid),
    .io_bus_response_bits_data(dmem88_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu89 ( // @[top.scala 635:21]
    .clock(cpu89_clock),
    .reset(cpu89_reset),
    .io_imem_address(cpu89_io_imem_address),
    .io_imem_instruction(cpu89_io_imem_instruction),
    .io_dmem_address(cpu89_io_dmem_address),
    .io_dmem_valid(cpu89_io_dmem_valid),
    .io_dmem_writedata(cpu89_io_dmem_writedata),
    .io_dmem_memread(cpu89_io_dmem_memread),
    .io_dmem_memwrite(cpu89_io_dmem_memwrite),
    .io_dmem_maskmode(cpu89_io_dmem_maskmode),
    .io_dmem_sext(cpu89_io_dmem_sext),
    .io_dmem_readdata(cpu89_io_dmem_readdata)
  );
  DualPortedCombinMemory mem89 ( // @[top.scala 636:21]
    .clock(mem89_clock),
    .reset(mem89_reset),
    .io_imem_request_bits_address(mem89_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem89_io_imem_response_bits_data),
    .io_dmem_request_valid(mem89_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem89_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem89_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem89_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem89_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem89_io_dmem_response_bits_data)
  );
  ICombinMemPort imem89 ( // @[top.scala 637:22]
    .io_pipeline_address(imem89_io_pipeline_address),
    .io_pipeline_instruction(imem89_io_pipeline_instruction),
    .io_bus_request_bits_address(imem89_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem89_io_bus_response_bits_data)
  );
  DCombinMemPort dmem89 ( // @[top.scala 638:22]
    .clock(dmem89_clock),
    .reset(dmem89_reset),
    .io_pipeline_address(dmem89_io_pipeline_address),
    .io_pipeline_valid(dmem89_io_pipeline_valid),
    .io_pipeline_writedata(dmem89_io_pipeline_writedata),
    .io_pipeline_memread(dmem89_io_pipeline_memread),
    .io_pipeline_memwrite(dmem89_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem89_io_pipeline_maskmode),
    .io_pipeline_sext(dmem89_io_pipeline_sext),
    .io_pipeline_readdata(dmem89_io_pipeline_readdata),
    .io_bus_request_valid(dmem89_io_bus_request_valid),
    .io_bus_request_bits_address(dmem89_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem89_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem89_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem89_io_bus_response_valid),
    .io_bus_response_bits_data(dmem89_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu90 ( // @[top.scala 642:21]
    .clock(cpu90_clock),
    .reset(cpu90_reset),
    .io_imem_address(cpu90_io_imem_address),
    .io_imem_instruction(cpu90_io_imem_instruction),
    .io_dmem_address(cpu90_io_dmem_address),
    .io_dmem_valid(cpu90_io_dmem_valid),
    .io_dmem_writedata(cpu90_io_dmem_writedata),
    .io_dmem_memread(cpu90_io_dmem_memread),
    .io_dmem_memwrite(cpu90_io_dmem_memwrite),
    .io_dmem_maskmode(cpu90_io_dmem_maskmode),
    .io_dmem_sext(cpu90_io_dmem_sext),
    .io_dmem_readdata(cpu90_io_dmem_readdata)
  );
  DualPortedCombinMemory mem90 ( // @[top.scala 643:21]
    .clock(mem90_clock),
    .reset(mem90_reset),
    .io_imem_request_bits_address(mem90_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem90_io_imem_response_bits_data),
    .io_dmem_request_valid(mem90_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem90_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem90_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem90_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem90_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem90_io_dmem_response_bits_data)
  );
  ICombinMemPort imem90 ( // @[top.scala 644:22]
    .io_pipeline_address(imem90_io_pipeline_address),
    .io_pipeline_instruction(imem90_io_pipeline_instruction),
    .io_bus_request_bits_address(imem90_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem90_io_bus_response_bits_data)
  );
  DCombinMemPort dmem90 ( // @[top.scala 645:22]
    .clock(dmem90_clock),
    .reset(dmem90_reset),
    .io_pipeline_address(dmem90_io_pipeline_address),
    .io_pipeline_valid(dmem90_io_pipeline_valid),
    .io_pipeline_writedata(dmem90_io_pipeline_writedata),
    .io_pipeline_memread(dmem90_io_pipeline_memread),
    .io_pipeline_memwrite(dmem90_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem90_io_pipeline_maskmode),
    .io_pipeline_sext(dmem90_io_pipeline_sext),
    .io_pipeline_readdata(dmem90_io_pipeline_readdata),
    .io_bus_request_valid(dmem90_io_bus_request_valid),
    .io_bus_request_bits_address(dmem90_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem90_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem90_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem90_io_bus_response_valid),
    .io_bus_response_bits_data(dmem90_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu91 ( // @[top.scala 649:21]
    .clock(cpu91_clock),
    .reset(cpu91_reset),
    .io_imem_address(cpu91_io_imem_address),
    .io_imem_instruction(cpu91_io_imem_instruction),
    .io_dmem_address(cpu91_io_dmem_address),
    .io_dmem_valid(cpu91_io_dmem_valid),
    .io_dmem_writedata(cpu91_io_dmem_writedata),
    .io_dmem_memread(cpu91_io_dmem_memread),
    .io_dmem_memwrite(cpu91_io_dmem_memwrite),
    .io_dmem_maskmode(cpu91_io_dmem_maskmode),
    .io_dmem_sext(cpu91_io_dmem_sext),
    .io_dmem_readdata(cpu91_io_dmem_readdata)
  );
  DualPortedCombinMemory mem91 ( // @[top.scala 650:21]
    .clock(mem91_clock),
    .reset(mem91_reset),
    .io_imem_request_bits_address(mem91_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem91_io_imem_response_bits_data),
    .io_dmem_request_valid(mem91_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem91_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem91_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem91_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem91_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem91_io_dmem_response_bits_data)
  );
  ICombinMemPort imem91 ( // @[top.scala 651:22]
    .io_pipeline_address(imem91_io_pipeline_address),
    .io_pipeline_instruction(imem91_io_pipeline_instruction),
    .io_bus_request_bits_address(imem91_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem91_io_bus_response_bits_data)
  );
  DCombinMemPort dmem91 ( // @[top.scala 652:22]
    .clock(dmem91_clock),
    .reset(dmem91_reset),
    .io_pipeline_address(dmem91_io_pipeline_address),
    .io_pipeline_valid(dmem91_io_pipeline_valid),
    .io_pipeline_writedata(dmem91_io_pipeline_writedata),
    .io_pipeline_memread(dmem91_io_pipeline_memread),
    .io_pipeline_memwrite(dmem91_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem91_io_pipeline_maskmode),
    .io_pipeline_sext(dmem91_io_pipeline_sext),
    .io_pipeline_readdata(dmem91_io_pipeline_readdata),
    .io_bus_request_valid(dmem91_io_bus_request_valid),
    .io_bus_request_bits_address(dmem91_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem91_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem91_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem91_io_bus_response_valid),
    .io_bus_response_bits_data(dmem91_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu92 ( // @[top.scala 656:21]
    .clock(cpu92_clock),
    .reset(cpu92_reset),
    .io_imem_address(cpu92_io_imem_address),
    .io_imem_instruction(cpu92_io_imem_instruction),
    .io_dmem_address(cpu92_io_dmem_address),
    .io_dmem_valid(cpu92_io_dmem_valid),
    .io_dmem_writedata(cpu92_io_dmem_writedata),
    .io_dmem_memread(cpu92_io_dmem_memread),
    .io_dmem_memwrite(cpu92_io_dmem_memwrite),
    .io_dmem_maskmode(cpu92_io_dmem_maskmode),
    .io_dmem_sext(cpu92_io_dmem_sext),
    .io_dmem_readdata(cpu92_io_dmem_readdata)
  );
  DualPortedCombinMemory mem92 ( // @[top.scala 657:21]
    .clock(mem92_clock),
    .reset(mem92_reset),
    .io_imem_request_bits_address(mem92_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem92_io_imem_response_bits_data),
    .io_dmem_request_valid(mem92_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem92_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem92_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem92_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem92_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem92_io_dmem_response_bits_data)
  );
  ICombinMemPort imem92 ( // @[top.scala 658:22]
    .io_pipeline_address(imem92_io_pipeline_address),
    .io_pipeline_instruction(imem92_io_pipeline_instruction),
    .io_bus_request_bits_address(imem92_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem92_io_bus_response_bits_data)
  );
  DCombinMemPort dmem92 ( // @[top.scala 659:22]
    .clock(dmem92_clock),
    .reset(dmem92_reset),
    .io_pipeline_address(dmem92_io_pipeline_address),
    .io_pipeline_valid(dmem92_io_pipeline_valid),
    .io_pipeline_writedata(dmem92_io_pipeline_writedata),
    .io_pipeline_memread(dmem92_io_pipeline_memread),
    .io_pipeline_memwrite(dmem92_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem92_io_pipeline_maskmode),
    .io_pipeline_sext(dmem92_io_pipeline_sext),
    .io_pipeline_readdata(dmem92_io_pipeline_readdata),
    .io_bus_request_valid(dmem92_io_bus_request_valid),
    .io_bus_request_bits_address(dmem92_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem92_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem92_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem92_io_bus_response_valid),
    .io_bus_response_bits_data(dmem92_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu93 ( // @[top.scala 663:21]
    .clock(cpu93_clock),
    .reset(cpu93_reset),
    .io_imem_address(cpu93_io_imem_address),
    .io_imem_instruction(cpu93_io_imem_instruction),
    .io_dmem_address(cpu93_io_dmem_address),
    .io_dmem_valid(cpu93_io_dmem_valid),
    .io_dmem_writedata(cpu93_io_dmem_writedata),
    .io_dmem_memread(cpu93_io_dmem_memread),
    .io_dmem_memwrite(cpu93_io_dmem_memwrite),
    .io_dmem_maskmode(cpu93_io_dmem_maskmode),
    .io_dmem_sext(cpu93_io_dmem_sext),
    .io_dmem_readdata(cpu93_io_dmem_readdata)
  );
  DualPortedCombinMemory mem93 ( // @[top.scala 664:21]
    .clock(mem93_clock),
    .reset(mem93_reset),
    .io_imem_request_bits_address(mem93_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem93_io_imem_response_bits_data),
    .io_dmem_request_valid(mem93_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem93_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem93_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem93_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem93_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem93_io_dmem_response_bits_data)
  );
  ICombinMemPort imem93 ( // @[top.scala 665:22]
    .io_pipeline_address(imem93_io_pipeline_address),
    .io_pipeline_instruction(imem93_io_pipeline_instruction),
    .io_bus_request_bits_address(imem93_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem93_io_bus_response_bits_data)
  );
  DCombinMemPort dmem93 ( // @[top.scala 666:22]
    .clock(dmem93_clock),
    .reset(dmem93_reset),
    .io_pipeline_address(dmem93_io_pipeline_address),
    .io_pipeline_valid(dmem93_io_pipeline_valid),
    .io_pipeline_writedata(dmem93_io_pipeline_writedata),
    .io_pipeline_memread(dmem93_io_pipeline_memread),
    .io_pipeline_memwrite(dmem93_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem93_io_pipeline_maskmode),
    .io_pipeline_sext(dmem93_io_pipeline_sext),
    .io_pipeline_readdata(dmem93_io_pipeline_readdata),
    .io_bus_request_valid(dmem93_io_bus_request_valid),
    .io_bus_request_bits_address(dmem93_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem93_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem93_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem93_io_bus_response_valid),
    .io_bus_response_bits_data(dmem93_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu94 ( // @[top.scala 670:21]
    .clock(cpu94_clock),
    .reset(cpu94_reset),
    .io_imem_address(cpu94_io_imem_address),
    .io_imem_instruction(cpu94_io_imem_instruction),
    .io_dmem_address(cpu94_io_dmem_address),
    .io_dmem_valid(cpu94_io_dmem_valid),
    .io_dmem_writedata(cpu94_io_dmem_writedata),
    .io_dmem_memread(cpu94_io_dmem_memread),
    .io_dmem_memwrite(cpu94_io_dmem_memwrite),
    .io_dmem_maskmode(cpu94_io_dmem_maskmode),
    .io_dmem_sext(cpu94_io_dmem_sext),
    .io_dmem_readdata(cpu94_io_dmem_readdata)
  );
  DualPortedCombinMemory mem94 ( // @[top.scala 671:21]
    .clock(mem94_clock),
    .reset(mem94_reset),
    .io_imem_request_bits_address(mem94_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem94_io_imem_response_bits_data),
    .io_dmem_request_valid(mem94_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem94_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem94_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem94_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem94_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem94_io_dmem_response_bits_data)
  );
  ICombinMemPort imem94 ( // @[top.scala 672:22]
    .io_pipeline_address(imem94_io_pipeline_address),
    .io_pipeline_instruction(imem94_io_pipeline_instruction),
    .io_bus_request_bits_address(imem94_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem94_io_bus_response_bits_data)
  );
  DCombinMemPort dmem94 ( // @[top.scala 673:22]
    .clock(dmem94_clock),
    .reset(dmem94_reset),
    .io_pipeline_address(dmem94_io_pipeline_address),
    .io_pipeline_valid(dmem94_io_pipeline_valid),
    .io_pipeline_writedata(dmem94_io_pipeline_writedata),
    .io_pipeline_memread(dmem94_io_pipeline_memread),
    .io_pipeline_memwrite(dmem94_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem94_io_pipeline_maskmode),
    .io_pipeline_sext(dmem94_io_pipeline_sext),
    .io_pipeline_readdata(dmem94_io_pipeline_readdata),
    .io_bus_request_valid(dmem94_io_bus_request_valid),
    .io_bus_request_bits_address(dmem94_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem94_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem94_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem94_io_bus_response_valid),
    .io_bus_response_bits_data(dmem94_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu95 ( // @[top.scala 677:21]
    .clock(cpu95_clock),
    .reset(cpu95_reset),
    .io_imem_address(cpu95_io_imem_address),
    .io_imem_instruction(cpu95_io_imem_instruction),
    .io_dmem_address(cpu95_io_dmem_address),
    .io_dmem_valid(cpu95_io_dmem_valid),
    .io_dmem_writedata(cpu95_io_dmem_writedata),
    .io_dmem_memread(cpu95_io_dmem_memread),
    .io_dmem_memwrite(cpu95_io_dmem_memwrite),
    .io_dmem_maskmode(cpu95_io_dmem_maskmode),
    .io_dmem_sext(cpu95_io_dmem_sext),
    .io_dmem_readdata(cpu95_io_dmem_readdata)
  );
  DualPortedCombinMemory mem95 ( // @[top.scala 678:21]
    .clock(mem95_clock),
    .reset(mem95_reset),
    .io_imem_request_bits_address(mem95_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem95_io_imem_response_bits_data),
    .io_dmem_request_valid(mem95_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem95_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem95_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem95_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem95_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem95_io_dmem_response_bits_data)
  );
  ICombinMemPort imem95 ( // @[top.scala 679:22]
    .io_pipeline_address(imem95_io_pipeline_address),
    .io_pipeline_instruction(imem95_io_pipeline_instruction),
    .io_bus_request_bits_address(imem95_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem95_io_bus_response_bits_data)
  );
  DCombinMemPort dmem95 ( // @[top.scala 680:22]
    .clock(dmem95_clock),
    .reset(dmem95_reset),
    .io_pipeline_address(dmem95_io_pipeline_address),
    .io_pipeline_valid(dmem95_io_pipeline_valid),
    .io_pipeline_writedata(dmem95_io_pipeline_writedata),
    .io_pipeline_memread(dmem95_io_pipeline_memread),
    .io_pipeline_memwrite(dmem95_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem95_io_pipeline_maskmode),
    .io_pipeline_sext(dmem95_io_pipeline_sext),
    .io_pipeline_readdata(dmem95_io_pipeline_readdata),
    .io_bus_request_valid(dmem95_io_bus_request_valid),
    .io_bus_request_bits_address(dmem95_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem95_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem95_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem95_io_bus_response_valid),
    .io_bus_response_bits_data(dmem95_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu96 ( // @[top.scala 684:21]
    .clock(cpu96_clock),
    .reset(cpu96_reset),
    .io_imem_address(cpu96_io_imem_address),
    .io_imem_instruction(cpu96_io_imem_instruction),
    .io_dmem_address(cpu96_io_dmem_address),
    .io_dmem_valid(cpu96_io_dmem_valid),
    .io_dmem_writedata(cpu96_io_dmem_writedata),
    .io_dmem_memread(cpu96_io_dmem_memread),
    .io_dmem_memwrite(cpu96_io_dmem_memwrite),
    .io_dmem_maskmode(cpu96_io_dmem_maskmode),
    .io_dmem_sext(cpu96_io_dmem_sext),
    .io_dmem_readdata(cpu96_io_dmem_readdata)
  );
  DualPortedCombinMemory mem96 ( // @[top.scala 685:21]
    .clock(mem96_clock),
    .reset(mem96_reset),
    .io_imem_request_bits_address(mem96_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem96_io_imem_response_bits_data),
    .io_dmem_request_valid(mem96_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem96_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem96_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem96_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem96_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem96_io_dmem_response_bits_data)
  );
  ICombinMemPort imem96 ( // @[top.scala 686:22]
    .io_pipeline_address(imem96_io_pipeline_address),
    .io_pipeline_instruction(imem96_io_pipeline_instruction),
    .io_bus_request_bits_address(imem96_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem96_io_bus_response_bits_data)
  );
  DCombinMemPort dmem96 ( // @[top.scala 687:22]
    .clock(dmem96_clock),
    .reset(dmem96_reset),
    .io_pipeline_address(dmem96_io_pipeline_address),
    .io_pipeline_valid(dmem96_io_pipeline_valid),
    .io_pipeline_writedata(dmem96_io_pipeline_writedata),
    .io_pipeline_memread(dmem96_io_pipeline_memread),
    .io_pipeline_memwrite(dmem96_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem96_io_pipeline_maskmode),
    .io_pipeline_sext(dmem96_io_pipeline_sext),
    .io_pipeline_readdata(dmem96_io_pipeline_readdata),
    .io_bus_request_valid(dmem96_io_bus_request_valid),
    .io_bus_request_bits_address(dmem96_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem96_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem96_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem96_io_bus_response_valid),
    .io_bus_response_bits_data(dmem96_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu97 ( // @[top.scala 691:21]
    .clock(cpu97_clock),
    .reset(cpu97_reset),
    .io_imem_address(cpu97_io_imem_address),
    .io_imem_instruction(cpu97_io_imem_instruction),
    .io_dmem_address(cpu97_io_dmem_address),
    .io_dmem_valid(cpu97_io_dmem_valid),
    .io_dmem_writedata(cpu97_io_dmem_writedata),
    .io_dmem_memread(cpu97_io_dmem_memread),
    .io_dmem_memwrite(cpu97_io_dmem_memwrite),
    .io_dmem_maskmode(cpu97_io_dmem_maskmode),
    .io_dmem_sext(cpu97_io_dmem_sext),
    .io_dmem_readdata(cpu97_io_dmem_readdata)
  );
  DualPortedCombinMemory mem97 ( // @[top.scala 692:21]
    .clock(mem97_clock),
    .reset(mem97_reset),
    .io_imem_request_bits_address(mem97_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem97_io_imem_response_bits_data),
    .io_dmem_request_valid(mem97_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem97_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem97_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem97_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem97_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem97_io_dmem_response_bits_data)
  );
  ICombinMemPort imem97 ( // @[top.scala 693:22]
    .io_pipeline_address(imem97_io_pipeline_address),
    .io_pipeline_instruction(imem97_io_pipeline_instruction),
    .io_bus_request_bits_address(imem97_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem97_io_bus_response_bits_data)
  );
  DCombinMemPort dmem97 ( // @[top.scala 694:22]
    .clock(dmem97_clock),
    .reset(dmem97_reset),
    .io_pipeline_address(dmem97_io_pipeline_address),
    .io_pipeline_valid(dmem97_io_pipeline_valid),
    .io_pipeline_writedata(dmem97_io_pipeline_writedata),
    .io_pipeline_memread(dmem97_io_pipeline_memread),
    .io_pipeline_memwrite(dmem97_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem97_io_pipeline_maskmode),
    .io_pipeline_sext(dmem97_io_pipeline_sext),
    .io_pipeline_readdata(dmem97_io_pipeline_readdata),
    .io_bus_request_valid(dmem97_io_bus_request_valid),
    .io_bus_request_bits_address(dmem97_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem97_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem97_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem97_io_bus_response_valid),
    .io_bus_response_bits_data(dmem97_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu98 ( // @[top.scala 698:21]
    .clock(cpu98_clock),
    .reset(cpu98_reset),
    .io_imem_address(cpu98_io_imem_address),
    .io_imem_instruction(cpu98_io_imem_instruction),
    .io_dmem_address(cpu98_io_dmem_address),
    .io_dmem_valid(cpu98_io_dmem_valid),
    .io_dmem_writedata(cpu98_io_dmem_writedata),
    .io_dmem_memread(cpu98_io_dmem_memread),
    .io_dmem_memwrite(cpu98_io_dmem_memwrite),
    .io_dmem_maskmode(cpu98_io_dmem_maskmode),
    .io_dmem_sext(cpu98_io_dmem_sext),
    .io_dmem_readdata(cpu98_io_dmem_readdata)
  );
  DualPortedCombinMemory mem98 ( // @[top.scala 699:21]
    .clock(mem98_clock),
    .reset(mem98_reset),
    .io_imem_request_bits_address(mem98_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem98_io_imem_response_bits_data),
    .io_dmem_request_valid(mem98_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem98_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem98_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem98_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem98_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem98_io_dmem_response_bits_data)
  );
  ICombinMemPort imem98 ( // @[top.scala 700:22]
    .io_pipeline_address(imem98_io_pipeline_address),
    .io_pipeline_instruction(imem98_io_pipeline_instruction),
    .io_bus_request_bits_address(imem98_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem98_io_bus_response_bits_data)
  );
  DCombinMemPort dmem98 ( // @[top.scala 701:22]
    .clock(dmem98_clock),
    .reset(dmem98_reset),
    .io_pipeline_address(dmem98_io_pipeline_address),
    .io_pipeline_valid(dmem98_io_pipeline_valid),
    .io_pipeline_writedata(dmem98_io_pipeline_writedata),
    .io_pipeline_memread(dmem98_io_pipeline_memread),
    .io_pipeline_memwrite(dmem98_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem98_io_pipeline_maskmode),
    .io_pipeline_sext(dmem98_io_pipeline_sext),
    .io_pipeline_readdata(dmem98_io_pipeline_readdata),
    .io_bus_request_valid(dmem98_io_bus_request_valid),
    .io_bus_request_bits_address(dmem98_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem98_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem98_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem98_io_bus_response_valid),
    .io_bus_response_bits_data(dmem98_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu99 ( // @[top.scala 705:21]
    .clock(cpu99_clock),
    .reset(cpu99_reset),
    .io_imem_address(cpu99_io_imem_address),
    .io_imem_instruction(cpu99_io_imem_instruction),
    .io_dmem_address(cpu99_io_dmem_address),
    .io_dmem_valid(cpu99_io_dmem_valid),
    .io_dmem_writedata(cpu99_io_dmem_writedata),
    .io_dmem_memread(cpu99_io_dmem_memread),
    .io_dmem_memwrite(cpu99_io_dmem_memwrite),
    .io_dmem_maskmode(cpu99_io_dmem_maskmode),
    .io_dmem_sext(cpu99_io_dmem_sext),
    .io_dmem_readdata(cpu99_io_dmem_readdata)
  );
  DualPortedCombinMemory mem99 ( // @[top.scala 706:21]
    .clock(mem99_clock),
    .reset(mem99_reset),
    .io_imem_request_bits_address(mem99_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem99_io_imem_response_bits_data),
    .io_dmem_request_valid(mem99_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem99_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem99_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem99_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem99_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem99_io_dmem_response_bits_data)
  );
  ICombinMemPort imem99 ( // @[top.scala 707:22]
    .io_pipeline_address(imem99_io_pipeline_address),
    .io_pipeline_instruction(imem99_io_pipeline_instruction),
    .io_bus_request_bits_address(imem99_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem99_io_bus_response_bits_data)
  );
  DCombinMemPort dmem99 ( // @[top.scala 708:22]
    .clock(dmem99_clock),
    .reset(dmem99_reset),
    .io_pipeline_address(dmem99_io_pipeline_address),
    .io_pipeline_valid(dmem99_io_pipeline_valid),
    .io_pipeline_writedata(dmem99_io_pipeline_writedata),
    .io_pipeline_memread(dmem99_io_pipeline_memread),
    .io_pipeline_memwrite(dmem99_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem99_io_pipeline_maskmode),
    .io_pipeline_sext(dmem99_io_pipeline_sext),
    .io_pipeline_readdata(dmem99_io_pipeline_readdata),
    .io_bus_request_valid(dmem99_io_bus_request_valid),
    .io_bus_request_bits_address(dmem99_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem99_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem99_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem99_io_bus_response_valid),
    .io_bus_response_bits_data(dmem99_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu100 ( // @[top.scala 712:22]
    .clock(cpu100_clock),
    .reset(cpu100_reset),
    .io_imem_address(cpu100_io_imem_address),
    .io_imem_instruction(cpu100_io_imem_instruction),
    .io_dmem_address(cpu100_io_dmem_address),
    .io_dmem_valid(cpu100_io_dmem_valid),
    .io_dmem_writedata(cpu100_io_dmem_writedata),
    .io_dmem_memread(cpu100_io_dmem_memread),
    .io_dmem_memwrite(cpu100_io_dmem_memwrite),
    .io_dmem_maskmode(cpu100_io_dmem_maskmode),
    .io_dmem_sext(cpu100_io_dmem_sext),
    .io_dmem_readdata(cpu100_io_dmem_readdata)
  );
  DualPortedCombinMemory mem100 ( // @[top.scala 713:22]
    .clock(mem100_clock),
    .reset(mem100_reset),
    .io_imem_request_bits_address(mem100_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem100_io_imem_response_bits_data),
    .io_dmem_request_valid(mem100_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem100_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem100_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem100_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem100_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem100_io_dmem_response_bits_data)
  );
  ICombinMemPort imem100 ( // @[top.scala 714:23]
    .io_pipeline_address(imem100_io_pipeline_address),
    .io_pipeline_instruction(imem100_io_pipeline_instruction),
    .io_bus_request_bits_address(imem100_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem100_io_bus_response_bits_data)
  );
  DCombinMemPort dmem100 ( // @[top.scala 715:23]
    .clock(dmem100_clock),
    .reset(dmem100_reset),
    .io_pipeline_address(dmem100_io_pipeline_address),
    .io_pipeline_valid(dmem100_io_pipeline_valid),
    .io_pipeline_writedata(dmem100_io_pipeline_writedata),
    .io_pipeline_memread(dmem100_io_pipeline_memread),
    .io_pipeline_memwrite(dmem100_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem100_io_pipeline_maskmode),
    .io_pipeline_sext(dmem100_io_pipeline_sext),
    .io_pipeline_readdata(dmem100_io_pipeline_readdata),
    .io_bus_request_valid(dmem100_io_bus_request_valid),
    .io_bus_request_bits_address(dmem100_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem100_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem100_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem100_io_bus_response_valid),
    .io_bus_response_bits_data(dmem100_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu101 ( // @[top.scala 719:22]
    .clock(cpu101_clock),
    .reset(cpu101_reset),
    .io_imem_address(cpu101_io_imem_address),
    .io_imem_instruction(cpu101_io_imem_instruction),
    .io_dmem_address(cpu101_io_dmem_address),
    .io_dmem_valid(cpu101_io_dmem_valid),
    .io_dmem_writedata(cpu101_io_dmem_writedata),
    .io_dmem_memread(cpu101_io_dmem_memread),
    .io_dmem_memwrite(cpu101_io_dmem_memwrite),
    .io_dmem_maskmode(cpu101_io_dmem_maskmode),
    .io_dmem_sext(cpu101_io_dmem_sext),
    .io_dmem_readdata(cpu101_io_dmem_readdata)
  );
  DualPortedCombinMemory mem101 ( // @[top.scala 720:22]
    .clock(mem101_clock),
    .reset(mem101_reset),
    .io_imem_request_bits_address(mem101_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem101_io_imem_response_bits_data),
    .io_dmem_request_valid(mem101_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem101_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem101_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem101_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem101_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem101_io_dmem_response_bits_data)
  );
  ICombinMemPort imem101 ( // @[top.scala 721:23]
    .io_pipeline_address(imem101_io_pipeline_address),
    .io_pipeline_instruction(imem101_io_pipeline_instruction),
    .io_bus_request_bits_address(imem101_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem101_io_bus_response_bits_data)
  );
  DCombinMemPort dmem101 ( // @[top.scala 722:23]
    .clock(dmem101_clock),
    .reset(dmem101_reset),
    .io_pipeline_address(dmem101_io_pipeline_address),
    .io_pipeline_valid(dmem101_io_pipeline_valid),
    .io_pipeline_writedata(dmem101_io_pipeline_writedata),
    .io_pipeline_memread(dmem101_io_pipeline_memread),
    .io_pipeline_memwrite(dmem101_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem101_io_pipeline_maskmode),
    .io_pipeline_sext(dmem101_io_pipeline_sext),
    .io_pipeline_readdata(dmem101_io_pipeline_readdata),
    .io_bus_request_valid(dmem101_io_bus_request_valid),
    .io_bus_request_bits_address(dmem101_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem101_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem101_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem101_io_bus_response_valid),
    .io_bus_response_bits_data(dmem101_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu102 ( // @[top.scala 726:22]
    .clock(cpu102_clock),
    .reset(cpu102_reset),
    .io_imem_address(cpu102_io_imem_address),
    .io_imem_instruction(cpu102_io_imem_instruction),
    .io_dmem_address(cpu102_io_dmem_address),
    .io_dmem_valid(cpu102_io_dmem_valid),
    .io_dmem_writedata(cpu102_io_dmem_writedata),
    .io_dmem_memread(cpu102_io_dmem_memread),
    .io_dmem_memwrite(cpu102_io_dmem_memwrite),
    .io_dmem_maskmode(cpu102_io_dmem_maskmode),
    .io_dmem_sext(cpu102_io_dmem_sext),
    .io_dmem_readdata(cpu102_io_dmem_readdata)
  );
  DualPortedCombinMemory mem102 ( // @[top.scala 727:22]
    .clock(mem102_clock),
    .reset(mem102_reset),
    .io_imem_request_bits_address(mem102_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem102_io_imem_response_bits_data),
    .io_dmem_request_valid(mem102_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem102_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem102_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem102_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem102_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem102_io_dmem_response_bits_data)
  );
  ICombinMemPort imem102 ( // @[top.scala 728:23]
    .io_pipeline_address(imem102_io_pipeline_address),
    .io_pipeline_instruction(imem102_io_pipeline_instruction),
    .io_bus_request_bits_address(imem102_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem102_io_bus_response_bits_data)
  );
  DCombinMemPort dmem102 ( // @[top.scala 729:23]
    .clock(dmem102_clock),
    .reset(dmem102_reset),
    .io_pipeline_address(dmem102_io_pipeline_address),
    .io_pipeline_valid(dmem102_io_pipeline_valid),
    .io_pipeline_writedata(dmem102_io_pipeline_writedata),
    .io_pipeline_memread(dmem102_io_pipeline_memread),
    .io_pipeline_memwrite(dmem102_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem102_io_pipeline_maskmode),
    .io_pipeline_sext(dmem102_io_pipeline_sext),
    .io_pipeline_readdata(dmem102_io_pipeline_readdata),
    .io_bus_request_valid(dmem102_io_bus_request_valid),
    .io_bus_request_bits_address(dmem102_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem102_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem102_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem102_io_bus_response_valid),
    .io_bus_response_bits_data(dmem102_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu103 ( // @[top.scala 733:22]
    .clock(cpu103_clock),
    .reset(cpu103_reset),
    .io_imem_address(cpu103_io_imem_address),
    .io_imem_instruction(cpu103_io_imem_instruction),
    .io_dmem_address(cpu103_io_dmem_address),
    .io_dmem_valid(cpu103_io_dmem_valid),
    .io_dmem_writedata(cpu103_io_dmem_writedata),
    .io_dmem_memread(cpu103_io_dmem_memread),
    .io_dmem_memwrite(cpu103_io_dmem_memwrite),
    .io_dmem_maskmode(cpu103_io_dmem_maskmode),
    .io_dmem_sext(cpu103_io_dmem_sext),
    .io_dmem_readdata(cpu103_io_dmem_readdata)
  );
  DualPortedCombinMemory mem103 ( // @[top.scala 734:22]
    .clock(mem103_clock),
    .reset(mem103_reset),
    .io_imem_request_bits_address(mem103_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem103_io_imem_response_bits_data),
    .io_dmem_request_valid(mem103_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem103_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem103_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem103_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem103_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem103_io_dmem_response_bits_data)
  );
  ICombinMemPort imem103 ( // @[top.scala 735:23]
    .io_pipeline_address(imem103_io_pipeline_address),
    .io_pipeline_instruction(imem103_io_pipeline_instruction),
    .io_bus_request_bits_address(imem103_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem103_io_bus_response_bits_data)
  );
  DCombinMemPort dmem103 ( // @[top.scala 736:23]
    .clock(dmem103_clock),
    .reset(dmem103_reset),
    .io_pipeline_address(dmem103_io_pipeline_address),
    .io_pipeline_valid(dmem103_io_pipeline_valid),
    .io_pipeline_writedata(dmem103_io_pipeline_writedata),
    .io_pipeline_memread(dmem103_io_pipeline_memread),
    .io_pipeline_memwrite(dmem103_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem103_io_pipeline_maskmode),
    .io_pipeline_sext(dmem103_io_pipeline_sext),
    .io_pipeline_readdata(dmem103_io_pipeline_readdata),
    .io_bus_request_valid(dmem103_io_bus_request_valid),
    .io_bus_request_bits_address(dmem103_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem103_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem103_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem103_io_bus_response_valid),
    .io_bus_response_bits_data(dmem103_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu104 ( // @[top.scala 740:22]
    .clock(cpu104_clock),
    .reset(cpu104_reset),
    .io_imem_address(cpu104_io_imem_address),
    .io_imem_instruction(cpu104_io_imem_instruction),
    .io_dmem_address(cpu104_io_dmem_address),
    .io_dmem_valid(cpu104_io_dmem_valid),
    .io_dmem_writedata(cpu104_io_dmem_writedata),
    .io_dmem_memread(cpu104_io_dmem_memread),
    .io_dmem_memwrite(cpu104_io_dmem_memwrite),
    .io_dmem_maskmode(cpu104_io_dmem_maskmode),
    .io_dmem_sext(cpu104_io_dmem_sext),
    .io_dmem_readdata(cpu104_io_dmem_readdata)
  );
  DualPortedCombinMemory mem104 ( // @[top.scala 741:22]
    .clock(mem104_clock),
    .reset(mem104_reset),
    .io_imem_request_bits_address(mem104_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem104_io_imem_response_bits_data),
    .io_dmem_request_valid(mem104_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem104_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem104_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem104_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem104_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem104_io_dmem_response_bits_data)
  );
  ICombinMemPort imem104 ( // @[top.scala 742:23]
    .io_pipeline_address(imem104_io_pipeline_address),
    .io_pipeline_instruction(imem104_io_pipeline_instruction),
    .io_bus_request_bits_address(imem104_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem104_io_bus_response_bits_data)
  );
  DCombinMemPort dmem104 ( // @[top.scala 743:23]
    .clock(dmem104_clock),
    .reset(dmem104_reset),
    .io_pipeline_address(dmem104_io_pipeline_address),
    .io_pipeline_valid(dmem104_io_pipeline_valid),
    .io_pipeline_writedata(dmem104_io_pipeline_writedata),
    .io_pipeline_memread(dmem104_io_pipeline_memread),
    .io_pipeline_memwrite(dmem104_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem104_io_pipeline_maskmode),
    .io_pipeline_sext(dmem104_io_pipeline_sext),
    .io_pipeline_readdata(dmem104_io_pipeline_readdata),
    .io_bus_request_valid(dmem104_io_bus_request_valid),
    .io_bus_request_bits_address(dmem104_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem104_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem104_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem104_io_bus_response_valid),
    .io_bus_response_bits_data(dmem104_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu105 ( // @[top.scala 747:22]
    .clock(cpu105_clock),
    .reset(cpu105_reset),
    .io_imem_address(cpu105_io_imem_address),
    .io_imem_instruction(cpu105_io_imem_instruction),
    .io_dmem_address(cpu105_io_dmem_address),
    .io_dmem_valid(cpu105_io_dmem_valid),
    .io_dmem_writedata(cpu105_io_dmem_writedata),
    .io_dmem_memread(cpu105_io_dmem_memread),
    .io_dmem_memwrite(cpu105_io_dmem_memwrite),
    .io_dmem_maskmode(cpu105_io_dmem_maskmode),
    .io_dmem_sext(cpu105_io_dmem_sext),
    .io_dmem_readdata(cpu105_io_dmem_readdata)
  );
  DualPortedCombinMemory mem105 ( // @[top.scala 748:22]
    .clock(mem105_clock),
    .reset(mem105_reset),
    .io_imem_request_bits_address(mem105_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem105_io_imem_response_bits_data),
    .io_dmem_request_valid(mem105_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem105_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem105_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem105_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem105_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem105_io_dmem_response_bits_data)
  );
  ICombinMemPort imem105 ( // @[top.scala 749:23]
    .io_pipeline_address(imem105_io_pipeline_address),
    .io_pipeline_instruction(imem105_io_pipeline_instruction),
    .io_bus_request_bits_address(imem105_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem105_io_bus_response_bits_data)
  );
  DCombinMemPort dmem105 ( // @[top.scala 750:23]
    .clock(dmem105_clock),
    .reset(dmem105_reset),
    .io_pipeline_address(dmem105_io_pipeline_address),
    .io_pipeline_valid(dmem105_io_pipeline_valid),
    .io_pipeline_writedata(dmem105_io_pipeline_writedata),
    .io_pipeline_memread(dmem105_io_pipeline_memread),
    .io_pipeline_memwrite(dmem105_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem105_io_pipeline_maskmode),
    .io_pipeline_sext(dmem105_io_pipeline_sext),
    .io_pipeline_readdata(dmem105_io_pipeline_readdata),
    .io_bus_request_valid(dmem105_io_bus_request_valid),
    .io_bus_request_bits_address(dmem105_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem105_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem105_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem105_io_bus_response_valid),
    .io_bus_response_bits_data(dmem105_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu106 ( // @[top.scala 754:22]
    .clock(cpu106_clock),
    .reset(cpu106_reset),
    .io_imem_address(cpu106_io_imem_address),
    .io_imem_instruction(cpu106_io_imem_instruction),
    .io_dmem_address(cpu106_io_dmem_address),
    .io_dmem_valid(cpu106_io_dmem_valid),
    .io_dmem_writedata(cpu106_io_dmem_writedata),
    .io_dmem_memread(cpu106_io_dmem_memread),
    .io_dmem_memwrite(cpu106_io_dmem_memwrite),
    .io_dmem_maskmode(cpu106_io_dmem_maskmode),
    .io_dmem_sext(cpu106_io_dmem_sext),
    .io_dmem_readdata(cpu106_io_dmem_readdata)
  );
  DualPortedCombinMemory mem106 ( // @[top.scala 755:22]
    .clock(mem106_clock),
    .reset(mem106_reset),
    .io_imem_request_bits_address(mem106_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem106_io_imem_response_bits_data),
    .io_dmem_request_valid(mem106_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem106_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem106_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem106_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem106_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem106_io_dmem_response_bits_data)
  );
  ICombinMemPort imem106 ( // @[top.scala 756:23]
    .io_pipeline_address(imem106_io_pipeline_address),
    .io_pipeline_instruction(imem106_io_pipeline_instruction),
    .io_bus_request_bits_address(imem106_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem106_io_bus_response_bits_data)
  );
  DCombinMemPort dmem106 ( // @[top.scala 757:23]
    .clock(dmem106_clock),
    .reset(dmem106_reset),
    .io_pipeline_address(dmem106_io_pipeline_address),
    .io_pipeline_valid(dmem106_io_pipeline_valid),
    .io_pipeline_writedata(dmem106_io_pipeline_writedata),
    .io_pipeline_memread(dmem106_io_pipeline_memread),
    .io_pipeline_memwrite(dmem106_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem106_io_pipeline_maskmode),
    .io_pipeline_sext(dmem106_io_pipeline_sext),
    .io_pipeline_readdata(dmem106_io_pipeline_readdata),
    .io_bus_request_valid(dmem106_io_bus_request_valid),
    .io_bus_request_bits_address(dmem106_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem106_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem106_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem106_io_bus_response_valid),
    .io_bus_response_bits_data(dmem106_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu107 ( // @[top.scala 761:22]
    .clock(cpu107_clock),
    .reset(cpu107_reset),
    .io_imem_address(cpu107_io_imem_address),
    .io_imem_instruction(cpu107_io_imem_instruction),
    .io_dmem_address(cpu107_io_dmem_address),
    .io_dmem_valid(cpu107_io_dmem_valid),
    .io_dmem_writedata(cpu107_io_dmem_writedata),
    .io_dmem_memread(cpu107_io_dmem_memread),
    .io_dmem_memwrite(cpu107_io_dmem_memwrite),
    .io_dmem_maskmode(cpu107_io_dmem_maskmode),
    .io_dmem_sext(cpu107_io_dmem_sext),
    .io_dmem_readdata(cpu107_io_dmem_readdata)
  );
  DualPortedCombinMemory mem107 ( // @[top.scala 762:22]
    .clock(mem107_clock),
    .reset(mem107_reset),
    .io_imem_request_bits_address(mem107_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem107_io_imem_response_bits_data),
    .io_dmem_request_valid(mem107_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem107_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem107_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem107_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem107_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem107_io_dmem_response_bits_data)
  );
  ICombinMemPort imem107 ( // @[top.scala 763:23]
    .io_pipeline_address(imem107_io_pipeline_address),
    .io_pipeline_instruction(imem107_io_pipeline_instruction),
    .io_bus_request_bits_address(imem107_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem107_io_bus_response_bits_data)
  );
  DCombinMemPort dmem107 ( // @[top.scala 764:23]
    .clock(dmem107_clock),
    .reset(dmem107_reset),
    .io_pipeline_address(dmem107_io_pipeline_address),
    .io_pipeline_valid(dmem107_io_pipeline_valid),
    .io_pipeline_writedata(dmem107_io_pipeline_writedata),
    .io_pipeline_memread(dmem107_io_pipeline_memread),
    .io_pipeline_memwrite(dmem107_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem107_io_pipeline_maskmode),
    .io_pipeline_sext(dmem107_io_pipeline_sext),
    .io_pipeline_readdata(dmem107_io_pipeline_readdata),
    .io_bus_request_valid(dmem107_io_bus_request_valid),
    .io_bus_request_bits_address(dmem107_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem107_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem107_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem107_io_bus_response_valid),
    .io_bus_response_bits_data(dmem107_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu108 ( // @[top.scala 768:22]
    .clock(cpu108_clock),
    .reset(cpu108_reset),
    .io_imem_address(cpu108_io_imem_address),
    .io_imem_instruction(cpu108_io_imem_instruction),
    .io_dmem_address(cpu108_io_dmem_address),
    .io_dmem_valid(cpu108_io_dmem_valid),
    .io_dmem_writedata(cpu108_io_dmem_writedata),
    .io_dmem_memread(cpu108_io_dmem_memread),
    .io_dmem_memwrite(cpu108_io_dmem_memwrite),
    .io_dmem_maskmode(cpu108_io_dmem_maskmode),
    .io_dmem_sext(cpu108_io_dmem_sext),
    .io_dmem_readdata(cpu108_io_dmem_readdata)
  );
  DualPortedCombinMemory mem108 ( // @[top.scala 769:22]
    .clock(mem108_clock),
    .reset(mem108_reset),
    .io_imem_request_bits_address(mem108_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem108_io_imem_response_bits_data),
    .io_dmem_request_valid(mem108_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem108_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem108_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem108_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem108_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem108_io_dmem_response_bits_data)
  );
  ICombinMemPort imem108 ( // @[top.scala 770:23]
    .io_pipeline_address(imem108_io_pipeline_address),
    .io_pipeline_instruction(imem108_io_pipeline_instruction),
    .io_bus_request_bits_address(imem108_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem108_io_bus_response_bits_data)
  );
  DCombinMemPort dmem108 ( // @[top.scala 771:23]
    .clock(dmem108_clock),
    .reset(dmem108_reset),
    .io_pipeline_address(dmem108_io_pipeline_address),
    .io_pipeline_valid(dmem108_io_pipeline_valid),
    .io_pipeline_writedata(dmem108_io_pipeline_writedata),
    .io_pipeline_memread(dmem108_io_pipeline_memread),
    .io_pipeline_memwrite(dmem108_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem108_io_pipeline_maskmode),
    .io_pipeline_sext(dmem108_io_pipeline_sext),
    .io_pipeline_readdata(dmem108_io_pipeline_readdata),
    .io_bus_request_valid(dmem108_io_bus_request_valid),
    .io_bus_request_bits_address(dmem108_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem108_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem108_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem108_io_bus_response_valid),
    .io_bus_response_bits_data(dmem108_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu109 ( // @[top.scala 775:22]
    .clock(cpu109_clock),
    .reset(cpu109_reset),
    .io_imem_address(cpu109_io_imem_address),
    .io_imem_instruction(cpu109_io_imem_instruction),
    .io_dmem_address(cpu109_io_dmem_address),
    .io_dmem_valid(cpu109_io_dmem_valid),
    .io_dmem_writedata(cpu109_io_dmem_writedata),
    .io_dmem_memread(cpu109_io_dmem_memread),
    .io_dmem_memwrite(cpu109_io_dmem_memwrite),
    .io_dmem_maskmode(cpu109_io_dmem_maskmode),
    .io_dmem_sext(cpu109_io_dmem_sext),
    .io_dmem_readdata(cpu109_io_dmem_readdata)
  );
  DualPortedCombinMemory mem109 ( // @[top.scala 776:22]
    .clock(mem109_clock),
    .reset(mem109_reset),
    .io_imem_request_bits_address(mem109_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem109_io_imem_response_bits_data),
    .io_dmem_request_valid(mem109_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem109_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem109_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem109_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem109_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem109_io_dmem_response_bits_data)
  );
  ICombinMemPort imem109 ( // @[top.scala 777:23]
    .io_pipeline_address(imem109_io_pipeline_address),
    .io_pipeline_instruction(imem109_io_pipeline_instruction),
    .io_bus_request_bits_address(imem109_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem109_io_bus_response_bits_data)
  );
  DCombinMemPort dmem109 ( // @[top.scala 778:23]
    .clock(dmem109_clock),
    .reset(dmem109_reset),
    .io_pipeline_address(dmem109_io_pipeline_address),
    .io_pipeline_valid(dmem109_io_pipeline_valid),
    .io_pipeline_writedata(dmem109_io_pipeline_writedata),
    .io_pipeline_memread(dmem109_io_pipeline_memread),
    .io_pipeline_memwrite(dmem109_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem109_io_pipeline_maskmode),
    .io_pipeline_sext(dmem109_io_pipeline_sext),
    .io_pipeline_readdata(dmem109_io_pipeline_readdata),
    .io_bus_request_valid(dmem109_io_bus_request_valid),
    .io_bus_request_bits_address(dmem109_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem109_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem109_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem109_io_bus_response_valid),
    .io_bus_response_bits_data(dmem109_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu110 ( // @[top.scala 782:22]
    .clock(cpu110_clock),
    .reset(cpu110_reset),
    .io_imem_address(cpu110_io_imem_address),
    .io_imem_instruction(cpu110_io_imem_instruction),
    .io_dmem_address(cpu110_io_dmem_address),
    .io_dmem_valid(cpu110_io_dmem_valid),
    .io_dmem_writedata(cpu110_io_dmem_writedata),
    .io_dmem_memread(cpu110_io_dmem_memread),
    .io_dmem_memwrite(cpu110_io_dmem_memwrite),
    .io_dmem_maskmode(cpu110_io_dmem_maskmode),
    .io_dmem_sext(cpu110_io_dmem_sext),
    .io_dmem_readdata(cpu110_io_dmem_readdata)
  );
  DualPortedCombinMemory mem110 ( // @[top.scala 783:22]
    .clock(mem110_clock),
    .reset(mem110_reset),
    .io_imem_request_bits_address(mem110_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem110_io_imem_response_bits_data),
    .io_dmem_request_valid(mem110_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem110_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem110_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem110_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem110_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem110_io_dmem_response_bits_data)
  );
  ICombinMemPort imem110 ( // @[top.scala 784:23]
    .io_pipeline_address(imem110_io_pipeline_address),
    .io_pipeline_instruction(imem110_io_pipeline_instruction),
    .io_bus_request_bits_address(imem110_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem110_io_bus_response_bits_data)
  );
  DCombinMemPort dmem110 ( // @[top.scala 785:23]
    .clock(dmem110_clock),
    .reset(dmem110_reset),
    .io_pipeline_address(dmem110_io_pipeline_address),
    .io_pipeline_valid(dmem110_io_pipeline_valid),
    .io_pipeline_writedata(dmem110_io_pipeline_writedata),
    .io_pipeline_memread(dmem110_io_pipeline_memread),
    .io_pipeline_memwrite(dmem110_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem110_io_pipeline_maskmode),
    .io_pipeline_sext(dmem110_io_pipeline_sext),
    .io_pipeline_readdata(dmem110_io_pipeline_readdata),
    .io_bus_request_valid(dmem110_io_bus_request_valid),
    .io_bus_request_bits_address(dmem110_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem110_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem110_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem110_io_bus_response_valid),
    .io_bus_response_bits_data(dmem110_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu111 ( // @[top.scala 789:22]
    .clock(cpu111_clock),
    .reset(cpu111_reset),
    .io_imem_address(cpu111_io_imem_address),
    .io_imem_instruction(cpu111_io_imem_instruction),
    .io_dmem_address(cpu111_io_dmem_address),
    .io_dmem_valid(cpu111_io_dmem_valid),
    .io_dmem_writedata(cpu111_io_dmem_writedata),
    .io_dmem_memread(cpu111_io_dmem_memread),
    .io_dmem_memwrite(cpu111_io_dmem_memwrite),
    .io_dmem_maskmode(cpu111_io_dmem_maskmode),
    .io_dmem_sext(cpu111_io_dmem_sext),
    .io_dmem_readdata(cpu111_io_dmem_readdata)
  );
  DualPortedCombinMemory mem111 ( // @[top.scala 790:22]
    .clock(mem111_clock),
    .reset(mem111_reset),
    .io_imem_request_bits_address(mem111_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem111_io_imem_response_bits_data),
    .io_dmem_request_valid(mem111_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem111_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem111_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem111_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem111_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem111_io_dmem_response_bits_data)
  );
  ICombinMemPort imem111 ( // @[top.scala 791:23]
    .io_pipeline_address(imem111_io_pipeline_address),
    .io_pipeline_instruction(imem111_io_pipeline_instruction),
    .io_bus_request_bits_address(imem111_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem111_io_bus_response_bits_data)
  );
  DCombinMemPort dmem111 ( // @[top.scala 792:23]
    .clock(dmem111_clock),
    .reset(dmem111_reset),
    .io_pipeline_address(dmem111_io_pipeline_address),
    .io_pipeline_valid(dmem111_io_pipeline_valid),
    .io_pipeline_writedata(dmem111_io_pipeline_writedata),
    .io_pipeline_memread(dmem111_io_pipeline_memread),
    .io_pipeline_memwrite(dmem111_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem111_io_pipeline_maskmode),
    .io_pipeline_sext(dmem111_io_pipeline_sext),
    .io_pipeline_readdata(dmem111_io_pipeline_readdata),
    .io_bus_request_valid(dmem111_io_bus_request_valid),
    .io_bus_request_bits_address(dmem111_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem111_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem111_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem111_io_bus_response_valid),
    .io_bus_response_bits_data(dmem111_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu112 ( // @[top.scala 796:22]
    .clock(cpu112_clock),
    .reset(cpu112_reset),
    .io_imem_address(cpu112_io_imem_address),
    .io_imem_instruction(cpu112_io_imem_instruction),
    .io_dmem_address(cpu112_io_dmem_address),
    .io_dmem_valid(cpu112_io_dmem_valid),
    .io_dmem_writedata(cpu112_io_dmem_writedata),
    .io_dmem_memread(cpu112_io_dmem_memread),
    .io_dmem_memwrite(cpu112_io_dmem_memwrite),
    .io_dmem_maskmode(cpu112_io_dmem_maskmode),
    .io_dmem_sext(cpu112_io_dmem_sext),
    .io_dmem_readdata(cpu112_io_dmem_readdata)
  );
  DualPortedCombinMemory mem112 ( // @[top.scala 797:22]
    .clock(mem112_clock),
    .reset(mem112_reset),
    .io_imem_request_bits_address(mem112_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem112_io_imem_response_bits_data),
    .io_dmem_request_valid(mem112_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem112_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem112_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem112_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem112_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem112_io_dmem_response_bits_data)
  );
  ICombinMemPort imem112 ( // @[top.scala 798:23]
    .io_pipeline_address(imem112_io_pipeline_address),
    .io_pipeline_instruction(imem112_io_pipeline_instruction),
    .io_bus_request_bits_address(imem112_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem112_io_bus_response_bits_data)
  );
  DCombinMemPort dmem112 ( // @[top.scala 799:23]
    .clock(dmem112_clock),
    .reset(dmem112_reset),
    .io_pipeline_address(dmem112_io_pipeline_address),
    .io_pipeline_valid(dmem112_io_pipeline_valid),
    .io_pipeline_writedata(dmem112_io_pipeline_writedata),
    .io_pipeline_memread(dmem112_io_pipeline_memread),
    .io_pipeline_memwrite(dmem112_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem112_io_pipeline_maskmode),
    .io_pipeline_sext(dmem112_io_pipeline_sext),
    .io_pipeline_readdata(dmem112_io_pipeline_readdata),
    .io_bus_request_valid(dmem112_io_bus_request_valid),
    .io_bus_request_bits_address(dmem112_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem112_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem112_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem112_io_bus_response_valid),
    .io_bus_response_bits_data(dmem112_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu113 ( // @[top.scala 803:22]
    .clock(cpu113_clock),
    .reset(cpu113_reset),
    .io_imem_address(cpu113_io_imem_address),
    .io_imem_instruction(cpu113_io_imem_instruction),
    .io_dmem_address(cpu113_io_dmem_address),
    .io_dmem_valid(cpu113_io_dmem_valid),
    .io_dmem_writedata(cpu113_io_dmem_writedata),
    .io_dmem_memread(cpu113_io_dmem_memread),
    .io_dmem_memwrite(cpu113_io_dmem_memwrite),
    .io_dmem_maskmode(cpu113_io_dmem_maskmode),
    .io_dmem_sext(cpu113_io_dmem_sext),
    .io_dmem_readdata(cpu113_io_dmem_readdata)
  );
  DualPortedCombinMemory mem113 ( // @[top.scala 804:22]
    .clock(mem113_clock),
    .reset(mem113_reset),
    .io_imem_request_bits_address(mem113_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem113_io_imem_response_bits_data),
    .io_dmem_request_valid(mem113_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem113_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem113_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem113_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem113_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem113_io_dmem_response_bits_data)
  );
  ICombinMemPort imem113 ( // @[top.scala 805:23]
    .io_pipeline_address(imem113_io_pipeline_address),
    .io_pipeline_instruction(imem113_io_pipeline_instruction),
    .io_bus_request_bits_address(imem113_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem113_io_bus_response_bits_data)
  );
  DCombinMemPort dmem113 ( // @[top.scala 806:23]
    .clock(dmem113_clock),
    .reset(dmem113_reset),
    .io_pipeline_address(dmem113_io_pipeline_address),
    .io_pipeline_valid(dmem113_io_pipeline_valid),
    .io_pipeline_writedata(dmem113_io_pipeline_writedata),
    .io_pipeline_memread(dmem113_io_pipeline_memread),
    .io_pipeline_memwrite(dmem113_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem113_io_pipeline_maskmode),
    .io_pipeline_sext(dmem113_io_pipeline_sext),
    .io_pipeline_readdata(dmem113_io_pipeline_readdata),
    .io_bus_request_valid(dmem113_io_bus_request_valid),
    .io_bus_request_bits_address(dmem113_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem113_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem113_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem113_io_bus_response_valid),
    .io_bus_response_bits_data(dmem113_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu114 ( // @[top.scala 810:22]
    .clock(cpu114_clock),
    .reset(cpu114_reset),
    .io_imem_address(cpu114_io_imem_address),
    .io_imem_instruction(cpu114_io_imem_instruction),
    .io_dmem_address(cpu114_io_dmem_address),
    .io_dmem_valid(cpu114_io_dmem_valid),
    .io_dmem_writedata(cpu114_io_dmem_writedata),
    .io_dmem_memread(cpu114_io_dmem_memread),
    .io_dmem_memwrite(cpu114_io_dmem_memwrite),
    .io_dmem_maskmode(cpu114_io_dmem_maskmode),
    .io_dmem_sext(cpu114_io_dmem_sext),
    .io_dmem_readdata(cpu114_io_dmem_readdata)
  );
  DualPortedCombinMemory mem114 ( // @[top.scala 811:22]
    .clock(mem114_clock),
    .reset(mem114_reset),
    .io_imem_request_bits_address(mem114_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem114_io_imem_response_bits_data),
    .io_dmem_request_valid(mem114_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem114_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem114_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem114_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem114_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem114_io_dmem_response_bits_data)
  );
  ICombinMemPort imem114 ( // @[top.scala 812:23]
    .io_pipeline_address(imem114_io_pipeline_address),
    .io_pipeline_instruction(imem114_io_pipeline_instruction),
    .io_bus_request_bits_address(imem114_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem114_io_bus_response_bits_data)
  );
  DCombinMemPort dmem114 ( // @[top.scala 813:23]
    .clock(dmem114_clock),
    .reset(dmem114_reset),
    .io_pipeline_address(dmem114_io_pipeline_address),
    .io_pipeline_valid(dmem114_io_pipeline_valid),
    .io_pipeline_writedata(dmem114_io_pipeline_writedata),
    .io_pipeline_memread(dmem114_io_pipeline_memread),
    .io_pipeline_memwrite(dmem114_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem114_io_pipeline_maskmode),
    .io_pipeline_sext(dmem114_io_pipeline_sext),
    .io_pipeline_readdata(dmem114_io_pipeline_readdata),
    .io_bus_request_valid(dmem114_io_bus_request_valid),
    .io_bus_request_bits_address(dmem114_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem114_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem114_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem114_io_bus_response_valid),
    .io_bus_response_bits_data(dmem114_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu115 ( // @[top.scala 817:22]
    .clock(cpu115_clock),
    .reset(cpu115_reset),
    .io_imem_address(cpu115_io_imem_address),
    .io_imem_instruction(cpu115_io_imem_instruction),
    .io_dmem_address(cpu115_io_dmem_address),
    .io_dmem_valid(cpu115_io_dmem_valid),
    .io_dmem_writedata(cpu115_io_dmem_writedata),
    .io_dmem_memread(cpu115_io_dmem_memread),
    .io_dmem_memwrite(cpu115_io_dmem_memwrite),
    .io_dmem_maskmode(cpu115_io_dmem_maskmode),
    .io_dmem_sext(cpu115_io_dmem_sext),
    .io_dmem_readdata(cpu115_io_dmem_readdata)
  );
  DualPortedCombinMemory mem115 ( // @[top.scala 818:22]
    .clock(mem115_clock),
    .reset(mem115_reset),
    .io_imem_request_bits_address(mem115_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem115_io_imem_response_bits_data),
    .io_dmem_request_valid(mem115_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem115_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem115_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem115_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem115_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem115_io_dmem_response_bits_data)
  );
  ICombinMemPort imem115 ( // @[top.scala 819:23]
    .io_pipeline_address(imem115_io_pipeline_address),
    .io_pipeline_instruction(imem115_io_pipeline_instruction),
    .io_bus_request_bits_address(imem115_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem115_io_bus_response_bits_data)
  );
  DCombinMemPort dmem115 ( // @[top.scala 820:23]
    .clock(dmem115_clock),
    .reset(dmem115_reset),
    .io_pipeline_address(dmem115_io_pipeline_address),
    .io_pipeline_valid(dmem115_io_pipeline_valid),
    .io_pipeline_writedata(dmem115_io_pipeline_writedata),
    .io_pipeline_memread(dmem115_io_pipeline_memread),
    .io_pipeline_memwrite(dmem115_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem115_io_pipeline_maskmode),
    .io_pipeline_sext(dmem115_io_pipeline_sext),
    .io_pipeline_readdata(dmem115_io_pipeline_readdata),
    .io_bus_request_valid(dmem115_io_bus_request_valid),
    .io_bus_request_bits_address(dmem115_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem115_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem115_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem115_io_bus_response_valid),
    .io_bus_response_bits_data(dmem115_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu116 ( // @[top.scala 824:22]
    .clock(cpu116_clock),
    .reset(cpu116_reset),
    .io_imem_address(cpu116_io_imem_address),
    .io_imem_instruction(cpu116_io_imem_instruction),
    .io_dmem_address(cpu116_io_dmem_address),
    .io_dmem_valid(cpu116_io_dmem_valid),
    .io_dmem_writedata(cpu116_io_dmem_writedata),
    .io_dmem_memread(cpu116_io_dmem_memread),
    .io_dmem_memwrite(cpu116_io_dmem_memwrite),
    .io_dmem_maskmode(cpu116_io_dmem_maskmode),
    .io_dmem_sext(cpu116_io_dmem_sext),
    .io_dmem_readdata(cpu116_io_dmem_readdata)
  );
  DualPortedCombinMemory mem116 ( // @[top.scala 825:22]
    .clock(mem116_clock),
    .reset(mem116_reset),
    .io_imem_request_bits_address(mem116_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem116_io_imem_response_bits_data),
    .io_dmem_request_valid(mem116_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem116_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem116_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem116_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem116_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem116_io_dmem_response_bits_data)
  );
  ICombinMemPort imem116 ( // @[top.scala 826:23]
    .io_pipeline_address(imem116_io_pipeline_address),
    .io_pipeline_instruction(imem116_io_pipeline_instruction),
    .io_bus_request_bits_address(imem116_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem116_io_bus_response_bits_data)
  );
  DCombinMemPort dmem116 ( // @[top.scala 827:23]
    .clock(dmem116_clock),
    .reset(dmem116_reset),
    .io_pipeline_address(dmem116_io_pipeline_address),
    .io_pipeline_valid(dmem116_io_pipeline_valid),
    .io_pipeline_writedata(dmem116_io_pipeline_writedata),
    .io_pipeline_memread(dmem116_io_pipeline_memread),
    .io_pipeline_memwrite(dmem116_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem116_io_pipeline_maskmode),
    .io_pipeline_sext(dmem116_io_pipeline_sext),
    .io_pipeline_readdata(dmem116_io_pipeline_readdata),
    .io_bus_request_valid(dmem116_io_bus_request_valid),
    .io_bus_request_bits_address(dmem116_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem116_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem116_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem116_io_bus_response_valid),
    .io_bus_response_bits_data(dmem116_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu117 ( // @[top.scala 831:22]
    .clock(cpu117_clock),
    .reset(cpu117_reset),
    .io_imem_address(cpu117_io_imem_address),
    .io_imem_instruction(cpu117_io_imem_instruction),
    .io_dmem_address(cpu117_io_dmem_address),
    .io_dmem_valid(cpu117_io_dmem_valid),
    .io_dmem_writedata(cpu117_io_dmem_writedata),
    .io_dmem_memread(cpu117_io_dmem_memread),
    .io_dmem_memwrite(cpu117_io_dmem_memwrite),
    .io_dmem_maskmode(cpu117_io_dmem_maskmode),
    .io_dmem_sext(cpu117_io_dmem_sext),
    .io_dmem_readdata(cpu117_io_dmem_readdata)
  );
  DualPortedCombinMemory mem117 ( // @[top.scala 832:22]
    .clock(mem117_clock),
    .reset(mem117_reset),
    .io_imem_request_bits_address(mem117_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem117_io_imem_response_bits_data),
    .io_dmem_request_valid(mem117_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem117_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem117_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem117_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem117_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem117_io_dmem_response_bits_data)
  );
  ICombinMemPort imem117 ( // @[top.scala 833:23]
    .io_pipeline_address(imem117_io_pipeline_address),
    .io_pipeline_instruction(imem117_io_pipeline_instruction),
    .io_bus_request_bits_address(imem117_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem117_io_bus_response_bits_data)
  );
  DCombinMemPort dmem117 ( // @[top.scala 834:23]
    .clock(dmem117_clock),
    .reset(dmem117_reset),
    .io_pipeline_address(dmem117_io_pipeline_address),
    .io_pipeline_valid(dmem117_io_pipeline_valid),
    .io_pipeline_writedata(dmem117_io_pipeline_writedata),
    .io_pipeline_memread(dmem117_io_pipeline_memread),
    .io_pipeline_memwrite(dmem117_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem117_io_pipeline_maskmode),
    .io_pipeline_sext(dmem117_io_pipeline_sext),
    .io_pipeline_readdata(dmem117_io_pipeline_readdata),
    .io_bus_request_valid(dmem117_io_bus_request_valid),
    .io_bus_request_bits_address(dmem117_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem117_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem117_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem117_io_bus_response_valid),
    .io_bus_response_bits_data(dmem117_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu118 ( // @[top.scala 838:22]
    .clock(cpu118_clock),
    .reset(cpu118_reset),
    .io_imem_address(cpu118_io_imem_address),
    .io_imem_instruction(cpu118_io_imem_instruction),
    .io_dmem_address(cpu118_io_dmem_address),
    .io_dmem_valid(cpu118_io_dmem_valid),
    .io_dmem_writedata(cpu118_io_dmem_writedata),
    .io_dmem_memread(cpu118_io_dmem_memread),
    .io_dmem_memwrite(cpu118_io_dmem_memwrite),
    .io_dmem_maskmode(cpu118_io_dmem_maskmode),
    .io_dmem_sext(cpu118_io_dmem_sext),
    .io_dmem_readdata(cpu118_io_dmem_readdata)
  );
  DualPortedCombinMemory mem118 ( // @[top.scala 839:22]
    .clock(mem118_clock),
    .reset(mem118_reset),
    .io_imem_request_bits_address(mem118_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem118_io_imem_response_bits_data),
    .io_dmem_request_valid(mem118_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem118_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem118_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem118_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem118_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem118_io_dmem_response_bits_data)
  );
  ICombinMemPort imem118 ( // @[top.scala 840:23]
    .io_pipeline_address(imem118_io_pipeline_address),
    .io_pipeline_instruction(imem118_io_pipeline_instruction),
    .io_bus_request_bits_address(imem118_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem118_io_bus_response_bits_data)
  );
  DCombinMemPort dmem118 ( // @[top.scala 841:23]
    .clock(dmem118_clock),
    .reset(dmem118_reset),
    .io_pipeline_address(dmem118_io_pipeline_address),
    .io_pipeline_valid(dmem118_io_pipeline_valid),
    .io_pipeline_writedata(dmem118_io_pipeline_writedata),
    .io_pipeline_memread(dmem118_io_pipeline_memread),
    .io_pipeline_memwrite(dmem118_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem118_io_pipeline_maskmode),
    .io_pipeline_sext(dmem118_io_pipeline_sext),
    .io_pipeline_readdata(dmem118_io_pipeline_readdata),
    .io_bus_request_valid(dmem118_io_bus_request_valid),
    .io_bus_request_bits_address(dmem118_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem118_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem118_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem118_io_bus_response_valid),
    .io_bus_response_bits_data(dmem118_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu119 ( // @[top.scala 845:22]
    .clock(cpu119_clock),
    .reset(cpu119_reset),
    .io_imem_address(cpu119_io_imem_address),
    .io_imem_instruction(cpu119_io_imem_instruction),
    .io_dmem_address(cpu119_io_dmem_address),
    .io_dmem_valid(cpu119_io_dmem_valid),
    .io_dmem_writedata(cpu119_io_dmem_writedata),
    .io_dmem_memread(cpu119_io_dmem_memread),
    .io_dmem_memwrite(cpu119_io_dmem_memwrite),
    .io_dmem_maskmode(cpu119_io_dmem_maskmode),
    .io_dmem_sext(cpu119_io_dmem_sext),
    .io_dmem_readdata(cpu119_io_dmem_readdata)
  );
  DualPortedCombinMemory mem119 ( // @[top.scala 846:22]
    .clock(mem119_clock),
    .reset(mem119_reset),
    .io_imem_request_bits_address(mem119_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem119_io_imem_response_bits_data),
    .io_dmem_request_valid(mem119_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem119_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem119_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem119_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem119_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem119_io_dmem_response_bits_data)
  );
  ICombinMemPort imem119 ( // @[top.scala 847:23]
    .io_pipeline_address(imem119_io_pipeline_address),
    .io_pipeline_instruction(imem119_io_pipeline_instruction),
    .io_bus_request_bits_address(imem119_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem119_io_bus_response_bits_data)
  );
  DCombinMemPort dmem119 ( // @[top.scala 848:23]
    .clock(dmem119_clock),
    .reset(dmem119_reset),
    .io_pipeline_address(dmem119_io_pipeline_address),
    .io_pipeline_valid(dmem119_io_pipeline_valid),
    .io_pipeline_writedata(dmem119_io_pipeline_writedata),
    .io_pipeline_memread(dmem119_io_pipeline_memread),
    .io_pipeline_memwrite(dmem119_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem119_io_pipeline_maskmode),
    .io_pipeline_sext(dmem119_io_pipeline_sext),
    .io_pipeline_readdata(dmem119_io_pipeline_readdata),
    .io_bus_request_valid(dmem119_io_bus_request_valid),
    .io_bus_request_bits_address(dmem119_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem119_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem119_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem119_io_bus_response_valid),
    .io_bus_response_bits_data(dmem119_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu120 ( // @[top.scala 852:22]
    .clock(cpu120_clock),
    .reset(cpu120_reset),
    .io_imem_address(cpu120_io_imem_address),
    .io_imem_instruction(cpu120_io_imem_instruction),
    .io_dmem_address(cpu120_io_dmem_address),
    .io_dmem_valid(cpu120_io_dmem_valid),
    .io_dmem_writedata(cpu120_io_dmem_writedata),
    .io_dmem_memread(cpu120_io_dmem_memread),
    .io_dmem_memwrite(cpu120_io_dmem_memwrite),
    .io_dmem_maskmode(cpu120_io_dmem_maskmode),
    .io_dmem_sext(cpu120_io_dmem_sext),
    .io_dmem_readdata(cpu120_io_dmem_readdata)
  );
  DualPortedCombinMemory mem120 ( // @[top.scala 853:22]
    .clock(mem120_clock),
    .reset(mem120_reset),
    .io_imem_request_bits_address(mem120_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem120_io_imem_response_bits_data),
    .io_dmem_request_valid(mem120_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem120_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem120_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem120_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem120_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem120_io_dmem_response_bits_data)
  );
  ICombinMemPort imem120 ( // @[top.scala 854:23]
    .io_pipeline_address(imem120_io_pipeline_address),
    .io_pipeline_instruction(imem120_io_pipeline_instruction),
    .io_bus_request_bits_address(imem120_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem120_io_bus_response_bits_data)
  );
  DCombinMemPort dmem120 ( // @[top.scala 855:23]
    .clock(dmem120_clock),
    .reset(dmem120_reset),
    .io_pipeline_address(dmem120_io_pipeline_address),
    .io_pipeline_valid(dmem120_io_pipeline_valid),
    .io_pipeline_writedata(dmem120_io_pipeline_writedata),
    .io_pipeline_memread(dmem120_io_pipeline_memread),
    .io_pipeline_memwrite(dmem120_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem120_io_pipeline_maskmode),
    .io_pipeline_sext(dmem120_io_pipeline_sext),
    .io_pipeline_readdata(dmem120_io_pipeline_readdata),
    .io_bus_request_valid(dmem120_io_bus_request_valid),
    .io_bus_request_bits_address(dmem120_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem120_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem120_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem120_io_bus_response_valid),
    .io_bus_response_bits_data(dmem120_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu121 ( // @[top.scala 859:22]
    .clock(cpu121_clock),
    .reset(cpu121_reset),
    .io_imem_address(cpu121_io_imem_address),
    .io_imem_instruction(cpu121_io_imem_instruction),
    .io_dmem_address(cpu121_io_dmem_address),
    .io_dmem_valid(cpu121_io_dmem_valid),
    .io_dmem_writedata(cpu121_io_dmem_writedata),
    .io_dmem_memread(cpu121_io_dmem_memread),
    .io_dmem_memwrite(cpu121_io_dmem_memwrite),
    .io_dmem_maskmode(cpu121_io_dmem_maskmode),
    .io_dmem_sext(cpu121_io_dmem_sext),
    .io_dmem_readdata(cpu121_io_dmem_readdata)
  );
  DualPortedCombinMemory mem121 ( // @[top.scala 860:22]
    .clock(mem121_clock),
    .reset(mem121_reset),
    .io_imem_request_bits_address(mem121_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem121_io_imem_response_bits_data),
    .io_dmem_request_valid(mem121_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem121_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem121_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem121_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem121_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem121_io_dmem_response_bits_data)
  );
  ICombinMemPort imem121 ( // @[top.scala 861:23]
    .io_pipeline_address(imem121_io_pipeline_address),
    .io_pipeline_instruction(imem121_io_pipeline_instruction),
    .io_bus_request_bits_address(imem121_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem121_io_bus_response_bits_data)
  );
  DCombinMemPort dmem121 ( // @[top.scala 862:23]
    .clock(dmem121_clock),
    .reset(dmem121_reset),
    .io_pipeline_address(dmem121_io_pipeline_address),
    .io_pipeline_valid(dmem121_io_pipeline_valid),
    .io_pipeline_writedata(dmem121_io_pipeline_writedata),
    .io_pipeline_memread(dmem121_io_pipeline_memread),
    .io_pipeline_memwrite(dmem121_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem121_io_pipeline_maskmode),
    .io_pipeline_sext(dmem121_io_pipeline_sext),
    .io_pipeline_readdata(dmem121_io_pipeline_readdata),
    .io_bus_request_valid(dmem121_io_bus_request_valid),
    .io_bus_request_bits_address(dmem121_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem121_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem121_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem121_io_bus_response_valid),
    .io_bus_response_bits_data(dmem121_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu122 ( // @[top.scala 866:22]
    .clock(cpu122_clock),
    .reset(cpu122_reset),
    .io_imem_address(cpu122_io_imem_address),
    .io_imem_instruction(cpu122_io_imem_instruction),
    .io_dmem_address(cpu122_io_dmem_address),
    .io_dmem_valid(cpu122_io_dmem_valid),
    .io_dmem_writedata(cpu122_io_dmem_writedata),
    .io_dmem_memread(cpu122_io_dmem_memread),
    .io_dmem_memwrite(cpu122_io_dmem_memwrite),
    .io_dmem_maskmode(cpu122_io_dmem_maskmode),
    .io_dmem_sext(cpu122_io_dmem_sext),
    .io_dmem_readdata(cpu122_io_dmem_readdata)
  );
  DualPortedCombinMemory mem122 ( // @[top.scala 867:22]
    .clock(mem122_clock),
    .reset(mem122_reset),
    .io_imem_request_bits_address(mem122_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem122_io_imem_response_bits_data),
    .io_dmem_request_valid(mem122_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem122_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem122_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem122_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem122_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem122_io_dmem_response_bits_data)
  );
  ICombinMemPort imem122 ( // @[top.scala 868:23]
    .io_pipeline_address(imem122_io_pipeline_address),
    .io_pipeline_instruction(imem122_io_pipeline_instruction),
    .io_bus_request_bits_address(imem122_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem122_io_bus_response_bits_data)
  );
  DCombinMemPort dmem122 ( // @[top.scala 869:23]
    .clock(dmem122_clock),
    .reset(dmem122_reset),
    .io_pipeline_address(dmem122_io_pipeline_address),
    .io_pipeline_valid(dmem122_io_pipeline_valid),
    .io_pipeline_writedata(dmem122_io_pipeline_writedata),
    .io_pipeline_memread(dmem122_io_pipeline_memread),
    .io_pipeline_memwrite(dmem122_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem122_io_pipeline_maskmode),
    .io_pipeline_sext(dmem122_io_pipeline_sext),
    .io_pipeline_readdata(dmem122_io_pipeline_readdata),
    .io_bus_request_valid(dmem122_io_bus_request_valid),
    .io_bus_request_bits_address(dmem122_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem122_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem122_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem122_io_bus_response_valid),
    .io_bus_response_bits_data(dmem122_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu123 ( // @[top.scala 873:22]
    .clock(cpu123_clock),
    .reset(cpu123_reset),
    .io_imem_address(cpu123_io_imem_address),
    .io_imem_instruction(cpu123_io_imem_instruction),
    .io_dmem_address(cpu123_io_dmem_address),
    .io_dmem_valid(cpu123_io_dmem_valid),
    .io_dmem_writedata(cpu123_io_dmem_writedata),
    .io_dmem_memread(cpu123_io_dmem_memread),
    .io_dmem_memwrite(cpu123_io_dmem_memwrite),
    .io_dmem_maskmode(cpu123_io_dmem_maskmode),
    .io_dmem_sext(cpu123_io_dmem_sext),
    .io_dmem_readdata(cpu123_io_dmem_readdata)
  );
  DualPortedCombinMemory mem123 ( // @[top.scala 874:22]
    .clock(mem123_clock),
    .reset(mem123_reset),
    .io_imem_request_bits_address(mem123_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem123_io_imem_response_bits_data),
    .io_dmem_request_valid(mem123_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem123_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem123_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem123_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem123_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem123_io_dmem_response_bits_data)
  );
  ICombinMemPort imem123 ( // @[top.scala 875:23]
    .io_pipeline_address(imem123_io_pipeline_address),
    .io_pipeline_instruction(imem123_io_pipeline_instruction),
    .io_bus_request_bits_address(imem123_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem123_io_bus_response_bits_data)
  );
  DCombinMemPort dmem123 ( // @[top.scala 876:23]
    .clock(dmem123_clock),
    .reset(dmem123_reset),
    .io_pipeline_address(dmem123_io_pipeline_address),
    .io_pipeline_valid(dmem123_io_pipeline_valid),
    .io_pipeline_writedata(dmem123_io_pipeline_writedata),
    .io_pipeline_memread(dmem123_io_pipeline_memread),
    .io_pipeline_memwrite(dmem123_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem123_io_pipeline_maskmode),
    .io_pipeline_sext(dmem123_io_pipeline_sext),
    .io_pipeline_readdata(dmem123_io_pipeline_readdata),
    .io_bus_request_valid(dmem123_io_bus_request_valid),
    .io_bus_request_bits_address(dmem123_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem123_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem123_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem123_io_bus_response_valid),
    .io_bus_response_bits_data(dmem123_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu124 ( // @[top.scala 880:22]
    .clock(cpu124_clock),
    .reset(cpu124_reset),
    .io_imem_address(cpu124_io_imem_address),
    .io_imem_instruction(cpu124_io_imem_instruction),
    .io_dmem_address(cpu124_io_dmem_address),
    .io_dmem_valid(cpu124_io_dmem_valid),
    .io_dmem_writedata(cpu124_io_dmem_writedata),
    .io_dmem_memread(cpu124_io_dmem_memread),
    .io_dmem_memwrite(cpu124_io_dmem_memwrite),
    .io_dmem_maskmode(cpu124_io_dmem_maskmode),
    .io_dmem_sext(cpu124_io_dmem_sext),
    .io_dmem_readdata(cpu124_io_dmem_readdata)
  );
  DualPortedCombinMemory mem124 ( // @[top.scala 881:22]
    .clock(mem124_clock),
    .reset(mem124_reset),
    .io_imem_request_bits_address(mem124_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem124_io_imem_response_bits_data),
    .io_dmem_request_valid(mem124_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem124_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem124_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem124_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem124_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem124_io_dmem_response_bits_data)
  );
  ICombinMemPort imem124 ( // @[top.scala 882:23]
    .io_pipeline_address(imem124_io_pipeline_address),
    .io_pipeline_instruction(imem124_io_pipeline_instruction),
    .io_bus_request_bits_address(imem124_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem124_io_bus_response_bits_data)
  );
  DCombinMemPort dmem124 ( // @[top.scala 883:23]
    .clock(dmem124_clock),
    .reset(dmem124_reset),
    .io_pipeline_address(dmem124_io_pipeline_address),
    .io_pipeline_valid(dmem124_io_pipeline_valid),
    .io_pipeline_writedata(dmem124_io_pipeline_writedata),
    .io_pipeline_memread(dmem124_io_pipeline_memread),
    .io_pipeline_memwrite(dmem124_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem124_io_pipeline_maskmode),
    .io_pipeline_sext(dmem124_io_pipeline_sext),
    .io_pipeline_readdata(dmem124_io_pipeline_readdata),
    .io_bus_request_valid(dmem124_io_bus_request_valid),
    .io_bus_request_bits_address(dmem124_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem124_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem124_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem124_io_bus_response_valid),
    .io_bus_response_bits_data(dmem124_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu125 ( // @[top.scala 887:22]
    .clock(cpu125_clock),
    .reset(cpu125_reset),
    .io_imem_address(cpu125_io_imem_address),
    .io_imem_instruction(cpu125_io_imem_instruction),
    .io_dmem_address(cpu125_io_dmem_address),
    .io_dmem_valid(cpu125_io_dmem_valid),
    .io_dmem_writedata(cpu125_io_dmem_writedata),
    .io_dmem_memread(cpu125_io_dmem_memread),
    .io_dmem_memwrite(cpu125_io_dmem_memwrite),
    .io_dmem_maskmode(cpu125_io_dmem_maskmode),
    .io_dmem_sext(cpu125_io_dmem_sext),
    .io_dmem_readdata(cpu125_io_dmem_readdata)
  );
  DualPortedCombinMemory mem125 ( // @[top.scala 888:22]
    .clock(mem125_clock),
    .reset(mem125_reset),
    .io_imem_request_bits_address(mem125_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem125_io_imem_response_bits_data),
    .io_dmem_request_valid(mem125_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem125_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem125_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem125_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem125_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem125_io_dmem_response_bits_data)
  );
  ICombinMemPort imem125 ( // @[top.scala 889:23]
    .io_pipeline_address(imem125_io_pipeline_address),
    .io_pipeline_instruction(imem125_io_pipeline_instruction),
    .io_bus_request_bits_address(imem125_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem125_io_bus_response_bits_data)
  );
  DCombinMemPort dmem125 ( // @[top.scala 890:23]
    .clock(dmem125_clock),
    .reset(dmem125_reset),
    .io_pipeline_address(dmem125_io_pipeline_address),
    .io_pipeline_valid(dmem125_io_pipeline_valid),
    .io_pipeline_writedata(dmem125_io_pipeline_writedata),
    .io_pipeline_memread(dmem125_io_pipeline_memread),
    .io_pipeline_memwrite(dmem125_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem125_io_pipeline_maskmode),
    .io_pipeline_sext(dmem125_io_pipeline_sext),
    .io_pipeline_readdata(dmem125_io_pipeline_readdata),
    .io_bus_request_valid(dmem125_io_bus_request_valid),
    .io_bus_request_bits_address(dmem125_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem125_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem125_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem125_io_bus_response_valid),
    .io_bus_response_bits_data(dmem125_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu126 ( // @[top.scala 894:22]
    .clock(cpu126_clock),
    .reset(cpu126_reset),
    .io_imem_address(cpu126_io_imem_address),
    .io_imem_instruction(cpu126_io_imem_instruction),
    .io_dmem_address(cpu126_io_dmem_address),
    .io_dmem_valid(cpu126_io_dmem_valid),
    .io_dmem_writedata(cpu126_io_dmem_writedata),
    .io_dmem_memread(cpu126_io_dmem_memread),
    .io_dmem_memwrite(cpu126_io_dmem_memwrite),
    .io_dmem_maskmode(cpu126_io_dmem_maskmode),
    .io_dmem_sext(cpu126_io_dmem_sext),
    .io_dmem_readdata(cpu126_io_dmem_readdata)
  );
  DualPortedCombinMemory mem126 ( // @[top.scala 895:22]
    .clock(mem126_clock),
    .reset(mem126_reset),
    .io_imem_request_bits_address(mem126_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem126_io_imem_response_bits_data),
    .io_dmem_request_valid(mem126_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem126_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem126_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem126_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem126_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem126_io_dmem_response_bits_data)
  );
  ICombinMemPort imem126 ( // @[top.scala 896:23]
    .io_pipeline_address(imem126_io_pipeline_address),
    .io_pipeline_instruction(imem126_io_pipeline_instruction),
    .io_bus_request_bits_address(imem126_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem126_io_bus_response_bits_data)
  );
  DCombinMemPort dmem126 ( // @[top.scala 897:23]
    .clock(dmem126_clock),
    .reset(dmem126_reset),
    .io_pipeline_address(dmem126_io_pipeline_address),
    .io_pipeline_valid(dmem126_io_pipeline_valid),
    .io_pipeline_writedata(dmem126_io_pipeline_writedata),
    .io_pipeline_memread(dmem126_io_pipeline_memread),
    .io_pipeline_memwrite(dmem126_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem126_io_pipeline_maskmode),
    .io_pipeline_sext(dmem126_io_pipeline_sext),
    .io_pipeline_readdata(dmem126_io_pipeline_readdata),
    .io_bus_request_valid(dmem126_io_bus_request_valid),
    .io_bus_request_bits_address(dmem126_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem126_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem126_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem126_io_bus_response_valid),
    .io_bus_response_bits_data(dmem126_io_bus_response_bits_data)
  );
  PipelinedCPUBP cpu127 ( // @[top.scala 901:22]
    .clock(cpu127_clock),
    .reset(cpu127_reset),
    .io_imem_address(cpu127_io_imem_address),
    .io_imem_instruction(cpu127_io_imem_instruction),
    .io_dmem_address(cpu127_io_dmem_address),
    .io_dmem_valid(cpu127_io_dmem_valid),
    .io_dmem_writedata(cpu127_io_dmem_writedata),
    .io_dmem_memread(cpu127_io_dmem_memread),
    .io_dmem_memwrite(cpu127_io_dmem_memwrite),
    .io_dmem_maskmode(cpu127_io_dmem_maskmode),
    .io_dmem_sext(cpu127_io_dmem_sext),
    .io_dmem_readdata(cpu127_io_dmem_readdata)
  );
  DualPortedCombinMemory mem127 ( // @[top.scala 902:22]
    .clock(mem127_clock),
    .reset(mem127_reset),
    .io_imem_request_bits_address(mem127_io_imem_request_bits_address),
    .io_imem_response_bits_data(mem127_io_imem_response_bits_data),
    .io_dmem_request_valid(mem127_io_dmem_request_valid),
    .io_dmem_request_bits_address(mem127_io_dmem_request_bits_address),
    .io_dmem_request_bits_writedata(mem127_io_dmem_request_bits_writedata),
    .io_dmem_request_bits_operation(mem127_io_dmem_request_bits_operation),
    .io_dmem_response_valid(mem127_io_dmem_response_valid),
    .io_dmem_response_bits_data(mem127_io_dmem_response_bits_data)
  );
  ICombinMemPort imem127 ( // @[top.scala 903:23]
    .io_pipeline_address(imem127_io_pipeline_address),
    .io_pipeline_instruction(imem127_io_pipeline_instruction),
    .io_bus_request_bits_address(imem127_io_bus_request_bits_address),
    .io_bus_response_bits_data(imem127_io_bus_response_bits_data)
  );
  DCombinMemPort dmem127 ( // @[top.scala 904:23]
    .clock(dmem127_clock),
    .reset(dmem127_reset),
    .io_pipeline_address(dmem127_io_pipeline_address),
    .io_pipeline_valid(dmem127_io_pipeline_valid),
    .io_pipeline_writedata(dmem127_io_pipeline_writedata),
    .io_pipeline_memread(dmem127_io_pipeline_memread),
    .io_pipeline_memwrite(dmem127_io_pipeline_memwrite),
    .io_pipeline_maskmode(dmem127_io_pipeline_maskmode),
    .io_pipeline_sext(dmem127_io_pipeline_sext),
    .io_pipeline_readdata(dmem127_io_pipeline_readdata),
    .io_bus_request_valid(dmem127_io_bus_request_valid),
    .io_bus_request_bits_address(dmem127_io_bus_request_bits_address),
    .io_bus_request_bits_writedata(dmem127_io_bus_request_bits_writedata),
    .io_bus_request_bits_operation(dmem127_io_bus_request_bits_operation),
    .io_bus_response_valid(dmem127_io_bus_response_valid),
    .io_bus_response_bits_data(dmem127_io_bus_response_bits_data)
  );
  assign io_success = 1'h0;
  assign cpu0_clock = clock;
  assign cpu0_reset = reset;
  assign cpu0_io_imem_instruction = imem0_io_pipeline_instruction; // @[top.scala 17:16]
  assign cpu0_io_dmem_readdata = dmem0_io_pipeline_readdata; // @[top.scala 18:16]
  assign mem0_clock = clock;
  assign mem0_reset = reset;
  assign mem0_io_imem_request_bits_address = imem0_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem0_io_dmem_request_valid = dmem0_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem0_io_dmem_request_bits_address = dmem0_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem0_io_dmem_request_bits_writedata = dmem0_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem0_io_dmem_request_bits_operation = dmem0_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem0_io_pipeline_address = cpu0_io_imem_address; // @[top.scala 17:16]
  assign imem0_io_bus_response_bits_data = mem0_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem0_clock = clock;
  assign dmem0_reset = reset;
  assign dmem0_io_pipeline_address = cpu0_io_dmem_address; // @[top.scala 18:16]
  assign dmem0_io_pipeline_valid = cpu0_io_dmem_valid; // @[top.scala 18:16]
  assign dmem0_io_pipeline_writedata = cpu0_io_dmem_writedata; // @[top.scala 18:16]
  assign dmem0_io_pipeline_memread = cpu0_io_dmem_memread; // @[top.scala 18:16]
  assign dmem0_io_pipeline_memwrite = cpu0_io_dmem_memwrite; // @[top.scala 18:16]
  assign dmem0_io_pipeline_maskmode = cpu0_io_dmem_maskmode; // @[top.scala 18:16]
  assign dmem0_io_pipeline_sext = cpu0_io_dmem_sext; // @[top.scala 18:16]
  assign dmem0_io_bus_response_valid = mem0_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem0_io_bus_response_bits_data = mem0_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu1_clock = clock;
  assign cpu1_reset = reset;
  assign cpu1_io_imem_instruction = imem1_io_pipeline_instruction; // @[top.scala 24:16]
  assign cpu1_io_dmem_readdata = dmem1_io_pipeline_readdata; // @[top.scala 25:16]
  assign mem1_clock = clock;
  assign mem1_reset = reset;
  assign mem1_io_imem_request_bits_address = imem1_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem1_io_dmem_request_valid = dmem1_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem1_io_dmem_request_bits_address = dmem1_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem1_io_dmem_request_bits_writedata = dmem1_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem1_io_dmem_request_bits_operation = dmem1_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem1_io_pipeline_address = cpu1_io_imem_address; // @[top.scala 24:16]
  assign imem1_io_bus_response_bits_data = mem1_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem1_clock = clock;
  assign dmem1_reset = reset;
  assign dmem1_io_pipeline_address = cpu1_io_dmem_address; // @[top.scala 25:16]
  assign dmem1_io_pipeline_valid = cpu1_io_dmem_valid; // @[top.scala 25:16]
  assign dmem1_io_pipeline_writedata = cpu1_io_dmem_writedata; // @[top.scala 25:16]
  assign dmem1_io_pipeline_memread = cpu1_io_dmem_memread; // @[top.scala 25:16]
  assign dmem1_io_pipeline_memwrite = cpu1_io_dmem_memwrite; // @[top.scala 25:16]
  assign dmem1_io_pipeline_maskmode = cpu1_io_dmem_maskmode; // @[top.scala 25:16]
  assign dmem1_io_pipeline_sext = cpu1_io_dmem_sext; // @[top.scala 25:16]
  assign dmem1_io_bus_response_valid = mem1_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem1_io_bus_response_bits_data = mem1_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu2_clock = clock;
  assign cpu2_reset = reset;
  assign cpu2_io_imem_instruction = imem2_io_pipeline_instruction; // @[top.scala 31:16]
  assign cpu2_io_dmem_readdata = dmem2_io_pipeline_readdata; // @[top.scala 32:16]
  assign mem2_clock = clock;
  assign mem2_reset = reset;
  assign mem2_io_imem_request_bits_address = imem2_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem2_io_dmem_request_valid = dmem2_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem2_io_dmem_request_bits_address = dmem2_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem2_io_dmem_request_bits_writedata = dmem2_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem2_io_dmem_request_bits_operation = dmem2_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem2_io_pipeline_address = cpu2_io_imem_address; // @[top.scala 31:16]
  assign imem2_io_bus_response_bits_data = mem2_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem2_clock = clock;
  assign dmem2_reset = reset;
  assign dmem2_io_pipeline_address = cpu2_io_dmem_address; // @[top.scala 32:16]
  assign dmem2_io_pipeline_valid = cpu2_io_dmem_valid; // @[top.scala 32:16]
  assign dmem2_io_pipeline_writedata = cpu2_io_dmem_writedata; // @[top.scala 32:16]
  assign dmem2_io_pipeline_memread = cpu2_io_dmem_memread; // @[top.scala 32:16]
  assign dmem2_io_pipeline_memwrite = cpu2_io_dmem_memwrite; // @[top.scala 32:16]
  assign dmem2_io_pipeline_maskmode = cpu2_io_dmem_maskmode; // @[top.scala 32:16]
  assign dmem2_io_pipeline_sext = cpu2_io_dmem_sext; // @[top.scala 32:16]
  assign dmem2_io_bus_response_valid = mem2_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem2_io_bus_response_bits_data = mem2_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu3_clock = clock;
  assign cpu3_reset = reset;
  assign cpu3_io_imem_instruction = imem3_io_pipeline_instruction; // @[top.scala 38:16]
  assign cpu3_io_dmem_readdata = dmem3_io_pipeline_readdata; // @[top.scala 39:16]
  assign mem3_clock = clock;
  assign mem3_reset = reset;
  assign mem3_io_imem_request_bits_address = imem3_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem3_io_dmem_request_valid = dmem3_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem3_io_dmem_request_bits_address = dmem3_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem3_io_dmem_request_bits_writedata = dmem3_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem3_io_dmem_request_bits_operation = dmem3_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem3_io_pipeline_address = cpu3_io_imem_address; // @[top.scala 38:16]
  assign imem3_io_bus_response_bits_data = mem3_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem3_clock = clock;
  assign dmem3_reset = reset;
  assign dmem3_io_pipeline_address = cpu3_io_dmem_address; // @[top.scala 39:16]
  assign dmem3_io_pipeline_valid = cpu3_io_dmem_valid; // @[top.scala 39:16]
  assign dmem3_io_pipeline_writedata = cpu3_io_dmem_writedata; // @[top.scala 39:16]
  assign dmem3_io_pipeline_memread = cpu3_io_dmem_memread; // @[top.scala 39:16]
  assign dmem3_io_pipeline_memwrite = cpu3_io_dmem_memwrite; // @[top.scala 39:16]
  assign dmem3_io_pipeline_maskmode = cpu3_io_dmem_maskmode; // @[top.scala 39:16]
  assign dmem3_io_pipeline_sext = cpu3_io_dmem_sext; // @[top.scala 39:16]
  assign dmem3_io_bus_response_valid = mem3_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem3_io_bus_response_bits_data = mem3_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu4_clock = clock;
  assign cpu4_reset = reset;
  assign cpu4_io_imem_instruction = imem4_io_pipeline_instruction; // @[top.scala 45:16]
  assign cpu4_io_dmem_readdata = dmem4_io_pipeline_readdata; // @[top.scala 46:16]
  assign mem4_clock = clock;
  assign mem4_reset = reset;
  assign mem4_io_imem_request_bits_address = imem4_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem4_io_dmem_request_valid = dmem4_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem4_io_dmem_request_bits_address = dmem4_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem4_io_dmem_request_bits_writedata = dmem4_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem4_io_dmem_request_bits_operation = dmem4_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem4_io_pipeline_address = cpu4_io_imem_address; // @[top.scala 45:16]
  assign imem4_io_bus_response_bits_data = mem4_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem4_clock = clock;
  assign dmem4_reset = reset;
  assign dmem4_io_pipeline_address = cpu4_io_dmem_address; // @[top.scala 46:16]
  assign dmem4_io_pipeline_valid = cpu4_io_dmem_valid; // @[top.scala 46:16]
  assign dmem4_io_pipeline_writedata = cpu4_io_dmem_writedata; // @[top.scala 46:16]
  assign dmem4_io_pipeline_memread = cpu4_io_dmem_memread; // @[top.scala 46:16]
  assign dmem4_io_pipeline_memwrite = cpu4_io_dmem_memwrite; // @[top.scala 46:16]
  assign dmem4_io_pipeline_maskmode = cpu4_io_dmem_maskmode; // @[top.scala 46:16]
  assign dmem4_io_pipeline_sext = cpu4_io_dmem_sext; // @[top.scala 46:16]
  assign dmem4_io_bus_response_valid = mem4_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem4_io_bus_response_bits_data = mem4_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu5_clock = clock;
  assign cpu5_reset = reset;
  assign cpu5_io_imem_instruction = imem5_io_pipeline_instruction; // @[top.scala 52:16]
  assign cpu5_io_dmem_readdata = dmem5_io_pipeline_readdata; // @[top.scala 53:16]
  assign mem5_clock = clock;
  assign mem5_reset = reset;
  assign mem5_io_imem_request_bits_address = imem5_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem5_io_dmem_request_valid = dmem5_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem5_io_dmem_request_bits_address = dmem5_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem5_io_dmem_request_bits_writedata = dmem5_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem5_io_dmem_request_bits_operation = dmem5_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem5_io_pipeline_address = cpu5_io_imem_address; // @[top.scala 52:16]
  assign imem5_io_bus_response_bits_data = mem5_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem5_clock = clock;
  assign dmem5_reset = reset;
  assign dmem5_io_pipeline_address = cpu5_io_dmem_address; // @[top.scala 53:16]
  assign dmem5_io_pipeline_valid = cpu5_io_dmem_valid; // @[top.scala 53:16]
  assign dmem5_io_pipeline_writedata = cpu5_io_dmem_writedata; // @[top.scala 53:16]
  assign dmem5_io_pipeline_memread = cpu5_io_dmem_memread; // @[top.scala 53:16]
  assign dmem5_io_pipeline_memwrite = cpu5_io_dmem_memwrite; // @[top.scala 53:16]
  assign dmem5_io_pipeline_maskmode = cpu5_io_dmem_maskmode; // @[top.scala 53:16]
  assign dmem5_io_pipeline_sext = cpu5_io_dmem_sext; // @[top.scala 53:16]
  assign dmem5_io_bus_response_valid = mem5_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem5_io_bus_response_bits_data = mem5_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu6_clock = clock;
  assign cpu6_reset = reset;
  assign cpu6_io_imem_instruction = imem6_io_pipeline_instruction; // @[top.scala 59:16]
  assign cpu6_io_dmem_readdata = dmem6_io_pipeline_readdata; // @[top.scala 60:16]
  assign mem6_clock = clock;
  assign mem6_reset = reset;
  assign mem6_io_imem_request_bits_address = imem6_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem6_io_dmem_request_valid = dmem6_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem6_io_dmem_request_bits_address = dmem6_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem6_io_dmem_request_bits_writedata = dmem6_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem6_io_dmem_request_bits_operation = dmem6_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem6_io_pipeline_address = cpu6_io_imem_address; // @[top.scala 59:16]
  assign imem6_io_bus_response_bits_data = mem6_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem6_clock = clock;
  assign dmem6_reset = reset;
  assign dmem6_io_pipeline_address = cpu6_io_dmem_address; // @[top.scala 60:16]
  assign dmem6_io_pipeline_valid = cpu6_io_dmem_valid; // @[top.scala 60:16]
  assign dmem6_io_pipeline_writedata = cpu6_io_dmem_writedata; // @[top.scala 60:16]
  assign dmem6_io_pipeline_memread = cpu6_io_dmem_memread; // @[top.scala 60:16]
  assign dmem6_io_pipeline_memwrite = cpu6_io_dmem_memwrite; // @[top.scala 60:16]
  assign dmem6_io_pipeline_maskmode = cpu6_io_dmem_maskmode; // @[top.scala 60:16]
  assign dmem6_io_pipeline_sext = cpu6_io_dmem_sext; // @[top.scala 60:16]
  assign dmem6_io_bus_response_valid = mem6_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem6_io_bus_response_bits_data = mem6_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu7_clock = clock;
  assign cpu7_reset = reset;
  assign cpu7_io_imem_instruction = imem7_io_pipeline_instruction; // @[top.scala 66:16]
  assign cpu7_io_dmem_readdata = dmem7_io_pipeline_readdata; // @[top.scala 67:16]
  assign mem7_clock = clock;
  assign mem7_reset = reset;
  assign mem7_io_imem_request_bits_address = imem7_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem7_io_dmem_request_valid = dmem7_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem7_io_dmem_request_bits_address = dmem7_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem7_io_dmem_request_bits_writedata = dmem7_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem7_io_dmem_request_bits_operation = dmem7_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem7_io_pipeline_address = cpu7_io_imem_address; // @[top.scala 66:16]
  assign imem7_io_bus_response_bits_data = mem7_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem7_clock = clock;
  assign dmem7_reset = reset;
  assign dmem7_io_pipeline_address = cpu7_io_dmem_address; // @[top.scala 67:16]
  assign dmem7_io_pipeline_valid = cpu7_io_dmem_valid; // @[top.scala 67:16]
  assign dmem7_io_pipeline_writedata = cpu7_io_dmem_writedata; // @[top.scala 67:16]
  assign dmem7_io_pipeline_memread = cpu7_io_dmem_memread; // @[top.scala 67:16]
  assign dmem7_io_pipeline_memwrite = cpu7_io_dmem_memwrite; // @[top.scala 67:16]
  assign dmem7_io_pipeline_maskmode = cpu7_io_dmem_maskmode; // @[top.scala 67:16]
  assign dmem7_io_pipeline_sext = cpu7_io_dmem_sext; // @[top.scala 67:16]
  assign dmem7_io_bus_response_valid = mem7_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem7_io_bus_response_bits_data = mem7_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu8_clock = clock;
  assign cpu8_reset = reset;
  assign cpu8_io_imem_instruction = imem8_io_pipeline_instruction; // @[top.scala 73:16]
  assign cpu8_io_dmem_readdata = dmem8_io_pipeline_readdata; // @[top.scala 74:16]
  assign mem8_clock = clock;
  assign mem8_reset = reset;
  assign mem8_io_imem_request_bits_address = imem8_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem8_io_dmem_request_valid = dmem8_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem8_io_dmem_request_bits_address = dmem8_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem8_io_dmem_request_bits_writedata = dmem8_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem8_io_dmem_request_bits_operation = dmem8_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem8_io_pipeline_address = cpu8_io_imem_address; // @[top.scala 73:16]
  assign imem8_io_bus_response_bits_data = mem8_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem8_clock = clock;
  assign dmem8_reset = reset;
  assign dmem8_io_pipeline_address = cpu8_io_dmem_address; // @[top.scala 74:16]
  assign dmem8_io_pipeline_valid = cpu8_io_dmem_valid; // @[top.scala 74:16]
  assign dmem8_io_pipeline_writedata = cpu8_io_dmem_writedata; // @[top.scala 74:16]
  assign dmem8_io_pipeline_memread = cpu8_io_dmem_memread; // @[top.scala 74:16]
  assign dmem8_io_pipeline_memwrite = cpu8_io_dmem_memwrite; // @[top.scala 74:16]
  assign dmem8_io_pipeline_maskmode = cpu8_io_dmem_maskmode; // @[top.scala 74:16]
  assign dmem8_io_pipeline_sext = cpu8_io_dmem_sext; // @[top.scala 74:16]
  assign dmem8_io_bus_response_valid = mem8_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem8_io_bus_response_bits_data = mem8_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu9_clock = clock;
  assign cpu9_reset = reset;
  assign cpu9_io_imem_instruction = imem9_io_pipeline_instruction; // @[top.scala 80:16]
  assign cpu9_io_dmem_readdata = dmem9_io_pipeline_readdata; // @[top.scala 81:16]
  assign mem9_clock = clock;
  assign mem9_reset = reset;
  assign mem9_io_imem_request_bits_address = imem9_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem9_io_dmem_request_valid = dmem9_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem9_io_dmem_request_bits_address = dmem9_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem9_io_dmem_request_bits_writedata = dmem9_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem9_io_dmem_request_bits_operation = dmem9_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem9_io_pipeline_address = cpu9_io_imem_address; // @[top.scala 80:16]
  assign imem9_io_bus_response_bits_data = mem9_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem9_clock = clock;
  assign dmem9_reset = reset;
  assign dmem9_io_pipeline_address = cpu9_io_dmem_address; // @[top.scala 81:16]
  assign dmem9_io_pipeline_valid = cpu9_io_dmem_valid; // @[top.scala 81:16]
  assign dmem9_io_pipeline_writedata = cpu9_io_dmem_writedata; // @[top.scala 81:16]
  assign dmem9_io_pipeline_memread = cpu9_io_dmem_memread; // @[top.scala 81:16]
  assign dmem9_io_pipeline_memwrite = cpu9_io_dmem_memwrite; // @[top.scala 81:16]
  assign dmem9_io_pipeline_maskmode = cpu9_io_dmem_maskmode; // @[top.scala 81:16]
  assign dmem9_io_pipeline_sext = cpu9_io_dmem_sext; // @[top.scala 81:16]
  assign dmem9_io_bus_response_valid = mem9_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem9_io_bus_response_bits_data = mem9_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu10_clock = clock;
  assign cpu10_reset = reset;
  assign cpu10_io_imem_instruction = imem10_io_pipeline_instruction; // @[top.scala 87:17]
  assign cpu10_io_dmem_readdata = dmem10_io_pipeline_readdata; // @[top.scala 88:17]
  assign mem10_clock = clock;
  assign mem10_reset = reset;
  assign mem10_io_imem_request_bits_address = imem10_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem10_io_dmem_request_valid = dmem10_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem10_io_dmem_request_bits_address = dmem10_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem10_io_dmem_request_bits_writedata = dmem10_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem10_io_dmem_request_bits_operation = dmem10_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem10_io_pipeline_address = cpu10_io_imem_address; // @[top.scala 87:17]
  assign imem10_io_bus_response_bits_data = mem10_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem10_clock = clock;
  assign dmem10_reset = reset;
  assign dmem10_io_pipeline_address = cpu10_io_dmem_address; // @[top.scala 88:17]
  assign dmem10_io_pipeline_valid = cpu10_io_dmem_valid; // @[top.scala 88:17]
  assign dmem10_io_pipeline_writedata = cpu10_io_dmem_writedata; // @[top.scala 88:17]
  assign dmem10_io_pipeline_memread = cpu10_io_dmem_memread; // @[top.scala 88:17]
  assign dmem10_io_pipeline_memwrite = cpu10_io_dmem_memwrite; // @[top.scala 88:17]
  assign dmem10_io_pipeline_maskmode = cpu10_io_dmem_maskmode; // @[top.scala 88:17]
  assign dmem10_io_pipeline_sext = cpu10_io_dmem_sext; // @[top.scala 88:17]
  assign dmem10_io_bus_response_valid = mem10_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem10_io_bus_response_bits_data = mem10_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu11_clock = clock;
  assign cpu11_reset = reset;
  assign cpu11_io_imem_instruction = imem11_io_pipeline_instruction; // @[top.scala 94:17]
  assign cpu11_io_dmem_readdata = dmem11_io_pipeline_readdata; // @[top.scala 95:17]
  assign mem11_clock = clock;
  assign mem11_reset = reset;
  assign mem11_io_imem_request_bits_address = imem11_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem11_io_dmem_request_valid = dmem11_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem11_io_dmem_request_bits_address = dmem11_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem11_io_dmem_request_bits_writedata = dmem11_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem11_io_dmem_request_bits_operation = dmem11_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem11_io_pipeline_address = cpu11_io_imem_address; // @[top.scala 94:17]
  assign imem11_io_bus_response_bits_data = mem11_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem11_clock = clock;
  assign dmem11_reset = reset;
  assign dmem11_io_pipeline_address = cpu11_io_dmem_address; // @[top.scala 95:17]
  assign dmem11_io_pipeline_valid = cpu11_io_dmem_valid; // @[top.scala 95:17]
  assign dmem11_io_pipeline_writedata = cpu11_io_dmem_writedata; // @[top.scala 95:17]
  assign dmem11_io_pipeline_memread = cpu11_io_dmem_memread; // @[top.scala 95:17]
  assign dmem11_io_pipeline_memwrite = cpu11_io_dmem_memwrite; // @[top.scala 95:17]
  assign dmem11_io_pipeline_maskmode = cpu11_io_dmem_maskmode; // @[top.scala 95:17]
  assign dmem11_io_pipeline_sext = cpu11_io_dmem_sext; // @[top.scala 95:17]
  assign dmem11_io_bus_response_valid = mem11_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem11_io_bus_response_bits_data = mem11_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu12_clock = clock;
  assign cpu12_reset = reset;
  assign cpu12_io_imem_instruction = imem12_io_pipeline_instruction; // @[top.scala 101:17]
  assign cpu12_io_dmem_readdata = dmem12_io_pipeline_readdata; // @[top.scala 102:17]
  assign mem12_clock = clock;
  assign mem12_reset = reset;
  assign mem12_io_imem_request_bits_address = imem12_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem12_io_dmem_request_valid = dmem12_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem12_io_dmem_request_bits_address = dmem12_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem12_io_dmem_request_bits_writedata = dmem12_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem12_io_dmem_request_bits_operation = dmem12_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem12_io_pipeline_address = cpu12_io_imem_address; // @[top.scala 101:17]
  assign imem12_io_bus_response_bits_data = mem12_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem12_clock = clock;
  assign dmem12_reset = reset;
  assign dmem12_io_pipeline_address = cpu12_io_dmem_address; // @[top.scala 102:17]
  assign dmem12_io_pipeline_valid = cpu12_io_dmem_valid; // @[top.scala 102:17]
  assign dmem12_io_pipeline_writedata = cpu12_io_dmem_writedata; // @[top.scala 102:17]
  assign dmem12_io_pipeline_memread = cpu12_io_dmem_memread; // @[top.scala 102:17]
  assign dmem12_io_pipeline_memwrite = cpu12_io_dmem_memwrite; // @[top.scala 102:17]
  assign dmem12_io_pipeline_maskmode = cpu12_io_dmem_maskmode; // @[top.scala 102:17]
  assign dmem12_io_pipeline_sext = cpu12_io_dmem_sext; // @[top.scala 102:17]
  assign dmem12_io_bus_response_valid = mem12_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem12_io_bus_response_bits_data = mem12_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu13_clock = clock;
  assign cpu13_reset = reset;
  assign cpu13_io_imem_instruction = imem13_io_pipeline_instruction; // @[top.scala 108:17]
  assign cpu13_io_dmem_readdata = dmem13_io_pipeline_readdata; // @[top.scala 109:17]
  assign mem13_clock = clock;
  assign mem13_reset = reset;
  assign mem13_io_imem_request_bits_address = imem13_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem13_io_dmem_request_valid = dmem13_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem13_io_dmem_request_bits_address = dmem13_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem13_io_dmem_request_bits_writedata = dmem13_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem13_io_dmem_request_bits_operation = dmem13_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem13_io_pipeline_address = cpu13_io_imem_address; // @[top.scala 108:17]
  assign imem13_io_bus_response_bits_data = mem13_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem13_clock = clock;
  assign dmem13_reset = reset;
  assign dmem13_io_pipeline_address = cpu13_io_dmem_address; // @[top.scala 109:17]
  assign dmem13_io_pipeline_valid = cpu13_io_dmem_valid; // @[top.scala 109:17]
  assign dmem13_io_pipeline_writedata = cpu13_io_dmem_writedata; // @[top.scala 109:17]
  assign dmem13_io_pipeline_memread = cpu13_io_dmem_memread; // @[top.scala 109:17]
  assign dmem13_io_pipeline_memwrite = cpu13_io_dmem_memwrite; // @[top.scala 109:17]
  assign dmem13_io_pipeline_maskmode = cpu13_io_dmem_maskmode; // @[top.scala 109:17]
  assign dmem13_io_pipeline_sext = cpu13_io_dmem_sext; // @[top.scala 109:17]
  assign dmem13_io_bus_response_valid = mem13_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem13_io_bus_response_bits_data = mem13_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu14_clock = clock;
  assign cpu14_reset = reset;
  assign cpu14_io_imem_instruction = imem14_io_pipeline_instruction; // @[top.scala 115:17]
  assign cpu14_io_dmem_readdata = dmem14_io_pipeline_readdata; // @[top.scala 116:17]
  assign mem14_clock = clock;
  assign mem14_reset = reset;
  assign mem14_io_imem_request_bits_address = imem14_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem14_io_dmem_request_valid = dmem14_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem14_io_dmem_request_bits_address = dmem14_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem14_io_dmem_request_bits_writedata = dmem14_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem14_io_dmem_request_bits_operation = dmem14_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem14_io_pipeline_address = cpu14_io_imem_address; // @[top.scala 115:17]
  assign imem14_io_bus_response_bits_data = mem14_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem14_clock = clock;
  assign dmem14_reset = reset;
  assign dmem14_io_pipeline_address = cpu14_io_dmem_address; // @[top.scala 116:17]
  assign dmem14_io_pipeline_valid = cpu14_io_dmem_valid; // @[top.scala 116:17]
  assign dmem14_io_pipeline_writedata = cpu14_io_dmem_writedata; // @[top.scala 116:17]
  assign dmem14_io_pipeline_memread = cpu14_io_dmem_memread; // @[top.scala 116:17]
  assign dmem14_io_pipeline_memwrite = cpu14_io_dmem_memwrite; // @[top.scala 116:17]
  assign dmem14_io_pipeline_maskmode = cpu14_io_dmem_maskmode; // @[top.scala 116:17]
  assign dmem14_io_pipeline_sext = cpu14_io_dmem_sext; // @[top.scala 116:17]
  assign dmem14_io_bus_response_valid = mem14_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem14_io_bus_response_bits_data = mem14_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu15_clock = clock;
  assign cpu15_reset = reset;
  assign cpu15_io_imem_instruction = imem15_io_pipeline_instruction; // @[top.scala 122:17]
  assign cpu15_io_dmem_readdata = dmem15_io_pipeline_readdata; // @[top.scala 123:17]
  assign mem15_clock = clock;
  assign mem15_reset = reset;
  assign mem15_io_imem_request_bits_address = imem15_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem15_io_dmem_request_valid = dmem15_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem15_io_dmem_request_bits_address = dmem15_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem15_io_dmem_request_bits_writedata = dmem15_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem15_io_dmem_request_bits_operation = dmem15_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem15_io_pipeline_address = cpu15_io_imem_address; // @[top.scala 122:17]
  assign imem15_io_bus_response_bits_data = mem15_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem15_clock = clock;
  assign dmem15_reset = reset;
  assign dmem15_io_pipeline_address = cpu15_io_dmem_address; // @[top.scala 123:17]
  assign dmem15_io_pipeline_valid = cpu15_io_dmem_valid; // @[top.scala 123:17]
  assign dmem15_io_pipeline_writedata = cpu15_io_dmem_writedata; // @[top.scala 123:17]
  assign dmem15_io_pipeline_memread = cpu15_io_dmem_memread; // @[top.scala 123:17]
  assign dmem15_io_pipeline_memwrite = cpu15_io_dmem_memwrite; // @[top.scala 123:17]
  assign dmem15_io_pipeline_maskmode = cpu15_io_dmem_maskmode; // @[top.scala 123:17]
  assign dmem15_io_pipeline_sext = cpu15_io_dmem_sext; // @[top.scala 123:17]
  assign dmem15_io_bus_response_valid = mem15_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem15_io_bus_response_bits_data = mem15_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu16_clock = clock;
  assign cpu16_reset = reset;
  assign cpu16_io_imem_instruction = imem16_io_pipeline_instruction; // @[top.scala 129:17]
  assign cpu16_io_dmem_readdata = dmem16_io_pipeline_readdata; // @[top.scala 130:17]
  assign mem16_clock = clock;
  assign mem16_reset = reset;
  assign mem16_io_imem_request_bits_address = imem16_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem16_io_dmem_request_valid = dmem16_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem16_io_dmem_request_bits_address = dmem16_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem16_io_dmem_request_bits_writedata = dmem16_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem16_io_dmem_request_bits_operation = dmem16_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem16_io_pipeline_address = cpu16_io_imem_address; // @[top.scala 129:17]
  assign imem16_io_bus_response_bits_data = mem16_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem16_clock = clock;
  assign dmem16_reset = reset;
  assign dmem16_io_pipeline_address = cpu16_io_dmem_address; // @[top.scala 130:17]
  assign dmem16_io_pipeline_valid = cpu16_io_dmem_valid; // @[top.scala 130:17]
  assign dmem16_io_pipeline_writedata = cpu16_io_dmem_writedata; // @[top.scala 130:17]
  assign dmem16_io_pipeline_memread = cpu16_io_dmem_memread; // @[top.scala 130:17]
  assign dmem16_io_pipeline_memwrite = cpu16_io_dmem_memwrite; // @[top.scala 130:17]
  assign dmem16_io_pipeline_maskmode = cpu16_io_dmem_maskmode; // @[top.scala 130:17]
  assign dmem16_io_pipeline_sext = cpu16_io_dmem_sext; // @[top.scala 130:17]
  assign dmem16_io_bus_response_valid = mem16_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem16_io_bus_response_bits_data = mem16_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu17_clock = clock;
  assign cpu17_reset = reset;
  assign cpu17_io_imem_instruction = imem17_io_pipeline_instruction; // @[top.scala 136:17]
  assign cpu17_io_dmem_readdata = dmem17_io_pipeline_readdata; // @[top.scala 137:17]
  assign mem17_clock = clock;
  assign mem17_reset = reset;
  assign mem17_io_imem_request_bits_address = imem17_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem17_io_dmem_request_valid = dmem17_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem17_io_dmem_request_bits_address = dmem17_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem17_io_dmem_request_bits_writedata = dmem17_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem17_io_dmem_request_bits_operation = dmem17_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem17_io_pipeline_address = cpu17_io_imem_address; // @[top.scala 136:17]
  assign imem17_io_bus_response_bits_data = mem17_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem17_clock = clock;
  assign dmem17_reset = reset;
  assign dmem17_io_pipeline_address = cpu17_io_dmem_address; // @[top.scala 137:17]
  assign dmem17_io_pipeline_valid = cpu17_io_dmem_valid; // @[top.scala 137:17]
  assign dmem17_io_pipeline_writedata = cpu17_io_dmem_writedata; // @[top.scala 137:17]
  assign dmem17_io_pipeline_memread = cpu17_io_dmem_memread; // @[top.scala 137:17]
  assign dmem17_io_pipeline_memwrite = cpu17_io_dmem_memwrite; // @[top.scala 137:17]
  assign dmem17_io_pipeline_maskmode = cpu17_io_dmem_maskmode; // @[top.scala 137:17]
  assign dmem17_io_pipeline_sext = cpu17_io_dmem_sext; // @[top.scala 137:17]
  assign dmem17_io_bus_response_valid = mem17_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem17_io_bus_response_bits_data = mem17_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu18_clock = clock;
  assign cpu18_reset = reset;
  assign cpu18_io_imem_instruction = imem18_io_pipeline_instruction; // @[top.scala 143:17]
  assign cpu18_io_dmem_readdata = dmem18_io_pipeline_readdata; // @[top.scala 144:17]
  assign mem18_clock = clock;
  assign mem18_reset = reset;
  assign mem18_io_imem_request_bits_address = imem18_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem18_io_dmem_request_valid = dmem18_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem18_io_dmem_request_bits_address = dmem18_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem18_io_dmem_request_bits_writedata = dmem18_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem18_io_dmem_request_bits_operation = dmem18_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem18_io_pipeline_address = cpu18_io_imem_address; // @[top.scala 143:17]
  assign imem18_io_bus_response_bits_data = mem18_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem18_clock = clock;
  assign dmem18_reset = reset;
  assign dmem18_io_pipeline_address = cpu18_io_dmem_address; // @[top.scala 144:17]
  assign dmem18_io_pipeline_valid = cpu18_io_dmem_valid; // @[top.scala 144:17]
  assign dmem18_io_pipeline_writedata = cpu18_io_dmem_writedata; // @[top.scala 144:17]
  assign dmem18_io_pipeline_memread = cpu18_io_dmem_memread; // @[top.scala 144:17]
  assign dmem18_io_pipeline_memwrite = cpu18_io_dmem_memwrite; // @[top.scala 144:17]
  assign dmem18_io_pipeline_maskmode = cpu18_io_dmem_maskmode; // @[top.scala 144:17]
  assign dmem18_io_pipeline_sext = cpu18_io_dmem_sext; // @[top.scala 144:17]
  assign dmem18_io_bus_response_valid = mem18_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem18_io_bus_response_bits_data = mem18_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu19_clock = clock;
  assign cpu19_reset = reset;
  assign cpu19_io_imem_instruction = imem19_io_pipeline_instruction; // @[top.scala 150:17]
  assign cpu19_io_dmem_readdata = dmem19_io_pipeline_readdata; // @[top.scala 151:17]
  assign mem19_clock = clock;
  assign mem19_reset = reset;
  assign mem19_io_imem_request_bits_address = imem19_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem19_io_dmem_request_valid = dmem19_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem19_io_dmem_request_bits_address = dmem19_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem19_io_dmem_request_bits_writedata = dmem19_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem19_io_dmem_request_bits_operation = dmem19_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem19_io_pipeline_address = cpu19_io_imem_address; // @[top.scala 150:17]
  assign imem19_io_bus_response_bits_data = mem19_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem19_clock = clock;
  assign dmem19_reset = reset;
  assign dmem19_io_pipeline_address = cpu19_io_dmem_address; // @[top.scala 151:17]
  assign dmem19_io_pipeline_valid = cpu19_io_dmem_valid; // @[top.scala 151:17]
  assign dmem19_io_pipeline_writedata = cpu19_io_dmem_writedata; // @[top.scala 151:17]
  assign dmem19_io_pipeline_memread = cpu19_io_dmem_memread; // @[top.scala 151:17]
  assign dmem19_io_pipeline_memwrite = cpu19_io_dmem_memwrite; // @[top.scala 151:17]
  assign dmem19_io_pipeline_maskmode = cpu19_io_dmem_maskmode; // @[top.scala 151:17]
  assign dmem19_io_pipeline_sext = cpu19_io_dmem_sext; // @[top.scala 151:17]
  assign dmem19_io_bus_response_valid = mem19_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem19_io_bus_response_bits_data = mem19_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu20_clock = clock;
  assign cpu20_reset = reset;
  assign cpu20_io_imem_instruction = imem20_io_pipeline_instruction; // @[top.scala 157:17]
  assign cpu20_io_dmem_readdata = dmem20_io_pipeline_readdata; // @[top.scala 158:17]
  assign mem20_clock = clock;
  assign mem20_reset = reset;
  assign mem20_io_imem_request_bits_address = imem20_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem20_io_dmem_request_valid = dmem20_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem20_io_dmem_request_bits_address = dmem20_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem20_io_dmem_request_bits_writedata = dmem20_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem20_io_dmem_request_bits_operation = dmem20_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem20_io_pipeline_address = cpu20_io_imem_address; // @[top.scala 157:17]
  assign imem20_io_bus_response_bits_data = mem20_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem20_clock = clock;
  assign dmem20_reset = reset;
  assign dmem20_io_pipeline_address = cpu20_io_dmem_address; // @[top.scala 158:17]
  assign dmem20_io_pipeline_valid = cpu20_io_dmem_valid; // @[top.scala 158:17]
  assign dmem20_io_pipeline_writedata = cpu20_io_dmem_writedata; // @[top.scala 158:17]
  assign dmem20_io_pipeline_memread = cpu20_io_dmem_memread; // @[top.scala 158:17]
  assign dmem20_io_pipeline_memwrite = cpu20_io_dmem_memwrite; // @[top.scala 158:17]
  assign dmem20_io_pipeline_maskmode = cpu20_io_dmem_maskmode; // @[top.scala 158:17]
  assign dmem20_io_pipeline_sext = cpu20_io_dmem_sext; // @[top.scala 158:17]
  assign dmem20_io_bus_response_valid = mem20_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem20_io_bus_response_bits_data = mem20_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu21_clock = clock;
  assign cpu21_reset = reset;
  assign cpu21_io_imem_instruction = imem21_io_pipeline_instruction; // @[top.scala 164:17]
  assign cpu21_io_dmem_readdata = dmem21_io_pipeline_readdata; // @[top.scala 165:17]
  assign mem21_clock = clock;
  assign mem21_reset = reset;
  assign mem21_io_imem_request_bits_address = imem21_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem21_io_dmem_request_valid = dmem21_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem21_io_dmem_request_bits_address = dmem21_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem21_io_dmem_request_bits_writedata = dmem21_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem21_io_dmem_request_bits_operation = dmem21_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem21_io_pipeline_address = cpu21_io_imem_address; // @[top.scala 164:17]
  assign imem21_io_bus_response_bits_data = mem21_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem21_clock = clock;
  assign dmem21_reset = reset;
  assign dmem21_io_pipeline_address = cpu21_io_dmem_address; // @[top.scala 165:17]
  assign dmem21_io_pipeline_valid = cpu21_io_dmem_valid; // @[top.scala 165:17]
  assign dmem21_io_pipeline_writedata = cpu21_io_dmem_writedata; // @[top.scala 165:17]
  assign dmem21_io_pipeline_memread = cpu21_io_dmem_memread; // @[top.scala 165:17]
  assign dmem21_io_pipeline_memwrite = cpu21_io_dmem_memwrite; // @[top.scala 165:17]
  assign dmem21_io_pipeline_maskmode = cpu21_io_dmem_maskmode; // @[top.scala 165:17]
  assign dmem21_io_pipeline_sext = cpu21_io_dmem_sext; // @[top.scala 165:17]
  assign dmem21_io_bus_response_valid = mem21_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem21_io_bus_response_bits_data = mem21_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu22_clock = clock;
  assign cpu22_reset = reset;
  assign cpu22_io_imem_instruction = imem22_io_pipeline_instruction; // @[top.scala 171:17]
  assign cpu22_io_dmem_readdata = dmem22_io_pipeline_readdata; // @[top.scala 172:17]
  assign mem22_clock = clock;
  assign mem22_reset = reset;
  assign mem22_io_imem_request_bits_address = imem22_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem22_io_dmem_request_valid = dmem22_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem22_io_dmem_request_bits_address = dmem22_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem22_io_dmem_request_bits_writedata = dmem22_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem22_io_dmem_request_bits_operation = dmem22_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem22_io_pipeline_address = cpu22_io_imem_address; // @[top.scala 171:17]
  assign imem22_io_bus_response_bits_data = mem22_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem22_clock = clock;
  assign dmem22_reset = reset;
  assign dmem22_io_pipeline_address = cpu22_io_dmem_address; // @[top.scala 172:17]
  assign dmem22_io_pipeline_valid = cpu22_io_dmem_valid; // @[top.scala 172:17]
  assign dmem22_io_pipeline_writedata = cpu22_io_dmem_writedata; // @[top.scala 172:17]
  assign dmem22_io_pipeline_memread = cpu22_io_dmem_memread; // @[top.scala 172:17]
  assign dmem22_io_pipeline_memwrite = cpu22_io_dmem_memwrite; // @[top.scala 172:17]
  assign dmem22_io_pipeline_maskmode = cpu22_io_dmem_maskmode; // @[top.scala 172:17]
  assign dmem22_io_pipeline_sext = cpu22_io_dmem_sext; // @[top.scala 172:17]
  assign dmem22_io_bus_response_valid = mem22_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem22_io_bus_response_bits_data = mem22_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu23_clock = clock;
  assign cpu23_reset = reset;
  assign cpu23_io_imem_instruction = imem23_io_pipeline_instruction; // @[top.scala 178:17]
  assign cpu23_io_dmem_readdata = dmem23_io_pipeline_readdata; // @[top.scala 179:17]
  assign mem23_clock = clock;
  assign mem23_reset = reset;
  assign mem23_io_imem_request_bits_address = imem23_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem23_io_dmem_request_valid = dmem23_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem23_io_dmem_request_bits_address = dmem23_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem23_io_dmem_request_bits_writedata = dmem23_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem23_io_dmem_request_bits_operation = dmem23_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem23_io_pipeline_address = cpu23_io_imem_address; // @[top.scala 178:17]
  assign imem23_io_bus_response_bits_data = mem23_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem23_clock = clock;
  assign dmem23_reset = reset;
  assign dmem23_io_pipeline_address = cpu23_io_dmem_address; // @[top.scala 179:17]
  assign dmem23_io_pipeline_valid = cpu23_io_dmem_valid; // @[top.scala 179:17]
  assign dmem23_io_pipeline_writedata = cpu23_io_dmem_writedata; // @[top.scala 179:17]
  assign dmem23_io_pipeline_memread = cpu23_io_dmem_memread; // @[top.scala 179:17]
  assign dmem23_io_pipeline_memwrite = cpu23_io_dmem_memwrite; // @[top.scala 179:17]
  assign dmem23_io_pipeline_maskmode = cpu23_io_dmem_maskmode; // @[top.scala 179:17]
  assign dmem23_io_pipeline_sext = cpu23_io_dmem_sext; // @[top.scala 179:17]
  assign dmem23_io_bus_response_valid = mem23_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem23_io_bus_response_bits_data = mem23_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu24_clock = clock;
  assign cpu24_reset = reset;
  assign cpu24_io_imem_instruction = imem24_io_pipeline_instruction; // @[top.scala 185:17]
  assign cpu24_io_dmem_readdata = dmem24_io_pipeline_readdata; // @[top.scala 186:17]
  assign mem24_clock = clock;
  assign mem24_reset = reset;
  assign mem24_io_imem_request_bits_address = imem24_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem24_io_dmem_request_valid = dmem24_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem24_io_dmem_request_bits_address = dmem24_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem24_io_dmem_request_bits_writedata = dmem24_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem24_io_dmem_request_bits_operation = dmem24_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem24_io_pipeline_address = cpu24_io_imem_address; // @[top.scala 185:17]
  assign imem24_io_bus_response_bits_data = mem24_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem24_clock = clock;
  assign dmem24_reset = reset;
  assign dmem24_io_pipeline_address = cpu24_io_dmem_address; // @[top.scala 186:17]
  assign dmem24_io_pipeline_valid = cpu24_io_dmem_valid; // @[top.scala 186:17]
  assign dmem24_io_pipeline_writedata = cpu24_io_dmem_writedata; // @[top.scala 186:17]
  assign dmem24_io_pipeline_memread = cpu24_io_dmem_memread; // @[top.scala 186:17]
  assign dmem24_io_pipeline_memwrite = cpu24_io_dmem_memwrite; // @[top.scala 186:17]
  assign dmem24_io_pipeline_maskmode = cpu24_io_dmem_maskmode; // @[top.scala 186:17]
  assign dmem24_io_pipeline_sext = cpu24_io_dmem_sext; // @[top.scala 186:17]
  assign dmem24_io_bus_response_valid = mem24_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem24_io_bus_response_bits_data = mem24_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu25_clock = clock;
  assign cpu25_reset = reset;
  assign cpu25_io_imem_instruction = imem25_io_pipeline_instruction; // @[top.scala 192:17]
  assign cpu25_io_dmem_readdata = dmem25_io_pipeline_readdata; // @[top.scala 193:17]
  assign mem25_clock = clock;
  assign mem25_reset = reset;
  assign mem25_io_imem_request_bits_address = imem25_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem25_io_dmem_request_valid = dmem25_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem25_io_dmem_request_bits_address = dmem25_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem25_io_dmem_request_bits_writedata = dmem25_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem25_io_dmem_request_bits_operation = dmem25_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem25_io_pipeline_address = cpu25_io_imem_address; // @[top.scala 192:17]
  assign imem25_io_bus_response_bits_data = mem25_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem25_clock = clock;
  assign dmem25_reset = reset;
  assign dmem25_io_pipeline_address = cpu25_io_dmem_address; // @[top.scala 193:17]
  assign dmem25_io_pipeline_valid = cpu25_io_dmem_valid; // @[top.scala 193:17]
  assign dmem25_io_pipeline_writedata = cpu25_io_dmem_writedata; // @[top.scala 193:17]
  assign dmem25_io_pipeline_memread = cpu25_io_dmem_memread; // @[top.scala 193:17]
  assign dmem25_io_pipeline_memwrite = cpu25_io_dmem_memwrite; // @[top.scala 193:17]
  assign dmem25_io_pipeline_maskmode = cpu25_io_dmem_maskmode; // @[top.scala 193:17]
  assign dmem25_io_pipeline_sext = cpu25_io_dmem_sext; // @[top.scala 193:17]
  assign dmem25_io_bus_response_valid = mem25_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem25_io_bus_response_bits_data = mem25_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu26_clock = clock;
  assign cpu26_reset = reset;
  assign cpu26_io_imem_instruction = imem26_io_pipeline_instruction; // @[top.scala 199:17]
  assign cpu26_io_dmem_readdata = dmem26_io_pipeline_readdata; // @[top.scala 200:17]
  assign mem26_clock = clock;
  assign mem26_reset = reset;
  assign mem26_io_imem_request_bits_address = imem26_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem26_io_dmem_request_valid = dmem26_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem26_io_dmem_request_bits_address = dmem26_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem26_io_dmem_request_bits_writedata = dmem26_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem26_io_dmem_request_bits_operation = dmem26_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem26_io_pipeline_address = cpu26_io_imem_address; // @[top.scala 199:17]
  assign imem26_io_bus_response_bits_data = mem26_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem26_clock = clock;
  assign dmem26_reset = reset;
  assign dmem26_io_pipeline_address = cpu26_io_dmem_address; // @[top.scala 200:17]
  assign dmem26_io_pipeline_valid = cpu26_io_dmem_valid; // @[top.scala 200:17]
  assign dmem26_io_pipeline_writedata = cpu26_io_dmem_writedata; // @[top.scala 200:17]
  assign dmem26_io_pipeline_memread = cpu26_io_dmem_memread; // @[top.scala 200:17]
  assign dmem26_io_pipeline_memwrite = cpu26_io_dmem_memwrite; // @[top.scala 200:17]
  assign dmem26_io_pipeline_maskmode = cpu26_io_dmem_maskmode; // @[top.scala 200:17]
  assign dmem26_io_pipeline_sext = cpu26_io_dmem_sext; // @[top.scala 200:17]
  assign dmem26_io_bus_response_valid = mem26_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem26_io_bus_response_bits_data = mem26_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu27_clock = clock;
  assign cpu27_reset = reset;
  assign cpu27_io_imem_instruction = imem27_io_pipeline_instruction; // @[top.scala 206:17]
  assign cpu27_io_dmem_readdata = dmem27_io_pipeline_readdata; // @[top.scala 207:17]
  assign mem27_clock = clock;
  assign mem27_reset = reset;
  assign mem27_io_imem_request_bits_address = imem27_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem27_io_dmem_request_valid = dmem27_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem27_io_dmem_request_bits_address = dmem27_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem27_io_dmem_request_bits_writedata = dmem27_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem27_io_dmem_request_bits_operation = dmem27_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem27_io_pipeline_address = cpu27_io_imem_address; // @[top.scala 206:17]
  assign imem27_io_bus_response_bits_data = mem27_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem27_clock = clock;
  assign dmem27_reset = reset;
  assign dmem27_io_pipeline_address = cpu27_io_dmem_address; // @[top.scala 207:17]
  assign dmem27_io_pipeline_valid = cpu27_io_dmem_valid; // @[top.scala 207:17]
  assign dmem27_io_pipeline_writedata = cpu27_io_dmem_writedata; // @[top.scala 207:17]
  assign dmem27_io_pipeline_memread = cpu27_io_dmem_memread; // @[top.scala 207:17]
  assign dmem27_io_pipeline_memwrite = cpu27_io_dmem_memwrite; // @[top.scala 207:17]
  assign dmem27_io_pipeline_maskmode = cpu27_io_dmem_maskmode; // @[top.scala 207:17]
  assign dmem27_io_pipeline_sext = cpu27_io_dmem_sext; // @[top.scala 207:17]
  assign dmem27_io_bus_response_valid = mem27_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem27_io_bus_response_bits_data = mem27_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu28_clock = clock;
  assign cpu28_reset = reset;
  assign cpu28_io_imem_instruction = imem28_io_pipeline_instruction; // @[top.scala 213:17]
  assign cpu28_io_dmem_readdata = dmem28_io_pipeline_readdata; // @[top.scala 214:17]
  assign mem28_clock = clock;
  assign mem28_reset = reset;
  assign mem28_io_imem_request_bits_address = imem28_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem28_io_dmem_request_valid = dmem28_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem28_io_dmem_request_bits_address = dmem28_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem28_io_dmem_request_bits_writedata = dmem28_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem28_io_dmem_request_bits_operation = dmem28_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem28_io_pipeline_address = cpu28_io_imem_address; // @[top.scala 213:17]
  assign imem28_io_bus_response_bits_data = mem28_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem28_clock = clock;
  assign dmem28_reset = reset;
  assign dmem28_io_pipeline_address = cpu28_io_dmem_address; // @[top.scala 214:17]
  assign dmem28_io_pipeline_valid = cpu28_io_dmem_valid; // @[top.scala 214:17]
  assign dmem28_io_pipeline_writedata = cpu28_io_dmem_writedata; // @[top.scala 214:17]
  assign dmem28_io_pipeline_memread = cpu28_io_dmem_memread; // @[top.scala 214:17]
  assign dmem28_io_pipeline_memwrite = cpu28_io_dmem_memwrite; // @[top.scala 214:17]
  assign dmem28_io_pipeline_maskmode = cpu28_io_dmem_maskmode; // @[top.scala 214:17]
  assign dmem28_io_pipeline_sext = cpu28_io_dmem_sext; // @[top.scala 214:17]
  assign dmem28_io_bus_response_valid = mem28_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem28_io_bus_response_bits_data = mem28_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu29_clock = clock;
  assign cpu29_reset = reset;
  assign cpu29_io_imem_instruction = imem29_io_pipeline_instruction; // @[top.scala 220:17]
  assign cpu29_io_dmem_readdata = dmem29_io_pipeline_readdata; // @[top.scala 221:17]
  assign mem29_clock = clock;
  assign mem29_reset = reset;
  assign mem29_io_imem_request_bits_address = imem29_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem29_io_dmem_request_valid = dmem29_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem29_io_dmem_request_bits_address = dmem29_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem29_io_dmem_request_bits_writedata = dmem29_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem29_io_dmem_request_bits_operation = dmem29_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem29_io_pipeline_address = cpu29_io_imem_address; // @[top.scala 220:17]
  assign imem29_io_bus_response_bits_data = mem29_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem29_clock = clock;
  assign dmem29_reset = reset;
  assign dmem29_io_pipeline_address = cpu29_io_dmem_address; // @[top.scala 221:17]
  assign dmem29_io_pipeline_valid = cpu29_io_dmem_valid; // @[top.scala 221:17]
  assign dmem29_io_pipeline_writedata = cpu29_io_dmem_writedata; // @[top.scala 221:17]
  assign dmem29_io_pipeline_memread = cpu29_io_dmem_memread; // @[top.scala 221:17]
  assign dmem29_io_pipeline_memwrite = cpu29_io_dmem_memwrite; // @[top.scala 221:17]
  assign dmem29_io_pipeline_maskmode = cpu29_io_dmem_maskmode; // @[top.scala 221:17]
  assign dmem29_io_pipeline_sext = cpu29_io_dmem_sext; // @[top.scala 221:17]
  assign dmem29_io_bus_response_valid = mem29_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem29_io_bus_response_bits_data = mem29_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu30_clock = clock;
  assign cpu30_reset = reset;
  assign cpu30_io_imem_instruction = imem30_io_pipeline_instruction; // @[top.scala 227:17]
  assign cpu30_io_dmem_readdata = dmem30_io_pipeline_readdata; // @[top.scala 228:17]
  assign mem30_clock = clock;
  assign mem30_reset = reset;
  assign mem30_io_imem_request_bits_address = imem30_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem30_io_dmem_request_valid = dmem30_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem30_io_dmem_request_bits_address = dmem30_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem30_io_dmem_request_bits_writedata = dmem30_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem30_io_dmem_request_bits_operation = dmem30_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem30_io_pipeline_address = cpu30_io_imem_address; // @[top.scala 227:17]
  assign imem30_io_bus_response_bits_data = mem30_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem30_clock = clock;
  assign dmem30_reset = reset;
  assign dmem30_io_pipeline_address = cpu30_io_dmem_address; // @[top.scala 228:17]
  assign dmem30_io_pipeline_valid = cpu30_io_dmem_valid; // @[top.scala 228:17]
  assign dmem30_io_pipeline_writedata = cpu30_io_dmem_writedata; // @[top.scala 228:17]
  assign dmem30_io_pipeline_memread = cpu30_io_dmem_memread; // @[top.scala 228:17]
  assign dmem30_io_pipeline_memwrite = cpu30_io_dmem_memwrite; // @[top.scala 228:17]
  assign dmem30_io_pipeline_maskmode = cpu30_io_dmem_maskmode; // @[top.scala 228:17]
  assign dmem30_io_pipeline_sext = cpu30_io_dmem_sext; // @[top.scala 228:17]
  assign dmem30_io_bus_response_valid = mem30_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem30_io_bus_response_bits_data = mem30_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu31_clock = clock;
  assign cpu31_reset = reset;
  assign cpu31_io_imem_instruction = imem31_io_pipeline_instruction; // @[top.scala 234:17]
  assign cpu31_io_dmem_readdata = dmem31_io_pipeline_readdata; // @[top.scala 235:17]
  assign mem31_clock = clock;
  assign mem31_reset = reset;
  assign mem31_io_imem_request_bits_address = imem31_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem31_io_dmem_request_valid = dmem31_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem31_io_dmem_request_bits_address = dmem31_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem31_io_dmem_request_bits_writedata = dmem31_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem31_io_dmem_request_bits_operation = dmem31_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem31_io_pipeline_address = cpu31_io_imem_address; // @[top.scala 234:17]
  assign imem31_io_bus_response_bits_data = mem31_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem31_clock = clock;
  assign dmem31_reset = reset;
  assign dmem31_io_pipeline_address = cpu31_io_dmem_address; // @[top.scala 235:17]
  assign dmem31_io_pipeline_valid = cpu31_io_dmem_valid; // @[top.scala 235:17]
  assign dmem31_io_pipeline_writedata = cpu31_io_dmem_writedata; // @[top.scala 235:17]
  assign dmem31_io_pipeline_memread = cpu31_io_dmem_memread; // @[top.scala 235:17]
  assign dmem31_io_pipeline_memwrite = cpu31_io_dmem_memwrite; // @[top.scala 235:17]
  assign dmem31_io_pipeline_maskmode = cpu31_io_dmem_maskmode; // @[top.scala 235:17]
  assign dmem31_io_pipeline_sext = cpu31_io_dmem_sext; // @[top.scala 235:17]
  assign dmem31_io_bus_response_valid = mem31_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem31_io_bus_response_bits_data = mem31_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu32_clock = clock;
  assign cpu32_reset = reset;
  assign cpu32_io_imem_instruction = imem32_io_pipeline_instruction; // @[top.scala 241:17]
  assign cpu32_io_dmem_readdata = dmem32_io_pipeline_readdata; // @[top.scala 242:17]
  assign mem32_clock = clock;
  assign mem32_reset = reset;
  assign mem32_io_imem_request_bits_address = imem32_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem32_io_dmem_request_valid = dmem32_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem32_io_dmem_request_bits_address = dmem32_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem32_io_dmem_request_bits_writedata = dmem32_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem32_io_dmem_request_bits_operation = dmem32_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem32_io_pipeline_address = cpu32_io_imem_address; // @[top.scala 241:17]
  assign imem32_io_bus_response_bits_data = mem32_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem32_clock = clock;
  assign dmem32_reset = reset;
  assign dmem32_io_pipeline_address = cpu32_io_dmem_address; // @[top.scala 242:17]
  assign dmem32_io_pipeline_valid = cpu32_io_dmem_valid; // @[top.scala 242:17]
  assign dmem32_io_pipeline_writedata = cpu32_io_dmem_writedata; // @[top.scala 242:17]
  assign dmem32_io_pipeline_memread = cpu32_io_dmem_memread; // @[top.scala 242:17]
  assign dmem32_io_pipeline_memwrite = cpu32_io_dmem_memwrite; // @[top.scala 242:17]
  assign dmem32_io_pipeline_maskmode = cpu32_io_dmem_maskmode; // @[top.scala 242:17]
  assign dmem32_io_pipeline_sext = cpu32_io_dmem_sext; // @[top.scala 242:17]
  assign dmem32_io_bus_response_valid = mem32_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem32_io_bus_response_bits_data = mem32_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu33_clock = clock;
  assign cpu33_reset = reset;
  assign cpu33_io_imem_instruction = imem33_io_pipeline_instruction; // @[top.scala 248:17]
  assign cpu33_io_dmem_readdata = dmem33_io_pipeline_readdata; // @[top.scala 249:17]
  assign mem33_clock = clock;
  assign mem33_reset = reset;
  assign mem33_io_imem_request_bits_address = imem33_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem33_io_dmem_request_valid = dmem33_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem33_io_dmem_request_bits_address = dmem33_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem33_io_dmem_request_bits_writedata = dmem33_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem33_io_dmem_request_bits_operation = dmem33_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem33_io_pipeline_address = cpu33_io_imem_address; // @[top.scala 248:17]
  assign imem33_io_bus_response_bits_data = mem33_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem33_clock = clock;
  assign dmem33_reset = reset;
  assign dmem33_io_pipeline_address = cpu33_io_dmem_address; // @[top.scala 249:17]
  assign dmem33_io_pipeline_valid = cpu33_io_dmem_valid; // @[top.scala 249:17]
  assign dmem33_io_pipeline_writedata = cpu33_io_dmem_writedata; // @[top.scala 249:17]
  assign dmem33_io_pipeline_memread = cpu33_io_dmem_memread; // @[top.scala 249:17]
  assign dmem33_io_pipeline_memwrite = cpu33_io_dmem_memwrite; // @[top.scala 249:17]
  assign dmem33_io_pipeline_maskmode = cpu33_io_dmem_maskmode; // @[top.scala 249:17]
  assign dmem33_io_pipeline_sext = cpu33_io_dmem_sext; // @[top.scala 249:17]
  assign dmem33_io_bus_response_valid = mem33_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem33_io_bus_response_bits_data = mem33_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu34_clock = clock;
  assign cpu34_reset = reset;
  assign cpu34_io_imem_instruction = imem34_io_pipeline_instruction; // @[top.scala 255:17]
  assign cpu34_io_dmem_readdata = dmem34_io_pipeline_readdata; // @[top.scala 256:17]
  assign mem34_clock = clock;
  assign mem34_reset = reset;
  assign mem34_io_imem_request_bits_address = imem34_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem34_io_dmem_request_valid = dmem34_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem34_io_dmem_request_bits_address = dmem34_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem34_io_dmem_request_bits_writedata = dmem34_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem34_io_dmem_request_bits_operation = dmem34_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem34_io_pipeline_address = cpu34_io_imem_address; // @[top.scala 255:17]
  assign imem34_io_bus_response_bits_data = mem34_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem34_clock = clock;
  assign dmem34_reset = reset;
  assign dmem34_io_pipeline_address = cpu34_io_dmem_address; // @[top.scala 256:17]
  assign dmem34_io_pipeline_valid = cpu34_io_dmem_valid; // @[top.scala 256:17]
  assign dmem34_io_pipeline_writedata = cpu34_io_dmem_writedata; // @[top.scala 256:17]
  assign dmem34_io_pipeline_memread = cpu34_io_dmem_memread; // @[top.scala 256:17]
  assign dmem34_io_pipeline_memwrite = cpu34_io_dmem_memwrite; // @[top.scala 256:17]
  assign dmem34_io_pipeline_maskmode = cpu34_io_dmem_maskmode; // @[top.scala 256:17]
  assign dmem34_io_pipeline_sext = cpu34_io_dmem_sext; // @[top.scala 256:17]
  assign dmem34_io_bus_response_valid = mem34_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem34_io_bus_response_bits_data = mem34_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu35_clock = clock;
  assign cpu35_reset = reset;
  assign cpu35_io_imem_instruction = imem35_io_pipeline_instruction; // @[top.scala 262:17]
  assign cpu35_io_dmem_readdata = dmem35_io_pipeline_readdata; // @[top.scala 263:17]
  assign mem35_clock = clock;
  assign mem35_reset = reset;
  assign mem35_io_imem_request_bits_address = imem35_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem35_io_dmem_request_valid = dmem35_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem35_io_dmem_request_bits_address = dmem35_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem35_io_dmem_request_bits_writedata = dmem35_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem35_io_dmem_request_bits_operation = dmem35_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem35_io_pipeline_address = cpu35_io_imem_address; // @[top.scala 262:17]
  assign imem35_io_bus_response_bits_data = mem35_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem35_clock = clock;
  assign dmem35_reset = reset;
  assign dmem35_io_pipeline_address = cpu35_io_dmem_address; // @[top.scala 263:17]
  assign dmem35_io_pipeline_valid = cpu35_io_dmem_valid; // @[top.scala 263:17]
  assign dmem35_io_pipeline_writedata = cpu35_io_dmem_writedata; // @[top.scala 263:17]
  assign dmem35_io_pipeline_memread = cpu35_io_dmem_memread; // @[top.scala 263:17]
  assign dmem35_io_pipeline_memwrite = cpu35_io_dmem_memwrite; // @[top.scala 263:17]
  assign dmem35_io_pipeline_maskmode = cpu35_io_dmem_maskmode; // @[top.scala 263:17]
  assign dmem35_io_pipeline_sext = cpu35_io_dmem_sext; // @[top.scala 263:17]
  assign dmem35_io_bus_response_valid = mem35_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem35_io_bus_response_bits_data = mem35_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu36_clock = clock;
  assign cpu36_reset = reset;
  assign cpu36_io_imem_instruction = imem36_io_pipeline_instruction; // @[top.scala 269:17]
  assign cpu36_io_dmem_readdata = dmem36_io_pipeline_readdata; // @[top.scala 270:17]
  assign mem36_clock = clock;
  assign mem36_reset = reset;
  assign mem36_io_imem_request_bits_address = imem36_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem36_io_dmem_request_valid = dmem36_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem36_io_dmem_request_bits_address = dmem36_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem36_io_dmem_request_bits_writedata = dmem36_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem36_io_dmem_request_bits_operation = dmem36_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem36_io_pipeline_address = cpu36_io_imem_address; // @[top.scala 269:17]
  assign imem36_io_bus_response_bits_data = mem36_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem36_clock = clock;
  assign dmem36_reset = reset;
  assign dmem36_io_pipeline_address = cpu36_io_dmem_address; // @[top.scala 270:17]
  assign dmem36_io_pipeline_valid = cpu36_io_dmem_valid; // @[top.scala 270:17]
  assign dmem36_io_pipeline_writedata = cpu36_io_dmem_writedata; // @[top.scala 270:17]
  assign dmem36_io_pipeline_memread = cpu36_io_dmem_memread; // @[top.scala 270:17]
  assign dmem36_io_pipeline_memwrite = cpu36_io_dmem_memwrite; // @[top.scala 270:17]
  assign dmem36_io_pipeline_maskmode = cpu36_io_dmem_maskmode; // @[top.scala 270:17]
  assign dmem36_io_pipeline_sext = cpu36_io_dmem_sext; // @[top.scala 270:17]
  assign dmem36_io_bus_response_valid = mem36_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem36_io_bus_response_bits_data = mem36_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu37_clock = clock;
  assign cpu37_reset = reset;
  assign cpu37_io_imem_instruction = imem37_io_pipeline_instruction; // @[top.scala 276:17]
  assign cpu37_io_dmem_readdata = dmem37_io_pipeline_readdata; // @[top.scala 277:17]
  assign mem37_clock = clock;
  assign mem37_reset = reset;
  assign mem37_io_imem_request_bits_address = imem37_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem37_io_dmem_request_valid = dmem37_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem37_io_dmem_request_bits_address = dmem37_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem37_io_dmem_request_bits_writedata = dmem37_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem37_io_dmem_request_bits_operation = dmem37_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem37_io_pipeline_address = cpu37_io_imem_address; // @[top.scala 276:17]
  assign imem37_io_bus_response_bits_data = mem37_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem37_clock = clock;
  assign dmem37_reset = reset;
  assign dmem37_io_pipeline_address = cpu37_io_dmem_address; // @[top.scala 277:17]
  assign dmem37_io_pipeline_valid = cpu37_io_dmem_valid; // @[top.scala 277:17]
  assign dmem37_io_pipeline_writedata = cpu37_io_dmem_writedata; // @[top.scala 277:17]
  assign dmem37_io_pipeline_memread = cpu37_io_dmem_memread; // @[top.scala 277:17]
  assign dmem37_io_pipeline_memwrite = cpu37_io_dmem_memwrite; // @[top.scala 277:17]
  assign dmem37_io_pipeline_maskmode = cpu37_io_dmem_maskmode; // @[top.scala 277:17]
  assign dmem37_io_pipeline_sext = cpu37_io_dmem_sext; // @[top.scala 277:17]
  assign dmem37_io_bus_response_valid = mem37_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem37_io_bus_response_bits_data = mem37_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu38_clock = clock;
  assign cpu38_reset = reset;
  assign cpu38_io_imem_instruction = imem38_io_pipeline_instruction; // @[top.scala 283:17]
  assign cpu38_io_dmem_readdata = dmem38_io_pipeline_readdata; // @[top.scala 284:17]
  assign mem38_clock = clock;
  assign mem38_reset = reset;
  assign mem38_io_imem_request_bits_address = imem38_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem38_io_dmem_request_valid = dmem38_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem38_io_dmem_request_bits_address = dmem38_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem38_io_dmem_request_bits_writedata = dmem38_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem38_io_dmem_request_bits_operation = dmem38_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem38_io_pipeline_address = cpu38_io_imem_address; // @[top.scala 283:17]
  assign imem38_io_bus_response_bits_data = mem38_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem38_clock = clock;
  assign dmem38_reset = reset;
  assign dmem38_io_pipeline_address = cpu38_io_dmem_address; // @[top.scala 284:17]
  assign dmem38_io_pipeline_valid = cpu38_io_dmem_valid; // @[top.scala 284:17]
  assign dmem38_io_pipeline_writedata = cpu38_io_dmem_writedata; // @[top.scala 284:17]
  assign dmem38_io_pipeline_memread = cpu38_io_dmem_memread; // @[top.scala 284:17]
  assign dmem38_io_pipeline_memwrite = cpu38_io_dmem_memwrite; // @[top.scala 284:17]
  assign dmem38_io_pipeline_maskmode = cpu38_io_dmem_maskmode; // @[top.scala 284:17]
  assign dmem38_io_pipeline_sext = cpu38_io_dmem_sext; // @[top.scala 284:17]
  assign dmem38_io_bus_response_valid = mem38_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem38_io_bus_response_bits_data = mem38_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu39_clock = clock;
  assign cpu39_reset = reset;
  assign cpu39_io_imem_instruction = imem39_io_pipeline_instruction; // @[top.scala 290:17]
  assign cpu39_io_dmem_readdata = dmem39_io_pipeline_readdata; // @[top.scala 291:17]
  assign mem39_clock = clock;
  assign mem39_reset = reset;
  assign mem39_io_imem_request_bits_address = imem39_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem39_io_dmem_request_valid = dmem39_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem39_io_dmem_request_bits_address = dmem39_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem39_io_dmem_request_bits_writedata = dmem39_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem39_io_dmem_request_bits_operation = dmem39_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem39_io_pipeline_address = cpu39_io_imem_address; // @[top.scala 290:17]
  assign imem39_io_bus_response_bits_data = mem39_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem39_clock = clock;
  assign dmem39_reset = reset;
  assign dmem39_io_pipeline_address = cpu39_io_dmem_address; // @[top.scala 291:17]
  assign dmem39_io_pipeline_valid = cpu39_io_dmem_valid; // @[top.scala 291:17]
  assign dmem39_io_pipeline_writedata = cpu39_io_dmem_writedata; // @[top.scala 291:17]
  assign dmem39_io_pipeline_memread = cpu39_io_dmem_memread; // @[top.scala 291:17]
  assign dmem39_io_pipeline_memwrite = cpu39_io_dmem_memwrite; // @[top.scala 291:17]
  assign dmem39_io_pipeline_maskmode = cpu39_io_dmem_maskmode; // @[top.scala 291:17]
  assign dmem39_io_pipeline_sext = cpu39_io_dmem_sext; // @[top.scala 291:17]
  assign dmem39_io_bus_response_valid = mem39_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem39_io_bus_response_bits_data = mem39_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu40_clock = clock;
  assign cpu40_reset = reset;
  assign cpu40_io_imem_instruction = imem40_io_pipeline_instruction; // @[top.scala 297:17]
  assign cpu40_io_dmem_readdata = dmem40_io_pipeline_readdata; // @[top.scala 298:17]
  assign mem40_clock = clock;
  assign mem40_reset = reset;
  assign mem40_io_imem_request_bits_address = imem40_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem40_io_dmem_request_valid = dmem40_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem40_io_dmem_request_bits_address = dmem40_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem40_io_dmem_request_bits_writedata = dmem40_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem40_io_dmem_request_bits_operation = dmem40_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem40_io_pipeline_address = cpu40_io_imem_address; // @[top.scala 297:17]
  assign imem40_io_bus_response_bits_data = mem40_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem40_clock = clock;
  assign dmem40_reset = reset;
  assign dmem40_io_pipeline_address = cpu40_io_dmem_address; // @[top.scala 298:17]
  assign dmem40_io_pipeline_valid = cpu40_io_dmem_valid; // @[top.scala 298:17]
  assign dmem40_io_pipeline_writedata = cpu40_io_dmem_writedata; // @[top.scala 298:17]
  assign dmem40_io_pipeline_memread = cpu40_io_dmem_memread; // @[top.scala 298:17]
  assign dmem40_io_pipeline_memwrite = cpu40_io_dmem_memwrite; // @[top.scala 298:17]
  assign dmem40_io_pipeline_maskmode = cpu40_io_dmem_maskmode; // @[top.scala 298:17]
  assign dmem40_io_pipeline_sext = cpu40_io_dmem_sext; // @[top.scala 298:17]
  assign dmem40_io_bus_response_valid = mem40_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem40_io_bus_response_bits_data = mem40_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu41_clock = clock;
  assign cpu41_reset = reset;
  assign cpu41_io_imem_instruction = imem41_io_pipeline_instruction; // @[top.scala 304:17]
  assign cpu41_io_dmem_readdata = dmem41_io_pipeline_readdata; // @[top.scala 305:17]
  assign mem41_clock = clock;
  assign mem41_reset = reset;
  assign mem41_io_imem_request_bits_address = imem41_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem41_io_dmem_request_valid = dmem41_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem41_io_dmem_request_bits_address = dmem41_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem41_io_dmem_request_bits_writedata = dmem41_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem41_io_dmem_request_bits_operation = dmem41_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem41_io_pipeline_address = cpu41_io_imem_address; // @[top.scala 304:17]
  assign imem41_io_bus_response_bits_data = mem41_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem41_clock = clock;
  assign dmem41_reset = reset;
  assign dmem41_io_pipeline_address = cpu41_io_dmem_address; // @[top.scala 305:17]
  assign dmem41_io_pipeline_valid = cpu41_io_dmem_valid; // @[top.scala 305:17]
  assign dmem41_io_pipeline_writedata = cpu41_io_dmem_writedata; // @[top.scala 305:17]
  assign dmem41_io_pipeline_memread = cpu41_io_dmem_memread; // @[top.scala 305:17]
  assign dmem41_io_pipeline_memwrite = cpu41_io_dmem_memwrite; // @[top.scala 305:17]
  assign dmem41_io_pipeline_maskmode = cpu41_io_dmem_maskmode; // @[top.scala 305:17]
  assign dmem41_io_pipeline_sext = cpu41_io_dmem_sext; // @[top.scala 305:17]
  assign dmem41_io_bus_response_valid = mem41_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem41_io_bus_response_bits_data = mem41_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu42_clock = clock;
  assign cpu42_reset = reset;
  assign cpu42_io_imem_instruction = imem42_io_pipeline_instruction; // @[top.scala 311:17]
  assign cpu42_io_dmem_readdata = dmem42_io_pipeline_readdata; // @[top.scala 312:17]
  assign mem42_clock = clock;
  assign mem42_reset = reset;
  assign mem42_io_imem_request_bits_address = imem42_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem42_io_dmem_request_valid = dmem42_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem42_io_dmem_request_bits_address = dmem42_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem42_io_dmem_request_bits_writedata = dmem42_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem42_io_dmem_request_bits_operation = dmem42_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem42_io_pipeline_address = cpu42_io_imem_address; // @[top.scala 311:17]
  assign imem42_io_bus_response_bits_data = mem42_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem42_clock = clock;
  assign dmem42_reset = reset;
  assign dmem42_io_pipeline_address = cpu42_io_dmem_address; // @[top.scala 312:17]
  assign dmem42_io_pipeline_valid = cpu42_io_dmem_valid; // @[top.scala 312:17]
  assign dmem42_io_pipeline_writedata = cpu42_io_dmem_writedata; // @[top.scala 312:17]
  assign dmem42_io_pipeline_memread = cpu42_io_dmem_memread; // @[top.scala 312:17]
  assign dmem42_io_pipeline_memwrite = cpu42_io_dmem_memwrite; // @[top.scala 312:17]
  assign dmem42_io_pipeline_maskmode = cpu42_io_dmem_maskmode; // @[top.scala 312:17]
  assign dmem42_io_pipeline_sext = cpu42_io_dmem_sext; // @[top.scala 312:17]
  assign dmem42_io_bus_response_valid = mem42_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem42_io_bus_response_bits_data = mem42_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu43_clock = clock;
  assign cpu43_reset = reset;
  assign cpu43_io_imem_instruction = imem43_io_pipeline_instruction; // @[top.scala 318:17]
  assign cpu43_io_dmem_readdata = dmem43_io_pipeline_readdata; // @[top.scala 319:17]
  assign mem43_clock = clock;
  assign mem43_reset = reset;
  assign mem43_io_imem_request_bits_address = imem43_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem43_io_dmem_request_valid = dmem43_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem43_io_dmem_request_bits_address = dmem43_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem43_io_dmem_request_bits_writedata = dmem43_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem43_io_dmem_request_bits_operation = dmem43_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem43_io_pipeline_address = cpu43_io_imem_address; // @[top.scala 318:17]
  assign imem43_io_bus_response_bits_data = mem43_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem43_clock = clock;
  assign dmem43_reset = reset;
  assign dmem43_io_pipeline_address = cpu43_io_dmem_address; // @[top.scala 319:17]
  assign dmem43_io_pipeline_valid = cpu43_io_dmem_valid; // @[top.scala 319:17]
  assign dmem43_io_pipeline_writedata = cpu43_io_dmem_writedata; // @[top.scala 319:17]
  assign dmem43_io_pipeline_memread = cpu43_io_dmem_memread; // @[top.scala 319:17]
  assign dmem43_io_pipeline_memwrite = cpu43_io_dmem_memwrite; // @[top.scala 319:17]
  assign dmem43_io_pipeline_maskmode = cpu43_io_dmem_maskmode; // @[top.scala 319:17]
  assign dmem43_io_pipeline_sext = cpu43_io_dmem_sext; // @[top.scala 319:17]
  assign dmem43_io_bus_response_valid = mem43_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem43_io_bus_response_bits_data = mem43_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu44_clock = clock;
  assign cpu44_reset = reset;
  assign cpu44_io_imem_instruction = imem44_io_pipeline_instruction; // @[top.scala 325:17]
  assign cpu44_io_dmem_readdata = dmem44_io_pipeline_readdata; // @[top.scala 326:17]
  assign mem44_clock = clock;
  assign mem44_reset = reset;
  assign mem44_io_imem_request_bits_address = imem44_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem44_io_dmem_request_valid = dmem44_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem44_io_dmem_request_bits_address = dmem44_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem44_io_dmem_request_bits_writedata = dmem44_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem44_io_dmem_request_bits_operation = dmem44_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem44_io_pipeline_address = cpu44_io_imem_address; // @[top.scala 325:17]
  assign imem44_io_bus_response_bits_data = mem44_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem44_clock = clock;
  assign dmem44_reset = reset;
  assign dmem44_io_pipeline_address = cpu44_io_dmem_address; // @[top.scala 326:17]
  assign dmem44_io_pipeline_valid = cpu44_io_dmem_valid; // @[top.scala 326:17]
  assign dmem44_io_pipeline_writedata = cpu44_io_dmem_writedata; // @[top.scala 326:17]
  assign dmem44_io_pipeline_memread = cpu44_io_dmem_memread; // @[top.scala 326:17]
  assign dmem44_io_pipeline_memwrite = cpu44_io_dmem_memwrite; // @[top.scala 326:17]
  assign dmem44_io_pipeline_maskmode = cpu44_io_dmem_maskmode; // @[top.scala 326:17]
  assign dmem44_io_pipeline_sext = cpu44_io_dmem_sext; // @[top.scala 326:17]
  assign dmem44_io_bus_response_valid = mem44_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem44_io_bus_response_bits_data = mem44_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu45_clock = clock;
  assign cpu45_reset = reset;
  assign cpu45_io_imem_instruction = imem45_io_pipeline_instruction; // @[top.scala 332:17]
  assign cpu45_io_dmem_readdata = dmem45_io_pipeline_readdata; // @[top.scala 333:17]
  assign mem45_clock = clock;
  assign mem45_reset = reset;
  assign mem45_io_imem_request_bits_address = imem45_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem45_io_dmem_request_valid = dmem45_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem45_io_dmem_request_bits_address = dmem45_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem45_io_dmem_request_bits_writedata = dmem45_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem45_io_dmem_request_bits_operation = dmem45_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem45_io_pipeline_address = cpu45_io_imem_address; // @[top.scala 332:17]
  assign imem45_io_bus_response_bits_data = mem45_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem45_clock = clock;
  assign dmem45_reset = reset;
  assign dmem45_io_pipeline_address = cpu45_io_dmem_address; // @[top.scala 333:17]
  assign dmem45_io_pipeline_valid = cpu45_io_dmem_valid; // @[top.scala 333:17]
  assign dmem45_io_pipeline_writedata = cpu45_io_dmem_writedata; // @[top.scala 333:17]
  assign dmem45_io_pipeline_memread = cpu45_io_dmem_memread; // @[top.scala 333:17]
  assign dmem45_io_pipeline_memwrite = cpu45_io_dmem_memwrite; // @[top.scala 333:17]
  assign dmem45_io_pipeline_maskmode = cpu45_io_dmem_maskmode; // @[top.scala 333:17]
  assign dmem45_io_pipeline_sext = cpu45_io_dmem_sext; // @[top.scala 333:17]
  assign dmem45_io_bus_response_valid = mem45_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem45_io_bus_response_bits_data = mem45_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu46_clock = clock;
  assign cpu46_reset = reset;
  assign cpu46_io_imem_instruction = imem46_io_pipeline_instruction; // @[top.scala 339:17]
  assign cpu46_io_dmem_readdata = dmem46_io_pipeline_readdata; // @[top.scala 340:17]
  assign mem46_clock = clock;
  assign mem46_reset = reset;
  assign mem46_io_imem_request_bits_address = imem46_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem46_io_dmem_request_valid = dmem46_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem46_io_dmem_request_bits_address = dmem46_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem46_io_dmem_request_bits_writedata = dmem46_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem46_io_dmem_request_bits_operation = dmem46_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem46_io_pipeline_address = cpu46_io_imem_address; // @[top.scala 339:17]
  assign imem46_io_bus_response_bits_data = mem46_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem46_clock = clock;
  assign dmem46_reset = reset;
  assign dmem46_io_pipeline_address = cpu46_io_dmem_address; // @[top.scala 340:17]
  assign dmem46_io_pipeline_valid = cpu46_io_dmem_valid; // @[top.scala 340:17]
  assign dmem46_io_pipeline_writedata = cpu46_io_dmem_writedata; // @[top.scala 340:17]
  assign dmem46_io_pipeline_memread = cpu46_io_dmem_memread; // @[top.scala 340:17]
  assign dmem46_io_pipeline_memwrite = cpu46_io_dmem_memwrite; // @[top.scala 340:17]
  assign dmem46_io_pipeline_maskmode = cpu46_io_dmem_maskmode; // @[top.scala 340:17]
  assign dmem46_io_pipeline_sext = cpu46_io_dmem_sext; // @[top.scala 340:17]
  assign dmem46_io_bus_response_valid = mem46_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem46_io_bus_response_bits_data = mem46_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu47_clock = clock;
  assign cpu47_reset = reset;
  assign cpu47_io_imem_instruction = imem47_io_pipeline_instruction; // @[top.scala 346:17]
  assign cpu47_io_dmem_readdata = dmem47_io_pipeline_readdata; // @[top.scala 347:17]
  assign mem47_clock = clock;
  assign mem47_reset = reset;
  assign mem47_io_imem_request_bits_address = imem47_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem47_io_dmem_request_valid = dmem47_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem47_io_dmem_request_bits_address = dmem47_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem47_io_dmem_request_bits_writedata = dmem47_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem47_io_dmem_request_bits_operation = dmem47_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem47_io_pipeline_address = cpu47_io_imem_address; // @[top.scala 346:17]
  assign imem47_io_bus_response_bits_data = mem47_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem47_clock = clock;
  assign dmem47_reset = reset;
  assign dmem47_io_pipeline_address = cpu47_io_dmem_address; // @[top.scala 347:17]
  assign dmem47_io_pipeline_valid = cpu47_io_dmem_valid; // @[top.scala 347:17]
  assign dmem47_io_pipeline_writedata = cpu47_io_dmem_writedata; // @[top.scala 347:17]
  assign dmem47_io_pipeline_memread = cpu47_io_dmem_memread; // @[top.scala 347:17]
  assign dmem47_io_pipeline_memwrite = cpu47_io_dmem_memwrite; // @[top.scala 347:17]
  assign dmem47_io_pipeline_maskmode = cpu47_io_dmem_maskmode; // @[top.scala 347:17]
  assign dmem47_io_pipeline_sext = cpu47_io_dmem_sext; // @[top.scala 347:17]
  assign dmem47_io_bus_response_valid = mem47_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem47_io_bus_response_bits_data = mem47_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu48_clock = clock;
  assign cpu48_reset = reset;
  assign cpu48_io_imem_instruction = imem48_io_pipeline_instruction; // @[top.scala 353:17]
  assign cpu48_io_dmem_readdata = dmem48_io_pipeline_readdata; // @[top.scala 354:17]
  assign mem48_clock = clock;
  assign mem48_reset = reset;
  assign mem48_io_imem_request_bits_address = imem48_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem48_io_dmem_request_valid = dmem48_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem48_io_dmem_request_bits_address = dmem48_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem48_io_dmem_request_bits_writedata = dmem48_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem48_io_dmem_request_bits_operation = dmem48_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem48_io_pipeline_address = cpu48_io_imem_address; // @[top.scala 353:17]
  assign imem48_io_bus_response_bits_data = mem48_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem48_clock = clock;
  assign dmem48_reset = reset;
  assign dmem48_io_pipeline_address = cpu48_io_dmem_address; // @[top.scala 354:17]
  assign dmem48_io_pipeline_valid = cpu48_io_dmem_valid; // @[top.scala 354:17]
  assign dmem48_io_pipeline_writedata = cpu48_io_dmem_writedata; // @[top.scala 354:17]
  assign dmem48_io_pipeline_memread = cpu48_io_dmem_memread; // @[top.scala 354:17]
  assign dmem48_io_pipeline_memwrite = cpu48_io_dmem_memwrite; // @[top.scala 354:17]
  assign dmem48_io_pipeline_maskmode = cpu48_io_dmem_maskmode; // @[top.scala 354:17]
  assign dmem48_io_pipeline_sext = cpu48_io_dmem_sext; // @[top.scala 354:17]
  assign dmem48_io_bus_response_valid = mem48_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem48_io_bus_response_bits_data = mem48_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu49_clock = clock;
  assign cpu49_reset = reset;
  assign cpu49_io_imem_instruction = imem49_io_pipeline_instruction; // @[top.scala 360:17]
  assign cpu49_io_dmem_readdata = dmem49_io_pipeline_readdata; // @[top.scala 361:17]
  assign mem49_clock = clock;
  assign mem49_reset = reset;
  assign mem49_io_imem_request_bits_address = imem49_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem49_io_dmem_request_valid = dmem49_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem49_io_dmem_request_bits_address = dmem49_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem49_io_dmem_request_bits_writedata = dmem49_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem49_io_dmem_request_bits_operation = dmem49_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem49_io_pipeline_address = cpu49_io_imem_address; // @[top.scala 360:17]
  assign imem49_io_bus_response_bits_data = mem49_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem49_clock = clock;
  assign dmem49_reset = reset;
  assign dmem49_io_pipeline_address = cpu49_io_dmem_address; // @[top.scala 361:17]
  assign dmem49_io_pipeline_valid = cpu49_io_dmem_valid; // @[top.scala 361:17]
  assign dmem49_io_pipeline_writedata = cpu49_io_dmem_writedata; // @[top.scala 361:17]
  assign dmem49_io_pipeline_memread = cpu49_io_dmem_memread; // @[top.scala 361:17]
  assign dmem49_io_pipeline_memwrite = cpu49_io_dmem_memwrite; // @[top.scala 361:17]
  assign dmem49_io_pipeline_maskmode = cpu49_io_dmem_maskmode; // @[top.scala 361:17]
  assign dmem49_io_pipeline_sext = cpu49_io_dmem_sext; // @[top.scala 361:17]
  assign dmem49_io_bus_response_valid = mem49_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem49_io_bus_response_bits_data = mem49_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu50_clock = clock;
  assign cpu50_reset = reset;
  assign cpu50_io_imem_instruction = imem50_io_pipeline_instruction; // @[top.scala 367:17]
  assign cpu50_io_dmem_readdata = dmem50_io_pipeline_readdata; // @[top.scala 368:17]
  assign mem50_clock = clock;
  assign mem50_reset = reset;
  assign mem50_io_imem_request_bits_address = imem50_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem50_io_dmem_request_valid = dmem50_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem50_io_dmem_request_bits_address = dmem50_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem50_io_dmem_request_bits_writedata = dmem50_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem50_io_dmem_request_bits_operation = dmem50_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem50_io_pipeline_address = cpu50_io_imem_address; // @[top.scala 367:17]
  assign imem50_io_bus_response_bits_data = mem50_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem50_clock = clock;
  assign dmem50_reset = reset;
  assign dmem50_io_pipeline_address = cpu50_io_dmem_address; // @[top.scala 368:17]
  assign dmem50_io_pipeline_valid = cpu50_io_dmem_valid; // @[top.scala 368:17]
  assign dmem50_io_pipeline_writedata = cpu50_io_dmem_writedata; // @[top.scala 368:17]
  assign dmem50_io_pipeline_memread = cpu50_io_dmem_memread; // @[top.scala 368:17]
  assign dmem50_io_pipeline_memwrite = cpu50_io_dmem_memwrite; // @[top.scala 368:17]
  assign dmem50_io_pipeline_maskmode = cpu50_io_dmem_maskmode; // @[top.scala 368:17]
  assign dmem50_io_pipeline_sext = cpu50_io_dmem_sext; // @[top.scala 368:17]
  assign dmem50_io_bus_response_valid = mem50_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem50_io_bus_response_bits_data = mem50_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu51_clock = clock;
  assign cpu51_reset = reset;
  assign cpu51_io_imem_instruction = imem51_io_pipeline_instruction; // @[top.scala 374:17]
  assign cpu51_io_dmem_readdata = dmem51_io_pipeline_readdata; // @[top.scala 375:17]
  assign mem51_clock = clock;
  assign mem51_reset = reset;
  assign mem51_io_imem_request_bits_address = imem51_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem51_io_dmem_request_valid = dmem51_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem51_io_dmem_request_bits_address = dmem51_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem51_io_dmem_request_bits_writedata = dmem51_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem51_io_dmem_request_bits_operation = dmem51_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem51_io_pipeline_address = cpu51_io_imem_address; // @[top.scala 374:17]
  assign imem51_io_bus_response_bits_data = mem51_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem51_clock = clock;
  assign dmem51_reset = reset;
  assign dmem51_io_pipeline_address = cpu51_io_dmem_address; // @[top.scala 375:17]
  assign dmem51_io_pipeline_valid = cpu51_io_dmem_valid; // @[top.scala 375:17]
  assign dmem51_io_pipeline_writedata = cpu51_io_dmem_writedata; // @[top.scala 375:17]
  assign dmem51_io_pipeline_memread = cpu51_io_dmem_memread; // @[top.scala 375:17]
  assign dmem51_io_pipeline_memwrite = cpu51_io_dmem_memwrite; // @[top.scala 375:17]
  assign dmem51_io_pipeline_maskmode = cpu51_io_dmem_maskmode; // @[top.scala 375:17]
  assign dmem51_io_pipeline_sext = cpu51_io_dmem_sext; // @[top.scala 375:17]
  assign dmem51_io_bus_response_valid = mem51_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem51_io_bus_response_bits_data = mem51_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu52_clock = clock;
  assign cpu52_reset = reset;
  assign cpu52_io_imem_instruction = imem52_io_pipeline_instruction; // @[top.scala 381:17]
  assign cpu52_io_dmem_readdata = dmem52_io_pipeline_readdata; // @[top.scala 382:17]
  assign mem52_clock = clock;
  assign mem52_reset = reset;
  assign mem52_io_imem_request_bits_address = imem52_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem52_io_dmem_request_valid = dmem52_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem52_io_dmem_request_bits_address = dmem52_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem52_io_dmem_request_bits_writedata = dmem52_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem52_io_dmem_request_bits_operation = dmem52_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem52_io_pipeline_address = cpu52_io_imem_address; // @[top.scala 381:17]
  assign imem52_io_bus_response_bits_data = mem52_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem52_clock = clock;
  assign dmem52_reset = reset;
  assign dmem52_io_pipeline_address = cpu52_io_dmem_address; // @[top.scala 382:17]
  assign dmem52_io_pipeline_valid = cpu52_io_dmem_valid; // @[top.scala 382:17]
  assign dmem52_io_pipeline_writedata = cpu52_io_dmem_writedata; // @[top.scala 382:17]
  assign dmem52_io_pipeline_memread = cpu52_io_dmem_memread; // @[top.scala 382:17]
  assign dmem52_io_pipeline_memwrite = cpu52_io_dmem_memwrite; // @[top.scala 382:17]
  assign dmem52_io_pipeline_maskmode = cpu52_io_dmem_maskmode; // @[top.scala 382:17]
  assign dmem52_io_pipeline_sext = cpu52_io_dmem_sext; // @[top.scala 382:17]
  assign dmem52_io_bus_response_valid = mem52_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem52_io_bus_response_bits_data = mem52_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu53_clock = clock;
  assign cpu53_reset = reset;
  assign cpu53_io_imem_instruction = imem53_io_pipeline_instruction; // @[top.scala 388:17]
  assign cpu53_io_dmem_readdata = dmem53_io_pipeline_readdata; // @[top.scala 389:17]
  assign mem53_clock = clock;
  assign mem53_reset = reset;
  assign mem53_io_imem_request_bits_address = imem53_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem53_io_dmem_request_valid = dmem53_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem53_io_dmem_request_bits_address = dmem53_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem53_io_dmem_request_bits_writedata = dmem53_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem53_io_dmem_request_bits_operation = dmem53_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem53_io_pipeline_address = cpu53_io_imem_address; // @[top.scala 388:17]
  assign imem53_io_bus_response_bits_data = mem53_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem53_clock = clock;
  assign dmem53_reset = reset;
  assign dmem53_io_pipeline_address = cpu53_io_dmem_address; // @[top.scala 389:17]
  assign dmem53_io_pipeline_valid = cpu53_io_dmem_valid; // @[top.scala 389:17]
  assign dmem53_io_pipeline_writedata = cpu53_io_dmem_writedata; // @[top.scala 389:17]
  assign dmem53_io_pipeline_memread = cpu53_io_dmem_memread; // @[top.scala 389:17]
  assign dmem53_io_pipeline_memwrite = cpu53_io_dmem_memwrite; // @[top.scala 389:17]
  assign dmem53_io_pipeline_maskmode = cpu53_io_dmem_maskmode; // @[top.scala 389:17]
  assign dmem53_io_pipeline_sext = cpu53_io_dmem_sext; // @[top.scala 389:17]
  assign dmem53_io_bus_response_valid = mem53_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem53_io_bus_response_bits_data = mem53_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu54_clock = clock;
  assign cpu54_reset = reset;
  assign cpu54_io_imem_instruction = imem54_io_pipeline_instruction; // @[top.scala 395:17]
  assign cpu54_io_dmem_readdata = dmem54_io_pipeline_readdata; // @[top.scala 396:17]
  assign mem54_clock = clock;
  assign mem54_reset = reset;
  assign mem54_io_imem_request_bits_address = imem54_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem54_io_dmem_request_valid = dmem54_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem54_io_dmem_request_bits_address = dmem54_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem54_io_dmem_request_bits_writedata = dmem54_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem54_io_dmem_request_bits_operation = dmem54_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem54_io_pipeline_address = cpu54_io_imem_address; // @[top.scala 395:17]
  assign imem54_io_bus_response_bits_data = mem54_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem54_clock = clock;
  assign dmem54_reset = reset;
  assign dmem54_io_pipeline_address = cpu54_io_dmem_address; // @[top.scala 396:17]
  assign dmem54_io_pipeline_valid = cpu54_io_dmem_valid; // @[top.scala 396:17]
  assign dmem54_io_pipeline_writedata = cpu54_io_dmem_writedata; // @[top.scala 396:17]
  assign dmem54_io_pipeline_memread = cpu54_io_dmem_memread; // @[top.scala 396:17]
  assign dmem54_io_pipeline_memwrite = cpu54_io_dmem_memwrite; // @[top.scala 396:17]
  assign dmem54_io_pipeline_maskmode = cpu54_io_dmem_maskmode; // @[top.scala 396:17]
  assign dmem54_io_pipeline_sext = cpu54_io_dmem_sext; // @[top.scala 396:17]
  assign dmem54_io_bus_response_valid = mem54_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem54_io_bus_response_bits_data = mem54_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu55_clock = clock;
  assign cpu55_reset = reset;
  assign cpu55_io_imem_instruction = imem55_io_pipeline_instruction; // @[top.scala 402:17]
  assign cpu55_io_dmem_readdata = dmem55_io_pipeline_readdata; // @[top.scala 403:17]
  assign mem55_clock = clock;
  assign mem55_reset = reset;
  assign mem55_io_imem_request_bits_address = imem55_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem55_io_dmem_request_valid = dmem55_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem55_io_dmem_request_bits_address = dmem55_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem55_io_dmem_request_bits_writedata = dmem55_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem55_io_dmem_request_bits_operation = dmem55_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem55_io_pipeline_address = cpu55_io_imem_address; // @[top.scala 402:17]
  assign imem55_io_bus_response_bits_data = mem55_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem55_clock = clock;
  assign dmem55_reset = reset;
  assign dmem55_io_pipeline_address = cpu55_io_dmem_address; // @[top.scala 403:17]
  assign dmem55_io_pipeline_valid = cpu55_io_dmem_valid; // @[top.scala 403:17]
  assign dmem55_io_pipeline_writedata = cpu55_io_dmem_writedata; // @[top.scala 403:17]
  assign dmem55_io_pipeline_memread = cpu55_io_dmem_memread; // @[top.scala 403:17]
  assign dmem55_io_pipeline_memwrite = cpu55_io_dmem_memwrite; // @[top.scala 403:17]
  assign dmem55_io_pipeline_maskmode = cpu55_io_dmem_maskmode; // @[top.scala 403:17]
  assign dmem55_io_pipeline_sext = cpu55_io_dmem_sext; // @[top.scala 403:17]
  assign dmem55_io_bus_response_valid = mem55_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem55_io_bus_response_bits_data = mem55_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu56_clock = clock;
  assign cpu56_reset = reset;
  assign cpu56_io_imem_instruction = imem56_io_pipeline_instruction; // @[top.scala 409:17]
  assign cpu56_io_dmem_readdata = dmem56_io_pipeline_readdata; // @[top.scala 410:17]
  assign mem56_clock = clock;
  assign mem56_reset = reset;
  assign mem56_io_imem_request_bits_address = imem56_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem56_io_dmem_request_valid = dmem56_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem56_io_dmem_request_bits_address = dmem56_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem56_io_dmem_request_bits_writedata = dmem56_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem56_io_dmem_request_bits_operation = dmem56_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem56_io_pipeline_address = cpu56_io_imem_address; // @[top.scala 409:17]
  assign imem56_io_bus_response_bits_data = mem56_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem56_clock = clock;
  assign dmem56_reset = reset;
  assign dmem56_io_pipeline_address = cpu56_io_dmem_address; // @[top.scala 410:17]
  assign dmem56_io_pipeline_valid = cpu56_io_dmem_valid; // @[top.scala 410:17]
  assign dmem56_io_pipeline_writedata = cpu56_io_dmem_writedata; // @[top.scala 410:17]
  assign dmem56_io_pipeline_memread = cpu56_io_dmem_memread; // @[top.scala 410:17]
  assign dmem56_io_pipeline_memwrite = cpu56_io_dmem_memwrite; // @[top.scala 410:17]
  assign dmem56_io_pipeline_maskmode = cpu56_io_dmem_maskmode; // @[top.scala 410:17]
  assign dmem56_io_pipeline_sext = cpu56_io_dmem_sext; // @[top.scala 410:17]
  assign dmem56_io_bus_response_valid = mem56_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem56_io_bus_response_bits_data = mem56_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu57_clock = clock;
  assign cpu57_reset = reset;
  assign cpu57_io_imem_instruction = imem57_io_pipeline_instruction; // @[top.scala 416:17]
  assign cpu57_io_dmem_readdata = dmem57_io_pipeline_readdata; // @[top.scala 417:17]
  assign mem57_clock = clock;
  assign mem57_reset = reset;
  assign mem57_io_imem_request_bits_address = imem57_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem57_io_dmem_request_valid = dmem57_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem57_io_dmem_request_bits_address = dmem57_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem57_io_dmem_request_bits_writedata = dmem57_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem57_io_dmem_request_bits_operation = dmem57_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem57_io_pipeline_address = cpu57_io_imem_address; // @[top.scala 416:17]
  assign imem57_io_bus_response_bits_data = mem57_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem57_clock = clock;
  assign dmem57_reset = reset;
  assign dmem57_io_pipeline_address = cpu57_io_dmem_address; // @[top.scala 417:17]
  assign dmem57_io_pipeline_valid = cpu57_io_dmem_valid; // @[top.scala 417:17]
  assign dmem57_io_pipeline_writedata = cpu57_io_dmem_writedata; // @[top.scala 417:17]
  assign dmem57_io_pipeline_memread = cpu57_io_dmem_memread; // @[top.scala 417:17]
  assign dmem57_io_pipeline_memwrite = cpu57_io_dmem_memwrite; // @[top.scala 417:17]
  assign dmem57_io_pipeline_maskmode = cpu57_io_dmem_maskmode; // @[top.scala 417:17]
  assign dmem57_io_pipeline_sext = cpu57_io_dmem_sext; // @[top.scala 417:17]
  assign dmem57_io_bus_response_valid = mem57_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem57_io_bus_response_bits_data = mem57_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu58_clock = clock;
  assign cpu58_reset = reset;
  assign cpu58_io_imem_instruction = imem58_io_pipeline_instruction; // @[top.scala 423:17]
  assign cpu58_io_dmem_readdata = dmem58_io_pipeline_readdata; // @[top.scala 424:17]
  assign mem58_clock = clock;
  assign mem58_reset = reset;
  assign mem58_io_imem_request_bits_address = imem58_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem58_io_dmem_request_valid = dmem58_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem58_io_dmem_request_bits_address = dmem58_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem58_io_dmem_request_bits_writedata = dmem58_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem58_io_dmem_request_bits_operation = dmem58_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem58_io_pipeline_address = cpu58_io_imem_address; // @[top.scala 423:17]
  assign imem58_io_bus_response_bits_data = mem58_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem58_clock = clock;
  assign dmem58_reset = reset;
  assign dmem58_io_pipeline_address = cpu58_io_dmem_address; // @[top.scala 424:17]
  assign dmem58_io_pipeline_valid = cpu58_io_dmem_valid; // @[top.scala 424:17]
  assign dmem58_io_pipeline_writedata = cpu58_io_dmem_writedata; // @[top.scala 424:17]
  assign dmem58_io_pipeline_memread = cpu58_io_dmem_memread; // @[top.scala 424:17]
  assign dmem58_io_pipeline_memwrite = cpu58_io_dmem_memwrite; // @[top.scala 424:17]
  assign dmem58_io_pipeline_maskmode = cpu58_io_dmem_maskmode; // @[top.scala 424:17]
  assign dmem58_io_pipeline_sext = cpu58_io_dmem_sext; // @[top.scala 424:17]
  assign dmem58_io_bus_response_valid = mem58_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem58_io_bus_response_bits_data = mem58_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu59_clock = clock;
  assign cpu59_reset = reset;
  assign cpu59_io_imem_instruction = imem59_io_pipeline_instruction; // @[top.scala 430:17]
  assign cpu59_io_dmem_readdata = dmem59_io_pipeline_readdata; // @[top.scala 431:17]
  assign mem59_clock = clock;
  assign mem59_reset = reset;
  assign mem59_io_imem_request_bits_address = imem59_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem59_io_dmem_request_valid = dmem59_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem59_io_dmem_request_bits_address = dmem59_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem59_io_dmem_request_bits_writedata = dmem59_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem59_io_dmem_request_bits_operation = dmem59_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem59_io_pipeline_address = cpu59_io_imem_address; // @[top.scala 430:17]
  assign imem59_io_bus_response_bits_data = mem59_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem59_clock = clock;
  assign dmem59_reset = reset;
  assign dmem59_io_pipeline_address = cpu59_io_dmem_address; // @[top.scala 431:17]
  assign dmem59_io_pipeline_valid = cpu59_io_dmem_valid; // @[top.scala 431:17]
  assign dmem59_io_pipeline_writedata = cpu59_io_dmem_writedata; // @[top.scala 431:17]
  assign dmem59_io_pipeline_memread = cpu59_io_dmem_memread; // @[top.scala 431:17]
  assign dmem59_io_pipeline_memwrite = cpu59_io_dmem_memwrite; // @[top.scala 431:17]
  assign dmem59_io_pipeline_maskmode = cpu59_io_dmem_maskmode; // @[top.scala 431:17]
  assign dmem59_io_pipeline_sext = cpu59_io_dmem_sext; // @[top.scala 431:17]
  assign dmem59_io_bus_response_valid = mem59_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem59_io_bus_response_bits_data = mem59_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu60_clock = clock;
  assign cpu60_reset = reset;
  assign cpu60_io_imem_instruction = imem60_io_pipeline_instruction; // @[top.scala 437:17]
  assign cpu60_io_dmem_readdata = dmem60_io_pipeline_readdata; // @[top.scala 438:17]
  assign mem60_clock = clock;
  assign mem60_reset = reset;
  assign mem60_io_imem_request_bits_address = imem60_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem60_io_dmem_request_valid = dmem60_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem60_io_dmem_request_bits_address = dmem60_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem60_io_dmem_request_bits_writedata = dmem60_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem60_io_dmem_request_bits_operation = dmem60_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem60_io_pipeline_address = cpu60_io_imem_address; // @[top.scala 437:17]
  assign imem60_io_bus_response_bits_data = mem60_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem60_clock = clock;
  assign dmem60_reset = reset;
  assign dmem60_io_pipeline_address = cpu60_io_dmem_address; // @[top.scala 438:17]
  assign dmem60_io_pipeline_valid = cpu60_io_dmem_valid; // @[top.scala 438:17]
  assign dmem60_io_pipeline_writedata = cpu60_io_dmem_writedata; // @[top.scala 438:17]
  assign dmem60_io_pipeline_memread = cpu60_io_dmem_memread; // @[top.scala 438:17]
  assign dmem60_io_pipeline_memwrite = cpu60_io_dmem_memwrite; // @[top.scala 438:17]
  assign dmem60_io_pipeline_maskmode = cpu60_io_dmem_maskmode; // @[top.scala 438:17]
  assign dmem60_io_pipeline_sext = cpu60_io_dmem_sext; // @[top.scala 438:17]
  assign dmem60_io_bus_response_valid = mem60_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem60_io_bus_response_bits_data = mem60_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu61_clock = clock;
  assign cpu61_reset = reset;
  assign cpu61_io_imem_instruction = imem61_io_pipeline_instruction; // @[top.scala 444:17]
  assign cpu61_io_dmem_readdata = dmem61_io_pipeline_readdata; // @[top.scala 445:17]
  assign mem61_clock = clock;
  assign mem61_reset = reset;
  assign mem61_io_imem_request_bits_address = imem61_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem61_io_dmem_request_valid = dmem61_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem61_io_dmem_request_bits_address = dmem61_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem61_io_dmem_request_bits_writedata = dmem61_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem61_io_dmem_request_bits_operation = dmem61_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem61_io_pipeline_address = cpu61_io_imem_address; // @[top.scala 444:17]
  assign imem61_io_bus_response_bits_data = mem61_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem61_clock = clock;
  assign dmem61_reset = reset;
  assign dmem61_io_pipeline_address = cpu61_io_dmem_address; // @[top.scala 445:17]
  assign dmem61_io_pipeline_valid = cpu61_io_dmem_valid; // @[top.scala 445:17]
  assign dmem61_io_pipeline_writedata = cpu61_io_dmem_writedata; // @[top.scala 445:17]
  assign dmem61_io_pipeline_memread = cpu61_io_dmem_memread; // @[top.scala 445:17]
  assign dmem61_io_pipeline_memwrite = cpu61_io_dmem_memwrite; // @[top.scala 445:17]
  assign dmem61_io_pipeline_maskmode = cpu61_io_dmem_maskmode; // @[top.scala 445:17]
  assign dmem61_io_pipeline_sext = cpu61_io_dmem_sext; // @[top.scala 445:17]
  assign dmem61_io_bus_response_valid = mem61_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem61_io_bus_response_bits_data = mem61_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu62_clock = clock;
  assign cpu62_reset = reset;
  assign cpu62_io_imem_instruction = imem62_io_pipeline_instruction; // @[top.scala 451:17]
  assign cpu62_io_dmem_readdata = dmem62_io_pipeline_readdata; // @[top.scala 452:17]
  assign mem62_clock = clock;
  assign mem62_reset = reset;
  assign mem62_io_imem_request_bits_address = imem62_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem62_io_dmem_request_valid = dmem62_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem62_io_dmem_request_bits_address = dmem62_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem62_io_dmem_request_bits_writedata = dmem62_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem62_io_dmem_request_bits_operation = dmem62_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem62_io_pipeline_address = cpu62_io_imem_address; // @[top.scala 451:17]
  assign imem62_io_bus_response_bits_data = mem62_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem62_clock = clock;
  assign dmem62_reset = reset;
  assign dmem62_io_pipeline_address = cpu62_io_dmem_address; // @[top.scala 452:17]
  assign dmem62_io_pipeline_valid = cpu62_io_dmem_valid; // @[top.scala 452:17]
  assign dmem62_io_pipeline_writedata = cpu62_io_dmem_writedata; // @[top.scala 452:17]
  assign dmem62_io_pipeline_memread = cpu62_io_dmem_memread; // @[top.scala 452:17]
  assign dmem62_io_pipeline_memwrite = cpu62_io_dmem_memwrite; // @[top.scala 452:17]
  assign dmem62_io_pipeline_maskmode = cpu62_io_dmem_maskmode; // @[top.scala 452:17]
  assign dmem62_io_pipeline_sext = cpu62_io_dmem_sext; // @[top.scala 452:17]
  assign dmem62_io_bus_response_valid = mem62_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem62_io_bus_response_bits_data = mem62_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu63_clock = clock;
  assign cpu63_reset = reset;
  assign cpu63_io_imem_instruction = imem63_io_pipeline_instruction; // @[top.scala 458:17]
  assign cpu63_io_dmem_readdata = dmem63_io_pipeline_readdata; // @[top.scala 459:17]
  assign mem63_clock = clock;
  assign mem63_reset = reset;
  assign mem63_io_imem_request_bits_address = imem63_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem63_io_dmem_request_valid = dmem63_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem63_io_dmem_request_bits_address = dmem63_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem63_io_dmem_request_bits_writedata = dmem63_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem63_io_dmem_request_bits_operation = dmem63_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem63_io_pipeline_address = cpu63_io_imem_address; // @[top.scala 458:17]
  assign imem63_io_bus_response_bits_data = mem63_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem63_clock = clock;
  assign dmem63_reset = reset;
  assign dmem63_io_pipeline_address = cpu63_io_dmem_address; // @[top.scala 459:17]
  assign dmem63_io_pipeline_valid = cpu63_io_dmem_valid; // @[top.scala 459:17]
  assign dmem63_io_pipeline_writedata = cpu63_io_dmem_writedata; // @[top.scala 459:17]
  assign dmem63_io_pipeline_memread = cpu63_io_dmem_memread; // @[top.scala 459:17]
  assign dmem63_io_pipeline_memwrite = cpu63_io_dmem_memwrite; // @[top.scala 459:17]
  assign dmem63_io_pipeline_maskmode = cpu63_io_dmem_maskmode; // @[top.scala 459:17]
  assign dmem63_io_pipeline_sext = cpu63_io_dmem_sext; // @[top.scala 459:17]
  assign dmem63_io_bus_response_valid = mem63_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem63_io_bus_response_bits_data = mem63_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu64_clock = clock;
  assign cpu64_reset = reset;
  assign cpu64_io_imem_instruction = imem64_io_pipeline_instruction; // @[top.scala 465:17]
  assign cpu64_io_dmem_readdata = dmem64_io_pipeline_readdata; // @[top.scala 466:17]
  assign mem64_clock = clock;
  assign mem64_reset = reset;
  assign mem64_io_imem_request_bits_address = imem64_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem64_io_dmem_request_valid = dmem64_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem64_io_dmem_request_bits_address = dmem64_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem64_io_dmem_request_bits_writedata = dmem64_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem64_io_dmem_request_bits_operation = dmem64_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem64_io_pipeline_address = cpu64_io_imem_address; // @[top.scala 465:17]
  assign imem64_io_bus_response_bits_data = mem64_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem64_clock = clock;
  assign dmem64_reset = reset;
  assign dmem64_io_pipeline_address = cpu64_io_dmem_address; // @[top.scala 466:17]
  assign dmem64_io_pipeline_valid = cpu64_io_dmem_valid; // @[top.scala 466:17]
  assign dmem64_io_pipeline_writedata = cpu64_io_dmem_writedata; // @[top.scala 466:17]
  assign dmem64_io_pipeline_memread = cpu64_io_dmem_memread; // @[top.scala 466:17]
  assign dmem64_io_pipeline_memwrite = cpu64_io_dmem_memwrite; // @[top.scala 466:17]
  assign dmem64_io_pipeline_maskmode = cpu64_io_dmem_maskmode; // @[top.scala 466:17]
  assign dmem64_io_pipeline_sext = cpu64_io_dmem_sext; // @[top.scala 466:17]
  assign dmem64_io_bus_response_valid = mem64_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem64_io_bus_response_bits_data = mem64_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu65_clock = clock;
  assign cpu65_reset = reset;
  assign cpu65_io_imem_instruction = imem65_io_pipeline_instruction; // @[top.scala 472:17]
  assign cpu65_io_dmem_readdata = dmem65_io_pipeline_readdata; // @[top.scala 473:17]
  assign mem65_clock = clock;
  assign mem65_reset = reset;
  assign mem65_io_imem_request_bits_address = imem65_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem65_io_dmem_request_valid = dmem65_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem65_io_dmem_request_bits_address = dmem65_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem65_io_dmem_request_bits_writedata = dmem65_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem65_io_dmem_request_bits_operation = dmem65_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem65_io_pipeline_address = cpu65_io_imem_address; // @[top.scala 472:17]
  assign imem65_io_bus_response_bits_data = mem65_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem65_clock = clock;
  assign dmem65_reset = reset;
  assign dmem65_io_pipeline_address = cpu65_io_dmem_address; // @[top.scala 473:17]
  assign dmem65_io_pipeline_valid = cpu65_io_dmem_valid; // @[top.scala 473:17]
  assign dmem65_io_pipeline_writedata = cpu65_io_dmem_writedata; // @[top.scala 473:17]
  assign dmem65_io_pipeline_memread = cpu65_io_dmem_memread; // @[top.scala 473:17]
  assign dmem65_io_pipeline_memwrite = cpu65_io_dmem_memwrite; // @[top.scala 473:17]
  assign dmem65_io_pipeline_maskmode = cpu65_io_dmem_maskmode; // @[top.scala 473:17]
  assign dmem65_io_pipeline_sext = cpu65_io_dmem_sext; // @[top.scala 473:17]
  assign dmem65_io_bus_response_valid = mem65_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem65_io_bus_response_bits_data = mem65_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu66_clock = clock;
  assign cpu66_reset = reset;
  assign cpu66_io_imem_instruction = imem66_io_pipeline_instruction; // @[top.scala 479:17]
  assign cpu66_io_dmem_readdata = dmem66_io_pipeline_readdata; // @[top.scala 480:17]
  assign mem66_clock = clock;
  assign mem66_reset = reset;
  assign mem66_io_imem_request_bits_address = imem66_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem66_io_dmem_request_valid = dmem66_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem66_io_dmem_request_bits_address = dmem66_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem66_io_dmem_request_bits_writedata = dmem66_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem66_io_dmem_request_bits_operation = dmem66_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem66_io_pipeline_address = cpu66_io_imem_address; // @[top.scala 479:17]
  assign imem66_io_bus_response_bits_data = mem66_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem66_clock = clock;
  assign dmem66_reset = reset;
  assign dmem66_io_pipeline_address = cpu66_io_dmem_address; // @[top.scala 480:17]
  assign dmem66_io_pipeline_valid = cpu66_io_dmem_valid; // @[top.scala 480:17]
  assign dmem66_io_pipeline_writedata = cpu66_io_dmem_writedata; // @[top.scala 480:17]
  assign dmem66_io_pipeline_memread = cpu66_io_dmem_memread; // @[top.scala 480:17]
  assign dmem66_io_pipeline_memwrite = cpu66_io_dmem_memwrite; // @[top.scala 480:17]
  assign dmem66_io_pipeline_maskmode = cpu66_io_dmem_maskmode; // @[top.scala 480:17]
  assign dmem66_io_pipeline_sext = cpu66_io_dmem_sext; // @[top.scala 480:17]
  assign dmem66_io_bus_response_valid = mem66_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem66_io_bus_response_bits_data = mem66_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu67_clock = clock;
  assign cpu67_reset = reset;
  assign cpu67_io_imem_instruction = imem67_io_pipeline_instruction; // @[top.scala 486:17]
  assign cpu67_io_dmem_readdata = dmem67_io_pipeline_readdata; // @[top.scala 487:17]
  assign mem67_clock = clock;
  assign mem67_reset = reset;
  assign mem67_io_imem_request_bits_address = imem67_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem67_io_dmem_request_valid = dmem67_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem67_io_dmem_request_bits_address = dmem67_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem67_io_dmem_request_bits_writedata = dmem67_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem67_io_dmem_request_bits_operation = dmem67_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem67_io_pipeline_address = cpu67_io_imem_address; // @[top.scala 486:17]
  assign imem67_io_bus_response_bits_data = mem67_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem67_clock = clock;
  assign dmem67_reset = reset;
  assign dmem67_io_pipeline_address = cpu67_io_dmem_address; // @[top.scala 487:17]
  assign dmem67_io_pipeline_valid = cpu67_io_dmem_valid; // @[top.scala 487:17]
  assign dmem67_io_pipeline_writedata = cpu67_io_dmem_writedata; // @[top.scala 487:17]
  assign dmem67_io_pipeline_memread = cpu67_io_dmem_memread; // @[top.scala 487:17]
  assign dmem67_io_pipeline_memwrite = cpu67_io_dmem_memwrite; // @[top.scala 487:17]
  assign dmem67_io_pipeline_maskmode = cpu67_io_dmem_maskmode; // @[top.scala 487:17]
  assign dmem67_io_pipeline_sext = cpu67_io_dmem_sext; // @[top.scala 487:17]
  assign dmem67_io_bus_response_valid = mem67_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem67_io_bus_response_bits_data = mem67_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu68_clock = clock;
  assign cpu68_reset = reset;
  assign cpu68_io_imem_instruction = imem68_io_pipeline_instruction; // @[top.scala 493:17]
  assign cpu68_io_dmem_readdata = dmem68_io_pipeline_readdata; // @[top.scala 494:17]
  assign mem68_clock = clock;
  assign mem68_reset = reset;
  assign mem68_io_imem_request_bits_address = imem68_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem68_io_dmem_request_valid = dmem68_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem68_io_dmem_request_bits_address = dmem68_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem68_io_dmem_request_bits_writedata = dmem68_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem68_io_dmem_request_bits_operation = dmem68_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem68_io_pipeline_address = cpu68_io_imem_address; // @[top.scala 493:17]
  assign imem68_io_bus_response_bits_data = mem68_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem68_clock = clock;
  assign dmem68_reset = reset;
  assign dmem68_io_pipeline_address = cpu68_io_dmem_address; // @[top.scala 494:17]
  assign dmem68_io_pipeline_valid = cpu68_io_dmem_valid; // @[top.scala 494:17]
  assign dmem68_io_pipeline_writedata = cpu68_io_dmem_writedata; // @[top.scala 494:17]
  assign dmem68_io_pipeline_memread = cpu68_io_dmem_memread; // @[top.scala 494:17]
  assign dmem68_io_pipeline_memwrite = cpu68_io_dmem_memwrite; // @[top.scala 494:17]
  assign dmem68_io_pipeline_maskmode = cpu68_io_dmem_maskmode; // @[top.scala 494:17]
  assign dmem68_io_pipeline_sext = cpu68_io_dmem_sext; // @[top.scala 494:17]
  assign dmem68_io_bus_response_valid = mem68_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem68_io_bus_response_bits_data = mem68_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu69_clock = clock;
  assign cpu69_reset = reset;
  assign cpu69_io_imem_instruction = imem69_io_pipeline_instruction; // @[top.scala 500:17]
  assign cpu69_io_dmem_readdata = dmem69_io_pipeline_readdata; // @[top.scala 501:17]
  assign mem69_clock = clock;
  assign mem69_reset = reset;
  assign mem69_io_imem_request_bits_address = imem69_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem69_io_dmem_request_valid = dmem69_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem69_io_dmem_request_bits_address = dmem69_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem69_io_dmem_request_bits_writedata = dmem69_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem69_io_dmem_request_bits_operation = dmem69_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem69_io_pipeline_address = cpu69_io_imem_address; // @[top.scala 500:17]
  assign imem69_io_bus_response_bits_data = mem69_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem69_clock = clock;
  assign dmem69_reset = reset;
  assign dmem69_io_pipeline_address = cpu69_io_dmem_address; // @[top.scala 501:17]
  assign dmem69_io_pipeline_valid = cpu69_io_dmem_valid; // @[top.scala 501:17]
  assign dmem69_io_pipeline_writedata = cpu69_io_dmem_writedata; // @[top.scala 501:17]
  assign dmem69_io_pipeline_memread = cpu69_io_dmem_memread; // @[top.scala 501:17]
  assign dmem69_io_pipeline_memwrite = cpu69_io_dmem_memwrite; // @[top.scala 501:17]
  assign dmem69_io_pipeline_maskmode = cpu69_io_dmem_maskmode; // @[top.scala 501:17]
  assign dmem69_io_pipeline_sext = cpu69_io_dmem_sext; // @[top.scala 501:17]
  assign dmem69_io_bus_response_valid = mem69_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem69_io_bus_response_bits_data = mem69_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu70_clock = clock;
  assign cpu70_reset = reset;
  assign cpu70_io_imem_instruction = imem70_io_pipeline_instruction; // @[top.scala 507:17]
  assign cpu70_io_dmem_readdata = dmem70_io_pipeline_readdata; // @[top.scala 508:17]
  assign mem70_clock = clock;
  assign mem70_reset = reset;
  assign mem70_io_imem_request_bits_address = imem70_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem70_io_dmem_request_valid = dmem70_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem70_io_dmem_request_bits_address = dmem70_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem70_io_dmem_request_bits_writedata = dmem70_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem70_io_dmem_request_bits_operation = dmem70_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem70_io_pipeline_address = cpu70_io_imem_address; // @[top.scala 507:17]
  assign imem70_io_bus_response_bits_data = mem70_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem70_clock = clock;
  assign dmem70_reset = reset;
  assign dmem70_io_pipeline_address = cpu70_io_dmem_address; // @[top.scala 508:17]
  assign dmem70_io_pipeline_valid = cpu70_io_dmem_valid; // @[top.scala 508:17]
  assign dmem70_io_pipeline_writedata = cpu70_io_dmem_writedata; // @[top.scala 508:17]
  assign dmem70_io_pipeline_memread = cpu70_io_dmem_memread; // @[top.scala 508:17]
  assign dmem70_io_pipeline_memwrite = cpu70_io_dmem_memwrite; // @[top.scala 508:17]
  assign dmem70_io_pipeline_maskmode = cpu70_io_dmem_maskmode; // @[top.scala 508:17]
  assign dmem70_io_pipeline_sext = cpu70_io_dmem_sext; // @[top.scala 508:17]
  assign dmem70_io_bus_response_valid = mem70_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem70_io_bus_response_bits_data = mem70_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu71_clock = clock;
  assign cpu71_reset = reset;
  assign cpu71_io_imem_instruction = imem71_io_pipeline_instruction; // @[top.scala 514:17]
  assign cpu71_io_dmem_readdata = dmem71_io_pipeline_readdata; // @[top.scala 515:17]
  assign mem71_clock = clock;
  assign mem71_reset = reset;
  assign mem71_io_imem_request_bits_address = imem71_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem71_io_dmem_request_valid = dmem71_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem71_io_dmem_request_bits_address = dmem71_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem71_io_dmem_request_bits_writedata = dmem71_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem71_io_dmem_request_bits_operation = dmem71_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem71_io_pipeline_address = cpu71_io_imem_address; // @[top.scala 514:17]
  assign imem71_io_bus_response_bits_data = mem71_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem71_clock = clock;
  assign dmem71_reset = reset;
  assign dmem71_io_pipeline_address = cpu71_io_dmem_address; // @[top.scala 515:17]
  assign dmem71_io_pipeline_valid = cpu71_io_dmem_valid; // @[top.scala 515:17]
  assign dmem71_io_pipeline_writedata = cpu71_io_dmem_writedata; // @[top.scala 515:17]
  assign dmem71_io_pipeline_memread = cpu71_io_dmem_memread; // @[top.scala 515:17]
  assign dmem71_io_pipeline_memwrite = cpu71_io_dmem_memwrite; // @[top.scala 515:17]
  assign dmem71_io_pipeline_maskmode = cpu71_io_dmem_maskmode; // @[top.scala 515:17]
  assign dmem71_io_pipeline_sext = cpu71_io_dmem_sext; // @[top.scala 515:17]
  assign dmem71_io_bus_response_valid = mem71_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem71_io_bus_response_bits_data = mem71_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu72_clock = clock;
  assign cpu72_reset = reset;
  assign cpu72_io_imem_instruction = imem72_io_pipeline_instruction; // @[top.scala 521:17]
  assign cpu72_io_dmem_readdata = dmem72_io_pipeline_readdata; // @[top.scala 522:17]
  assign mem72_clock = clock;
  assign mem72_reset = reset;
  assign mem72_io_imem_request_bits_address = imem72_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem72_io_dmem_request_valid = dmem72_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem72_io_dmem_request_bits_address = dmem72_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem72_io_dmem_request_bits_writedata = dmem72_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem72_io_dmem_request_bits_operation = dmem72_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem72_io_pipeline_address = cpu72_io_imem_address; // @[top.scala 521:17]
  assign imem72_io_bus_response_bits_data = mem72_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem72_clock = clock;
  assign dmem72_reset = reset;
  assign dmem72_io_pipeline_address = cpu72_io_dmem_address; // @[top.scala 522:17]
  assign dmem72_io_pipeline_valid = cpu72_io_dmem_valid; // @[top.scala 522:17]
  assign dmem72_io_pipeline_writedata = cpu72_io_dmem_writedata; // @[top.scala 522:17]
  assign dmem72_io_pipeline_memread = cpu72_io_dmem_memread; // @[top.scala 522:17]
  assign dmem72_io_pipeline_memwrite = cpu72_io_dmem_memwrite; // @[top.scala 522:17]
  assign dmem72_io_pipeline_maskmode = cpu72_io_dmem_maskmode; // @[top.scala 522:17]
  assign dmem72_io_pipeline_sext = cpu72_io_dmem_sext; // @[top.scala 522:17]
  assign dmem72_io_bus_response_valid = mem72_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem72_io_bus_response_bits_data = mem72_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu73_clock = clock;
  assign cpu73_reset = reset;
  assign cpu73_io_imem_instruction = imem73_io_pipeline_instruction; // @[top.scala 528:17]
  assign cpu73_io_dmem_readdata = dmem73_io_pipeline_readdata; // @[top.scala 529:17]
  assign mem73_clock = clock;
  assign mem73_reset = reset;
  assign mem73_io_imem_request_bits_address = imem73_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem73_io_dmem_request_valid = dmem73_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem73_io_dmem_request_bits_address = dmem73_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem73_io_dmem_request_bits_writedata = dmem73_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem73_io_dmem_request_bits_operation = dmem73_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem73_io_pipeline_address = cpu73_io_imem_address; // @[top.scala 528:17]
  assign imem73_io_bus_response_bits_data = mem73_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem73_clock = clock;
  assign dmem73_reset = reset;
  assign dmem73_io_pipeline_address = cpu73_io_dmem_address; // @[top.scala 529:17]
  assign dmem73_io_pipeline_valid = cpu73_io_dmem_valid; // @[top.scala 529:17]
  assign dmem73_io_pipeline_writedata = cpu73_io_dmem_writedata; // @[top.scala 529:17]
  assign dmem73_io_pipeline_memread = cpu73_io_dmem_memread; // @[top.scala 529:17]
  assign dmem73_io_pipeline_memwrite = cpu73_io_dmem_memwrite; // @[top.scala 529:17]
  assign dmem73_io_pipeline_maskmode = cpu73_io_dmem_maskmode; // @[top.scala 529:17]
  assign dmem73_io_pipeline_sext = cpu73_io_dmem_sext; // @[top.scala 529:17]
  assign dmem73_io_bus_response_valid = mem73_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem73_io_bus_response_bits_data = mem73_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu74_clock = clock;
  assign cpu74_reset = reset;
  assign cpu74_io_imem_instruction = imem74_io_pipeline_instruction; // @[top.scala 535:17]
  assign cpu74_io_dmem_readdata = dmem74_io_pipeline_readdata; // @[top.scala 536:17]
  assign mem74_clock = clock;
  assign mem74_reset = reset;
  assign mem74_io_imem_request_bits_address = imem74_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem74_io_dmem_request_valid = dmem74_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem74_io_dmem_request_bits_address = dmem74_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem74_io_dmem_request_bits_writedata = dmem74_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem74_io_dmem_request_bits_operation = dmem74_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem74_io_pipeline_address = cpu74_io_imem_address; // @[top.scala 535:17]
  assign imem74_io_bus_response_bits_data = mem74_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem74_clock = clock;
  assign dmem74_reset = reset;
  assign dmem74_io_pipeline_address = cpu74_io_dmem_address; // @[top.scala 536:17]
  assign dmem74_io_pipeline_valid = cpu74_io_dmem_valid; // @[top.scala 536:17]
  assign dmem74_io_pipeline_writedata = cpu74_io_dmem_writedata; // @[top.scala 536:17]
  assign dmem74_io_pipeline_memread = cpu74_io_dmem_memread; // @[top.scala 536:17]
  assign dmem74_io_pipeline_memwrite = cpu74_io_dmem_memwrite; // @[top.scala 536:17]
  assign dmem74_io_pipeline_maskmode = cpu74_io_dmem_maskmode; // @[top.scala 536:17]
  assign dmem74_io_pipeline_sext = cpu74_io_dmem_sext; // @[top.scala 536:17]
  assign dmem74_io_bus_response_valid = mem74_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem74_io_bus_response_bits_data = mem74_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu75_clock = clock;
  assign cpu75_reset = reset;
  assign cpu75_io_imem_instruction = imem75_io_pipeline_instruction; // @[top.scala 542:17]
  assign cpu75_io_dmem_readdata = dmem75_io_pipeline_readdata; // @[top.scala 543:17]
  assign mem75_clock = clock;
  assign mem75_reset = reset;
  assign mem75_io_imem_request_bits_address = imem75_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem75_io_dmem_request_valid = dmem75_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem75_io_dmem_request_bits_address = dmem75_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem75_io_dmem_request_bits_writedata = dmem75_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem75_io_dmem_request_bits_operation = dmem75_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem75_io_pipeline_address = cpu75_io_imem_address; // @[top.scala 542:17]
  assign imem75_io_bus_response_bits_data = mem75_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem75_clock = clock;
  assign dmem75_reset = reset;
  assign dmem75_io_pipeline_address = cpu75_io_dmem_address; // @[top.scala 543:17]
  assign dmem75_io_pipeline_valid = cpu75_io_dmem_valid; // @[top.scala 543:17]
  assign dmem75_io_pipeline_writedata = cpu75_io_dmem_writedata; // @[top.scala 543:17]
  assign dmem75_io_pipeline_memread = cpu75_io_dmem_memread; // @[top.scala 543:17]
  assign dmem75_io_pipeline_memwrite = cpu75_io_dmem_memwrite; // @[top.scala 543:17]
  assign dmem75_io_pipeline_maskmode = cpu75_io_dmem_maskmode; // @[top.scala 543:17]
  assign dmem75_io_pipeline_sext = cpu75_io_dmem_sext; // @[top.scala 543:17]
  assign dmem75_io_bus_response_valid = mem75_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem75_io_bus_response_bits_data = mem75_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu76_clock = clock;
  assign cpu76_reset = reset;
  assign cpu76_io_imem_instruction = imem76_io_pipeline_instruction; // @[top.scala 549:17]
  assign cpu76_io_dmem_readdata = dmem76_io_pipeline_readdata; // @[top.scala 550:17]
  assign mem76_clock = clock;
  assign mem76_reset = reset;
  assign mem76_io_imem_request_bits_address = imem76_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem76_io_dmem_request_valid = dmem76_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem76_io_dmem_request_bits_address = dmem76_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem76_io_dmem_request_bits_writedata = dmem76_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem76_io_dmem_request_bits_operation = dmem76_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem76_io_pipeline_address = cpu76_io_imem_address; // @[top.scala 549:17]
  assign imem76_io_bus_response_bits_data = mem76_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem76_clock = clock;
  assign dmem76_reset = reset;
  assign dmem76_io_pipeline_address = cpu76_io_dmem_address; // @[top.scala 550:17]
  assign dmem76_io_pipeline_valid = cpu76_io_dmem_valid; // @[top.scala 550:17]
  assign dmem76_io_pipeline_writedata = cpu76_io_dmem_writedata; // @[top.scala 550:17]
  assign dmem76_io_pipeline_memread = cpu76_io_dmem_memread; // @[top.scala 550:17]
  assign dmem76_io_pipeline_memwrite = cpu76_io_dmem_memwrite; // @[top.scala 550:17]
  assign dmem76_io_pipeline_maskmode = cpu76_io_dmem_maskmode; // @[top.scala 550:17]
  assign dmem76_io_pipeline_sext = cpu76_io_dmem_sext; // @[top.scala 550:17]
  assign dmem76_io_bus_response_valid = mem76_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem76_io_bus_response_bits_data = mem76_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu77_clock = clock;
  assign cpu77_reset = reset;
  assign cpu77_io_imem_instruction = imem77_io_pipeline_instruction; // @[top.scala 556:17]
  assign cpu77_io_dmem_readdata = dmem77_io_pipeline_readdata; // @[top.scala 557:17]
  assign mem77_clock = clock;
  assign mem77_reset = reset;
  assign mem77_io_imem_request_bits_address = imem77_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem77_io_dmem_request_valid = dmem77_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem77_io_dmem_request_bits_address = dmem77_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem77_io_dmem_request_bits_writedata = dmem77_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem77_io_dmem_request_bits_operation = dmem77_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem77_io_pipeline_address = cpu77_io_imem_address; // @[top.scala 556:17]
  assign imem77_io_bus_response_bits_data = mem77_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem77_clock = clock;
  assign dmem77_reset = reset;
  assign dmem77_io_pipeline_address = cpu77_io_dmem_address; // @[top.scala 557:17]
  assign dmem77_io_pipeline_valid = cpu77_io_dmem_valid; // @[top.scala 557:17]
  assign dmem77_io_pipeline_writedata = cpu77_io_dmem_writedata; // @[top.scala 557:17]
  assign dmem77_io_pipeline_memread = cpu77_io_dmem_memread; // @[top.scala 557:17]
  assign dmem77_io_pipeline_memwrite = cpu77_io_dmem_memwrite; // @[top.scala 557:17]
  assign dmem77_io_pipeline_maskmode = cpu77_io_dmem_maskmode; // @[top.scala 557:17]
  assign dmem77_io_pipeline_sext = cpu77_io_dmem_sext; // @[top.scala 557:17]
  assign dmem77_io_bus_response_valid = mem77_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem77_io_bus_response_bits_data = mem77_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu78_clock = clock;
  assign cpu78_reset = reset;
  assign cpu78_io_imem_instruction = imem78_io_pipeline_instruction; // @[top.scala 563:17]
  assign cpu78_io_dmem_readdata = dmem78_io_pipeline_readdata; // @[top.scala 564:17]
  assign mem78_clock = clock;
  assign mem78_reset = reset;
  assign mem78_io_imem_request_bits_address = imem78_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem78_io_dmem_request_valid = dmem78_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem78_io_dmem_request_bits_address = dmem78_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem78_io_dmem_request_bits_writedata = dmem78_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem78_io_dmem_request_bits_operation = dmem78_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem78_io_pipeline_address = cpu78_io_imem_address; // @[top.scala 563:17]
  assign imem78_io_bus_response_bits_data = mem78_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem78_clock = clock;
  assign dmem78_reset = reset;
  assign dmem78_io_pipeline_address = cpu78_io_dmem_address; // @[top.scala 564:17]
  assign dmem78_io_pipeline_valid = cpu78_io_dmem_valid; // @[top.scala 564:17]
  assign dmem78_io_pipeline_writedata = cpu78_io_dmem_writedata; // @[top.scala 564:17]
  assign dmem78_io_pipeline_memread = cpu78_io_dmem_memread; // @[top.scala 564:17]
  assign dmem78_io_pipeline_memwrite = cpu78_io_dmem_memwrite; // @[top.scala 564:17]
  assign dmem78_io_pipeline_maskmode = cpu78_io_dmem_maskmode; // @[top.scala 564:17]
  assign dmem78_io_pipeline_sext = cpu78_io_dmem_sext; // @[top.scala 564:17]
  assign dmem78_io_bus_response_valid = mem78_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem78_io_bus_response_bits_data = mem78_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu79_clock = clock;
  assign cpu79_reset = reset;
  assign cpu79_io_imem_instruction = imem79_io_pipeline_instruction; // @[top.scala 570:17]
  assign cpu79_io_dmem_readdata = dmem79_io_pipeline_readdata; // @[top.scala 571:17]
  assign mem79_clock = clock;
  assign mem79_reset = reset;
  assign mem79_io_imem_request_bits_address = imem79_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem79_io_dmem_request_valid = dmem79_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem79_io_dmem_request_bits_address = dmem79_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem79_io_dmem_request_bits_writedata = dmem79_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem79_io_dmem_request_bits_operation = dmem79_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem79_io_pipeline_address = cpu79_io_imem_address; // @[top.scala 570:17]
  assign imem79_io_bus_response_bits_data = mem79_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem79_clock = clock;
  assign dmem79_reset = reset;
  assign dmem79_io_pipeline_address = cpu79_io_dmem_address; // @[top.scala 571:17]
  assign dmem79_io_pipeline_valid = cpu79_io_dmem_valid; // @[top.scala 571:17]
  assign dmem79_io_pipeline_writedata = cpu79_io_dmem_writedata; // @[top.scala 571:17]
  assign dmem79_io_pipeline_memread = cpu79_io_dmem_memread; // @[top.scala 571:17]
  assign dmem79_io_pipeline_memwrite = cpu79_io_dmem_memwrite; // @[top.scala 571:17]
  assign dmem79_io_pipeline_maskmode = cpu79_io_dmem_maskmode; // @[top.scala 571:17]
  assign dmem79_io_pipeline_sext = cpu79_io_dmem_sext; // @[top.scala 571:17]
  assign dmem79_io_bus_response_valid = mem79_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem79_io_bus_response_bits_data = mem79_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu80_clock = clock;
  assign cpu80_reset = reset;
  assign cpu80_io_imem_instruction = imem80_io_pipeline_instruction; // @[top.scala 577:17]
  assign cpu80_io_dmem_readdata = dmem80_io_pipeline_readdata; // @[top.scala 578:17]
  assign mem80_clock = clock;
  assign mem80_reset = reset;
  assign mem80_io_imem_request_bits_address = imem80_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem80_io_dmem_request_valid = dmem80_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem80_io_dmem_request_bits_address = dmem80_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem80_io_dmem_request_bits_writedata = dmem80_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem80_io_dmem_request_bits_operation = dmem80_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem80_io_pipeline_address = cpu80_io_imem_address; // @[top.scala 577:17]
  assign imem80_io_bus_response_bits_data = mem80_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem80_clock = clock;
  assign dmem80_reset = reset;
  assign dmem80_io_pipeline_address = cpu80_io_dmem_address; // @[top.scala 578:17]
  assign dmem80_io_pipeline_valid = cpu80_io_dmem_valid; // @[top.scala 578:17]
  assign dmem80_io_pipeline_writedata = cpu80_io_dmem_writedata; // @[top.scala 578:17]
  assign dmem80_io_pipeline_memread = cpu80_io_dmem_memread; // @[top.scala 578:17]
  assign dmem80_io_pipeline_memwrite = cpu80_io_dmem_memwrite; // @[top.scala 578:17]
  assign dmem80_io_pipeline_maskmode = cpu80_io_dmem_maskmode; // @[top.scala 578:17]
  assign dmem80_io_pipeline_sext = cpu80_io_dmem_sext; // @[top.scala 578:17]
  assign dmem80_io_bus_response_valid = mem80_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem80_io_bus_response_bits_data = mem80_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu81_clock = clock;
  assign cpu81_reset = reset;
  assign cpu81_io_imem_instruction = imem81_io_pipeline_instruction; // @[top.scala 584:17]
  assign cpu81_io_dmem_readdata = dmem81_io_pipeline_readdata; // @[top.scala 585:17]
  assign mem81_clock = clock;
  assign mem81_reset = reset;
  assign mem81_io_imem_request_bits_address = imem81_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem81_io_dmem_request_valid = dmem81_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem81_io_dmem_request_bits_address = dmem81_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem81_io_dmem_request_bits_writedata = dmem81_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem81_io_dmem_request_bits_operation = dmem81_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem81_io_pipeline_address = cpu81_io_imem_address; // @[top.scala 584:17]
  assign imem81_io_bus_response_bits_data = mem81_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem81_clock = clock;
  assign dmem81_reset = reset;
  assign dmem81_io_pipeline_address = cpu81_io_dmem_address; // @[top.scala 585:17]
  assign dmem81_io_pipeline_valid = cpu81_io_dmem_valid; // @[top.scala 585:17]
  assign dmem81_io_pipeline_writedata = cpu81_io_dmem_writedata; // @[top.scala 585:17]
  assign dmem81_io_pipeline_memread = cpu81_io_dmem_memread; // @[top.scala 585:17]
  assign dmem81_io_pipeline_memwrite = cpu81_io_dmem_memwrite; // @[top.scala 585:17]
  assign dmem81_io_pipeline_maskmode = cpu81_io_dmem_maskmode; // @[top.scala 585:17]
  assign dmem81_io_pipeline_sext = cpu81_io_dmem_sext; // @[top.scala 585:17]
  assign dmem81_io_bus_response_valid = mem81_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem81_io_bus_response_bits_data = mem81_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu82_clock = clock;
  assign cpu82_reset = reset;
  assign cpu82_io_imem_instruction = imem82_io_pipeline_instruction; // @[top.scala 591:17]
  assign cpu82_io_dmem_readdata = dmem82_io_pipeline_readdata; // @[top.scala 592:17]
  assign mem82_clock = clock;
  assign mem82_reset = reset;
  assign mem82_io_imem_request_bits_address = imem82_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem82_io_dmem_request_valid = dmem82_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem82_io_dmem_request_bits_address = dmem82_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem82_io_dmem_request_bits_writedata = dmem82_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem82_io_dmem_request_bits_operation = dmem82_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem82_io_pipeline_address = cpu82_io_imem_address; // @[top.scala 591:17]
  assign imem82_io_bus_response_bits_data = mem82_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem82_clock = clock;
  assign dmem82_reset = reset;
  assign dmem82_io_pipeline_address = cpu82_io_dmem_address; // @[top.scala 592:17]
  assign dmem82_io_pipeline_valid = cpu82_io_dmem_valid; // @[top.scala 592:17]
  assign dmem82_io_pipeline_writedata = cpu82_io_dmem_writedata; // @[top.scala 592:17]
  assign dmem82_io_pipeline_memread = cpu82_io_dmem_memread; // @[top.scala 592:17]
  assign dmem82_io_pipeline_memwrite = cpu82_io_dmem_memwrite; // @[top.scala 592:17]
  assign dmem82_io_pipeline_maskmode = cpu82_io_dmem_maskmode; // @[top.scala 592:17]
  assign dmem82_io_pipeline_sext = cpu82_io_dmem_sext; // @[top.scala 592:17]
  assign dmem82_io_bus_response_valid = mem82_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem82_io_bus_response_bits_data = mem82_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu83_clock = clock;
  assign cpu83_reset = reset;
  assign cpu83_io_imem_instruction = imem83_io_pipeline_instruction; // @[top.scala 598:17]
  assign cpu83_io_dmem_readdata = dmem83_io_pipeline_readdata; // @[top.scala 599:17]
  assign mem83_clock = clock;
  assign mem83_reset = reset;
  assign mem83_io_imem_request_bits_address = imem83_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem83_io_dmem_request_valid = dmem83_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem83_io_dmem_request_bits_address = dmem83_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem83_io_dmem_request_bits_writedata = dmem83_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem83_io_dmem_request_bits_operation = dmem83_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem83_io_pipeline_address = cpu83_io_imem_address; // @[top.scala 598:17]
  assign imem83_io_bus_response_bits_data = mem83_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem83_clock = clock;
  assign dmem83_reset = reset;
  assign dmem83_io_pipeline_address = cpu83_io_dmem_address; // @[top.scala 599:17]
  assign dmem83_io_pipeline_valid = cpu83_io_dmem_valid; // @[top.scala 599:17]
  assign dmem83_io_pipeline_writedata = cpu83_io_dmem_writedata; // @[top.scala 599:17]
  assign dmem83_io_pipeline_memread = cpu83_io_dmem_memread; // @[top.scala 599:17]
  assign dmem83_io_pipeline_memwrite = cpu83_io_dmem_memwrite; // @[top.scala 599:17]
  assign dmem83_io_pipeline_maskmode = cpu83_io_dmem_maskmode; // @[top.scala 599:17]
  assign dmem83_io_pipeline_sext = cpu83_io_dmem_sext; // @[top.scala 599:17]
  assign dmem83_io_bus_response_valid = mem83_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem83_io_bus_response_bits_data = mem83_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu84_clock = clock;
  assign cpu84_reset = reset;
  assign cpu84_io_imem_instruction = imem84_io_pipeline_instruction; // @[top.scala 605:17]
  assign cpu84_io_dmem_readdata = dmem84_io_pipeline_readdata; // @[top.scala 606:17]
  assign mem84_clock = clock;
  assign mem84_reset = reset;
  assign mem84_io_imem_request_bits_address = imem84_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem84_io_dmem_request_valid = dmem84_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem84_io_dmem_request_bits_address = dmem84_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem84_io_dmem_request_bits_writedata = dmem84_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem84_io_dmem_request_bits_operation = dmem84_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem84_io_pipeline_address = cpu84_io_imem_address; // @[top.scala 605:17]
  assign imem84_io_bus_response_bits_data = mem84_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem84_clock = clock;
  assign dmem84_reset = reset;
  assign dmem84_io_pipeline_address = cpu84_io_dmem_address; // @[top.scala 606:17]
  assign dmem84_io_pipeline_valid = cpu84_io_dmem_valid; // @[top.scala 606:17]
  assign dmem84_io_pipeline_writedata = cpu84_io_dmem_writedata; // @[top.scala 606:17]
  assign dmem84_io_pipeline_memread = cpu84_io_dmem_memread; // @[top.scala 606:17]
  assign dmem84_io_pipeline_memwrite = cpu84_io_dmem_memwrite; // @[top.scala 606:17]
  assign dmem84_io_pipeline_maskmode = cpu84_io_dmem_maskmode; // @[top.scala 606:17]
  assign dmem84_io_pipeline_sext = cpu84_io_dmem_sext; // @[top.scala 606:17]
  assign dmem84_io_bus_response_valid = mem84_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem84_io_bus_response_bits_data = mem84_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu85_clock = clock;
  assign cpu85_reset = reset;
  assign cpu85_io_imem_instruction = imem85_io_pipeline_instruction; // @[top.scala 612:17]
  assign cpu85_io_dmem_readdata = dmem85_io_pipeline_readdata; // @[top.scala 613:17]
  assign mem85_clock = clock;
  assign mem85_reset = reset;
  assign mem85_io_imem_request_bits_address = imem85_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem85_io_dmem_request_valid = dmem85_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem85_io_dmem_request_bits_address = dmem85_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem85_io_dmem_request_bits_writedata = dmem85_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem85_io_dmem_request_bits_operation = dmem85_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem85_io_pipeline_address = cpu85_io_imem_address; // @[top.scala 612:17]
  assign imem85_io_bus_response_bits_data = mem85_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem85_clock = clock;
  assign dmem85_reset = reset;
  assign dmem85_io_pipeline_address = cpu85_io_dmem_address; // @[top.scala 613:17]
  assign dmem85_io_pipeline_valid = cpu85_io_dmem_valid; // @[top.scala 613:17]
  assign dmem85_io_pipeline_writedata = cpu85_io_dmem_writedata; // @[top.scala 613:17]
  assign dmem85_io_pipeline_memread = cpu85_io_dmem_memread; // @[top.scala 613:17]
  assign dmem85_io_pipeline_memwrite = cpu85_io_dmem_memwrite; // @[top.scala 613:17]
  assign dmem85_io_pipeline_maskmode = cpu85_io_dmem_maskmode; // @[top.scala 613:17]
  assign dmem85_io_pipeline_sext = cpu85_io_dmem_sext; // @[top.scala 613:17]
  assign dmem85_io_bus_response_valid = mem85_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem85_io_bus_response_bits_data = mem85_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu86_clock = clock;
  assign cpu86_reset = reset;
  assign cpu86_io_imem_instruction = imem86_io_pipeline_instruction; // @[top.scala 619:17]
  assign cpu86_io_dmem_readdata = dmem86_io_pipeline_readdata; // @[top.scala 620:17]
  assign mem86_clock = clock;
  assign mem86_reset = reset;
  assign mem86_io_imem_request_bits_address = imem86_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem86_io_dmem_request_valid = dmem86_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem86_io_dmem_request_bits_address = dmem86_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem86_io_dmem_request_bits_writedata = dmem86_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem86_io_dmem_request_bits_operation = dmem86_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem86_io_pipeline_address = cpu86_io_imem_address; // @[top.scala 619:17]
  assign imem86_io_bus_response_bits_data = mem86_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem86_clock = clock;
  assign dmem86_reset = reset;
  assign dmem86_io_pipeline_address = cpu86_io_dmem_address; // @[top.scala 620:17]
  assign dmem86_io_pipeline_valid = cpu86_io_dmem_valid; // @[top.scala 620:17]
  assign dmem86_io_pipeline_writedata = cpu86_io_dmem_writedata; // @[top.scala 620:17]
  assign dmem86_io_pipeline_memread = cpu86_io_dmem_memread; // @[top.scala 620:17]
  assign dmem86_io_pipeline_memwrite = cpu86_io_dmem_memwrite; // @[top.scala 620:17]
  assign dmem86_io_pipeline_maskmode = cpu86_io_dmem_maskmode; // @[top.scala 620:17]
  assign dmem86_io_pipeline_sext = cpu86_io_dmem_sext; // @[top.scala 620:17]
  assign dmem86_io_bus_response_valid = mem86_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem86_io_bus_response_bits_data = mem86_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu87_clock = clock;
  assign cpu87_reset = reset;
  assign cpu87_io_imem_instruction = imem87_io_pipeline_instruction; // @[top.scala 626:17]
  assign cpu87_io_dmem_readdata = dmem87_io_pipeline_readdata; // @[top.scala 627:17]
  assign mem87_clock = clock;
  assign mem87_reset = reset;
  assign mem87_io_imem_request_bits_address = imem87_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem87_io_dmem_request_valid = dmem87_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem87_io_dmem_request_bits_address = dmem87_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem87_io_dmem_request_bits_writedata = dmem87_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem87_io_dmem_request_bits_operation = dmem87_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem87_io_pipeline_address = cpu87_io_imem_address; // @[top.scala 626:17]
  assign imem87_io_bus_response_bits_data = mem87_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem87_clock = clock;
  assign dmem87_reset = reset;
  assign dmem87_io_pipeline_address = cpu87_io_dmem_address; // @[top.scala 627:17]
  assign dmem87_io_pipeline_valid = cpu87_io_dmem_valid; // @[top.scala 627:17]
  assign dmem87_io_pipeline_writedata = cpu87_io_dmem_writedata; // @[top.scala 627:17]
  assign dmem87_io_pipeline_memread = cpu87_io_dmem_memread; // @[top.scala 627:17]
  assign dmem87_io_pipeline_memwrite = cpu87_io_dmem_memwrite; // @[top.scala 627:17]
  assign dmem87_io_pipeline_maskmode = cpu87_io_dmem_maskmode; // @[top.scala 627:17]
  assign dmem87_io_pipeline_sext = cpu87_io_dmem_sext; // @[top.scala 627:17]
  assign dmem87_io_bus_response_valid = mem87_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem87_io_bus_response_bits_data = mem87_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu88_clock = clock;
  assign cpu88_reset = reset;
  assign cpu88_io_imem_instruction = imem88_io_pipeline_instruction; // @[top.scala 633:17]
  assign cpu88_io_dmem_readdata = dmem88_io_pipeline_readdata; // @[top.scala 634:17]
  assign mem88_clock = clock;
  assign mem88_reset = reset;
  assign mem88_io_imem_request_bits_address = imem88_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem88_io_dmem_request_valid = dmem88_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem88_io_dmem_request_bits_address = dmem88_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem88_io_dmem_request_bits_writedata = dmem88_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem88_io_dmem_request_bits_operation = dmem88_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem88_io_pipeline_address = cpu88_io_imem_address; // @[top.scala 633:17]
  assign imem88_io_bus_response_bits_data = mem88_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem88_clock = clock;
  assign dmem88_reset = reset;
  assign dmem88_io_pipeline_address = cpu88_io_dmem_address; // @[top.scala 634:17]
  assign dmem88_io_pipeline_valid = cpu88_io_dmem_valid; // @[top.scala 634:17]
  assign dmem88_io_pipeline_writedata = cpu88_io_dmem_writedata; // @[top.scala 634:17]
  assign dmem88_io_pipeline_memread = cpu88_io_dmem_memread; // @[top.scala 634:17]
  assign dmem88_io_pipeline_memwrite = cpu88_io_dmem_memwrite; // @[top.scala 634:17]
  assign dmem88_io_pipeline_maskmode = cpu88_io_dmem_maskmode; // @[top.scala 634:17]
  assign dmem88_io_pipeline_sext = cpu88_io_dmem_sext; // @[top.scala 634:17]
  assign dmem88_io_bus_response_valid = mem88_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem88_io_bus_response_bits_data = mem88_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu89_clock = clock;
  assign cpu89_reset = reset;
  assign cpu89_io_imem_instruction = imem89_io_pipeline_instruction; // @[top.scala 640:17]
  assign cpu89_io_dmem_readdata = dmem89_io_pipeline_readdata; // @[top.scala 641:17]
  assign mem89_clock = clock;
  assign mem89_reset = reset;
  assign mem89_io_imem_request_bits_address = imem89_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem89_io_dmem_request_valid = dmem89_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem89_io_dmem_request_bits_address = dmem89_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem89_io_dmem_request_bits_writedata = dmem89_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem89_io_dmem_request_bits_operation = dmem89_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem89_io_pipeline_address = cpu89_io_imem_address; // @[top.scala 640:17]
  assign imem89_io_bus_response_bits_data = mem89_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem89_clock = clock;
  assign dmem89_reset = reset;
  assign dmem89_io_pipeline_address = cpu89_io_dmem_address; // @[top.scala 641:17]
  assign dmem89_io_pipeline_valid = cpu89_io_dmem_valid; // @[top.scala 641:17]
  assign dmem89_io_pipeline_writedata = cpu89_io_dmem_writedata; // @[top.scala 641:17]
  assign dmem89_io_pipeline_memread = cpu89_io_dmem_memread; // @[top.scala 641:17]
  assign dmem89_io_pipeline_memwrite = cpu89_io_dmem_memwrite; // @[top.scala 641:17]
  assign dmem89_io_pipeline_maskmode = cpu89_io_dmem_maskmode; // @[top.scala 641:17]
  assign dmem89_io_pipeline_sext = cpu89_io_dmem_sext; // @[top.scala 641:17]
  assign dmem89_io_bus_response_valid = mem89_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem89_io_bus_response_bits_data = mem89_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu90_clock = clock;
  assign cpu90_reset = reset;
  assign cpu90_io_imem_instruction = imem90_io_pipeline_instruction; // @[top.scala 647:17]
  assign cpu90_io_dmem_readdata = dmem90_io_pipeline_readdata; // @[top.scala 648:17]
  assign mem90_clock = clock;
  assign mem90_reset = reset;
  assign mem90_io_imem_request_bits_address = imem90_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem90_io_dmem_request_valid = dmem90_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem90_io_dmem_request_bits_address = dmem90_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem90_io_dmem_request_bits_writedata = dmem90_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem90_io_dmem_request_bits_operation = dmem90_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem90_io_pipeline_address = cpu90_io_imem_address; // @[top.scala 647:17]
  assign imem90_io_bus_response_bits_data = mem90_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem90_clock = clock;
  assign dmem90_reset = reset;
  assign dmem90_io_pipeline_address = cpu90_io_dmem_address; // @[top.scala 648:17]
  assign dmem90_io_pipeline_valid = cpu90_io_dmem_valid; // @[top.scala 648:17]
  assign dmem90_io_pipeline_writedata = cpu90_io_dmem_writedata; // @[top.scala 648:17]
  assign dmem90_io_pipeline_memread = cpu90_io_dmem_memread; // @[top.scala 648:17]
  assign dmem90_io_pipeline_memwrite = cpu90_io_dmem_memwrite; // @[top.scala 648:17]
  assign dmem90_io_pipeline_maskmode = cpu90_io_dmem_maskmode; // @[top.scala 648:17]
  assign dmem90_io_pipeline_sext = cpu90_io_dmem_sext; // @[top.scala 648:17]
  assign dmem90_io_bus_response_valid = mem90_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem90_io_bus_response_bits_data = mem90_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu91_clock = clock;
  assign cpu91_reset = reset;
  assign cpu91_io_imem_instruction = imem91_io_pipeline_instruction; // @[top.scala 654:17]
  assign cpu91_io_dmem_readdata = dmem91_io_pipeline_readdata; // @[top.scala 655:17]
  assign mem91_clock = clock;
  assign mem91_reset = reset;
  assign mem91_io_imem_request_bits_address = imem91_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem91_io_dmem_request_valid = dmem91_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem91_io_dmem_request_bits_address = dmem91_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem91_io_dmem_request_bits_writedata = dmem91_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem91_io_dmem_request_bits_operation = dmem91_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem91_io_pipeline_address = cpu91_io_imem_address; // @[top.scala 654:17]
  assign imem91_io_bus_response_bits_data = mem91_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem91_clock = clock;
  assign dmem91_reset = reset;
  assign dmem91_io_pipeline_address = cpu91_io_dmem_address; // @[top.scala 655:17]
  assign dmem91_io_pipeline_valid = cpu91_io_dmem_valid; // @[top.scala 655:17]
  assign dmem91_io_pipeline_writedata = cpu91_io_dmem_writedata; // @[top.scala 655:17]
  assign dmem91_io_pipeline_memread = cpu91_io_dmem_memread; // @[top.scala 655:17]
  assign dmem91_io_pipeline_memwrite = cpu91_io_dmem_memwrite; // @[top.scala 655:17]
  assign dmem91_io_pipeline_maskmode = cpu91_io_dmem_maskmode; // @[top.scala 655:17]
  assign dmem91_io_pipeline_sext = cpu91_io_dmem_sext; // @[top.scala 655:17]
  assign dmem91_io_bus_response_valid = mem91_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem91_io_bus_response_bits_data = mem91_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu92_clock = clock;
  assign cpu92_reset = reset;
  assign cpu92_io_imem_instruction = imem92_io_pipeline_instruction; // @[top.scala 661:17]
  assign cpu92_io_dmem_readdata = dmem92_io_pipeline_readdata; // @[top.scala 662:17]
  assign mem92_clock = clock;
  assign mem92_reset = reset;
  assign mem92_io_imem_request_bits_address = imem92_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem92_io_dmem_request_valid = dmem92_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem92_io_dmem_request_bits_address = dmem92_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem92_io_dmem_request_bits_writedata = dmem92_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem92_io_dmem_request_bits_operation = dmem92_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem92_io_pipeline_address = cpu92_io_imem_address; // @[top.scala 661:17]
  assign imem92_io_bus_response_bits_data = mem92_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem92_clock = clock;
  assign dmem92_reset = reset;
  assign dmem92_io_pipeline_address = cpu92_io_dmem_address; // @[top.scala 662:17]
  assign dmem92_io_pipeline_valid = cpu92_io_dmem_valid; // @[top.scala 662:17]
  assign dmem92_io_pipeline_writedata = cpu92_io_dmem_writedata; // @[top.scala 662:17]
  assign dmem92_io_pipeline_memread = cpu92_io_dmem_memread; // @[top.scala 662:17]
  assign dmem92_io_pipeline_memwrite = cpu92_io_dmem_memwrite; // @[top.scala 662:17]
  assign dmem92_io_pipeline_maskmode = cpu92_io_dmem_maskmode; // @[top.scala 662:17]
  assign dmem92_io_pipeline_sext = cpu92_io_dmem_sext; // @[top.scala 662:17]
  assign dmem92_io_bus_response_valid = mem92_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem92_io_bus_response_bits_data = mem92_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu93_clock = clock;
  assign cpu93_reset = reset;
  assign cpu93_io_imem_instruction = imem93_io_pipeline_instruction; // @[top.scala 668:17]
  assign cpu93_io_dmem_readdata = dmem93_io_pipeline_readdata; // @[top.scala 669:17]
  assign mem93_clock = clock;
  assign mem93_reset = reset;
  assign mem93_io_imem_request_bits_address = imem93_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem93_io_dmem_request_valid = dmem93_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem93_io_dmem_request_bits_address = dmem93_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem93_io_dmem_request_bits_writedata = dmem93_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem93_io_dmem_request_bits_operation = dmem93_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem93_io_pipeline_address = cpu93_io_imem_address; // @[top.scala 668:17]
  assign imem93_io_bus_response_bits_data = mem93_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem93_clock = clock;
  assign dmem93_reset = reset;
  assign dmem93_io_pipeline_address = cpu93_io_dmem_address; // @[top.scala 669:17]
  assign dmem93_io_pipeline_valid = cpu93_io_dmem_valid; // @[top.scala 669:17]
  assign dmem93_io_pipeline_writedata = cpu93_io_dmem_writedata; // @[top.scala 669:17]
  assign dmem93_io_pipeline_memread = cpu93_io_dmem_memread; // @[top.scala 669:17]
  assign dmem93_io_pipeline_memwrite = cpu93_io_dmem_memwrite; // @[top.scala 669:17]
  assign dmem93_io_pipeline_maskmode = cpu93_io_dmem_maskmode; // @[top.scala 669:17]
  assign dmem93_io_pipeline_sext = cpu93_io_dmem_sext; // @[top.scala 669:17]
  assign dmem93_io_bus_response_valid = mem93_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem93_io_bus_response_bits_data = mem93_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu94_clock = clock;
  assign cpu94_reset = reset;
  assign cpu94_io_imem_instruction = imem94_io_pipeline_instruction; // @[top.scala 675:17]
  assign cpu94_io_dmem_readdata = dmem94_io_pipeline_readdata; // @[top.scala 676:17]
  assign mem94_clock = clock;
  assign mem94_reset = reset;
  assign mem94_io_imem_request_bits_address = imem94_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem94_io_dmem_request_valid = dmem94_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem94_io_dmem_request_bits_address = dmem94_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem94_io_dmem_request_bits_writedata = dmem94_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem94_io_dmem_request_bits_operation = dmem94_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem94_io_pipeline_address = cpu94_io_imem_address; // @[top.scala 675:17]
  assign imem94_io_bus_response_bits_data = mem94_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem94_clock = clock;
  assign dmem94_reset = reset;
  assign dmem94_io_pipeline_address = cpu94_io_dmem_address; // @[top.scala 676:17]
  assign dmem94_io_pipeline_valid = cpu94_io_dmem_valid; // @[top.scala 676:17]
  assign dmem94_io_pipeline_writedata = cpu94_io_dmem_writedata; // @[top.scala 676:17]
  assign dmem94_io_pipeline_memread = cpu94_io_dmem_memread; // @[top.scala 676:17]
  assign dmem94_io_pipeline_memwrite = cpu94_io_dmem_memwrite; // @[top.scala 676:17]
  assign dmem94_io_pipeline_maskmode = cpu94_io_dmem_maskmode; // @[top.scala 676:17]
  assign dmem94_io_pipeline_sext = cpu94_io_dmem_sext; // @[top.scala 676:17]
  assign dmem94_io_bus_response_valid = mem94_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem94_io_bus_response_bits_data = mem94_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu95_clock = clock;
  assign cpu95_reset = reset;
  assign cpu95_io_imem_instruction = imem95_io_pipeline_instruction; // @[top.scala 682:17]
  assign cpu95_io_dmem_readdata = dmem95_io_pipeline_readdata; // @[top.scala 683:17]
  assign mem95_clock = clock;
  assign mem95_reset = reset;
  assign mem95_io_imem_request_bits_address = imem95_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem95_io_dmem_request_valid = dmem95_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem95_io_dmem_request_bits_address = dmem95_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem95_io_dmem_request_bits_writedata = dmem95_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem95_io_dmem_request_bits_operation = dmem95_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem95_io_pipeline_address = cpu95_io_imem_address; // @[top.scala 682:17]
  assign imem95_io_bus_response_bits_data = mem95_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem95_clock = clock;
  assign dmem95_reset = reset;
  assign dmem95_io_pipeline_address = cpu95_io_dmem_address; // @[top.scala 683:17]
  assign dmem95_io_pipeline_valid = cpu95_io_dmem_valid; // @[top.scala 683:17]
  assign dmem95_io_pipeline_writedata = cpu95_io_dmem_writedata; // @[top.scala 683:17]
  assign dmem95_io_pipeline_memread = cpu95_io_dmem_memread; // @[top.scala 683:17]
  assign dmem95_io_pipeline_memwrite = cpu95_io_dmem_memwrite; // @[top.scala 683:17]
  assign dmem95_io_pipeline_maskmode = cpu95_io_dmem_maskmode; // @[top.scala 683:17]
  assign dmem95_io_pipeline_sext = cpu95_io_dmem_sext; // @[top.scala 683:17]
  assign dmem95_io_bus_response_valid = mem95_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem95_io_bus_response_bits_data = mem95_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu96_clock = clock;
  assign cpu96_reset = reset;
  assign cpu96_io_imem_instruction = imem96_io_pipeline_instruction; // @[top.scala 689:17]
  assign cpu96_io_dmem_readdata = dmem96_io_pipeline_readdata; // @[top.scala 690:17]
  assign mem96_clock = clock;
  assign mem96_reset = reset;
  assign mem96_io_imem_request_bits_address = imem96_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem96_io_dmem_request_valid = dmem96_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem96_io_dmem_request_bits_address = dmem96_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem96_io_dmem_request_bits_writedata = dmem96_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem96_io_dmem_request_bits_operation = dmem96_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem96_io_pipeline_address = cpu96_io_imem_address; // @[top.scala 689:17]
  assign imem96_io_bus_response_bits_data = mem96_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem96_clock = clock;
  assign dmem96_reset = reset;
  assign dmem96_io_pipeline_address = cpu96_io_dmem_address; // @[top.scala 690:17]
  assign dmem96_io_pipeline_valid = cpu96_io_dmem_valid; // @[top.scala 690:17]
  assign dmem96_io_pipeline_writedata = cpu96_io_dmem_writedata; // @[top.scala 690:17]
  assign dmem96_io_pipeline_memread = cpu96_io_dmem_memread; // @[top.scala 690:17]
  assign dmem96_io_pipeline_memwrite = cpu96_io_dmem_memwrite; // @[top.scala 690:17]
  assign dmem96_io_pipeline_maskmode = cpu96_io_dmem_maskmode; // @[top.scala 690:17]
  assign dmem96_io_pipeline_sext = cpu96_io_dmem_sext; // @[top.scala 690:17]
  assign dmem96_io_bus_response_valid = mem96_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem96_io_bus_response_bits_data = mem96_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu97_clock = clock;
  assign cpu97_reset = reset;
  assign cpu97_io_imem_instruction = imem97_io_pipeline_instruction; // @[top.scala 696:17]
  assign cpu97_io_dmem_readdata = dmem97_io_pipeline_readdata; // @[top.scala 697:17]
  assign mem97_clock = clock;
  assign mem97_reset = reset;
  assign mem97_io_imem_request_bits_address = imem97_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem97_io_dmem_request_valid = dmem97_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem97_io_dmem_request_bits_address = dmem97_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem97_io_dmem_request_bits_writedata = dmem97_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem97_io_dmem_request_bits_operation = dmem97_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem97_io_pipeline_address = cpu97_io_imem_address; // @[top.scala 696:17]
  assign imem97_io_bus_response_bits_data = mem97_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem97_clock = clock;
  assign dmem97_reset = reset;
  assign dmem97_io_pipeline_address = cpu97_io_dmem_address; // @[top.scala 697:17]
  assign dmem97_io_pipeline_valid = cpu97_io_dmem_valid; // @[top.scala 697:17]
  assign dmem97_io_pipeline_writedata = cpu97_io_dmem_writedata; // @[top.scala 697:17]
  assign dmem97_io_pipeline_memread = cpu97_io_dmem_memread; // @[top.scala 697:17]
  assign dmem97_io_pipeline_memwrite = cpu97_io_dmem_memwrite; // @[top.scala 697:17]
  assign dmem97_io_pipeline_maskmode = cpu97_io_dmem_maskmode; // @[top.scala 697:17]
  assign dmem97_io_pipeline_sext = cpu97_io_dmem_sext; // @[top.scala 697:17]
  assign dmem97_io_bus_response_valid = mem97_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem97_io_bus_response_bits_data = mem97_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu98_clock = clock;
  assign cpu98_reset = reset;
  assign cpu98_io_imem_instruction = imem98_io_pipeline_instruction; // @[top.scala 703:17]
  assign cpu98_io_dmem_readdata = dmem98_io_pipeline_readdata; // @[top.scala 704:17]
  assign mem98_clock = clock;
  assign mem98_reset = reset;
  assign mem98_io_imem_request_bits_address = imem98_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem98_io_dmem_request_valid = dmem98_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem98_io_dmem_request_bits_address = dmem98_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem98_io_dmem_request_bits_writedata = dmem98_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem98_io_dmem_request_bits_operation = dmem98_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem98_io_pipeline_address = cpu98_io_imem_address; // @[top.scala 703:17]
  assign imem98_io_bus_response_bits_data = mem98_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem98_clock = clock;
  assign dmem98_reset = reset;
  assign dmem98_io_pipeline_address = cpu98_io_dmem_address; // @[top.scala 704:17]
  assign dmem98_io_pipeline_valid = cpu98_io_dmem_valid; // @[top.scala 704:17]
  assign dmem98_io_pipeline_writedata = cpu98_io_dmem_writedata; // @[top.scala 704:17]
  assign dmem98_io_pipeline_memread = cpu98_io_dmem_memread; // @[top.scala 704:17]
  assign dmem98_io_pipeline_memwrite = cpu98_io_dmem_memwrite; // @[top.scala 704:17]
  assign dmem98_io_pipeline_maskmode = cpu98_io_dmem_maskmode; // @[top.scala 704:17]
  assign dmem98_io_pipeline_sext = cpu98_io_dmem_sext; // @[top.scala 704:17]
  assign dmem98_io_bus_response_valid = mem98_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem98_io_bus_response_bits_data = mem98_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu99_clock = clock;
  assign cpu99_reset = reset;
  assign cpu99_io_imem_instruction = imem99_io_pipeline_instruction; // @[top.scala 710:17]
  assign cpu99_io_dmem_readdata = dmem99_io_pipeline_readdata; // @[top.scala 711:17]
  assign mem99_clock = clock;
  assign mem99_reset = reset;
  assign mem99_io_imem_request_bits_address = imem99_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem99_io_dmem_request_valid = dmem99_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem99_io_dmem_request_bits_address = dmem99_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem99_io_dmem_request_bits_writedata = dmem99_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem99_io_dmem_request_bits_operation = dmem99_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem99_io_pipeline_address = cpu99_io_imem_address; // @[top.scala 710:17]
  assign imem99_io_bus_response_bits_data = mem99_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem99_clock = clock;
  assign dmem99_reset = reset;
  assign dmem99_io_pipeline_address = cpu99_io_dmem_address; // @[top.scala 711:17]
  assign dmem99_io_pipeline_valid = cpu99_io_dmem_valid; // @[top.scala 711:17]
  assign dmem99_io_pipeline_writedata = cpu99_io_dmem_writedata; // @[top.scala 711:17]
  assign dmem99_io_pipeline_memread = cpu99_io_dmem_memread; // @[top.scala 711:17]
  assign dmem99_io_pipeline_memwrite = cpu99_io_dmem_memwrite; // @[top.scala 711:17]
  assign dmem99_io_pipeline_maskmode = cpu99_io_dmem_maskmode; // @[top.scala 711:17]
  assign dmem99_io_pipeline_sext = cpu99_io_dmem_sext; // @[top.scala 711:17]
  assign dmem99_io_bus_response_valid = mem99_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem99_io_bus_response_bits_data = mem99_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu100_clock = clock;
  assign cpu100_reset = reset;
  assign cpu100_io_imem_instruction = imem100_io_pipeline_instruction; // @[top.scala 717:18]
  assign cpu100_io_dmem_readdata = dmem100_io_pipeline_readdata; // @[top.scala 718:18]
  assign mem100_clock = clock;
  assign mem100_reset = reset;
  assign mem100_io_imem_request_bits_address = imem100_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem100_io_dmem_request_valid = dmem100_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem100_io_dmem_request_bits_address = dmem100_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem100_io_dmem_request_bits_writedata = dmem100_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem100_io_dmem_request_bits_operation = dmem100_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem100_io_pipeline_address = cpu100_io_imem_address; // @[top.scala 717:18]
  assign imem100_io_bus_response_bits_data = mem100_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem100_clock = clock;
  assign dmem100_reset = reset;
  assign dmem100_io_pipeline_address = cpu100_io_dmem_address; // @[top.scala 718:18]
  assign dmem100_io_pipeline_valid = cpu100_io_dmem_valid; // @[top.scala 718:18]
  assign dmem100_io_pipeline_writedata = cpu100_io_dmem_writedata; // @[top.scala 718:18]
  assign dmem100_io_pipeline_memread = cpu100_io_dmem_memread; // @[top.scala 718:18]
  assign dmem100_io_pipeline_memwrite = cpu100_io_dmem_memwrite; // @[top.scala 718:18]
  assign dmem100_io_pipeline_maskmode = cpu100_io_dmem_maskmode; // @[top.scala 718:18]
  assign dmem100_io_pipeline_sext = cpu100_io_dmem_sext; // @[top.scala 718:18]
  assign dmem100_io_bus_response_valid = mem100_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem100_io_bus_response_bits_data = mem100_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu101_clock = clock;
  assign cpu101_reset = reset;
  assign cpu101_io_imem_instruction = imem101_io_pipeline_instruction; // @[top.scala 724:18]
  assign cpu101_io_dmem_readdata = dmem101_io_pipeline_readdata; // @[top.scala 725:18]
  assign mem101_clock = clock;
  assign mem101_reset = reset;
  assign mem101_io_imem_request_bits_address = imem101_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem101_io_dmem_request_valid = dmem101_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem101_io_dmem_request_bits_address = dmem101_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem101_io_dmem_request_bits_writedata = dmem101_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem101_io_dmem_request_bits_operation = dmem101_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem101_io_pipeline_address = cpu101_io_imem_address; // @[top.scala 724:18]
  assign imem101_io_bus_response_bits_data = mem101_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem101_clock = clock;
  assign dmem101_reset = reset;
  assign dmem101_io_pipeline_address = cpu101_io_dmem_address; // @[top.scala 725:18]
  assign dmem101_io_pipeline_valid = cpu101_io_dmem_valid; // @[top.scala 725:18]
  assign dmem101_io_pipeline_writedata = cpu101_io_dmem_writedata; // @[top.scala 725:18]
  assign dmem101_io_pipeline_memread = cpu101_io_dmem_memread; // @[top.scala 725:18]
  assign dmem101_io_pipeline_memwrite = cpu101_io_dmem_memwrite; // @[top.scala 725:18]
  assign dmem101_io_pipeline_maskmode = cpu101_io_dmem_maskmode; // @[top.scala 725:18]
  assign dmem101_io_pipeline_sext = cpu101_io_dmem_sext; // @[top.scala 725:18]
  assign dmem101_io_bus_response_valid = mem101_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem101_io_bus_response_bits_data = mem101_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu102_clock = clock;
  assign cpu102_reset = reset;
  assign cpu102_io_imem_instruction = imem102_io_pipeline_instruction; // @[top.scala 731:18]
  assign cpu102_io_dmem_readdata = dmem102_io_pipeline_readdata; // @[top.scala 732:18]
  assign mem102_clock = clock;
  assign mem102_reset = reset;
  assign mem102_io_imem_request_bits_address = imem102_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem102_io_dmem_request_valid = dmem102_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem102_io_dmem_request_bits_address = dmem102_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem102_io_dmem_request_bits_writedata = dmem102_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem102_io_dmem_request_bits_operation = dmem102_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem102_io_pipeline_address = cpu102_io_imem_address; // @[top.scala 731:18]
  assign imem102_io_bus_response_bits_data = mem102_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem102_clock = clock;
  assign dmem102_reset = reset;
  assign dmem102_io_pipeline_address = cpu102_io_dmem_address; // @[top.scala 732:18]
  assign dmem102_io_pipeline_valid = cpu102_io_dmem_valid; // @[top.scala 732:18]
  assign dmem102_io_pipeline_writedata = cpu102_io_dmem_writedata; // @[top.scala 732:18]
  assign dmem102_io_pipeline_memread = cpu102_io_dmem_memread; // @[top.scala 732:18]
  assign dmem102_io_pipeline_memwrite = cpu102_io_dmem_memwrite; // @[top.scala 732:18]
  assign dmem102_io_pipeline_maskmode = cpu102_io_dmem_maskmode; // @[top.scala 732:18]
  assign dmem102_io_pipeline_sext = cpu102_io_dmem_sext; // @[top.scala 732:18]
  assign dmem102_io_bus_response_valid = mem102_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem102_io_bus_response_bits_data = mem102_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu103_clock = clock;
  assign cpu103_reset = reset;
  assign cpu103_io_imem_instruction = imem103_io_pipeline_instruction; // @[top.scala 738:18]
  assign cpu103_io_dmem_readdata = dmem103_io_pipeline_readdata; // @[top.scala 739:18]
  assign mem103_clock = clock;
  assign mem103_reset = reset;
  assign mem103_io_imem_request_bits_address = imem103_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem103_io_dmem_request_valid = dmem103_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem103_io_dmem_request_bits_address = dmem103_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem103_io_dmem_request_bits_writedata = dmem103_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem103_io_dmem_request_bits_operation = dmem103_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem103_io_pipeline_address = cpu103_io_imem_address; // @[top.scala 738:18]
  assign imem103_io_bus_response_bits_data = mem103_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem103_clock = clock;
  assign dmem103_reset = reset;
  assign dmem103_io_pipeline_address = cpu103_io_dmem_address; // @[top.scala 739:18]
  assign dmem103_io_pipeline_valid = cpu103_io_dmem_valid; // @[top.scala 739:18]
  assign dmem103_io_pipeline_writedata = cpu103_io_dmem_writedata; // @[top.scala 739:18]
  assign dmem103_io_pipeline_memread = cpu103_io_dmem_memread; // @[top.scala 739:18]
  assign dmem103_io_pipeline_memwrite = cpu103_io_dmem_memwrite; // @[top.scala 739:18]
  assign dmem103_io_pipeline_maskmode = cpu103_io_dmem_maskmode; // @[top.scala 739:18]
  assign dmem103_io_pipeline_sext = cpu103_io_dmem_sext; // @[top.scala 739:18]
  assign dmem103_io_bus_response_valid = mem103_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem103_io_bus_response_bits_data = mem103_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu104_clock = clock;
  assign cpu104_reset = reset;
  assign cpu104_io_imem_instruction = imem104_io_pipeline_instruction; // @[top.scala 745:18]
  assign cpu104_io_dmem_readdata = dmem104_io_pipeline_readdata; // @[top.scala 746:18]
  assign mem104_clock = clock;
  assign mem104_reset = reset;
  assign mem104_io_imem_request_bits_address = imem104_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem104_io_dmem_request_valid = dmem104_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem104_io_dmem_request_bits_address = dmem104_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem104_io_dmem_request_bits_writedata = dmem104_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem104_io_dmem_request_bits_operation = dmem104_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem104_io_pipeline_address = cpu104_io_imem_address; // @[top.scala 745:18]
  assign imem104_io_bus_response_bits_data = mem104_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem104_clock = clock;
  assign dmem104_reset = reset;
  assign dmem104_io_pipeline_address = cpu104_io_dmem_address; // @[top.scala 746:18]
  assign dmem104_io_pipeline_valid = cpu104_io_dmem_valid; // @[top.scala 746:18]
  assign dmem104_io_pipeline_writedata = cpu104_io_dmem_writedata; // @[top.scala 746:18]
  assign dmem104_io_pipeline_memread = cpu104_io_dmem_memread; // @[top.scala 746:18]
  assign dmem104_io_pipeline_memwrite = cpu104_io_dmem_memwrite; // @[top.scala 746:18]
  assign dmem104_io_pipeline_maskmode = cpu104_io_dmem_maskmode; // @[top.scala 746:18]
  assign dmem104_io_pipeline_sext = cpu104_io_dmem_sext; // @[top.scala 746:18]
  assign dmem104_io_bus_response_valid = mem104_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem104_io_bus_response_bits_data = mem104_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu105_clock = clock;
  assign cpu105_reset = reset;
  assign cpu105_io_imem_instruction = imem105_io_pipeline_instruction; // @[top.scala 752:18]
  assign cpu105_io_dmem_readdata = dmem105_io_pipeline_readdata; // @[top.scala 753:18]
  assign mem105_clock = clock;
  assign mem105_reset = reset;
  assign mem105_io_imem_request_bits_address = imem105_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem105_io_dmem_request_valid = dmem105_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem105_io_dmem_request_bits_address = dmem105_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem105_io_dmem_request_bits_writedata = dmem105_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem105_io_dmem_request_bits_operation = dmem105_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem105_io_pipeline_address = cpu105_io_imem_address; // @[top.scala 752:18]
  assign imem105_io_bus_response_bits_data = mem105_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem105_clock = clock;
  assign dmem105_reset = reset;
  assign dmem105_io_pipeline_address = cpu105_io_dmem_address; // @[top.scala 753:18]
  assign dmem105_io_pipeline_valid = cpu105_io_dmem_valid; // @[top.scala 753:18]
  assign dmem105_io_pipeline_writedata = cpu105_io_dmem_writedata; // @[top.scala 753:18]
  assign dmem105_io_pipeline_memread = cpu105_io_dmem_memread; // @[top.scala 753:18]
  assign dmem105_io_pipeline_memwrite = cpu105_io_dmem_memwrite; // @[top.scala 753:18]
  assign dmem105_io_pipeline_maskmode = cpu105_io_dmem_maskmode; // @[top.scala 753:18]
  assign dmem105_io_pipeline_sext = cpu105_io_dmem_sext; // @[top.scala 753:18]
  assign dmem105_io_bus_response_valid = mem105_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem105_io_bus_response_bits_data = mem105_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu106_clock = clock;
  assign cpu106_reset = reset;
  assign cpu106_io_imem_instruction = imem106_io_pipeline_instruction; // @[top.scala 759:18]
  assign cpu106_io_dmem_readdata = dmem106_io_pipeline_readdata; // @[top.scala 760:18]
  assign mem106_clock = clock;
  assign mem106_reset = reset;
  assign mem106_io_imem_request_bits_address = imem106_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem106_io_dmem_request_valid = dmem106_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem106_io_dmem_request_bits_address = dmem106_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem106_io_dmem_request_bits_writedata = dmem106_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem106_io_dmem_request_bits_operation = dmem106_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem106_io_pipeline_address = cpu106_io_imem_address; // @[top.scala 759:18]
  assign imem106_io_bus_response_bits_data = mem106_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem106_clock = clock;
  assign dmem106_reset = reset;
  assign dmem106_io_pipeline_address = cpu106_io_dmem_address; // @[top.scala 760:18]
  assign dmem106_io_pipeline_valid = cpu106_io_dmem_valid; // @[top.scala 760:18]
  assign dmem106_io_pipeline_writedata = cpu106_io_dmem_writedata; // @[top.scala 760:18]
  assign dmem106_io_pipeline_memread = cpu106_io_dmem_memread; // @[top.scala 760:18]
  assign dmem106_io_pipeline_memwrite = cpu106_io_dmem_memwrite; // @[top.scala 760:18]
  assign dmem106_io_pipeline_maskmode = cpu106_io_dmem_maskmode; // @[top.scala 760:18]
  assign dmem106_io_pipeline_sext = cpu106_io_dmem_sext; // @[top.scala 760:18]
  assign dmem106_io_bus_response_valid = mem106_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem106_io_bus_response_bits_data = mem106_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu107_clock = clock;
  assign cpu107_reset = reset;
  assign cpu107_io_imem_instruction = imem107_io_pipeline_instruction; // @[top.scala 766:18]
  assign cpu107_io_dmem_readdata = dmem107_io_pipeline_readdata; // @[top.scala 767:18]
  assign mem107_clock = clock;
  assign mem107_reset = reset;
  assign mem107_io_imem_request_bits_address = imem107_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem107_io_dmem_request_valid = dmem107_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem107_io_dmem_request_bits_address = dmem107_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem107_io_dmem_request_bits_writedata = dmem107_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem107_io_dmem_request_bits_operation = dmem107_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem107_io_pipeline_address = cpu107_io_imem_address; // @[top.scala 766:18]
  assign imem107_io_bus_response_bits_data = mem107_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem107_clock = clock;
  assign dmem107_reset = reset;
  assign dmem107_io_pipeline_address = cpu107_io_dmem_address; // @[top.scala 767:18]
  assign dmem107_io_pipeline_valid = cpu107_io_dmem_valid; // @[top.scala 767:18]
  assign dmem107_io_pipeline_writedata = cpu107_io_dmem_writedata; // @[top.scala 767:18]
  assign dmem107_io_pipeline_memread = cpu107_io_dmem_memread; // @[top.scala 767:18]
  assign dmem107_io_pipeline_memwrite = cpu107_io_dmem_memwrite; // @[top.scala 767:18]
  assign dmem107_io_pipeline_maskmode = cpu107_io_dmem_maskmode; // @[top.scala 767:18]
  assign dmem107_io_pipeline_sext = cpu107_io_dmem_sext; // @[top.scala 767:18]
  assign dmem107_io_bus_response_valid = mem107_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem107_io_bus_response_bits_data = mem107_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu108_clock = clock;
  assign cpu108_reset = reset;
  assign cpu108_io_imem_instruction = imem108_io_pipeline_instruction; // @[top.scala 773:18]
  assign cpu108_io_dmem_readdata = dmem108_io_pipeline_readdata; // @[top.scala 774:18]
  assign mem108_clock = clock;
  assign mem108_reset = reset;
  assign mem108_io_imem_request_bits_address = imem108_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem108_io_dmem_request_valid = dmem108_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem108_io_dmem_request_bits_address = dmem108_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem108_io_dmem_request_bits_writedata = dmem108_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem108_io_dmem_request_bits_operation = dmem108_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem108_io_pipeline_address = cpu108_io_imem_address; // @[top.scala 773:18]
  assign imem108_io_bus_response_bits_data = mem108_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem108_clock = clock;
  assign dmem108_reset = reset;
  assign dmem108_io_pipeline_address = cpu108_io_dmem_address; // @[top.scala 774:18]
  assign dmem108_io_pipeline_valid = cpu108_io_dmem_valid; // @[top.scala 774:18]
  assign dmem108_io_pipeline_writedata = cpu108_io_dmem_writedata; // @[top.scala 774:18]
  assign dmem108_io_pipeline_memread = cpu108_io_dmem_memread; // @[top.scala 774:18]
  assign dmem108_io_pipeline_memwrite = cpu108_io_dmem_memwrite; // @[top.scala 774:18]
  assign dmem108_io_pipeline_maskmode = cpu108_io_dmem_maskmode; // @[top.scala 774:18]
  assign dmem108_io_pipeline_sext = cpu108_io_dmem_sext; // @[top.scala 774:18]
  assign dmem108_io_bus_response_valid = mem108_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem108_io_bus_response_bits_data = mem108_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu109_clock = clock;
  assign cpu109_reset = reset;
  assign cpu109_io_imem_instruction = imem109_io_pipeline_instruction; // @[top.scala 780:18]
  assign cpu109_io_dmem_readdata = dmem109_io_pipeline_readdata; // @[top.scala 781:18]
  assign mem109_clock = clock;
  assign mem109_reset = reset;
  assign mem109_io_imem_request_bits_address = imem109_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem109_io_dmem_request_valid = dmem109_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem109_io_dmem_request_bits_address = dmem109_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem109_io_dmem_request_bits_writedata = dmem109_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem109_io_dmem_request_bits_operation = dmem109_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem109_io_pipeline_address = cpu109_io_imem_address; // @[top.scala 780:18]
  assign imem109_io_bus_response_bits_data = mem109_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem109_clock = clock;
  assign dmem109_reset = reset;
  assign dmem109_io_pipeline_address = cpu109_io_dmem_address; // @[top.scala 781:18]
  assign dmem109_io_pipeline_valid = cpu109_io_dmem_valid; // @[top.scala 781:18]
  assign dmem109_io_pipeline_writedata = cpu109_io_dmem_writedata; // @[top.scala 781:18]
  assign dmem109_io_pipeline_memread = cpu109_io_dmem_memread; // @[top.scala 781:18]
  assign dmem109_io_pipeline_memwrite = cpu109_io_dmem_memwrite; // @[top.scala 781:18]
  assign dmem109_io_pipeline_maskmode = cpu109_io_dmem_maskmode; // @[top.scala 781:18]
  assign dmem109_io_pipeline_sext = cpu109_io_dmem_sext; // @[top.scala 781:18]
  assign dmem109_io_bus_response_valid = mem109_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem109_io_bus_response_bits_data = mem109_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu110_clock = clock;
  assign cpu110_reset = reset;
  assign cpu110_io_imem_instruction = imem110_io_pipeline_instruction; // @[top.scala 787:18]
  assign cpu110_io_dmem_readdata = dmem110_io_pipeline_readdata; // @[top.scala 788:18]
  assign mem110_clock = clock;
  assign mem110_reset = reset;
  assign mem110_io_imem_request_bits_address = imem110_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem110_io_dmem_request_valid = dmem110_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem110_io_dmem_request_bits_address = dmem110_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem110_io_dmem_request_bits_writedata = dmem110_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem110_io_dmem_request_bits_operation = dmem110_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem110_io_pipeline_address = cpu110_io_imem_address; // @[top.scala 787:18]
  assign imem110_io_bus_response_bits_data = mem110_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem110_clock = clock;
  assign dmem110_reset = reset;
  assign dmem110_io_pipeline_address = cpu110_io_dmem_address; // @[top.scala 788:18]
  assign dmem110_io_pipeline_valid = cpu110_io_dmem_valid; // @[top.scala 788:18]
  assign dmem110_io_pipeline_writedata = cpu110_io_dmem_writedata; // @[top.scala 788:18]
  assign dmem110_io_pipeline_memread = cpu110_io_dmem_memread; // @[top.scala 788:18]
  assign dmem110_io_pipeline_memwrite = cpu110_io_dmem_memwrite; // @[top.scala 788:18]
  assign dmem110_io_pipeline_maskmode = cpu110_io_dmem_maskmode; // @[top.scala 788:18]
  assign dmem110_io_pipeline_sext = cpu110_io_dmem_sext; // @[top.scala 788:18]
  assign dmem110_io_bus_response_valid = mem110_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem110_io_bus_response_bits_data = mem110_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu111_clock = clock;
  assign cpu111_reset = reset;
  assign cpu111_io_imem_instruction = imem111_io_pipeline_instruction; // @[top.scala 794:18]
  assign cpu111_io_dmem_readdata = dmem111_io_pipeline_readdata; // @[top.scala 795:18]
  assign mem111_clock = clock;
  assign mem111_reset = reset;
  assign mem111_io_imem_request_bits_address = imem111_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem111_io_dmem_request_valid = dmem111_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem111_io_dmem_request_bits_address = dmem111_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem111_io_dmem_request_bits_writedata = dmem111_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem111_io_dmem_request_bits_operation = dmem111_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem111_io_pipeline_address = cpu111_io_imem_address; // @[top.scala 794:18]
  assign imem111_io_bus_response_bits_data = mem111_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem111_clock = clock;
  assign dmem111_reset = reset;
  assign dmem111_io_pipeline_address = cpu111_io_dmem_address; // @[top.scala 795:18]
  assign dmem111_io_pipeline_valid = cpu111_io_dmem_valid; // @[top.scala 795:18]
  assign dmem111_io_pipeline_writedata = cpu111_io_dmem_writedata; // @[top.scala 795:18]
  assign dmem111_io_pipeline_memread = cpu111_io_dmem_memread; // @[top.scala 795:18]
  assign dmem111_io_pipeline_memwrite = cpu111_io_dmem_memwrite; // @[top.scala 795:18]
  assign dmem111_io_pipeline_maskmode = cpu111_io_dmem_maskmode; // @[top.scala 795:18]
  assign dmem111_io_pipeline_sext = cpu111_io_dmem_sext; // @[top.scala 795:18]
  assign dmem111_io_bus_response_valid = mem111_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem111_io_bus_response_bits_data = mem111_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu112_clock = clock;
  assign cpu112_reset = reset;
  assign cpu112_io_imem_instruction = imem112_io_pipeline_instruction; // @[top.scala 801:18]
  assign cpu112_io_dmem_readdata = dmem112_io_pipeline_readdata; // @[top.scala 802:18]
  assign mem112_clock = clock;
  assign mem112_reset = reset;
  assign mem112_io_imem_request_bits_address = imem112_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem112_io_dmem_request_valid = dmem112_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem112_io_dmem_request_bits_address = dmem112_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem112_io_dmem_request_bits_writedata = dmem112_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem112_io_dmem_request_bits_operation = dmem112_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem112_io_pipeline_address = cpu112_io_imem_address; // @[top.scala 801:18]
  assign imem112_io_bus_response_bits_data = mem112_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem112_clock = clock;
  assign dmem112_reset = reset;
  assign dmem112_io_pipeline_address = cpu112_io_dmem_address; // @[top.scala 802:18]
  assign dmem112_io_pipeline_valid = cpu112_io_dmem_valid; // @[top.scala 802:18]
  assign dmem112_io_pipeline_writedata = cpu112_io_dmem_writedata; // @[top.scala 802:18]
  assign dmem112_io_pipeline_memread = cpu112_io_dmem_memread; // @[top.scala 802:18]
  assign dmem112_io_pipeline_memwrite = cpu112_io_dmem_memwrite; // @[top.scala 802:18]
  assign dmem112_io_pipeline_maskmode = cpu112_io_dmem_maskmode; // @[top.scala 802:18]
  assign dmem112_io_pipeline_sext = cpu112_io_dmem_sext; // @[top.scala 802:18]
  assign dmem112_io_bus_response_valid = mem112_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem112_io_bus_response_bits_data = mem112_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu113_clock = clock;
  assign cpu113_reset = reset;
  assign cpu113_io_imem_instruction = imem113_io_pipeline_instruction; // @[top.scala 808:18]
  assign cpu113_io_dmem_readdata = dmem113_io_pipeline_readdata; // @[top.scala 809:18]
  assign mem113_clock = clock;
  assign mem113_reset = reset;
  assign mem113_io_imem_request_bits_address = imem113_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem113_io_dmem_request_valid = dmem113_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem113_io_dmem_request_bits_address = dmem113_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem113_io_dmem_request_bits_writedata = dmem113_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem113_io_dmem_request_bits_operation = dmem113_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem113_io_pipeline_address = cpu113_io_imem_address; // @[top.scala 808:18]
  assign imem113_io_bus_response_bits_data = mem113_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem113_clock = clock;
  assign dmem113_reset = reset;
  assign dmem113_io_pipeline_address = cpu113_io_dmem_address; // @[top.scala 809:18]
  assign dmem113_io_pipeline_valid = cpu113_io_dmem_valid; // @[top.scala 809:18]
  assign dmem113_io_pipeline_writedata = cpu113_io_dmem_writedata; // @[top.scala 809:18]
  assign dmem113_io_pipeline_memread = cpu113_io_dmem_memread; // @[top.scala 809:18]
  assign dmem113_io_pipeline_memwrite = cpu113_io_dmem_memwrite; // @[top.scala 809:18]
  assign dmem113_io_pipeline_maskmode = cpu113_io_dmem_maskmode; // @[top.scala 809:18]
  assign dmem113_io_pipeline_sext = cpu113_io_dmem_sext; // @[top.scala 809:18]
  assign dmem113_io_bus_response_valid = mem113_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem113_io_bus_response_bits_data = mem113_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu114_clock = clock;
  assign cpu114_reset = reset;
  assign cpu114_io_imem_instruction = imem114_io_pipeline_instruction; // @[top.scala 815:18]
  assign cpu114_io_dmem_readdata = dmem114_io_pipeline_readdata; // @[top.scala 816:18]
  assign mem114_clock = clock;
  assign mem114_reset = reset;
  assign mem114_io_imem_request_bits_address = imem114_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem114_io_dmem_request_valid = dmem114_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem114_io_dmem_request_bits_address = dmem114_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem114_io_dmem_request_bits_writedata = dmem114_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem114_io_dmem_request_bits_operation = dmem114_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem114_io_pipeline_address = cpu114_io_imem_address; // @[top.scala 815:18]
  assign imem114_io_bus_response_bits_data = mem114_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem114_clock = clock;
  assign dmem114_reset = reset;
  assign dmem114_io_pipeline_address = cpu114_io_dmem_address; // @[top.scala 816:18]
  assign dmem114_io_pipeline_valid = cpu114_io_dmem_valid; // @[top.scala 816:18]
  assign dmem114_io_pipeline_writedata = cpu114_io_dmem_writedata; // @[top.scala 816:18]
  assign dmem114_io_pipeline_memread = cpu114_io_dmem_memread; // @[top.scala 816:18]
  assign dmem114_io_pipeline_memwrite = cpu114_io_dmem_memwrite; // @[top.scala 816:18]
  assign dmem114_io_pipeline_maskmode = cpu114_io_dmem_maskmode; // @[top.scala 816:18]
  assign dmem114_io_pipeline_sext = cpu114_io_dmem_sext; // @[top.scala 816:18]
  assign dmem114_io_bus_response_valid = mem114_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem114_io_bus_response_bits_data = mem114_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu115_clock = clock;
  assign cpu115_reset = reset;
  assign cpu115_io_imem_instruction = imem115_io_pipeline_instruction; // @[top.scala 822:18]
  assign cpu115_io_dmem_readdata = dmem115_io_pipeline_readdata; // @[top.scala 823:18]
  assign mem115_clock = clock;
  assign mem115_reset = reset;
  assign mem115_io_imem_request_bits_address = imem115_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem115_io_dmem_request_valid = dmem115_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem115_io_dmem_request_bits_address = dmem115_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem115_io_dmem_request_bits_writedata = dmem115_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem115_io_dmem_request_bits_operation = dmem115_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem115_io_pipeline_address = cpu115_io_imem_address; // @[top.scala 822:18]
  assign imem115_io_bus_response_bits_data = mem115_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem115_clock = clock;
  assign dmem115_reset = reset;
  assign dmem115_io_pipeline_address = cpu115_io_dmem_address; // @[top.scala 823:18]
  assign dmem115_io_pipeline_valid = cpu115_io_dmem_valid; // @[top.scala 823:18]
  assign dmem115_io_pipeline_writedata = cpu115_io_dmem_writedata; // @[top.scala 823:18]
  assign dmem115_io_pipeline_memread = cpu115_io_dmem_memread; // @[top.scala 823:18]
  assign dmem115_io_pipeline_memwrite = cpu115_io_dmem_memwrite; // @[top.scala 823:18]
  assign dmem115_io_pipeline_maskmode = cpu115_io_dmem_maskmode; // @[top.scala 823:18]
  assign dmem115_io_pipeline_sext = cpu115_io_dmem_sext; // @[top.scala 823:18]
  assign dmem115_io_bus_response_valid = mem115_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem115_io_bus_response_bits_data = mem115_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu116_clock = clock;
  assign cpu116_reset = reset;
  assign cpu116_io_imem_instruction = imem116_io_pipeline_instruction; // @[top.scala 829:18]
  assign cpu116_io_dmem_readdata = dmem116_io_pipeline_readdata; // @[top.scala 830:18]
  assign mem116_clock = clock;
  assign mem116_reset = reset;
  assign mem116_io_imem_request_bits_address = imem116_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem116_io_dmem_request_valid = dmem116_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem116_io_dmem_request_bits_address = dmem116_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem116_io_dmem_request_bits_writedata = dmem116_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem116_io_dmem_request_bits_operation = dmem116_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem116_io_pipeline_address = cpu116_io_imem_address; // @[top.scala 829:18]
  assign imem116_io_bus_response_bits_data = mem116_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem116_clock = clock;
  assign dmem116_reset = reset;
  assign dmem116_io_pipeline_address = cpu116_io_dmem_address; // @[top.scala 830:18]
  assign dmem116_io_pipeline_valid = cpu116_io_dmem_valid; // @[top.scala 830:18]
  assign dmem116_io_pipeline_writedata = cpu116_io_dmem_writedata; // @[top.scala 830:18]
  assign dmem116_io_pipeline_memread = cpu116_io_dmem_memread; // @[top.scala 830:18]
  assign dmem116_io_pipeline_memwrite = cpu116_io_dmem_memwrite; // @[top.scala 830:18]
  assign dmem116_io_pipeline_maskmode = cpu116_io_dmem_maskmode; // @[top.scala 830:18]
  assign dmem116_io_pipeline_sext = cpu116_io_dmem_sext; // @[top.scala 830:18]
  assign dmem116_io_bus_response_valid = mem116_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem116_io_bus_response_bits_data = mem116_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu117_clock = clock;
  assign cpu117_reset = reset;
  assign cpu117_io_imem_instruction = imem117_io_pipeline_instruction; // @[top.scala 836:18]
  assign cpu117_io_dmem_readdata = dmem117_io_pipeline_readdata; // @[top.scala 837:18]
  assign mem117_clock = clock;
  assign mem117_reset = reset;
  assign mem117_io_imem_request_bits_address = imem117_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem117_io_dmem_request_valid = dmem117_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem117_io_dmem_request_bits_address = dmem117_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem117_io_dmem_request_bits_writedata = dmem117_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem117_io_dmem_request_bits_operation = dmem117_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem117_io_pipeline_address = cpu117_io_imem_address; // @[top.scala 836:18]
  assign imem117_io_bus_response_bits_data = mem117_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem117_clock = clock;
  assign dmem117_reset = reset;
  assign dmem117_io_pipeline_address = cpu117_io_dmem_address; // @[top.scala 837:18]
  assign dmem117_io_pipeline_valid = cpu117_io_dmem_valid; // @[top.scala 837:18]
  assign dmem117_io_pipeline_writedata = cpu117_io_dmem_writedata; // @[top.scala 837:18]
  assign dmem117_io_pipeline_memread = cpu117_io_dmem_memread; // @[top.scala 837:18]
  assign dmem117_io_pipeline_memwrite = cpu117_io_dmem_memwrite; // @[top.scala 837:18]
  assign dmem117_io_pipeline_maskmode = cpu117_io_dmem_maskmode; // @[top.scala 837:18]
  assign dmem117_io_pipeline_sext = cpu117_io_dmem_sext; // @[top.scala 837:18]
  assign dmem117_io_bus_response_valid = mem117_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem117_io_bus_response_bits_data = mem117_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu118_clock = clock;
  assign cpu118_reset = reset;
  assign cpu118_io_imem_instruction = imem118_io_pipeline_instruction; // @[top.scala 843:18]
  assign cpu118_io_dmem_readdata = dmem118_io_pipeline_readdata; // @[top.scala 844:18]
  assign mem118_clock = clock;
  assign mem118_reset = reset;
  assign mem118_io_imem_request_bits_address = imem118_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem118_io_dmem_request_valid = dmem118_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem118_io_dmem_request_bits_address = dmem118_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem118_io_dmem_request_bits_writedata = dmem118_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem118_io_dmem_request_bits_operation = dmem118_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem118_io_pipeline_address = cpu118_io_imem_address; // @[top.scala 843:18]
  assign imem118_io_bus_response_bits_data = mem118_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem118_clock = clock;
  assign dmem118_reset = reset;
  assign dmem118_io_pipeline_address = cpu118_io_dmem_address; // @[top.scala 844:18]
  assign dmem118_io_pipeline_valid = cpu118_io_dmem_valid; // @[top.scala 844:18]
  assign dmem118_io_pipeline_writedata = cpu118_io_dmem_writedata; // @[top.scala 844:18]
  assign dmem118_io_pipeline_memread = cpu118_io_dmem_memread; // @[top.scala 844:18]
  assign dmem118_io_pipeline_memwrite = cpu118_io_dmem_memwrite; // @[top.scala 844:18]
  assign dmem118_io_pipeline_maskmode = cpu118_io_dmem_maskmode; // @[top.scala 844:18]
  assign dmem118_io_pipeline_sext = cpu118_io_dmem_sext; // @[top.scala 844:18]
  assign dmem118_io_bus_response_valid = mem118_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem118_io_bus_response_bits_data = mem118_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu119_clock = clock;
  assign cpu119_reset = reset;
  assign cpu119_io_imem_instruction = imem119_io_pipeline_instruction; // @[top.scala 850:18]
  assign cpu119_io_dmem_readdata = dmem119_io_pipeline_readdata; // @[top.scala 851:18]
  assign mem119_clock = clock;
  assign mem119_reset = reset;
  assign mem119_io_imem_request_bits_address = imem119_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem119_io_dmem_request_valid = dmem119_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem119_io_dmem_request_bits_address = dmem119_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem119_io_dmem_request_bits_writedata = dmem119_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem119_io_dmem_request_bits_operation = dmem119_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem119_io_pipeline_address = cpu119_io_imem_address; // @[top.scala 850:18]
  assign imem119_io_bus_response_bits_data = mem119_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem119_clock = clock;
  assign dmem119_reset = reset;
  assign dmem119_io_pipeline_address = cpu119_io_dmem_address; // @[top.scala 851:18]
  assign dmem119_io_pipeline_valid = cpu119_io_dmem_valid; // @[top.scala 851:18]
  assign dmem119_io_pipeline_writedata = cpu119_io_dmem_writedata; // @[top.scala 851:18]
  assign dmem119_io_pipeline_memread = cpu119_io_dmem_memread; // @[top.scala 851:18]
  assign dmem119_io_pipeline_memwrite = cpu119_io_dmem_memwrite; // @[top.scala 851:18]
  assign dmem119_io_pipeline_maskmode = cpu119_io_dmem_maskmode; // @[top.scala 851:18]
  assign dmem119_io_pipeline_sext = cpu119_io_dmem_sext; // @[top.scala 851:18]
  assign dmem119_io_bus_response_valid = mem119_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem119_io_bus_response_bits_data = mem119_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu120_clock = clock;
  assign cpu120_reset = reset;
  assign cpu120_io_imem_instruction = imem120_io_pipeline_instruction; // @[top.scala 857:18]
  assign cpu120_io_dmem_readdata = dmem120_io_pipeline_readdata; // @[top.scala 858:18]
  assign mem120_clock = clock;
  assign mem120_reset = reset;
  assign mem120_io_imem_request_bits_address = imem120_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem120_io_dmem_request_valid = dmem120_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem120_io_dmem_request_bits_address = dmem120_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem120_io_dmem_request_bits_writedata = dmem120_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem120_io_dmem_request_bits_operation = dmem120_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem120_io_pipeline_address = cpu120_io_imem_address; // @[top.scala 857:18]
  assign imem120_io_bus_response_bits_data = mem120_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem120_clock = clock;
  assign dmem120_reset = reset;
  assign dmem120_io_pipeline_address = cpu120_io_dmem_address; // @[top.scala 858:18]
  assign dmem120_io_pipeline_valid = cpu120_io_dmem_valid; // @[top.scala 858:18]
  assign dmem120_io_pipeline_writedata = cpu120_io_dmem_writedata; // @[top.scala 858:18]
  assign dmem120_io_pipeline_memread = cpu120_io_dmem_memread; // @[top.scala 858:18]
  assign dmem120_io_pipeline_memwrite = cpu120_io_dmem_memwrite; // @[top.scala 858:18]
  assign dmem120_io_pipeline_maskmode = cpu120_io_dmem_maskmode; // @[top.scala 858:18]
  assign dmem120_io_pipeline_sext = cpu120_io_dmem_sext; // @[top.scala 858:18]
  assign dmem120_io_bus_response_valid = mem120_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem120_io_bus_response_bits_data = mem120_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu121_clock = clock;
  assign cpu121_reset = reset;
  assign cpu121_io_imem_instruction = imem121_io_pipeline_instruction; // @[top.scala 864:18]
  assign cpu121_io_dmem_readdata = dmem121_io_pipeline_readdata; // @[top.scala 865:18]
  assign mem121_clock = clock;
  assign mem121_reset = reset;
  assign mem121_io_imem_request_bits_address = imem121_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem121_io_dmem_request_valid = dmem121_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem121_io_dmem_request_bits_address = dmem121_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem121_io_dmem_request_bits_writedata = dmem121_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem121_io_dmem_request_bits_operation = dmem121_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem121_io_pipeline_address = cpu121_io_imem_address; // @[top.scala 864:18]
  assign imem121_io_bus_response_bits_data = mem121_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem121_clock = clock;
  assign dmem121_reset = reset;
  assign dmem121_io_pipeline_address = cpu121_io_dmem_address; // @[top.scala 865:18]
  assign dmem121_io_pipeline_valid = cpu121_io_dmem_valid; // @[top.scala 865:18]
  assign dmem121_io_pipeline_writedata = cpu121_io_dmem_writedata; // @[top.scala 865:18]
  assign dmem121_io_pipeline_memread = cpu121_io_dmem_memread; // @[top.scala 865:18]
  assign dmem121_io_pipeline_memwrite = cpu121_io_dmem_memwrite; // @[top.scala 865:18]
  assign dmem121_io_pipeline_maskmode = cpu121_io_dmem_maskmode; // @[top.scala 865:18]
  assign dmem121_io_pipeline_sext = cpu121_io_dmem_sext; // @[top.scala 865:18]
  assign dmem121_io_bus_response_valid = mem121_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem121_io_bus_response_bits_data = mem121_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu122_clock = clock;
  assign cpu122_reset = reset;
  assign cpu122_io_imem_instruction = imem122_io_pipeline_instruction; // @[top.scala 871:18]
  assign cpu122_io_dmem_readdata = dmem122_io_pipeline_readdata; // @[top.scala 872:18]
  assign mem122_clock = clock;
  assign mem122_reset = reset;
  assign mem122_io_imem_request_bits_address = imem122_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem122_io_dmem_request_valid = dmem122_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem122_io_dmem_request_bits_address = dmem122_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem122_io_dmem_request_bits_writedata = dmem122_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem122_io_dmem_request_bits_operation = dmem122_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem122_io_pipeline_address = cpu122_io_imem_address; // @[top.scala 871:18]
  assign imem122_io_bus_response_bits_data = mem122_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem122_clock = clock;
  assign dmem122_reset = reset;
  assign dmem122_io_pipeline_address = cpu122_io_dmem_address; // @[top.scala 872:18]
  assign dmem122_io_pipeline_valid = cpu122_io_dmem_valid; // @[top.scala 872:18]
  assign dmem122_io_pipeline_writedata = cpu122_io_dmem_writedata; // @[top.scala 872:18]
  assign dmem122_io_pipeline_memread = cpu122_io_dmem_memread; // @[top.scala 872:18]
  assign dmem122_io_pipeline_memwrite = cpu122_io_dmem_memwrite; // @[top.scala 872:18]
  assign dmem122_io_pipeline_maskmode = cpu122_io_dmem_maskmode; // @[top.scala 872:18]
  assign dmem122_io_pipeline_sext = cpu122_io_dmem_sext; // @[top.scala 872:18]
  assign dmem122_io_bus_response_valid = mem122_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem122_io_bus_response_bits_data = mem122_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu123_clock = clock;
  assign cpu123_reset = reset;
  assign cpu123_io_imem_instruction = imem123_io_pipeline_instruction; // @[top.scala 878:18]
  assign cpu123_io_dmem_readdata = dmem123_io_pipeline_readdata; // @[top.scala 879:18]
  assign mem123_clock = clock;
  assign mem123_reset = reset;
  assign mem123_io_imem_request_bits_address = imem123_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem123_io_dmem_request_valid = dmem123_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem123_io_dmem_request_bits_address = dmem123_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem123_io_dmem_request_bits_writedata = dmem123_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem123_io_dmem_request_bits_operation = dmem123_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem123_io_pipeline_address = cpu123_io_imem_address; // @[top.scala 878:18]
  assign imem123_io_bus_response_bits_data = mem123_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem123_clock = clock;
  assign dmem123_reset = reset;
  assign dmem123_io_pipeline_address = cpu123_io_dmem_address; // @[top.scala 879:18]
  assign dmem123_io_pipeline_valid = cpu123_io_dmem_valid; // @[top.scala 879:18]
  assign dmem123_io_pipeline_writedata = cpu123_io_dmem_writedata; // @[top.scala 879:18]
  assign dmem123_io_pipeline_memread = cpu123_io_dmem_memread; // @[top.scala 879:18]
  assign dmem123_io_pipeline_memwrite = cpu123_io_dmem_memwrite; // @[top.scala 879:18]
  assign dmem123_io_pipeline_maskmode = cpu123_io_dmem_maskmode; // @[top.scala 879:18]
  assign dmem123_io_pipeline_sext = cpu123_io_dmem_sext; // @[top.scala 879:18]
  assign dmem123_io_bus_response_valid = mem123_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem123_io_bus_response_bits_data = mem123_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu124_clock = clock;
  assign cpu124_reset = reset;
  assign cpu124_io_imem_instruction = imem124_io_pipeline_instruction; // @[top.scala 885:18]
  assign cpu124_io_dmem_readdata = dmem124_io_pipeline_readdata; // @[top.scala 886:18]
  assign mem124_clock = clock;
  assign mem124_reset = reset;
  assign mem124_io_imem_request_bits_address = imem124_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem124_io_dmem_request_valid = dmem124_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem124_io_dmem_request_bits_address = dmem124_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem124_io_dmem_request_bits_writedata = dmem124_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem124_io_dmem_request_bits_operation = dmem124_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem124_io_pipeline_address = cpu124_io_imem_address; // @[top.scala 885:18]
  assign imem124_io_bus_response_bits_data = mem124_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem124_clock = clock;
  assign dmem124_reset = reset;
  assign dmem124_io_pipeline_address = cpu124_io_dmem_address; // @[top.scala 886:18]
  assign dmem124_io_pipeline_valid = cpu124_io_dmem_valid; // @[top.scala 886:18]
  assign dmem124_io_pipeline_writedata = cpu124_io_dmem_writedata; // @[top.scala 886:18]
  assign dmem124_io_pipeline_memread = cpu124_io_dmem_memread; // @[top.scala 886:18]
  assign dmem124_io_pipeline_memwrite = cpu124_io_dmem_memwrite; // @[top.scala 886:18]
  assign dmem124_io_pipeline_maskmode = cpu124_io_dmem_maskmode; // @[top.scala 886:18]
  assign dmem124_io_pipeline_sext = cpu124_io_dmem_sext; // @[top.scala 886:18]
  assign dmem124_io_bus_response_valid = mem124_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem124_io_bus_response_bits_data = mem124_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu125_clock = clock;
  assign cpu125_reset = reset;
  assign cpu125_io_imem_instruction = imem125_io_pipeline_instruction; // @[top.scala 892:18]
  assign cpu125_io_dmem_readdata = dmem125_io_pipeline_readdata; // @[top.scala 893:18]
  assign mem125_clock = clock;
  assign mem125_reset = reset;
  assign mem125_io_imem_request_bits_address = imem125_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem125_io_dmem_request_valid = dmem125_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem125_io_dmem_request_bits_address = dmem125_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem125_io_dmem_request_bits_writedata = dmem125_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem125_io_dmem_request_bits_operation = dmem125_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem125_io_pipeline_address = cpu125_io_imem_address; // @[top.scala 892:18]
  assign imem125_io_bus_response_bits_data = mem125_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem125_clock = clock;
  assign dmem125_reset = reset;
  assign dmem125_io_pipeline_address = cpu125_io_dmem_address; // @[top.scala 893:18]
  assign dmem125_io_pipeline_valid = cpu125_io_dmem_valid; // @[top.scala 893:18]
  assign dmem125_io_pipeline_writedata = cpu125_io_dmem_writedata; // @[top.scala 893:18]
  assign dmem125_io_pipeline_memread = cpu125_io_dmem_memread; // @[top.scala 893:18]
  assign dmem125_io_pipeline_memwrite = cpu125_io_dmem_memwrite; // @[top.scala 893:18]
  assign dmem125_io_pipeline_maskmode = cpu125_io_dmem_maskmode; // @[top.scala 893:18]
  assign dmem125_io_pipeline_sext = cpu125_io_dmem_sext; // @[top.scala 893:18]
  assign dmem125_io_bus_response_valid = mem125_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem125_io_bus_response_bits_data = mem125_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu126_clock = clock;
  assign cpu126_reset = reset;
  assign cpu126_io_imem_instruction = imem126_io_pipeline_instruction; // @[top.scala 899:18]
  assign cpu126_io_dmem_readdata = dmem126_io_pipeline_readdata; // @[top.scala 900:18]
  assign mem126_clock = clock;
  assign mem126_reset = reset;
  assign mem126_io_imem_request_bits_address = imem126_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem126_io_dmem_request_valid = dmem126_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem126_io_dmem_request_bits_address = dmem126_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem126_io_dmem_request_bits_writedata = dmem126_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem126_io_dmem_request_bits_operation = dmem126_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem126_io_pipeline_address = cpu126_io_imem_address; // @[top.scala 899:18]
  assign imem126_io_bus_response_bits_data = mem126_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem126_clock = clock;
  assign dmem126_reset = reset;
  assign dmem126_io_pipeline_address = cpu126_io_dmem_address; // @[top.scala 900:18]
  assign dmem126_io_pipeline_valid = cpu126_io_dmem_valid; // @[top.scala 900:18]
  assign dmem126_io_pipeline_writedata = cpu126_io_dmem_writedata; // @[top.scala 900:18]
  assign dmem126_io_pipeline_memread = cpu126_io_dmem_memread; // @[top.scala 900:18]
  assign dmem126_io_pipeline_memwrite = cpu126_io_dmem_memwrite; // @[top.scala 900:18]
  assign dmem126_io_pipeline_maskmode = cpu126_io_dmem_maskmode; // @[top.scala 900:18]
  assign dmem126_io_pipeline_sext = cpu126_io_dmem_sext; // @[top.scala 900:18]
  assign dmem126_io_bus_response_valid = mem126_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem126_io_bus_response_bits_data = mem126_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
  assign cpu127_clock = clock;
  assign cpu127_reset = reset;
  assign cpu127_io_imem_instruction = imem127_io_pipeline_instruction; // @[top.scala 906:18]
  assign cpu127_io_dmem_readdata = dmem127_io_pipeline_readdata; // @[top.scala 907:18]
  assign mem127_clock = clock;
  assign mem127_reset = reset;
  assign mem127_io_imem_request_bits_address = imem127_io_bus_request_bits_address; // @[base-memory-components.scala 16:26]
  assign mem127_io_dmem_request_valid = dmem127_io_bus_request_valid; // @[base-memory-components.scala 19:26]
  assign mem127_io_dmem_request_bits_address = dmem127_io_bus_request_bits_address; // @[base-memory-components.scala 19:26]
  assign mem127_io_dmem_request_bits_writedata = dmem127_io_bus_request_bits_writedata; // @[base-memory-components.scala 19:26]
  assign mem127_io_dmem_request_bits_operation = dmem127_io_bus_request_bits_operation; // @[base-memory-components.scala 19:26]
  assign imem127_io_pipeline_address = cpu127_io_imem_address; // @[top.scala 906:18]
  assign imem127_io_bus_response_bits_data = mem127_io_imem_response_bits_data; // @[base-memory-components.scala 17:26]
  assign dmem127_clock = clock;
  assign dmem127_reset = reset;
  assign dmem127_io_pipeline_address = cpu127_io_dmem_address; // @[top.scala 907:18]
  assign dmem127_io_pipeline_valid = cpu127_io_dmem_valid; // @[top.scala 907:18]
  assign dmem127_io_pipeline_writedata = cpu127_io_dmem_writedata; // @[top.scala 907:18]
  assign dmem127_io_pipeline_memread = cpu127_io_dmem_memread; // @[top.scala 907:18]
  assign dmem127_io_pipeline_memwrite = cpu127_io_dmem_memwrite; // @[top.scala 907:18]
  assign dmem127_io_pipeline_maskmode = cpu127_io_dmem_maskmode; // @[top.scala 907:18]
  assign dmem127_io_pipeline_sext = cpu127_io_dmem_sext; // @[top.scala 907:18]
  assign dmem127_io_bus_response_valid = mem127_io_dmem_response_valid; // @[base-memory-components.scala 20:26]
  assign dmem127_io_bus_response_bits_data = mem127_io_dmem_response_bits_data; // @[base-memory-components.scala 20:26]
endmodule
