`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Rob(
  input         clock,
  input         reset,
  input         io_enq_valids_0,
  input         io_enq_valids_1,
  input  [39:0] io_enq_uops_0_pc,
  input  [7:0]  io_enq_uops_0_br_mask,
  input  [6:0]  io_enq_uops_0_rob_idx,
  input  [5:0]  io_enq_uops_0_brob_idx,
  input  [6:0]  io_enq_uops_0_pdst,
  input  [6:0]  io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_is_fence,
  input         io_enq_uops_0_is_fencei,
  input         io_enq_uops_0_is_store,
  input         io_enq_uops_0_is_load,
  input         io_enq_uops_0_is_sys_pc2epc,
  input         io_enq_uops_0_is_unique,
  input         io_enq_uops_0_flush_on_commit,
  input  [5:0]  io_enq_uops_0_ldst,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input         io_enq_uops_0_fp_val,
  input  [7:0]  io_enq_uops_1_br_mask,
  input  [6:0]  io_enq_uops_1_rob_idx,
  input  [6:0]  io_enq_uops_1_pdst,
  input  [6:0]  io_enq_uops_1_stale_pdst,
  input         io_enq_uops_1_exception,
  input  [63:0] io_enq_uops_1_exc_cause,
  input         io_enq_uops_1_is_fence,
  input         io_enq_uops_1_is_fencei,
  input         io_enq_uops_1_is_store,
  input         io_enq_uops_1_is_load,
  input         io_enq_uops_1_is_sys_pc2epc,
  input         io_enq_uops_1_is_unique,
  input         io_enq_uops_1_flush_on_commit,
  input  [5:0]  io_enq_uops_1_ldst,
  input         io_enq_uops_1_ldst_val,
  input  [1:0]  io_enq_uops_1_dst_rtype,
  input         io_enq_uops_1_fp_val,
  input         io_enq_has_br_or_jalr_in_packet,
  input         io_enq_partial_stall,
  input         io_enq_new_packet,
  output [6:0]  io_curr_rob_tail,
  input         io_brinfo_valid,
  input         io_brinfo_mispredict,
  input  [7:0]  io_brinfo_mask,
  input  [6:0]  io_brinfo_rob_idx,
  input  [6:0]  io_get_pc_rob_idx,
  output [39:0] io_get_pc_curr_pc,
  output [5:0]  io_get_pc_curr_brob_idx,
  output        io_get_pc_next_val,
  output [39:0] io_get_pc_next_pc,
  input         io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_rob_idx,
  input  [6:0]  io_wb_resps_0_bits_uop_pdst,
  input         io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_rob_idx,
  input  [6:0]  io_wb_resps_1_bits_uop_pdst,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_rob_idx,
  input  [6:0]  io_wb_resps_2_bits_uop_pdst,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_rob_idx,
  input  [6:0]  io_wb_resps_3_bits_uop_pdst,
  input         io_wb_resps_4_valid,
  input  [6:0]  io_wb_resps_4_bits_uop_rob_idx,
  input  [6:0]  io_wb_resps_4_bits_uop_pdst,
  input         io_lsu_clr_bsy_valid_0,
  input         io_lsu_clr_bsy_valid_1,
  input  [6:0]  io_lsu_clr_bsy_rob_idx_0,
  input  [6:0]  io_lsu_clr_bsy_rob_idx_1,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_rob_idx,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_1_valid,
  input  [6:0]  io_fflags_1_bits_uop_rob_idx,
  input  [4:0]  io_fflags_1_bits_flags,
  input         io_lxcpt_valid,
  input  [7:0]  io_lxcpt_bits_uop_br_mask,
  input  [6:0]  io_lxcpt_bits_uop_rob_idx,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_bxcpt_valid,
  input  [7:0]  io_bxcpt_bits_uop_br_mask,
  input  [6:0]  io_bxcpt_bits_uop_rob_idx,
  input  [39:0] io_bxcpt_bits_badvaddr,
  output        io_commit_valids_0,
  output        io_commit_valids_1,
  output [6:0]  io_commit_uops_0_pdst,
  output [6:0]  io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_is_fencei,
  output        io_commit_uops_0_is_store,
  output        io_commit_uops_0_is_load,
  output        io_commit_uops_0_is_sys_pc2epc,
  output        io_commit_uops_0_flush_on_commit,
  output [5:0]  io_commit_uops_0_ldst,
  output [1:0]  io_commit_uops_0_dst_rtype,
  output        io_commit_uops_0_fp_val,
  output [6:0]  io_commit_uops_1_pdst,
  output [6:0]  io_commit_uops_1_stale_pdst,
  output        io_commit_uops_1_is_fencei,
  output        io_commit_uops_1_is_store,
  output        io_commit_uops_1_is_load,
  output        io_commit_uops_1_is_sys_pc2epc,
  output        io_commit_uops_1_flush_on_commit,
  output [5:0]  io_commit_uops_1_ldst,
  output [1:0]  io_commit_uops_1_dst_rtype,
  output        io_commit_uops_1_fp_val,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output        io_commit_rbk_valids_0,
  output        io_commit_rbk_valids_1,
  output        io_commit_st_mask_0,
  output        io_commit_st_mask_1,
  output        io_commit_ld_mask_0,
  output        io_commit_ld_mask_1,
  output        io_com_load_is_at_rob_head,
  output        io_com_xcpt_valid,
  output [63:0] io_com_xcpt_bits_pc,
  output [63:0] io_com_xcpt_bits_cause,
  output [63:0] io_com_xcpt_bits_badvaddr,
  input         io_csr_eret,
  input  [39:0] io_csr_evec,
  input         io_csr_stall,
  output        io_flush_valid,
  output [63:0] io_flush_bits_pc,
  output        io_clear_brob,
  output        io_empty,
  output        io_ready,
  output        io_brob_deallocate_valid,
  output [5:0]  io_brob_deallocate_bits_brob_idx
);
  reg [1:0] rob_state;
  reg [31:0] _RAND_0;
  reg [5:0] rob_head;
  reg [31:0] _RAND_1;
  reg [5:0] rob_tail;
  reg [31:0] _RAND_2;
  wire [6:0] _GEN_421;
  wire [6:0] rob_tail_idx;
  wire  will_commit_0;
  wire  will_commit_1;
  wire  can_commit_0;
  wire  can_commit_1;
  wire  can_throw_exception_0;
  wire  can_throw_exception_1;
  wire  rob_head_vals_0;
  wire  rob_head_vals_1;
  wire  rob_head_is_store_0;
  wire  rob_head_is_store_1;
  wire  rob_head_is_load_0;
  wire  rob_head_is_load_1;
  wire [4:0] rob_head_fflags_0;
  wire [4:0] rob_head_fflags_1;
  wire  rob_getpc_next_vals_0;
  wire  rob_getpc_next_vals_1;
  wire  rob_getpc_curr_vals_0;
  wire  rob_getpc_curr_vals_1;
  wire  exception_thrown;
  reg  r_xcpt_val;
  reg [31:0] _RAND_3;
  reg [7:0] r_xcpt_uop_br_mask;
  reg [31:0] _RAND_4;
  reg [6:0] r_xcpt_uop_rob_idx;
  reg [31:0] _RAND_5;
  reg [63:0] r_xcpt_uop_exc_cause;
  reg [63:0] _RAND_6;
  reg [63:0] r_xcpt_badvaddr;
  reg [63:0] _RAND_7;
  reg [36:0] _T_2772 [0:19];
  reg [63:0] _RAND_8;
  wire [36:0] _T_2772__T_2805_data;
  wire [4:0] _T_2772__T_2805_addr;
  reg [63:0] _RAND_9;
  wire [36:0] _T_2772__T_8084_data;
  wire [4:0] _T_2772__T_8084_addr;
  reg [63:0] _RAND_10;
  wire [36:0] _T_2772__T_2788_data;
  wire [4:0] _T_2772__T_2788_addr;
  wire  _T_2772__T_2788_mask;
  wire  _T_2772__T_2788_en;
  wire [36:0] _GEN_112;
  reg [36:0] _T_2775 [0:19];
  reg [63:0] _RAND_11;
  wire [36:0] _T_2775__T_2811_data;
  wire [4:0] _T_2775__T_2811_addr;
  reg [63:0] _RAND_12;
  wire [36:0] _T_2775__T_8091_data;
  wire [4:0] _T_2775__T_8091_addr;
  reg [63:0] _RAND_13;
  wire [36:0] _T_2775__T_2784_data;
  wire [4:0] _T_2775__T_2784_addr;
  wire  _T_2775__T_2784_mask;
  wire  _T_2775__T_2784_en;
  wire  _T_2776;
  wire [39:0] _T_2779;
  wire  _T_2780;
  wire [5:0] _T_2782;
  wire [4:0] _T_2783;
  wire [4:0] _T_2787;
  wire  _GEN_553;
  wire  _GEN_557;
  wire  _GEN_561;
  wire [6:0] _T_2790;
  wire  _T_2791;
  wire [6:0] _T_2793;
  wire  _T_2795;
  wire [7:0] _T_2798;
  wire [6:0] _T_2799;
  wire [6:0] _T_2800;
  wire [6:0] _T_2803;
  wire [4:0] _T_2804;
  wire [39:0] _GEN_423;
  wire [39:0] _T_2807;
  wire [4:0] _T_2810;
  wire [39:0] _GEN_424;
  wire [39:0] _T_2813;
  wire [63:0] _T_2815;
  wire [63:0] _T_2817;
  wire [39:0] _T_2819;
  wire [39:0] _T_2821;
  wire [39:0] _T_2822;
  wire  _T_2823;
  wire [23:0] _T_2827;
  wire [63:0] curr_row_pc;
  wire [39:0] _T_2828;
  wire  _T_2829;
  wire [23:0] _T_2833;
  wire [63:0] next_row_pc;
  wire  _T_2834;
  wire [2:0] _T_2836;
  wire [63:0] _GEN_428;
  wire [64:0] _T_2837;
  wire [63:0] _T_2838;
  wire [1:0] _T_2841;
  wire  curr_idx;
  wire  curr_row_next_pc_val;
  wire  _GEN_0;
  wire  _GEN_563;
  wire  _T_2846;
  wire [2:0] _T_2848;
  wire [63:0] _GEN_429;
  wire [64:0] _T_2849;
  wire [63:0] curr_row_next_pc;
  wire [1:0] _T_2850;
  wire  _T_2851;
  wire  next_bank_idx;
  wire  rob_pc_hob_next_val;
  wire [1:0] _T_2855;
  wire  _T_2856;
  wire  bypass_next_bank_idx;
  wire [39:0] _T_2860;
  wire [39:0] _T_2862;
  wire [39:0] _T_2863;
  wire [39:0] _T_2864;
  wire [2:0] _T_2866;
  wire [39:0] _GEN_436;
  wire [40:0] _T_2867;
  wire [39:0] bypass_next_pc;
  wire  _T_2869;
  wire  _T_2870;
  wire [2:0] _T_2872;
  wire [63:0] _GEN_437;
  wire [64:0] _T_2873;
  wire [63:0] _T_2874;
  wire [63:0] _T_2875;
  wire [63:0] _T_2876;
  wire  finished_committing_row;
  reg  r_partial_row;
  reg [31:0] _RAND_14;
  reg [5:0] row_metadata_brob_idx [0:39];
  reg [31:0] _RAND_15;
  wire [5:0] row_metadata_brob_idx__T_2896_data;
  wire [5:0] row_metadata_brob_idx__T_2896_addr;
  reg [31:0] _RAND_16;
  wire [5:0] row_metadata_brob_idx__T_2900_data;
  wire [5:0] row_metadata_brob_idx__T_2900_addr;
  reg [31:0] _RAND_17;
  wire [5:0] row_metadata_brob_idx__T_2886_data;
  wire [5:0] row_metadata_brob_idx__T_2886_addr;
  wire  row_metadata_brob_idx__T_2886_mask;
  wire  row_metadata_brob_idx__T_2886_en;
  reg  row_metadata_has_brorjalr [0:39];
  reg [31:0] _RAND_18;
  wire  row_metadata_has_brorjalr__T_2894_data;
  wire [5:0] row_metadata_has_brorjalr__T_2894_addr;
  reg [31:0] _RAND_19;
  wire  row_metadata_has_brorjalr__T_2887_data;
  wire [5:0] row_metadata_has_brorjalr__T_2887_addr;
  wire  row_metadata_has_brorjalr__T_2887_mask;
  wire  row_metadata_has_brorjalr__T_2887_en;
  wire  row_metadata_has_brorjalr__T_2892_data;
  wire [5:0] row_metadata_has_brorjalr__T_2892_addr;
  wire  row_metadata_has_brorjalr__T_2892_mask;
  wire  row_metadata_has_brorjalr__T_2892_en;
  wire  _T_2885;
  wire  _T_2890;
  wire  _T_2891;
  wire  _GEN_564;
  wire  _GEN_570;
  wire  _T_2895;
  wire [5:0] _T_2899;
  wire  _T_2901;
  wire  _T_2902;
  wire  _T_2903;
  reg  _T_3073_0;
  reg [31:0] _RAND_20;
  reg  _T_3073_1;
  reg [31:0] _RAND_21;
  reg  _T_3073_2;
  reg [31:0] _RAND_22;
  reg  _T_3073_3;
  reg [31:0] _RAND_23;
  reg  _T_3073_4;
  reg [31:0] _RAND_24;
  reg  _T_3073_5;
  reg [31:0] _RAND_25;
  reg  _T_3073_6;
  reg [31:0] _RAND_26;
  reg  _T_3073_7;
  reg [31:0] _RAND_27;
  reg  _T_3073_8;
  reg [31:0] _RAND_28;
  reg  _T_3073_9;
  reg [31:0] _RAND_29;
  reg  _T_3073_10;
  reg [31:0] _RAND_30;
  reg  _T_3073_11;
  reg [31:0] _RAND_31;
  reg  _T_3073_12;
  reg [31:0] _RAND_32;
  reg  _T_3073_13;
  reg [31:0] _RAND_33;
  reg  _T_3073_14;
  reg [31:0] _RAND_34;
  reg  _T_3073_15;
  reg [31:0] _RAND_35;
  reg  _T_3073_16;
  reg [31:0] _RAND_36;
  reg  _T_3073_17;
  reg [31:0] _RAND_37;
  reg  _T_3073_18;
  reg [31:0] _RAND_38;
  reg  _T_3073_19;
  reg [31:0] _RAND_39;
  reg  _T_3073_20;
  reg [31:0] _RAND_40;
  reg  _T_3073_21;
  reg [31:0] _RAND_41;
  reg  _T_3073_22;
  reg [31:0] _RAND_42;
  reg  _T_3073_23;
  reg [31:0] _RAND_43;
  reg  _T_3073_24;
  reg [31:0] _RAND_44;
  reg  _T_3073_25;
  reg [31:0] _RAND_45;
  reg  _T_3073_26;
  reg [31:0] _RAND_46;
  reg  _T_3073_27;
  reg [31:0] _RAND_47;
  reg  _T_3073_28;
  reg [31:0] _RAND_48;
  reg  _T_3073_29;
  reg [31:0] _RAND_49;
  reg  _T_3073_30;
  reg [31:0] _RAND_50;
  reg  _T_3073_31;
  reg [31:0] _RAND_51;
  reg  _T_3073_32;
  reg [31:0] _RAND_52;
  reg  _T_3073_33;
  reg [31:0] _RAND_53;
  reg  _T_3073_34;
  reg [31:0] _RAND_54;
  reg  _T_3073_35;
  reg [31:0] _RAND_55;
  reg  _T_3073_36;
  reg [31:0] _RAND_56;
  reg  _T_3073_37;
  reg [31:0] _RAND_57;
  reg  _T_3073_38;
  reg [31:0] _RAND_58;
  reg  _T_3073_39;
  reg [31:0] _RAND_59;
  reg  _T_3200 [0:39];
  reg [31:0] _RAND_60;
  wire  _T_3200__T_3877_data;
  wire [5:0] _T_3200__T_3877_addr;
  reg [31:0] _RAND_61;
  wire  _T_3200__T_3904_data;
  wire [5:0] _T_3200__T_3904_addr;
  reg [31:0] _RAND_62;
  wire  _T_3200__T_4017_data;
  wire [5:0] _T_3200__T_4017_addr;
  reg [31:0] _RAND_63;
  wire  _T_3200__T_5128_data;
  wire [5:0] _T_3200__T_5128_addr;
  reg [31:0] _RAND_64;
  wire  _T_3200__T_5205_data;
  wire [5:0] _T_3200__T_5205_addr;
  reg [31:0] _RAND_65;
  wire  _T_3200__T_5282_data;
  wire [5:0] _T_3200__T_5282_addr;
  reg [31:0] _RAND_66;
  wire  _T_3200__T_5359_data;
  wire [5:0] _T_3200__T_5359_addr;
  reg [31:0] _RAND_67;
  wire  _T_3200__T_5436_data;
  wire [5:0] _T_3200__T_5436_addr;
  reg [31:0] _RAND_68;
  wire  _T_3200__T_3753_data;
  wire [5:0] _T_3200__T_3753_addr;
  wire  _T_3200__T_3753_mask;
  wire  _T_3200__T_3753_en;
  wire  _T_3200__T_3819_data;
  wire [5:0] _T_3200__T_3819_addr;
  wire  _T_3200__T_3819_mask;
  wire  _T_3200__T_3819_en;
  wire  _T_3200__T_3828_data;
  wire [5:0] _T_3200__T_3828_addr;
  wire  _T_3200__T_3828_mask;
  wire  _T_3200__T_3828_en;
  wire  _T_3200__T_3837_data;
  wire [5:0] _T_3200__T_3837_addr;
  wire  _T_3200__T_3837_mask;
  wire  _T_3200__T_3837_en;
  wire  _T_3200__T_3846_data;
  wire [5:0] _T_3200__T_3846_addr;
  wire  _T_3200__T_3846_mask;
  wire  _T_3200__T_3846_en;
  wire  _T_3200__T_3855_data;
  wire [5:0] _T_3200__T_3855_addr;
  wire  _T_3200__T_3855_mask;
  wire  _T_3200__T_3855_en;
  wire  _T_3200__T_3864_data;
  wire [5:0] _T_3200__T_3864_addr;
  wire  _T_3200__T_3864_mask;
  wire  _T_3200__T_3864_en;
  wire  _T_3200__T_3891_data;
  wire [5:0] _T_3200__T_3891_addr;
  wire  _T_3200__T_3891_mask;
  wire  _T_3200__T_3891_en;
  reg [7:0] _T_3372_0_br_mask;
  reg [31:0] _RAND_69;
  reg [6:0] _T_3372_0_pdst;
  reg [31:0] _RAND_70;
  reg [6:0] _T_3372_0_stale_pdst;
  reg [31:0] _RAND_71;
  reg  _T_3372_0_is_fencei;
  reg [31:0] _RAND_72;
  reg  _T_3372_0_is_store;
  reg [31:0] _RAND_73;
  reg  _T_3372_0_is_load;
  reg [31:0] _RAND_74;
  reg  _T_3372_0_is_sys_pc2epc;
  reg [31:0] _RAND_75;
  reg  _T_3372_0_flush_on_commit;
  reg [31:0] _RAND_76;
  reg [5:0] _T_3372_0_ldst;
  reg [31:0] _RAND_77;
  reg  _T_3372_0_ldst_val;
  reg [31:0] _RAND_78;
  reg [1:0] _T_3372_0_dst_rtype;
  reg [31:0] _RAND_79;
  reg  _T_3372_0_fp_val;
  reg [31:0] _RAND_80;
  reg [7:0] _T_3372_1_br_mask;
  reg [31:0] _RAND_81;
  reg [6:0] _T_3372_1_pdst;
  reg [31:0] _RAND_82;
  reg [6:0] _T_3372_1_stale_pdst;
  reg [31:0] _RAND_83;
  reg  _T_3372_1_is_fencei;
  reg [31:0] _RAND_84;
  reg  _T_3372_1_is_store;
  reg [31:0] _RAND_85;
  reg  _T_3372_1_is_load;
  reg [31:0] _RAND_86;
  reg  _T_3372_1_is_sys_pc2epc;
  reg [31:0] _RAND_87;
  reg  _T_3372_1_flush_on_commit;
  reg [31:0] _RAND_88;
  reg [5:0] _T_3372_1_ldst;
  reg [31:0] _RAND_89;
  reg  _T_3372_1_ldst_val;
  reg [31:0] _RAND_90;
  reg [1:0] _T_3372_1_dst_rtype;
  reg [31:0] _RAND_91;
  reg  _T_3372_1_fp_val;
  reg [31:0] _RAND_92;
  reg [7:0] _T_3372_2_br_mask;
  reg [31:0] _RAND_93;
  reg [6:0] _T_3372_2_pdst;
  reg [31:0] _RAND_94;
  reg [6:0] _T_3372_2_stale_pdst;
  reg [31:0] _RAND_95;
  reg  _T_3372_2_is_fencei;
  reg [31:0] _RAND_96;
  reg  _T_3372_2_is_store;
  reg [31:0] _RAND_97;
  reg  _T_3372_2_is_load;
  reg [31:0] _RAND_98;
  reg  _T_3372_2_is_sys_pc2epc;
  reg [31:0] _RAND_99;
  reg  _T_3372_2_flush_on_commit;
  reg [31:0] _RAND_100;
  reg [5:0] _T_3372_2_ldst;
  reg [31:0] _RAND_101;
  reg  _T_3372_2_ldst_val;
  reg [31:0] _RAND_102;
  reg [1:0] _T_3372_2_dst_rtype;
  reg [31:0] _RAND_103;
  reg  _T_3372_2_fp_val;
  reg [31:0] _RAND_104;
  reg [7:0] _T_3372_3_br_mask;
  reg [31:0] _RAND_105;
  reg [6:0] _T_3372_3_pdst;
  reg [31:0] _RAND_106;
  reg [6:0] _T_3372_3_stale_pdst;
  reg [31:0] _RAND_107;
  reg  _T_3372_3_is_fencei;
  reg [31:0] _RAND_108;
  reg  _T_3372_3_is_store;
  reg [31:0] _RAND_109;
  reg  _T_3372_3_is_load;
  reg [31:0] _RAND_110;
  reg  _T_3372_3_is_sys_pc2epc;
  reg [31:0] _RAND_111;
  reg  _T_3372_3_flush_on_commit;
  reg [31:0] _RAND_112;
  reg [5:0] _T_3372_3_ldst;
  reg [31:0] _RAND_113;
  reg  _T_3372_3_ldst_val;
  reg [31:0] _RAND_114;
  reg [1:0] _T_3372_3_dst_rtype;
  reg [31:0] _RAND_115;
  reg  _T_3372_3_fp_val;
  reg [31:0] _RAND_116;
  reg [7:0] _T_3372_4_br_mask;
  reg [31:0] _RAND_117;
  reg [6:0] _T_3372_4_pdst;
  reg [31:0] _RAND_118;
  reg [6:0] _T_3372_4_stale_pdst;
  reg [31:0] _RAND_119;
  reg  _T_3372_4_is_fencei;
  reg [31:0] _RAND_120;
  reg  _T_3372_4_is_store;
  reg [31:0] _RAND_121;
  reg  _T_3372_4_is_load;
  reg [31:0] _RAND_122;
  reg  _T_3372_4_is_sys_pc2epc;
  reg [31:0] _RAND_123;
  reg  _T_3372_4_flush_on_commit;
  reg [31:0] _RAND_124;
  reg [5:0] _T_3372_4_ldst;
  reg [31:0] _RAND_125;
  reg  _T_3372_4_ldst_val;
  reg [31:0] _RAND_126;
  reg [1:0] _T_3372_4_dst_rtype;
  reg [31:0] _RAND_127;
  reg  _T_3372_4_fp_val;
  reg [31:0] _RAND_128;
  reg [7:0] _T_3372_5_br_mask;
  reg [31:0] _RAND_129;
  reg [6:0] _T_3372_5_pdst;
  reg [31:0] _RAND_130;
  reg [6:0] _T_3372_5_stale_pdst;
  reg [31:0] _RAND_131;
  reg  _T_3372_5_is_fencei;
  reg [31:0] _RAND_132;
  reg  _T_3372_5_is_store;
  reg [31:0] _RAND_133;
  reg  _T_3372_5_is_load;
  reg [31:0] _RAND_134;
  reg  _T_3372_5_is_sys_pc2epc;
  reg [31:0] _RAND_135;
  reg  _T_3372_5_flush_on_commit;
  reg [31:0] _RAND_136;
  reg [5:0] _T_3372_5_ldst;
  reg [31:0] _RAND_137;
  reg  _T_3372_5_ldst_val;
  reg [31:0] _RAND_138;
  reg [1:0] _T_3372_5_dst_rtype;
  reg [31:0] _RAND_139;
  reg  _T_3372_5_fp_val;
  reg [31:0] _RAND_140;
  reg [7:0] _T_3372_6_br_mask;
  reg [31:0] _RAND_141;
  reg [6:0] _T_3372_6_pdst;
  reg [31:0] _RAND_142;
  reg [6:0] _T_3372_6_stale_pdst;
  reg [31:0] _RAND_143;
  reg  _T_3372_6_is_fencei;
  reg [31:0] _RAND_144;
  reg  _T_3372_6_is_store;
  reg [31:0] _RAND_145;
  reg  _T_3372_6_is_load;
  reg [31:0] _RAND_146;
  reg  _T_3372_6_is_sys_pc2epc;
  reg [31:0] _RAND_147;
  reg  _T_3372_6_flush_on_commit;
  reg [31:0] _RAND_148;
  reg [5:0] _T_3372_6_ldst;
  reg [31:0] _RAND_149;
  reg  _T_3372_6_ldst_val;
  reg [31:0] _RAND_150;
  reg [1:0] _T_3372_6_dst_rtype;
  reg [31:0] _RAND_151;
  reg  _T_3372_6_fp_val;
  reg [31:0] _RAND_152;
  reg [7:0] _T_3372_7_br_mask;
  reg [31:0] _RAND_153;
  reg [6:0] _T_3372_7_pdst;
  reg [31:0] _RAND_154;
  reg [6:0] _T_3372_7_stale_pdst;
  reg [31:0] _RAND_155;
  reg  _T_3372_7_is_fencei;
  reg [31:0] _RAND_156;
  reg  _T_3372_7_is_store;
  reg [31:0] _RAND_157;
  reg  _T_3372_7_is_load;
  reg [31:0] _RAND_158;
  reg  _T_3372_7_is_sys_pc2epc;
  reg [31:0] _RAND_159;
  reg  _T_3372_7_flush_on_commit;
  reg [31:0] _RAND_160;
  reg [5:0] _T_3372_7_ldst;
  reg [31:0] _RAND_161;
  reg  _T_3372_7_ldst_val;
  reg [31:0] _RAND_162;
  reg [1:0] _T_3372_7_dst_rtype;
  reg [31:0] _RAND_163;
  reg  _T_3372_7_fp_val;
  reg [31:0] _RAND_164;
  reg [7:0] _T_3372_8_br_mask;
  reg [31:0] _RAND_165;
  reg [6:0] _T_3372_8_pdst;
  reg [31:0] _RAND_166;
  reg [6:0] _T_3372_8_stale_pdst;
  reg [31:0] _RAND_167;
  reg  _T_3372_8_is_fencei;
  reg [31:0] _RAND_168;
  reg  _T_3372_8_is_store;
  reg [31:0] _RAND_169;
  reg  _T_3372_8_is_load;
  reg [31:0] _RAND_170;
  reg  _T_3372_8_is_sys_pc2epc;
  reg [31:0] _RAND_171;
  reg  _T_3372_8_flush_on_commit;
  reg [31:0] _RAND_172;
  reg [5:0] _T_3372_8_ldst;
  reg [31:0] _RAND_173;
  reg  _T_3372_8_ldst_val;
  reg [31:0] _RAND_174;
  reg [1:0] _T_3372_8_dst_rtype;
  reg [31:0] _RAND_175;
  reg  _T_3372_8_fp_val;
  reg [31:0] _RAND_176;
  reg [7:0] _T_3372_9_br_mask;
  reg [31:0] _RAND_177;
  reg [6:0] _T_3372_9_pdst;
  reg [31:0] _RAND_178;
  reg [6:0] _T_3372_9_stale_pdst;
  reg [31:0] _RAND_179;
  reg  _T_3372_9_is_fencei;
  reg [31:0] _RAND_180;
  reg  _T_3372_9_is_store;
  reg [31:0] _RAND_181;
  reg  _T_3372_9_is_load;
  reg [31:0] _RAND_182;
  reg  _T_3372_9_is_sys_pc2epc;
  reg [31:0] _RAND_183;
  reg  _T_3372_9_flush_on_commit;
  reg [31:0] _RAND_184;
  reg [5:0] _T_3372_9_ldst;
  reg [31:0] _RAND_185;
  reg  _T_3372_9_ldst_val;
  reg [31:0] _RAND_186;
  reg [1:0] _T_3372_9_dst_rtype;
  reg [31:0] _RAND_187;
  reg  _T_3372_9_fp_val;
  reg [31:0] _RAND_188;
  reg [7:0] _T_3372_10_br_mask;
  reg [31:0] _RAND_189;
  reg [6:0] _T_3372_10_pdst;
  reg [31:0] _RAND_190;
  reg [6:0] _T_3372_10_stale_pdst;
  reg [31:0] _RAND_191;
  reg  _T_3372_10_is_fencei;
  reg [31:0] _RAND_192;
  reg  _T_3372_10_is_store;
  reg [31:0] _RAND_193;
  reg  _T_3372_10_is_load;
  reg [31:0] _RAND_194;
  reg  _T_3372_10_is_sys_pc2epc;
  reg [31:0] _RAND_195;
  reg  _T_3372_10_flush_on_commit;
  reg [31:0] _RAND_196;
  reg [5:0] _T_3372_10_ldst;
  reg [31:0] _RAND_197;
  reg  _T_3372_10_ldst_val;
  reg [31:0] _RAND_198;
  reg [1:0] _T_3372_10_dst_rtype;
  reg [31:0] _RAND_199;
  reg  _T_3372_10_fp_val;
  reg [31:0] _RAND_200;
  reg [7:0] _T_3372_11_br_mask;
  reg [31:0] _RAND_201;
  reg [6:0] _T_3372_11_pdst;
  reg [31:0] _RAND_202;
  reg [6:0] _T_3372_11_stale_pdst;
  reg [31:0] _RAND_203;
  reg  _T_3372_11_is_fencei;
  reg [31:0] _RAND_204;
  reg  _T_3372_11_is_store;
  reg [31:0] _RAND_205;
  reg  _T_3372_11_is_load;
  reg [31:0] _RAND_206;
  reg  _T_3372_11_is_sys_pc2epc;
  reg [31:0] _RAND_207;
  reg  _T_3372_11_flush_on_commit;
  reg [31:0] _RAND_208;
  reg [5:0] _T_3372_11_ldst;
  reg [31:0] _RAND_209;
  reg  _T_3372_11_ldst_val;
  reg [31:0] _RAND_210;
  reg [1:0] _T_3372_11_dst_rtype;
  reg [31:0] _RAND_211;
  reg  _T_3372_11_fp_val;
  reg [31:0] _RAND_212;
  reg [7:0] _T_3372_12_br_mask;
  reg [31:0] _RAND_213;
  reg [6:0] _T_3372_12_pdst;
  reg [31:0] _RAND_214;
  reg [6:0] _T_3372_12_stale_pdst;
  reg [31:0] _RAND_215;
  reg  _T_3372_12_is_fencei;
  reg [31:0] _RAND_216;
  reg  _T_3372_12_is_store;
  reg [31:0] _RAND_217;
  reg  _T_3372_12_is_load;
  reg [31:0] _RAND_218;
  reg  _T_3372_12_is_sys_pc2epc;
  reg [31:0] _RAND_219;
  reg  _T_3372_12_flush_on_commit;
  reg [31:0] _RAND_220;
  reg [5:0] _T_3372_12_ldst;
  reg [31:0] _RAND_221;
  reg  _T_3372_12_ldst_val;
  reg [31:0] _RAND_222;
  reg [1:0] _T_3372_12_dst_rtype;
  reg [31:0] _RAND_223;
  reg  _T_3372_12_fp_val;
  reg [31:0] _RAND_224;
  reg [7:0] _T_3372_13_br_mask;
  reg [31:0] _RAND_225;
  reg [6:0] _T_3372_13_pdst;
  reg [31:0] _RAND_226;
  reg [6:0] _T_3372_13_stale_pdst;
  reg [31:0] _RAND_227;
  reg  _T_3372_13_is_fencei;
  reg [31:0] _RAND_228;
  reg  _T_3372_13_is_store;
  reg [31:0] _RAND_229;
  reg  _T_3372_13_is_load;
  reg [31:0] _RAND_230;
  reg  _T_3372_13_is_sys_pc2epc;
  reg [31:0] _RAND_231;
  reg  _T_3372_13_flush_on_commit;
  reg [31:0] _RAND_232;
  reg [5:0] _T_3372_13_ldst;
  reg [31:0] _RAND_233;
  reg  _T_3372_13_ldst_val;
  reg [31:0] _RAND_234;
  reg [1:0] _T_3372_13_dst_rtype;
  reg [31:0] _RAND_235;
  reg  _T_3372_13_fp_val;
  reg [31:0] _RAND_236;
  reg [7:0] _T_3372_14_br_mask;
  reg [31:0] _RAND_237;
  reg [6:0] _T_3372_14_pdst;
  reg [31:0] _RAND_238;
  reg [6:0] _T_3372_14_stale_pdst;
  reg [31:0] _RAND_239;
  reg  _T_3372_14_is_fencei;
  reg [31:0] _RAND_240;
  reg  _T_3372_14_is_store;
  reg [31:0] _RAND_241;
  reg  _T_3372_14_is_load;
  reg [31:0] _RAND_242;
  reg  _T_3372_14_is_sys_pc2epc;
  reg [31:0] _RAND_243;
  reg  _T_3372_14_flush_on_commit;
  reg [31:0] _RAND_244;
  reg [5:0] _T_3372_14_ldst;
  reg [31:0] _RAND_245;
  reg  _T_3372_14_ldst_val;
  reg [31:0] _RAND_246;
  reg [1:0] _T_3372_14_dst_rtype;
  reg [31:0] _RAND_247;
  reg  _T_3372_14_fp_val;
  reg [31:0] _RAND_248;
  reg [7:0] _T_3372_15_br_mask;
  reg [31:0] _RAND_249;
  reg [6:0] _T_3372_15_pdst;
  reg [31:0] _RAND_250;
  reg [6:0] _T_3372_15_stale_pdst;
  reg [31:0] _RAND_251;
  reg  _T_3372_15_is_fencei;
  reg [31:0] _RAND_252;
  reg  _T_3372_15_is_store;
  reg [31:0] _RAND_253;
  reg  _T_3372_15_is_load;
  reg [31:0] _RAND_254;
  reg  _T_3372_15_is_sys_pc2epc;
  reg [31:0] _RAND_255;
  reg  _T_3372_15_flush_on_commit;
  reg [31:0] _RAND_256;
  reg [5:0] _T_3372_15_ldst;
  reg [31:0] _RAND_257;
  reg  _T_3372_15_ldst_val;
  reg [31:0] _RAND_258;
  reg [1:0] _T_3372_15_dst_rtype;
  reg [31:0] _RAND_259;
  reg  _T_3372_15_fp_val;
  reg [31:0] _RAND_260;
  reg [7:0] _T_3372_16_br_mask;
  reg [31:0] _RAND_261;
  reg [6:0] _T_3372_16_pdst;
  reg [31:0] _RAND_262;
  reg [6:0] _T_3372_16_stale_pdst;
  reg [31:0] _RAND_263;
  reg  _T_3372_16_is_fencei;
  reg [31:0] _RAND_264;
  reg  _T_3372_16_is_store;
  reg [31:0] _RAND_265;
  reg  _T_3372_16_is_load;
  reg [31:0] _RAND_266;
  reg  _T_3372_16_is_sys_pc2epc;
  reg [31:0] _RAND_267;
  reg  _T_3372_16_flush_on_commit;
  reg [31:0] _RAND_268;
  reg [5:0] _T_3372_16_ldst;
  reg [31:0] _RAND_269;
  reg  _T_3372_16_ldst_val;
  reg [31:0] _RAND_270;
  reg [1:0] _T_3372_16_dst_rtype;
  reg [31:0] _RAND_271;
  reg  _T_3372_16_fp_val;
  reg [31:0] _RAND_272;
  reg [7:0] _T_3372_17_br_mask;
  reg [31:0] _RAND_273;
  reg [6:0] _T_3372_17_pdst;
  reg [31:0] _RAND_274;
  reg [6:0] _T_3372_17_stale_pdst;
  reg [31:0] _RAND_275;
  reg  _T_3372_17_is_fencei;
  reg [31:0] _RAND_276;
  reg  _T_3372_17_is_store;
  reg [31:0] _RAND_277;
  reg  _T_3372_17_is_load;
  reg [31:0] _RAND_278;
  reg  _T_3372_17_is_sys_pc2epc;
  reg [31:0] _RAND_279;
  reg  _T_3372_17_flush_on_commit;
  reg [31:0] _RAND_280;
  reg [5:0] _T_3372_17_ldst;
  reg [31:0] _RAND_281;
  reg  _T_3372_17_ldst_val;
  reg [31:0] _RAND_282;
  reg [1:0] _T_3372_17_dst_rtype;
  reg [31:0] _RAND_283;
  reg  _T_3372_17_fp_val;
  reg [31:0] _RAND_284;
  reg [7:0] _T_3372_18_br_mask;
  reg [31:0] _RAND_285;
  reg [6:0] _T_3372_18_pdst;
  reg [31:0] _RAND_286;
  reg [6:0] _T_3372_18_stale_pdst;
  reg [31:0] _RAND_287;
  reg  _T_3372_18_is_fencei;
  reg [31:0] _RAND_288;
  reg  _T_3372_18_is_store;
  reg [31:0] _RAND_289;
  reg  _T_3372_18_is_load;
  reg [31:0] _RAND_290;
  reg  _T_3372_18_is_sys_pc2epc;
  reg [31:0] _RAND_291;
  reg  _T_3372_18_flush_on_commit;
  reg [31:0] _RAND_292;
  reg [5:0] _T_3372_18_ldst;
  reg [31:0] _RAND_293;
  reg  _T_3372_18_ldst_val;
  reg [31:0] _RAND_294;
  reg [1:0] _T_3372_18_dst_rtype;
  reg [31:0] _RAND_295;
  reg  _T_3372_18_fp_val;
  reg [31:0] _RAND_296;
  reg [7:0] _T_3372_19_br_mask;
  reg [31:0] _RAND_297;
  reg [6:0] _T_3372_19_pdst;
  reg [31:0] _RAND_298;
  reg [6:0] _T_3372_19_stale_pdst;
  reg [31:0] _RAND_299;
  reg  _T_3372_19_is_fencei;
  reg [31:0] _RAND_300;
  reg  _T_3372_19_is_store;
  reg [31:0] _RAND_301;
  reg  _T_3372_19_is_load;
  reg [31:0] _RAND_302;
  reg  _T_3372_19_is_sys_pc2epc;
  reg [31:0] _RAND_303;
  reg  _T_3372_19_flush_on_commit;
  reg [31:0] _RAND_304;
  reg [5:0] _T_3372_19_ldst;
  reg [31:0] _RAND_305;
  reg  _T_3372_19_ldst_val;
  reg [31:0] _RAND_306;
  reg [1:0] _T_3372_19_dst_rtype;
  reg [31:0] _RAND_307;
  reg  _T_3372_19_fp_val;
  reg [31:0] _RAND_308;
  reg [7:0] _T_3372_20_br_mask;
  reg [31:0] _RAND_309;
  reg [6:0] _T_3372_20_pdst;
  reg [31:0] _RAND_310;
  reg [6:0] _T_3372_20_stale_pdst;
  reg [31:0] _RAND_311;
  reg  _T_3372_20_is_fencei;
  reg [31:0] _RAND_312;
  reg  _T_3372_20_is_store;
  reg [31:0] _RAND_313;
  reg  _T_3372_20_is_load;
  reg [31:0] _RAND_314;
  reg  _T_3372_20_is_sys_pc2epc;
  reg [31:0] _RAND_315;
  reg  _T_3372_20_flush_on_commit;
  reg [31:0] _RAND_316;
  reg [5:0] _T_3372_20_ldst;
  reg [31:0] _RAND_317;
  reg  _T_3372_20_ldst_val;
  reg [31:0] _RAND_318;
  reg [1:0] _T_3372_20_dst_rtype;
  reg [31:0] _RAND_319;
  reg  _T_3372_20_fp_val;
  reg [31:0] _RAND_320;
  reg [7:0] _T_3372_21_br_mask;
  reg [31:0] _RAND_321;
  reg [6:0] _T_3372_21_pdst;
  reg [31:0] _RAND_322;
  reg [6:0] _T_3372_21_stale_pdst;
  reg [31:0] _RAND_323;
  reg  _T_3372_21_is_fencei;
  reg [31:0] _RAND_324;
  reg  _T_3372_21_is_store;
  reg [31:0] _RAND_325;
  reg  _T_3372_21_is_load;
  reg [31:0] _RAND_326;
  reg  _T_3372_21_is_sys_pc2epc;
  reg [31:0] _RAND_327;
  reg  _T_3372_21_flush_on_commit;
  reg [31:0] _RAND_328;
  reg [5:0] _T_3372_21_ldst;
  reg [31:0] _RAND_329;
  reg  _T_3372_21_ldst_val;
  reg [31:0] _RAND_330;
  reg [1:0] _T_3372_21_dst_rtype;
  reg [31:0] _RAND_331;
  reg  _T_3372_21_fp_val;
  reg [31:0] _RAND_332;
  reg [7:0] _T_3372_22_br_mask;
  reg [31:0] _RAND_333;
  reg [6:0] _T_3372_22_pdst;
  reg [31:0] _RAND_334;
  reg [6:0] _T_3372_22_stale_pdst;
  reg [31:0] _RAND_335;
  reg  _T_3372_22_is_fencei;
  reg [31:0] _RAND_336;
  reg  _T_3372_22_is_store;
  reg [31:0] _RAND_337;
  reg  _T_3372_22_is_load;
  reg [31:0] _RAND_338;
  reg  _T_3372_22_is_sys_pc2epc;
  reg [31:0] _RAND_339;
  reg  _T_3372_22_flush_on_commit;
  reg [31:0] _RAND_340;
  reg [5:0] _T_3372_22_ldst;
  reg [31:0] _RAND_341;
  reg  _T_3372_22_ldst_val;
  reg [31:0] _RAND_342;
  reg [1:0] _T_3372_22_dst_rtype;
  reg [31:0] _RAND_343;
  reg  _T_3372_22_fp_val;
  reg [31:0] _RAND_344;
  reg [7:0] _T_3372_23_br_mask;
  reg [31:0] _RAND_345;
  reg [6:0] _T_3372_23_pdst;
  reg [31:0] _RAND_346;
  reg [6:0] _T_3372_23_stale_pdst;
  reg [31:0] _RAND_347;
  reg  _T_3372_23_is_fencei;
  reg [31:0] _RAND_348;
  reg  _T_3372_23_is_store;
  reg [31:0] _RAND_349;
  reg  _T_3372_23_is_load;
  reg [31:0] _RAND_350;
  reg  _T_3372_23_is_sys_pc2epc;
  reg [31:0] _RAND_351;
  reg  _T_3372_23_flush_on_commit;
  reg [31:0] _RAND_352;
  reg [5:0] _T_3372_23_ldst;
  reg [31:0] _RAND_353;
  reg  _T_3372_23_ldst_val;
  reg [31:0] _RAND_354;
  reg [1:0] _T_3372_23_dst_rtype;
  reg [31:0] _RAND_355;
  reg  _T_3372_23_fp_val;
  reg [31:0] _RAND_356;
  reg [7:0] _T_3372_24_br_mask;
  reg [31:0] _RAND_357;
  reg [6:0] _T_3372_24_pdst;
  reg [31:0] _RAND_358;
  reg [6:0] _T_3372_24_stale_pdst;
  reg [31:0] _RAND_359;
  reg  _T_3372_24_is_fencei;
  reg [31:0] _RAND_360;
  reg  _T_3372_24_is_store;
  reg [31:0] _RAND_361;
  reg  _T_3372_24_is_load;
  reg [31:0] _RAND_362;
  reg  _T_3372_24_is_sys_pc2epc;
  reg [31:0] _RAND_363;
  reg  _T_3372_24_flush_on_commit;
  reg [31:0] _RAND_364;
  reg [5:0] _T_3372_24_ldst;
  reg [31:0] _RAND_365;
  reg  _T_3372_24_ldst_val;
  reg [31:0] _RAND_366;
  reg [1:0] _T_3372_24_dst_rtype;
  reg [31:0] _RAND_367;
  reg  _T_3372_24_fp_val;
  reg [31:0] _RAND_368;
  reg [7:0] _T_3372_25_br_mask;
  reg [31:0] _RAND_369;
  reg [6:0] _T_3372_25_pdst;
  reg [31:0] _RAND_370;
  reg [6:0] _T_3372_25_stale_pdst;
  reg [31:0] _RAND_371;
  reg  _T_3372_25_is_fencei;
  reg [31:0] _RAND_372;
  reg  _T_3372_25_is_store;
  reg [31:0] _RAND_373;
  reg  _T_3372_25_is_load;
  reg [31:0] _RAND_374;
  reg  _T_3372_25_is_sys_pc2epc;
  reg [31:0] _RAND_375;
  reg  _T_3372_25_flush_on_commit;
  reg [31:0] _RAND_376;
  reg [5:0] _T_3372_25_ldst;
  reg [31:0] _RAND_377;
  reg  _T_3372_25_ldst_val;
  reg [31:0] _RAND_378;
  reg [1:0] _T_3372_25_dst_rtype;
  reg [31:0] _RAND_379;
  reg  _T_3372_25_fp_val;
  reg [31:0] _RAND_380;
  reg [7:0] _T_3372_26_br_mask;
  reg [31:0] _RAND_381;
  reg [6:0] _T_3372_26_pdst;
  reg [31:0] _RAND_382;
  reg [6:0] _T_3372_26_stale_pdst;
  reg [31:0] _RAND_383;
  reg  _T_3372_26_is_fencei;
  reg [31:0] _RAND_384;
  reg  _T_3372_26_is_store;
  reg [31:0] _RAND_385;
  reg  _T_3372_26_is_load;
  reg [31:0] _RAND_386;
  reg  _T_3372_26_is_sys_pc2epc;
  reg [31:0] _RAND_387;
  reg  _T_3372_26_flush_on_commit;
  reg [31:0] _RAND_388;
  reg [5:0] _T_3372_26_ldst;
  reg [31:0] _RAND_389;
  reg  _T_3372_26_ldst_val;
  reg [31:0] _RAND_390;
  reg [1:0] _T_3372_26_dst_rtype;
  reg [31:0] _RAND_391;
  reg  _T_3372_26_fp_val;
  reg [31:0] _RAND_392;
  reg [7:0] _T_3372_27_br_mask;
  reg [31:0] _RAND_393;
  reg [6:0] _T_3372_27_pdst;
  reg [31:0] _RAND_394;
  reg [6:0] _T_3372_27_stale_pdst;
  reg [31:0] _RAND_395;
  reg  _T_3372_27_is_fencei;
  reg [31:0] _RAND_396;
  reg  _T_3372_27_is_store;
  reg [31:0] _RAND_397;
  reg  _T_3372_27_is_load;
  reg [31:0] _RAND_398;
  reg  _T_3372_27_is_sys_pc2epc;
  reg [31:0] _RAND_399;
  reg  _T_3372_27_flush_on_commit;
  reg [31:0] _RAND_400;
  reg [5:0] _T_3372_27_ldst;
  reg [31:0] _RAND_401;
  reg  _T_3372_27_ldst_val;
  reg [31:0] _RAND_402;
  reg [1:0] _T_3372_27_dst_rtype;
  reg [31:0] _RAND_403;
  reg  _T_3372_27_fp_val;
  reg [31:0] _RAND_404;
  reg [7:0] _T_3372_28_br_mask;
  reg [31:0] _RAND_405;
  reg [6:0] _T_3372_28_pdst;
  reg [31:0] _RAND_406;
  reg [6:0] _T_3372_28_stale_pdst;
  reg [31:0] _RAND_407;
  reg  _T_3372_28_is_fencei;
  reg [31:0] _RAND_408;
  reg  _T_3372_28_is_store;
  reg [31:0] _RAND_409;
  reg  _T_3372_28_is_load;
  reg [31:0] _RAND_410;
  reg  _T_3372_28_is_sys_pc2epc;
  reg [31:0] _RAND_411;
  reg  _T_3372_28_flush_on_commit;
  reg [31:0] _RAND_412;
  reg [5:0] _T_3372_28_ldst;
  reg [31:0] _RAND_413;
  reg  _T_3372_28_ldst_val;
  reg [31:0] _RAND_414;
  reg [1:0] _T_3372_28_dst_rtype;
  reg [31:0] _RAND_415;
  reg  _T_3372_28_fp_val;
  reg [31:0] _RAND_416;
  reg [7:0] _T_3372_29_br_mask;
  reg [31:0] _RAND_417;
  reg [6:0] _T_3372_29_pdst;
  reg [31:0] _RAND_418;
  reg [6:0] _T_3372_29_stale_pdst;
  reg [31:0] _RAND_419;
  reg  _T_3372_29_is_fencei;
  reg [31:0] _RAND_420;
  reg  _T_3372_29_is_store;
  reg [31:0] _RAND_421;
  reg  _T_3372_29_is_load;
  reg [31:0] _RAND_422;
  reg  _T_3372_29_is_sys_pc2epc;
  reg [31:0] _RAND_423;
  reg  _T_3372_29_flush_on_commit;
  reg [31:0] _RAND_424;
  reg [5:0] _T_3372_29_ldst;
  reg [31:0] _RAND_425;
  reg  _T_3372_29_ldst_val;
  reg [31:0] _RAND_426;
  reg [1:0] _T_3372_29_dst_rtype;
  reg [31:0] _RAND_427;
  reg  _T_3372_29_fp_val;
  reg [31:0] _RAND_428;
  reg [7:0] _T_3372_30_br_mask;
  reg [31:0] _RAND_429;
  reg [6:0] _T_3372_30_pdst;
  reg [31:0] _RAND_430;
  reg [6:0] _T_3372_30_stale_pdst;
  reg [31:0] _RAND_431;
  reg  _T_3372_30_is_fencei;
  reg [31:0] _RAND_432;
  reg  _T_3372_30_is_store;
  reg [31:0] _RAND_433;
  reg  _T_3372_30_is_load;
  reg [31:0] _RAND_434;
  reg  _T_3372_30_is_sys_pc2epc;
  reg [31:0] _RAND_435;
  reg  _T_3372_30_flush_on_commit;
  reg [31:0] _RAND_436;
  reg [5:0] _T_3372_30_ldst;
  reg [31:0] _RAND_437;
  reg  _T_3372_30_ldst_val;
  reg [31:0] _RAND_438;
  reg [1:0] _T_3372_30_dst_rtype;
  reg [31:0] _RAND_439;
  reg  _T_3372_30_fp_val;
  reg [31:0] _RAND_440;
  reg [7:0] _T_3372_31_br_mask;
  reg [31:0] _RAND_441;
  reg [6:0] _T_3372_31_pdst;
  reg [31:0] _RAND_442;
  reg [6:0] _T_3372_31_stale_pdst;
  reg [31:0] _RAND_443;
  reg  _T_3372_31_is_fencei;
  reg [31:0] _RAND_444;
  reg  _T_3372_31_is_store;
  reg [31:0] _RAND_445;
  reg  _T_3372_31_is_load;
  reg [31:0] _RAND_446;
  reg  _T_3372_31_is_sys_pc2epc;
  reg [31:0] _RAND_447;
  reg  _T_3372_31_flush_on_commit;
  reg [31:0] _RAND_448;
  reg [5:0] _T_3372_31_ldst;
  reg [31:0] _RAND_449;
  reg  _T_3372_31_ldst_val;
  reg [31:0] _RAND_450;
  reg [1:0] _T_3372_31_dst_rtype;
  reg [31:0] _RAND_451;
  reg  _T_3372_31_fp_val;
  reg [31:0] _RAND_452;
  reg [7:0] _T_3372_32_br_mask;
  reg [31:0] _RAND_453;
  reg [6:0] _T_3372_32_pdst;
  reg [31:0] _RAND_454;
  reg [6:0] _T_3372_32_stale_pdst;
  reg [31:0] _RAND_455;
  reg  _T_3372_32_is_fencei;
  reg [31:0] _RAND_456;
  reg  _T_3372_32_is_store;
  reg [31:0] _RAND_457;
  reg  _T_3372_32_is_load;
  reg [31:0] _RAND_458;
  reg  _T_3372_32_is_sys_pc2epc;
  reg [31:0] _RAND_459;
  reg  _T_3372_32_flush_on_commit;
  reg [31:0] _RAND_460;
  reg [5:0] _T_3372_32_ldst;
  reg [31:0] _RAND_461;
  reg  _T_3372_32_ldst_val;
  reg [31:0] _RAND_462;
  reg [1:0] _T_3372_32_dst_rtype;
  reg [31:0] _RAND_463;
  reg  _T_3372_32_fp_val;
  reg [31:0] _RAND_464;
  reg [7:0] _T_3372_33_br_mask;
  reg [31:0] _RAND_465;
  reg [6:0] _T_3372_33_pdst;
  reg [31:0] _RAND_466;
  reg [6:0] _T_3372_33_stale_pdst;
  reg [31:0] _RAND_467;
  reg  _T_3372_33_is_fencei;
  reg [31:0] _RAND_468;
  reg  _T_3372_33_is_store;
  reg [31:0] _RAND_469;
  reg  _T_3372_33_is_load;
  reg [31:0] _RAND_470;
  reg  _T_3372_33_is_sys_pc2epc;
  reg [31:0] _RAND_471;
  reg  _T_3372_33_flush_on_commit;
  reg [31:0] _RAND_472;
  reg [5:0] _T_3372_33_ldst;
  reg [31:0] _RAND_473;
  reg  _T_3372_33_ldst_val;
  reg [31:0] _RAND_474;
  reg [1:0] _T_3372_33_dst_rtype;
  reg [31:0] _RAND_475;
  reg  _T_3372_33_fp_val;
  reg [31:0] _RAND_476;
  reg [7:0] _T_3372_34_br_mask;
  reg [31:0] _RAND_477;
  reg [6:0] _T_3372_34_pdst;
  reg [31:0] _RAND_478;
  reg [6:0] _T_3372_34_stale_pdst;
  reg [31:0] _RAND_479;
  reg  _T_3372_34_is_fencei;
  reg [31:0] _RAND_480;
  reg  _T_3372_34_is_store;
  reg [31:0] _RAND_481;
  reg  _T_3372_34_is_load;
  reg [31:0] _RAND_482;
  reg  _T_3372_34_is_sys_pc2epc;
  reg [31:0] _RAND_483;
  reg  _T_3372_34_flush_on_commit;
  reg [31:0] _RAND_484;
  reg [5:0] _T_3372_34_ldst;
  reg [31:0] _RAND_485;
  reg  _T_3372_34_ldst_val;
  reg [31:0] _RAND_486;
  reg [1:0] _T_3372_34_dst_rtype;
  reg [31:0] _RAND_487;
  reg  _T_3372_34_fp_val;
  reg [31:0] _RAND_488;
  reg [7:0] _T_3372_35_br_mask;
  reg [31:0] _RAND_489;
  reg [6:0] _T_3372_35_pdst;
  reg [31:0] _RAND_490;
  reg [6:0] _T_3372_35_stale_pdst;
  reg [31:0] _RAND_491;
  reg  _T_3372_35_is_fencei;
  reg [31:0] _RAND_492;
  reg  _T_3372_35_is_store;
  reg [31:0] _RAND_493;
  reg  _T_3372_35_is_load;
  reg [31:0] _RAND_494;
  reg  _T_3372_35_is_sys_pc2epc;
  reg [31:0] _RAND_495;
  reg  _T_3372_35_flush_on_commit;
  reg [31:0] _RAND_496;
  reg [5:0] _T_3372_35_ldst;
  reg [31:0] _RAND_497;
  reg  _T_3372_35_ldst_val;
  reg [31:0] _RAND_498;
  reg [1:0] _T_3372_35_dst_rtype;
  reg [31:0] _RAND_499;
  reg  _T_3372_35_fp_val;
  reg [31:0] _RAND_500;
  reg [7:0] _T_3372_36_br_mask;
  reg [31:0] _RAND_501;
  reg [6:0] _T_3372_36_pdst;
  reg [31:0] _RAND_502;
  reg [6:0] _T_3372_36_stale_pdst;
  reg [31:0] _RAND_503;
  reg  _T_3372_36_is_fencei;
  reg [31:0] _RAND_504;
  reg  _T_3372_36_is_store;
  reg [31:0] _RAND_505;
  reg  _T_3372_36_is_load;
  reg [31:0] _RAND_506;
  reg  _T_3372_36_is_sys_pc2epc;
  reg [31:0] _RAND_507;
  reg  _T_3372_36_flush_on_commit;
  reg [31:0] _RAND_508;
  reg [5:0] _T_3372_36_ldst;
  reg [31:0] _RAND_509;
  reg  _T_3372_36_ldst_val;
  reg [31:0] _RAND_510;
  reg [1:0] _T_3372_36_dst_rtype;
  reg [31:0] _RAND_511;
  reg  _T_3372_36_fp_val;
  reg [31:0] _RAND_512;
  reg [7:0] _T_3372_37_br_mask;
  reg [31:0] _RAND_513;
  reg [6:0] _T_3372_37_pdst;
  reg [31:0] _RAND_514;
  reg [6:0] _T_3372_37_stale_pdst;
  reg [31:0] _RAND_515;
  reg  _T_3372_37_is_fencei;
  reg [31:0] _RAND_516;
  reg  _T_3372_37_is_store;
  reg [31:0] _RAND_517;
  reg  _T_3372_37_is_load;
  reg [31:0] _RAND_518;
  reg  _T_3372_37_is_sys_pc2epc;
  reg [31:0] _RAND_519;
  reg  _T_3372_37_flush_on_commit;
  reg [31:0] _RAND_520;
  reg [5:0] _T_3372_37_ldst;
  reg [31:0] _RAND_521;
  reg  _T_3372_37_ldst_val;
  reg [31:0] _RAND_522;
  reg [1:0] _T_3372_37_dst_rtype;
  reg [31:0] _RAND_523;
  reg  _T_3372_37_fp_val;
  reg [31:0] _RAND_524;
  reg [7:0] _T_3372_38_br_mask;
  reg [31:0] _RAND_525;
  reg [6:0] _T_3372_38_pdst;
  reg [31:0] _RAND_526;
  reg [6:0] _T_3372_38_stale_pdst;
  reg [31:0] _RAND_527;
  reg  _T_3372_38_is_fencei;
  reg [31:0] _RAND_528;
  reg  _T_3372_38_is_store;
  reg [31:0] _RAND_529;
  reg  _T_3372_38_is_load;
  reg [31:0] _RAND_530;
  reg  _T_3372_38_is_sys_pc2epc;
  reg [31:0] _RAND_531;
  reg  _T_3372_38_flush_on_commit;
  reg [31:0] _RAND_532;
  reg [5:0] _T_3372_38_ldst;
  reg [31:0] _RAND_533;
  reg  _T_3372_38_ldst_val;
  reg [31:0] _RAND_534;
  reg [1:0] _T_3372_38_dst_rtype;
  reg [31:0] _RAND_535;
  reg  _T_3372_38_fp_val;
  reg [31:0] _RAND_536;
  reg [7:0] _T_3372_39_br_mask;
  reg [31:0] _RAND_537;
  reg [6:0] _T_3372_39_pdst;
  reg [31:0] _RAND_538;
  reg [6:0] _T_3372_39_stale_pdst;
  reg [31:0] _RAND_539;
  reg  _T_3372_39_is_fencei;
  reg [31:0] _RAND_540;
  reg  _T_3372_39_is_store;
  reg [31:0] _RAND_541;
  reg  _T_3372_39_is_load;
  reg [31:0] _RAND_542;
  reg  _T_3372_39_is_sys_pc2epc;
  reg [31:0] _RAND_543;
  reg  _T_3372_39_flush_on_commit;
  reg [31:0] _RAND_544;
  reg [5:0] _T_3372_39_ldst;
  reg [31:0] _RAND_545;
  reg  _T_3372_39_ldst_val;
  reg [31:0] _RAND_546;
  reg [1:0] _T_3372_39_dst_rtype;
  reg [31:0] _RAND_547;
  reg  _T_3372_39_fp_val;
  reg [31:0] _RAND_548;
  reg  _T_3745 [0:39];
  reg [31:0] _RAND_549;
  wire  _T_3745__T_4012_data;
  wire [5:0] _T_3745__T_4012_addr;
  reg [31:0] _RAND_550;
  wire  _T_3745__T_3768_data;
  wire [5:0] _T_3745__T_3768_addr;
  wire  _T_3745__T_3768_mask;
  wire  _T_3745__T_3768_en;
  wire  _T_3745__T_3998_data;
  wire [5:0] _T_3745__T_3998_addr;
  wire  _T_3745__T_3998_mask;
  wire  _T_3745__T_3998_en;
  wire  _T_3745__T_4007_data;
  wire [5:0] _T_3745__T_4007_addr;
  wire  _T_3745__T_4007_mask;
  wire  _T_3745__T_4007_en;
  wire  _T_3745__T_4088_data;
  wire [5:0] _T_3745__T_4088_addr;
  wire  _T_3745__T_4088_mask;
  wire  _T_3745__T_4088_en;
  reg [4:0] _T_3748 [0:39];
  reg [31:0] _RAND_551;
  wire [4:0] _T_3748__T_5017_data;
  wire [5:0] _T_3748__T_5017_addr;
  reg [31:0] _RAND_552;
  wire [4:0] _T_3748__T_3769_data;
  wire [5:0] _T_3748__T_3769_addr;
  wire  _T_3748__T_3769_mask;
  wire  _T_3748__T_3769_en;
  wire [4:0] _T_3748__T_3982_data;
  wire [5:0] _T_3748__T_3982_addr;
  wire  _T_3748__T_3982_mask;
  wire  _T_3748__T_3982_en;
  wire [4:0] _T_3748__T_3990_data;
  wire [5:0] _T_3748__T_3990_addr;
  wire  _T_3748__T_3990_mask;
  wire  _T_3748__T_3990_en;
  wire  _GEN_575;
  wire  _GEN_576;
  wire  _GEN_577;
  wire  _GEN_578;
  wire  _GEN_579;
  wire  _GEN_580;
  wire  _GEN_581;
  wire  _GEN_582;
  wire  _GEN_583;
  wire  _GEN_584;
  wire  _GEN_585;
  wire  _GEN_586;
  wire  _GEN_587;
  wire  _GEN_588;
  wire  _GEN_589;
  wire  _GEN_590;
  wire  _GEN_591;
  wire  _GEN_592;
  wire  _GEN_593;
  wire  _GEN_594;
  wire  _GEN_595;
  wire  _GEN_596;
  wire  _GEN_597;
  wire  _GEN_598;
  wire  _GEN_599;
  wire  _GEN_600;
  wire  _GEN_601;
  wire  _GEN_602;
  wire  _GEN_603;
  wire  _GEN_604;
  wire  _GEN_605;
  wire  _GEN_606;
  wire  _GEN_607;
  wire  _GEN_608;
  wire  _GEN_609;
  wire  _GEN_610;
  wire  _GEN_611;
  wire  _GEN_612;
  wire  _GEN_613;
  wire  _GEN_614;
  wire  _T_3755;
  wire  _T_3757;
  wire  _T_3758;
  wire [7:0] _GEN_26;
  wire [7:0] _GEN_1575;
  wire [7:0] _GEN_1576;
  wire [7:0] _GEN_1577;
  wire [7:0] _GEN_1578;
  wire [7:0] _GEN_1579;
  wire [7:0] _GEN_1580;
  wire [7:0] _GEN_1581;
  wire [7:0] _GEN_1582;
  wire [7:0] _GEN_1583;
  wire [7:0] _GEN_1584;
  wire [7:0] _GEN_1585;
  wire [7:0] _GEN_1586;
  wire [7:0] _GEN_1587;
  wire [7:0] _GEN_1588;
  wire [7:0] _GEN_1589;
  wire [7:0] _GEN_1590;
  wire [7:0] _GEN_1591;
  wire [7:0] _GEN_1592;
  wire [7:0] _GEN_1593;
  wire [7:0] _GEN_1594;
  wire [7:0] _GEN_1595;
  wire [7:0] _GEN_1596;
  wire [7:0] _GEN_1597;
  wire [7:0] _GEN_1598;
  wire [7:0] _GEN_1599;
  wire [7:0] _GEN_1600;
  wire [7:0] _GEN_1601;
  wire [7:0] _GEN_1602;
  wire [7:0] _GEN_1603;
  wire [7:0] _GEN_1604;
  wire [7:0] _GEN_1605;
  wire [7:0] _GEN_1606;
  wire [7:0] _GEN_1607;
  wire [7:0] _GEN_1608;
  wire [7:0] _GEN_1609;
  wire [7:0] _GEN_1610;
  wire [7:0] _GEN_1611;
  wire [7:0] _GEN_1612;
  wire [7:0] _GEN_1613;
  wire [7:0] _GEN_1614;
  wire [6:0] _GEN_54;
  wire [6:0] _GEN_2695;
  wire [6:0] _GEN_2696;
  wire [6:0] _GEN_2697;
  wire [6:0] _GEN_2698;
  wire [6:0] _GEN_2699;
  wire [6:0] _GEN_2700;
  wire [6:0] _GEN_2701;
  wire [6:0] _GEN_2702;
  wire [6:0] _GEN_2703;
  wire [6:0] _GEN_2704;
  wire [6:0] _GEN_2705;
  wire [6:0] _GEN_2706;
  wire [6:0] _GEN_2707;
  wire [6:0] _GEN_2708;
  wire [6:0] _GEN_2709;
  wire [6:0] _GEN_2710;
  wire [6:0] _GEN_2711;
  wire [6:0] _GEN_2712;
  wire [6:0] _GEN_2713;
  wire [6:0] _GEN_2714;
  wire [6:0] _GEN_2715;
  wire [6:0] _GEN_2716;
  wire [6:0] _GEN_2717;
  wire [6:0] _GEN_2718;
  wire [6:0] _GEN_2719;
  wire [6:0] _GEN_2720;
  wire [6:0] _GEN_2721;
  wire [6:0] _GEN_2722;
  wire [6:0] _GEN_2723;
  wire [6:0] _GEN_2724;
  wire [6:0] _GEN_2725;
  wire [6:0] _GEN_2726;
  wire [6:0] _GEN_2727;
  wire [6:0] _GEN_2728;
  wire [6:0] _GEN_2729;
  wire [6:0] _GEN_2730;
  wire [6:0] _GEN_2731;
  wire [6:0] _GEN_2732;
  wire [6:0] _GEN_2733;
  wire [6:0] _GEN_2734;
  wire [6:0] _GEN_61;
  wire [6:0] _GEN_2975;
  wire [6:0] _GEN_2976;
  wire [6:0] _GEN_2977;
  wire [6:0] _GEN_2978;
  wire [6:0] _GEN_2979;
  wire [6:0] _GEN_2980;
  wire [6:0] _GEN_2981;
  wire [6:0] _GEN_2982;
  wire [6:0] _GEN_2983;
  wire [6:0] _GEN_2984;
  wire [6:0] _GEN_2985;
  wire [6:0] _GEN_2986;
  wire [6:0] _GEN_2987;
  wire [6:0] _GEN_2988;
  wire [6:0] _GEN_2989;
  wire [6:0] _GEN_2990;
  wire [6:0] _GEN_2991;
  wire [6:0] _GEN_2992;
  wire [6:0] _GEN_2993;
  wire [6:0] _GEN_2994;
  wire [6:0] _GEN_2995;
  wire [6:0] _GEN_2996;
  wire [6:0] _GEN_2997;
  wire [6:0] _GEN_2998;
  wire [6:0] _GEN_2999;
  wire [6:0] _GEN_3000;
  wire [6:0] _GEN_3001;
  wire [6:0] _GEN_3002;
  wire [6:0] _GEN_3003;
  wire [6:0] _GEN_3004;
  wire [6:0] _GEN_3005;
  wire [6:0] _GEN_3006;
  wire [6:0] _GEN_3007;
  wire [6:0] _GEN_3008;
  wire [6:0] _GEN_3009;
  wire [6:0] _GEN_3010;
  wire [6:0] _GEN_3011;
  wire [6:0] _GEN_3012;
  wire [6:0] _GEN_3013;
  wire [6:0] _GEN_3014;
  wire  _GEN_68;
  wire  _GEN_3255;
  wire  _GEN_3256;
  wire  _GEN_3257;
  wire  _GEN_3258;
  wire  _GEN_3259;
  wire  _GEN_3260;
  wire  _GEN_3261;
  wire  _GEN_3262;
  wire  _GEN_3263;
  wire  _GEN_3264;
  wire  _GEN_3265;
  wire  _GEN_3266;
  wire  _GEN_3267;
  wire  _GEN_3268;
  wire  _GEN_3269;
  wire  _GEN_3270;
  wire  _GEN_3271;
  wire  _GEN_3272;
  wire  _GEN_3273;
  wire  _GEN_3274;
  wire  _GEN_3275;
  wire  _GEN_3276;
  wire  _GEN_3277;
  wire  _GEN_3278;
  wire  _GEN_3279;
  wire  _GEN_3280;
  wire  _GEN_3281;
  wire  _GEN_3282;
  wire  _GEN_3283;
  wire  _GEN_3284;
  wire  _GEN_3285;
  wire  _GEN_3286;
  wire  _GEN_3287;
  wire  _GEN_3288;
  wire  _GEN_3289;
  wire  _GEN_3290;
  wire  _GEN_3291;
  wire  _GEN_3292;
  wire  _GEN_3293;
  wire  _GEN_3294;
  wire  _GEN_69;
  wire  _GEN_3295;
  wire  _GEN_3296;
  wire  _GEN_3297;
  wire  _GEN_3298;
  wire  _GEN_3299;
  wire  _GEN_3300;
  wire  _GEN_3301;
  wire  _GEN_3302;
  wire  _GEN_3303;
  wire  _GEN_3304;
  wire  _GEN_3305;
  wire  _GEN_3306;
  wire  _GEN_3307;
  wire  _GEN_3308;
  wire  _GEN_3309;
  wire  _GEN_3310;
  wire  _GEN_3311;
  wire  _GEN_3312;
  wire  _GEN_3313;
  wire  _GEN_3314;
  wire  _GEN_3315;
  wire  _GEN_3316;
  wire  _GEN_3317;
  wire  _GEN_3318;
  wire  _GEN_3319;
  wire  _GEN_3320;
  wire  _GEN_3321;
  wire  _GEN_3322;
  wire  _GEN_3323;
  wire  _GEN_3324;
  wire  _GEN_3325;
  wire  _GEN_3326;
  wire  _GEN_3327;
  wire  _GEN_3328;
  wire  _GEN_3329;
  wire  _GEN_3330;
  wire  _GEN_3331;
  wire  _GEN_3332;
  wire  _GEN_3333;
  wire  _GEN_3334;
  wire  _GEN_71;
  wire  _GEN_3375;
  wire  _GEN_3376;
  wire  _GEN_3377;
  wire  _GEN_3378;
  wire  _GEN_3379;
  wire  _GEN_3380;
  wire  _GEN_3381;
  wire  _GEN_3382;
  wire  _GEN_3383;
  wire  _GEN_3384;
  wire  _GEN_3385;
  wire  _GEN_3386;
  wire  _GEN_3387;
  wire  _GEN_3388;
  wire  _GEN_3389;
  wire  _GEN_3390;
  wire  _GEN_3391;
  wire  _GEN_3392;
  wire  _GEN_3393;
  wire  _GEN_3394;
  wire  _GEN_3395;
  wire  _GEN_3396;
  wire  _GEN_3397;
  wire  _GEN_3398;
  wire  _GEN_3399;
  wire  _GEN_3400;
  wire  _GEN_3401;
  wire  _GEN_3402;
  wire  _GEN_3403;
  wire  _GEN_3404;
  wire  _GEN_3405;
  wire  _GEN_3406;
  wire  _GEN_3407;
  wire  _GEN_3408;
  wire  _GEN_3409;
  wire  _GEN_3410;
  wire  _GEN_3411;
  wire  _GEN_3412;
  wire  _GEN_3413;
  wire  _GEN_3414;
  wire  _GEN_72;
  wire  _GEN_3415;
  wire  _GEN_3416;
  wire  _GEN_3417;
  wire  _GEN_3418;
  wire  _GEN_3419;
  wire  _GEN_3420;
  wire  _GEN_3421;
  wire  _GEN_3422;
  wire  _GEN_3423;
  wire  _GEN_3424;
  wire  _GEN_3425;
  wire  _GEN_3426;
  wire  _GEN_3427;
  wire  _GEN_3428;
  wire  _GEN_3429;
  wire  _GEN_3430;
  wire  _GEN_3431;
  wire  _GEN_3432;
  wire  _GEN_3433;
  wire  _GEN_3434;
  wire  _GEN_3435;
  wire  _GEN_3436;
  wire  _GEN_3437;
  wire  _GEN_3438;
  wire  _GEN_3439;
  wire  _GEN_3440;
  wire  _GEN_3441;
  wire  _GEN_3442;
  wire  _GEN_3443;
  wire  _GEN_3444;
  wire  _GEN_3445;
  wire  _GEN_3446;
  wire  _GEN_3447;
  wire  _GEN_3448;
  wire  _GEN_3449;
  wire  _GEN_3450;
  wire  _GEN_3451;
  wire  _GEN_3452;
  wire  _GEN_3453;
  wire  _GEN_3454;
  wire  _GEN_74;
  wire  _GEN_3495;
  wire  _GEN_3496;
  wire  _GEN_3497;
  wire  _GEN_3498;
  wire  _GEN_3499;
  wire  _GEN_3500;
  wire  _GEN_3501;
  wire  _GEN_3502;
  wire  _GEN_3503;
  wire  _GEN_3504;
  wire  _GEN_3505;
  wire  _GEN_3506;
  wire  _GEN_3507;
  wire  _GEN_3508;
  wire  _GEN_3509;
  wire  _GEN_3510;
  wire  _GEN_3511;
  wire  _GEN_3512;
  wire  _GEN_3513;
  wire  _GEN_3514;
  wire  _GEN_3515;
  wire  _GEN_3516;
  wire  _GEN_3517;
  wire  _GEN_3518;
  wire  _GEN_3519;
  wire  _GEN_3520;
  wire  _GEN_3521;
  wire  _GEN_3522;
  wire  _GEN_3523;
  wire  _GEN_3524;
  wire  _GEN_3525;
  wire  _GEN_3526;
  wire  _GEN_3527;
  wire  _GEN_3528;
  wire  _GEN_3529;
  wire  _GEN_3530;
  wire  _GEN_3531;
  wire  _GEN_3532;
  wire  _GEN_3533;
  wire  _GEN_3534;
  wire [5:0] _GEN_75;
  wire [5:0] _GEN_3535;
  wire [5:0] _GEN_3536;
  wire [5:0] _GEN_3537;
  wire [5:0] _GEN_3538;
  wire [5:0] _GEN_3539;
  wire [5:0] _GEN_3540;
  wire [5:0] _GEN_3541;
  wire [5:0] _GEN_3542;
  wire [5:0] _GEN_3543;
  wire [5:0] _GEN_3544;
  wire [5:0] _GEN_3545;
  wire [5:0] _GEN_3546;
  wire [5:0] _GEN_3547;
  wire [5:0] _GEN_3548;
  wire [5:0] _GEN_3549;
  wire [5:0] _GEN_3550;
  wire [5:0] _GEN_3551;
  wire [5:0] _GEN_3552;
  wire [5:0] _GEN_3553;
  wire [5:0] _GEN_3554;
  wire [5:0] _GEN_3555;
  wire [5:0] _GEN_3556;
  wire [5:0] _GEN_3557;
  wire [5:0] _GEN_3558;
  wire [5:0] _GEN_3559;
  wire [5:0] _GEN_3560;
  wire [5:0] _GEN_3561;
  wire [5:0] _GEN_3562;
  wire [5:0] _GEN_3563;
  wire [5:0] _GEN_3564;
  wire [5:0] _GEN_3565;
  wire [5:0] _GEN_3566;
  wire [5:0] _GEN_3567;
  wire [5:0] _GEN_3568;
  wire [5:0] _GEN_3569;
  wire [5:0] _GEN_3570;
  wire [5:0] _GEN_3571;
  wire [5:0] _GEN_3572;
  wire [5:0] _GEN_3573;
  wire [5:0] _GEN_3574;
  wire  _GEN_79;
  wire  _GEN_3695;
  wire  _GEN_3696;
  wire  _GEN_3697;
  wire  _GEN_3698;
  wire  _GEN_3699;
  wire  _GEN_3700;
  wire  _GEN_3701;
  wire  _GEN_3702;
  wire  _GEN_3703;
  wire  _GEN_3704;
  wire  _GEN_3705;
  wire  _GEN_3706;
  wire  _GEN_3707;
  wire  _GEN_3708;
  wire  _GEN_3709;
  wire  _GEN_3710;
  wire  _GEN_3711;
  wire  _GEN_3712;
  wire  _GEN_3713;
  wire  _GEN_3714;
  wire  _GEN_3715;
  wire  _GEN_3716;
  wire  _GEN_3717;
  wire  _GEN_3718;
  wire  _GEN_3719;
  wire  _GEN_3720;
  wire  _GEN_3721;
  wire  _GEN_3722;
  wire  _GEN_3723;
  wire  _GEN_3724;
  wire  _GEN_3725;
  wire  _GEN_3726;
  wire  _GEN_3727;
  wire  _GEN_3728;
  wire  _GEN_3729;
  wire  _GEN_3730;
  wire  _GEN_3731;
  wire  _GEN_3732;
  wire  _GEN_3733;
  wire  _GEN_3734;
  wire [1:0] _GEN_80;
  wire [1:0] _GEN_3735;
  wire [1:0] _GEN_3736;
  wire [1:0] _GEN_3737;
  wire [1:0] _GEN_3738;
  wire [1:0] _GEN_3739;
  wire [1:0] _GEN_3740;
  wire [1:0] _GEN_3741;
  wire [1:0] _GEN_3742;
  wire [1:0] _GEN_3743;
  wire [1:0] _GEN_3744;
  wire [1:0] _GEN_3745;
  wire [1:0] _GEN_3746;
  wire [1:0] _GEN_3747;
  wire [1:0] _GEN_3748;
  wire [1:0] _GEN_3749;
  wire [1:0] _GEN_3750;
  wire [1:0] _GEN_3751;
  wire [1:0] _GEN_3752;
  wire [1:0] _GEN_3753;
  wire [1:0] _GEN_3754;
  wire [1:0] _GEN_3755;
  wire [1:0] _GEN_3756;
  wire [1:0] _GEN_3757;
  wire [1:0] _GEN_3758;
  wire [1:0] _GEN_3759;
  wire [1:0] _GEN_3760;
  wire [1:0] _GEN_3761;
  wire [1:0] _GEN_3762;
  wire [1:0] _GEN_3763;
  wire [1:0] _GEN_3764;
  wire [1:0] _GEN_3765;
  wire [1:0] _GEN_3766;
  wire [1:0] _GEN_3767;
  wire [1:0] _GEN_3768;
  wire [1:0] _GEN_3769;
  wire [1:0] _GEN_3770;
  wire [1:0] _GEN_3771;
  wire [1:0] _GEN_3772;
  wire [1:0] _GEN_3773;
  wire [1:0] _GEN_3774;
  wire  _GEN_84;
  wire  _GEN_3895;
  wire  _GEN_3896;
  wire  _GEN_3897;
  wire  _GEN_3898;
  wire  _GEN_3899;
  wire  _GEN_3900;
  wire  _GEN_3901;
  wire  _GEN_3902;
  wire  _GEN_3903;
  wire  _GEN_3904;
  wire  _GEN_3905;
  wire  _GEN_3906;
  wire  _GEN_3907;
  wire  _GEN_3908;
  wire  _GEN_3909;
  wire  _GEN_3910;
  wire  _GEN_3911;
  wire  _GEN_3912;
  wire  _GEN_3913;
  wire  _GEN_3914;
  wire  _GEN_3915;
  wire  _GEN_3916;
  wire  _GEN_3917;
  wire  _GEN_3918;
  wire  _GEN_3919;
  wire  _GEN_3920;
  wire  _GEN_3921;
  wire  _GEN_3922;
  wire  _GEN_3923;
  wire  _GEN_3924;
  wire  _GEN_3925;
  wire  _GEN_3926;
  wire  _GEN_3927;
  wire  _GEN_3928;
  wire  _GEN_3929;
  wire  _GEN_3930;
  wire  _GEN_3931;
  wire  _GEN_3932;
  wire  _GEN_3933;
  wire  _GEN_3934;
  wire  _GEN_93;
  wire  _GEN_4255;
  wire  _GEN_4256;
  wire  _GEN_4257;
  wire  _GEN_4258;
  wire  _GEN_4259;
  wire  _GEN_4260;
  wire  _GEN_4261;
  wire  _GEN_4262;
  wire  _GEN_4263;
  wire  _GEN_4264;
  wire  _GEN_4265;
  wire  _GEN_4266;
  wire  _GEN_4267;
  wire  _GEN_4268;
  wire  _GEN_4269;
  wire  _GEN_4270;
  wire  _GEN_4271;
  wire  _GEN_4272;
  wire  _GEN_4273;
  wire  _GEN_4274;
  wire  _GEN_4275;
  wire  _GEN_4276;
  wire  _GEN_4277;
  wire  _GEN_4278;
  wire  _GEN_4279;
  wire  _GEN_4280;
  wire  _GEN_4281;
  wire  _GEN_4282;
  wire  _GEN_4283;
  wire  _GEN_4284;
  wire  _GEN_4285;
  wire  _GEN_4286;
  wire  _GEN_4287;
  wire  _GEN_4288;
  wire  _GEN_4289;
  wire  _GEN_4290;
  wire  _GEN_4291;
  wire  _GEN_4292;
  wire  _GEN_4293;
  wire  _T_3785;
  wire  _T_3787;
  wire  _T_3789;
  wire [5:0] _T_3790;
  wire  _T_3791;
  wire  _T_3793;
  wire  _T_3795;
  wire  _GEN_4374;
  wire  _GEN_4375;
  wire  _GEN_4376;
  wire  _GEN_4377;
  wire  _GEN_4378;
  wire  _GEN_4379;
  wire  _GEN_4380;
  wire  _GEN_4381;
  wire  _GEN_4382;
  wire  _GEN_4383;
  wire  _GEN_4384;
  wire  _GEN_4385;
  wire  _GEN_4386;
  wire  _GEN_4387;
  wire  _GEN_4388;
  wire  _GEN_4389;
  wire  _GEN_4390;
  wire  _GEN_4391;
  wire  _GEN_4392;
  wire  _GEN_4393;
  wire  _GEN_4394;
  wire  _GEN_4395;
  wire  _GEN_4396;
  wire  _GEN_4397;
  wire  _GEN_4398;
  wire  _GEN_4399;
  wire  _GEN_4400;
  wire  _GEN_4401;
  wire  _GEN_4402;
  wire  _GEN_4403;
  wire  _GEN_4404;
  wire  _GEN_4405;
  wire  _GEN_4406;
  wire  _GEN_4407;
  wire  _GEN_4408;
  wire  _GEN_4409;
  wire  _GEN_4410;
  wire  _GEN_4411;
  wire  _GEN_4412;
  wire  _GEN_4413;
  wire [7:0] _GEN_5378;
  wire [7:0] _GEN_5379;
  wire [7:0] _GEN_5380;
  wire [7:0] _GEN_5381;
  wire [7:0] _GEN_5382;
  wire [7:0] _GEN_5383;
  wire [7:0] _GEN_5384;
  wire [7:0] _GEN_5385;
  wire [7:0] _GEN_5386;
  wire [7:0] _GEN_5387;
  wire [7:0] _GEN_5388;
  wire [7:0] _GEN_5389;
  wire [7:0] _GEN_5390;
  wire [7:0] _GEN_5391;
  wire [7:0] _GEN_5392;
  wire [7:0] _GEN_5393;
  wire [7:0] _GEN_5394;
  wire [7:0] _GEN_5395;
  wire [7:0] _GEN_5396;
  wire [7:0] _GEN_5397;
  wire [7:0] _GEN_5398;
  wire [7:0] _GEN_5399;
  wire [7:0] _GEN_5400;
  wire [7:0] _GEN_5401;
  wire [7:0] _GEN_5402;
  wire [7:0] _GEN_5403;
  wire [7:0] _GEN_5404;
  wire [7:0] _GEN_5405;
  wire [7:0] _GEN_5406;
  wire [7:0] _GEN_5407;
  wire [7:0] _GEN_5408;
  wire [7:0] _GEN_5409;
  wire [7:0] _GEN_5410;
  wire [7:0] _GEN_5411;
  wire [7:0] _GEN_5412;
  wire [7:0] _GEN_5413;
  wire [7:0] _GEN_5414;
  wire [7:0] _GEN_5415;
  wire [7:0] _GEN_5416;
  wire [7:0] _GEN_5417;
  wire [6:0] _GEN_6498;
  wire [6:0] _GEN_6499;
  wire [6:0] _GEN_6500;
  wire [6:0] _GEN_6501;
  wire [6:0] _GEN_6502;
  wire [6:0] _GEN_6503;
  wire [6:0] _GEN_6504;
  wire [6:0] _GEN_6505;
  wire [6:0] _GEN_6506;
  wire [6:0] _GEN_6507;
  wire [6:0] _GEN_6508;
  wire [6:0] _GEN_6509;
  wire [6:0] _GEN_6510;
  wire [6:0] _GEN_6511;
  wire [6:0] _GEN_6512;
  wire [6:0] _GEN_6513;
  wire [6:0] _GEN_6514;
  wire [6:0] _GEN_6515;
  wire [6:0] _GEN_6516;
  wire [6:0] _GEN_6517;
  wire [6:0] _GEN_6518;
  wire [6:0] _GEN_6519;
  wire [6:0] _GEN_6520;
  wire [6:0] _GEN_6521;
  wire [6:0] _GEN_6522;
  wire [6:0] _GEN_6523;
  wire [6:0] _GEN_6524;
  wire [6:0] _GEN_6525;
  wire [6:0] _GEN_6526;
  wire [6:0] _GEN_6527;
  wire [6:0] _GEN_6528;
  wire [6:0] _GEN_6529;
  wire [6:0] _GEN_6530;
  wire [6:0] _GEN_6531;
  wire [6:0] _GEN_6532;
  wire [6:0] _GEN_6533;
  wire [6:0] _GEN_6534;
  wire [6:0] _GEN_6535;
  wire [6:0] _GEN_6536;
  wire [6:0] _GEN_6537;
  wire [6:0] _GEN_6778;
  wire [6:0] _GEN_6779;
  wire [6:0] _GEN_6780;
  wire [6:0] _GEN_6781;
  wire [6:0] _GEN_6782;
  wire [6:0] _GEN_6783;
  wire [6:0] _GEN_6784;
  wire [6:0] _GEN_6785;
  wire [6:0] _GEN_6786;
  wire [6:0] _GEN_6787;
  wire [6:0] _GEN_6788;
  wire [6:0] _GEN_6789;
  wire [6:0] _GEN_6790;
  wire [6:0] _GEN_6791;
  wire [6:0] _GEN_6792;
  wire [6:0] _GEN_6793;
  wire [6:0] _GEN_6794;
  wire [6:0] _GEN_6795;
  wire [6:0] _GEN_6796;
  wire [6:0] _GEN_6797;
  wire [6:0] _GEN_6798;
  wire [6:0] _GEN_6799;
  wire [6:0] _GEN_6800;
  wire [6:0] _GEN_6801;
  wire [6:0] _GEN_6802;
  wire [6:0] _GEN_6803;
  wire [6:0] _GEN_6804;
  wire [6:0] _GEN_6805;
  wire [6:0] _GEN_6806;
  wire [6:0] _GEN_6807;
  wire [6:0] _GEN_6808;
  wire [6:0] _GEN_6809;
  wire [6:0] _GEN_6810;
  wire [6:0] _GEN_6811;
  wire [6:0] _GEN_6812;
  wire [6:0] _GEN_6813;
  wire [6:0] _GEN_6814;
  wire [6:0] _GEN_6815;
  wire [6:0] _GEN_6816;
  wire [6:0] _GEN_6817;
  wire  _GEN_7058;
  wire  _GEN_7059;
  wire  _GEN_7060;
  wire  _GEN_7061;
  wire  _GEN_7062;
  wire  _GEN_7063;
  wire  _GEN_7064;
  wire  _GEN_7065;
  wire  _GEN_7066;
  wire  _GEN_7067;
  wire  _GEN_7068;
  wire  _GEN_7069;
  wire  _GEN_7070;
  wire  _GEN_7071;
  wire  _GEN_7072;
  wire  _GEN_7073;
  wire  _GEN_7074;
  wire  _GEN_7075;
  wire  _GEN_7076;
  wire  _GEN_7077;
  wire  _GEN_7078;
  wire  _GEN_7079;
  wire  _GEN_7080;
  wire  _GEN_7081;
  wire  _GEN_7082;
  wire  _GEN_7083;
  wire  _GEN_7084;
  wire  _GEN_7085;
  wire  _GEN_7086;
  wire  _GEN_7087;
  wire  _GEN_7088;
  wire  _GEN_7089;
  wire  _GEN_7090;
  wire  _GEN_7091;
  wire  _GEN_7092;
  wire  _GEN_7093;
  wire  _GEN_7094;
  wire  _GEN_7095;
  wire  _GEN_7096;
  wire  _GEN_7097;
  wire  _GEN_7098;
  wire  _GEN_7099;
  wire  _GEN_7100;
  wire  _GEN_7101;
  wire  _GEN_7102;
  wire  _GEN_7103;
  wire  _GEN_7104;
  wire  _GEN_7105;
  wire  _GEN_7106;
  wire  _GEN_7107;
  wire  _GEN_7108;
  wire  _GEN_7109;
  wire  _GEN_7110;
  wire  _GEN_7111;
  wire  _GEN_7112;
  wire  _GEN_7113;
  wire  _GEN_7114;
  wire  _GEN_7115;
  wire  _GEN_7116;
  wire  _GEN_7117;
  wire  _GEN_7118;
  wire  _GEN_7119;
  wire  _GEN_7120;
  wire  _GEN_7121;
  wire  _GEN_7122;
  wire  _GEN_7123;
  wire  _GEN_7124;
  wire  _GEN_7125;
  wire  _GEN_7126;
  wire  _GEN_7127;
  wire  _GEN_7128;
  wire  _GEN_7129;
  wire  _GEN_7130;
  wire  _GEN_7131;
  wire  _GEN_7132;
  wire  _GEN_7133;
  wire  _GEN_7134;
  wire  _GEN_7135;
  wire  _GEN_7136;
  wire  _GEN_7137;
  wire  _GEN_7178;
  wire  _GEN_7179;
  wire  _GEN_7180;
  wire  _GEN_7181;
  wire  _GEN_7182;
  wire  _GEN_7183;
  wire  _GEN_7184;
  wire  _GEN_7185;
  wire  _GEN_7186;
  wire  _GEN_7187;
  wire  _GEN_7188;
  wire  _GEN_7189;
  wire  _GEN_7190;
  wire  _GEN_7191;
  wire  _GEN_7192;
  wire  _GEN_7193;
  wire  _GEN_7194;
  wire  _GEN_7195;
  wire  _GEN_7196;
  wire  _GEN_7197;
  wire  _GEN_7198;
  wire  _GEN_7199;
  wire  _GEN_7200;
  wire  _GEN_7201;
  wire  _GEN_7202;
  wire  _GEN_7203;
  wire  _GEN_7204;
  wire  _GEN_7205;
  wire  _GEN_7206;
  wire  _GEN_7207;
  wire  _GEN_7208;
  wire  _GEN_7209;
  wire  _GEN_7210;
  wire  _GEN_7211;
  wire  _GEN_7212;
  wire  _GEN_7213;
  wire  _GEN_7214;
  wire  _GEN_7215;
  wire  _GEN_7216;
  wire  _GEN_7217;
  wire  _GEN_7218;
  wire  _GEN_7219;
  wire  _GEN_7220;
  wire  _GEN_7221;
  wire  _GEN_7222;
  wire  _GEN_7223;
  wire  _GEN_7224;
  wire  _GEN_7225;
  wire  _GEN_7226;
  wire  _GEN_7227;
  wire  _GEN_7228;
  wire  _GEN_7229;
  wire  _GEN_7230;
  wire  _GEN_7231;
  wire  _GEN_7232;
  wire  _GEN_7233;
  wire  _GEN_7234;
  wire  _GEN_7235;
  wire  _GEN_7236;
  wire  _GEN_7237;
  wire  _GEN_7238;
  wire  _GEN_7239;
  wire  _GEN_7240;
  wire  _GEN_7241;
  wire  _GEN_7242;
  wire  _GEN_7243;
  wire  _GEN_7244;
  wire  _GEN_7245;
  wire  _GEN_7246;
  wire  _GEN_7247;
  wire  _GEN_7248;
  wire  _GEN_7249;
  wire  _GEN_7250;
  wire  _GEN_7251;
  wire  _GEN_7252;
  wire  _GEN_7253;
  wire  _GEN_7254;
  wire  _GEN_7255;
  wire  _GEN_7256;
  wire  _GEN_7257;
  wire  _GEN_7298;
  wire  _GEN_7299;
  wire  _GEN_7300;
  wire  _GEN_7301;
  wire  _GEN_7302;
  wire  _GEN_7303;
  wire  _GEN_7304;
  wire  _GEN_7305;
  wire  _GEN_7306;
  wire  _GEN_7307;
  wire  _GEN_7308;
  wire  _GEN_7309;
  wire  _GEN_7310;
  wire  _GEN_7311;
  wire  _GEN_7312;
  wire  _GEN_7313;
  wire  _GEN_7314;
  wire  _GEN_7315;
  wire  _GEN_7316;
  wire  _GEN_7317;
  wire  _GEN_7318;
  wire  _GEN_7319;
  wire  _GEN_7320;
  wire  _GEN_7321;
  wire  _GEN_7322;
  wire  _GEN_7323;
  wire  _GEN_7324;
  wire  _GEN_7325;
  wire  _GEN_7326;
  wire  _GEN_7327;
  wire  _GEN_7328;
  wire  _GEN_7329;
  wire  _GEN_7330;
  wire  _GEN_7331;
  wire  _GEN_7332;
  wire  _GEN_7333;
  wire  _GEN_7334;
  wire  _GEN_7335;
  wire  _GEN_7336;
  wire  _GEN_7337;
  wire [5:0] _GEN_7338;
  wire [5:0] _GEN_7339;
  wire [5:0] _GEN_7340;
  wire [5:0] _GEN_7341;
  wire [5:0] _GEN_7342;
  wire [5:0] _GEN_7343;
  wire [5:0] _GEN_7344;
  wire [5:0] _GEN_7345;
  wire [5:0] _GEN_7346;
  wire [5:0] _GEN_7347;
  wire [5:0] _GEN_7348;
  wire [5:0] _GEN_7349;
  wire [5:0] _GEN_7350;
  wire [5:0] _GEN_7351;
  wire [5:0] _GEN_7352;
  wire [5:0] _GEN_7353;
  wire [5:0] _GEN_7354;
  wire [5:0] _GEN_7355;
  wire [5:0] _GEN_7356;
  wire [5:0] _GEN_7357;
  wire [5:0] _GEN_7358;
  wire [5:0] _GEN_7359;
  wire [5:0] _GEN_7360;
  wire [5:0] _GEN_7361;
  wire [5:0] _GEN_7362;
  wire [5:0] _GEN_7363;
  wire [5:0] _GEN_7364;
  wire [5:0] _GEN_7365;
  wire [5:0] _GEN_7366;
  wire [5:0] _GEN_7367;
  wire [5:0] _GEN_7368;
  wire [5:0] _GEN_7369;
  wire [5:0] _GEN_7370;
  wire [5:0] _GEN_7371;
  wire [5:0] _GEN_7372;
  wire [5:0] _GEN_7373;
  wire [5:0] _GEN_7374;
  wire [5:0] _GEN_7375;
  wire [5:0] _GEN_7376;
  wire [5:0] _GEN_7377;
  wire  _GEN_7498;
  wire  _GEN_7499;
  wire  _GEN_7500;
  wire  _GEN_7501;
  wire  _GEN_7502;
  wire  _GEN_7503;
  wire  _GEN_7504;
  wire  _GEN_7505;
  wire  _GEN_7506;
  wire  _GEN_7507;
  wire  _GEN_7508;
  wire  _GEN_7509;
  wire  _GEN_7510;
  wire  _GEN_7511;
  wire  _GEN_7512;
  wire  _GEN_7513;
  wire  _GEN_7514;
  wire  _GEN_7515;
  wire  _GEN_7516;
  wire  _GEN_7517;
  wire  _GEN_7518;
  wire  _GEN_7519;
  wire  _GEN_7520;
  wire  _GEN_7521;
  wire  _GEN_7522;
  wire  _GEN_7523;
  wire  _GEN_7524;
  wire  _GEN_7525;
  wire  _GEN_7526;
  wire  _GEN_7527;
  wire  _GEN_7528;
  wire  _GEN_7529;
  wire  _GEN_7530;
  wire  _GEN_7531;
  wire  _GEN_7532;
  wire  _GEN_7533;
  wire  _GEN_7534;
  wire  _GEN_7535;
  wire  _GEN_7536;
  wire  _GEN_7537;
  wire [1:0] _GEN_7538;
  wire [1:0] _GEN_7539;
  wire [1:0] _GEN_7540;
  wire [1:0] _GEN_7541;
  wire [1:0] _GEN_7542;
  wire [1:0] _GEN_7543;
  wire [1:0] _GEN_7544;
  wire [1:0] _GEN_7545;
  wire [1:0] _GEN_7546;
  wire [1:0] _GEN_7547;
  wire [1:0] _GEN_7548;
  wire [1:0] _GEN_7549;
  wire [1:0] _GEN_7550;
  wire [1:0] _GEN_7551;
  wire [1:0] _GEN_7552;
  wire [1:0] _GEN_7553;
  wire [1:0] _GEN_7554;
  wire [1:0] _GEN_7555;
  wire [1:0] _GEN_7556;
  wire [1:0] _GEN_7557;
  wire [1:0] _GEN_7558;
  wire [1:0] _GEN_7559;
  wire [1:0] _GEN_7560;
  wire [1:0] _GEN_7561;
  wire [1:0] _GEN_7562;
  wire [1:0] _GEN_7563;
  wire [1:0] _GEN_7564;
  wire [1:0] _GEN_7565;
  wire [1:0] _GEN_7566;
  wire [1:0] _GEN_7567;
  wire [1:0] _GEN_7568;
  wire [1:0] _GEN_7569;
  wire [1:0] _GEN_7570;
  wire [1:0] _GEN_7571;
  wire [1:0] _GEN_7572;
  wire [1:0] _GEN_7573;
  wire [1:0] _GEN_7574;
  wire [1:0] _GEN_7575;
  wire [1:0] _GEN_7576;
  wire [1:0] _GEN_7577;
  wire  _GEN_7698;
  wire  _GEN_7699;
  wire  _GEN_7700;
  wire  _GEN_7701;
  wire  _GEN_7702;
  wire  _GEN_7703;
  wire  _GEN_7704;
  wire  _GEN_7705;
  wire  _GEN_7706;
  wire  _GEN_7707;
  wire  _GEN_7708;
  wire  _GEN_7709;
  wire  _GEN_7710;
  wire  _GEN_7711;
  wire  _GEN_7712;
  wire  _GEN_7713;
  wire  _GEN_7714;
  wire  _GEN_7715;
  wire  _GEN_7716;
  wire  _GEN_7717;
  wire  _GEN_7718;
  wire  _GEN_7719;
  wire  _GEN_7720;
  wire  _GEN_7721;
  wire  _GEN_7722;
  wire  _GEN_7723;
  wire  _GEN_7724;
  wire  _GEN_7725;
  wire  _GEN_7726;
  wire  _GEN_7727;
  wire  _GEN_7728;
  wire  _GEN_7729;
  wire  _GEN_7730;
  wire  _GEN_7731;
  wire  _GEN_7732;
  wire  _GEN_7733;
  wire  _GEN_7734;
  wire  _GEN_7735;
  wire  _GEN_7736;
  wire  _GEN_7737;
  wire [6:0] _T_3813;
  wire  _T_3814;
  wire  _T_3816;
  wire  _T_3817;
  wire [5:0] _T_3818;
  wire [6:0] _T_3822;
  wire  _T_3823;
  wire  _T_3825;
  wire  _T_3826;
  wire [5:0] _T_3827;
  wire [6:0] _T_3831;
  wire  _T_3832;
  wire  _T_3834;
  wire  _T_3835;
  wire [5:0] _T_3836;
  wire [6:0] _T_3840;
  wire  _T_3841;
  wire  _T_3843;
  wire  _T_3844;
  wire [5:0] _T_3845;
  wire [6:0] _T_3849;
  wire  _T_3850;
  wire  _T_3852;
  wire  _T_3853;
  wire [5:0] _T_3854;
  wire  _T_3857;
  wire  _T_3859;
  wire  _T_3860;
  wire [6:0] _T_3862;
  wire [5:0] _T_3863;
  wire  _GEN_96;
  wire  _GEN_8040;
  wire  _GEN_8041;
  wire  _GEN_8042;
  wire  _GEN_8043;
  wire  _GEN_8044;
  wire  _GEN_8045;
  wire  _GEN_8046;
  wire  _GEN_8047;
  wire  _GEN_8048;
  wire  _GEN_8049;
  wire  _GEN_8050;
  wire  _GEN_8051;
  wire  _GEN_8052;
  wire  _GEN_8053;
  wire  _GEN_8054;
  wire  _GEN_8055;
  wire  _GEN_8056;
  wire  _GEN_8057;
  wire  _GEN_8058;
  wire  _GEN_8059;
  wire  _GEN_8060;
  wire  _GEN_8061;
  wire  _GEN_8062;
  wire  _GEN_8063;
  wire  _GEN_8064;
  wire  _GEN_8065;
  wire  _GEN_8066;
  wire  _GEN_8067;
  wire  _GEN_8068;
  wire  _GEN_8069;
  wire  _GEN_8070;
  wire  _GEN_8071;
  wire  _GEN_8072;
  wire  _GEN_8073;
  wire  _GEN_8074;
  wire  _GEN_8075;
  wire  _GEN_8076;
  wire  _GEN_8077;
  wire  _GEN_8078;
  wire  _T_3873;
  wire  _T_3875;
  wire [5:0] _T_3876;
  wire  _T_3879;
  wire  _T_3881;
  wire  _T_3883;
  wire  _T_3884;
  wire  _T_3886;
  wire  _T_3887;
  wire [6:0] _T_3889;
  wire [5:0] _T_3890;
  wire  _GEN_97;
  wire  _GEN_8084;
  wire  _GEN_8085;
  wire  _GEN_8086;
  wire  _GEN_8087;
  wire  _GEN_8088;
  wire  _GEN_8089;
  wire  _GEN_8090;
  wire  _GEN_8091;
  wire  _GEN_8092;
  wire  _GEN_8093;
  wire  _GEN_8094;
  wire  _GEN_8095;
  wire  _GEN_8096;
  wire  _GEN_8097;
  wire  _GEN_8098;
  wire  _GEN_8099;
  wire  _GEN_8100;
  wire  _GEN_8101;
  wire  _GEN_8102;
  wire  _GEN_8103;
  wire  _GEN_8104;
  wire  _GEN_8105;
  wire  _GEN_8106;
  wire  _GEN_8107;
  wire  _GEN_8108;
  wire  _GEN_8109;
  wire  _GEN_8110;
  wire  _GEN_8111;
  wire  _GEN_8112;
  wire  _GEN_8113;
  wire  _GEN_8114;
  wire  _GEN_8115;
  wire  _GEN_8116;
  wire  _GEN_8117;
  wire  _GEN_8118;
  wire  _GEN_8119;
  wire  _GEN_8120;
  wire  _GEN_8121;
  wire  _GEN_8122;
  wire  _T_3900;
  wire  _T_3902;
  wire [5:0] _T_3903;
  wire  _T_3906;
  wire  _T_3908;
  wire  _T_3910;
  wire [6:0] _T_3916;
  wire  _T_3975;
  wire  _T_3977;
  wire  _T_3978;
  wire [6:0] _T_3980;
  wire [5:0] _T_3981;
  wire  _T_3983;
  wire  _T_3985;
  wire  _T_3986;
  wire [6:0] _T_3988;
  wire [5:0] _T_3989;
  wire  _T_3991;
  wire  _T_3993;
  wire  _T_3994;
  wire [6:0] _T_3996;
  wire [5:0] _T_3997;
  wire  _T_4000;
  wire  _T_4002;
  wire  _T_4003;
  wire [6:0] _T_4005;
  wire [5:0] _T_4006;
  wire  _GEN_103;
  wire  _GEN_8544;
  wire  _GEN_8545;
  wire  _GEN_8546;
  wire  _GEN_8547;
  wire  _GEN_8548;
  wire  _GEN_8549;
  wire  _GEN_8550;
  wire  _GEN_8551;
  wire  _GEN_8552;
  wire  _GEN_8553;
  wire  _GEN_8554;
  wire  _GEN_8555;
  wire  _GEN_8556;
  wire  _GEN_8557;
  wire  _GEN_8558;
  wire  _GEN_8559;
  wire  _GEN_8560;
  wire  _GEN_8561;
  wire  _GEN_8562;
  wire  _GEN_8563;
  wire  _GEN_8564;
  wire  _GEN_8565;
  wire  _GEN_8566;
  wire  _GEN_8567;
  wire  _GEN_8568;
  wire  _GEN_8569;
  wire  _GEN_8570;
  wire  _GEN_8571;
  wire  _GEN_8572;
  wire  _GEN_8573;
  wire  _GEN_8574;
  wire  _GEN_8575;
  wire  _GEN_8576;
  wire  _GEN_8577;
  wire  _GEN_8578;
  wire  _GEN_8579;
  wire  _GEN_8580;
  wire  _GEN_8581;
  wire  _GEN_8582;
  wire  _T_4013;
  wire  _T_4019;
  wire  _GEN_104;
  wire  _T_4020;
  wire  _T_4022;
  wire  _T_4023;
  wire [5:0] _T_4025;
  wire  _T_4026;
  wire [5:0] _GEN_8583;
  wire [6:0] _GEN_8636;
  wire [6:0] _GEN_8643;
  wire  _GEN_8650;
  wire  _GEN_8651;
  wire  _GEN_8653;
  wire  _GEN_8654;
  wire  _GEN_8656;
  wire [5:0] _GEN_8657;
  wire [1:0] _GEN_8662;
  wire  _GEN_8666;
  wire [6:0] _GEN_8726;
  wire [6:0] _GEN_8733;
  wire  _GEN_8740;
  wire  _GEN_8741;
  wire  _GEN_8743;
  wire  _GEN_8744;
  wire  _GEN_8746;
  wire [5:0] _GEN_8747;
  wire [1:0] _GEN_8752;
  wire  _GEN_8756;
  wire [6:0] _GEN_8816;
  wire [6:0] _GEN_8823;
  wire  _GEN_8830;
  wire  _GEN_8831;
  wire  _GEN_8833;
  wire  _GEN_8834;
  wire  _GEN_8836;
  wire [5:0] _GEN_8837;
  wire [1:0] _GEN_8842;
  wire  _GEN_8846;
  wire [6:0] _GEN_8906;
  wire [6:0] _GEN_8913;
  wire  _GEN_8920;
  wire  _GEN_8921;
  wire  _GEN_8923;
  wire  _GEN_8924;
  wire  _GEN_8926;
  wire [5:0] _GEN_8927;
  wire [1:0] _GEN_8932;
  wire  _GEN_8936;
  wire [6:0] _GEN_8996;
  wire [6:0] _GEN_9003;
  wire  _GEN_9010;
  wire  _GEN_9011;
  wire  _GEN_9013;
  wire  _GEN_9014;
  wire  _GEN_9016;
  wire [5:0] _GEN_9017;
  wire [1:0] _GEN_9022;
  wire  _GEN_9026;
  wire [6:0] _GEN_9086;
  wire [6:0] _GEN_9093;
  wire  _GEN_9100;
  wire  _GEN_9101;
  wire  _GEN_9103;
  wire  _GEN_9104;
  wire  _GEN_9106;
  wire [5:0] _GEN_9107;
  wire [1:0] _GEN_9112;
  wire  _GEN_9116;
  wire [6:0] _GEN_9176;
  wire [6:0] _GEN_9183;
  wire  _GEN_9190;
  wire  _GEN_9191;
  wire  _GEN_9193;
  wire  _GEN_9194;
  wire  _GEN_9196;
  wire [5:0] _GEN_9197;
  wire [1:0] _GEN_9202;
  wire  _GEN_9206;
  wire [6:0] _GEN_9266;
  wire [6:0] _GEN_9273;
  wire  _GEN_9280;
  wire  _GEN_9281;
  wire  _GEN_9283;
  wire  _GEN_9284;
  wire  _GEN_9286;
  wire [5:0] _GEN_9287;
  wire [1:0] _GEN_9292;
  wire  _GEN_9296;
  wire [6:0] _GEN_9356;
  wire [6:0] _GEN_9363;
  wire  _GEN_9370;
  wire  _GEN_9371;
  wire  _GEN_9373;
  wire  _GEN_9374;
  wire  _GEN_9376;
  wire [5:0] _GEN_9377;
  wire [1:0] _GEN_9382;
  wire  _GEN_9386;
  wire [6:0] _GEN_9446;
  wire [6:0] _GEN_9453;
  wire  _GEN_9460;
  wire  _GEN_9461;
  wire  _GEN_9463;
  wire  _GEN_9464;
  wire  _GEN_9466;
  wire [5:0] _GEN_9467;
  wire [1:0] _GEN_9472;
  wire  _GEN_9476;
  wire [6:0] _GEN_9536;
  wire [6:0] _GEN_9543;
  wire  _GEN_9550;
  wire  _GEN_9551;
  wire  _GEN_9553;
  wire  _GEN_9554;
  wire  _GEN_9556;
  wire [5:0] _GEN_9557;
  wire [1:0] _GEN_9562;
  wire  _GEN_9566;
  wire [6:0] _GEN_9626;
  wire [6:0] _GEN_9633;
  wire  _GEN_9640;
  wire  _GEN_9641;
  wire  _GEN_9643;
  wire  _GEN_9644;
  wire  _GEN_9646;
  wire [5:0] _GEN_9647;
  wire [1:0] _GEN_9652;
  wire  _GEN_9656;
  wire [6:0] _GEN_9716;
  wire [6:0] _GEN_9723;
  wire  _GEN_9730;
  wire  _GEN_9731;
  wire  _GEN_9733;
  wire  _GEN_9734;
  wire  _GEN_9736;
  wire [5:0] _GEN_9737;
  wire [1:0] _GEN_9742;
  wire  _GEN_9746;
  wire [6:0] _GEN_9806;
  wire [6:0] _GEN_9813;
  wire  _GEN_9820;
  wire  _GEN_9821;
  wire  _GEN_9823;
  wire  _GEN_9824;
  wire  _GEN_9826;
  wire [5:0] _GEN_9827;
  wire [1:0] _GEN_9832;
  wire  _GEN_9836;
  wire [6:0] _GEN_9896;
  wire [6:0] _GEN_9903;
  wire  _GEN_9910;
  wire  _GEN_9911;
  wire  _GEN_9913;
  wire  _GEN_9914;
  wire  _GEN_9916;
  wire [5:0] _GEN_9917;
  wire [1:0] _GEN_9922;
  wire  _GEN_9926;
  wire [6:0] _GEN_9986;
  wire [6:0] _GEN_9993;
  wire  _GEN_10000;
  wire  _GEN_10001;
  wire  _GEN_10003;
  wire  _GEN_10004;
  wire  _GEN_10006;
  wire [5:0] _GEN_10007;
  wire [1:0] _GEN_10012;
  wire  _GEN_10016;
  wire [6:0] _GEN_10076;
  wire [6:0] _GEN_10083;
  wire  _GEN_10090;
  wire  _GEN_10091;
  wire  _GEN_10093;
  wire  _GEN_10094;
  wire  _GEN_10096;
  wire [5:0] _GEN_10097;
  wire [1:0] _GEN_10102;
  wire  _GEN_10106;
  wire [6:0] _GEN_10166;
  wire [6:0] _GEN_10173;
  wire  _GEN_10180;
  wire  _GEN_10181;
  wire  _GEN_10183;
  wire  _GEN_10184;
  wire  _GEN_10186;
  wire [5:0] _GEN_10187;
  wire [1:0] _GEN_10192;
  wire  _GEN_10196;
  wire [6:0] _GEN_10256;
  wire [6:0] _GEN_10263;
  wire  _GEN_10270;
  wire  _GEN_10271;
  wire  _GEN_10273;
  wire  _GEN_10274;
  wire  _GEN_10276;
  wire [5:0] _GEN_10277;
  wire [1:0] _GEN_10282;
  wire  _GEN_10286;
  wire [6:0] _GEN_10346;
  wire [6:0] _GEN_10353;
  wire  _GEN_10360;
  wire  _GEN_10361;
  wire  _GEN_10363;
  wire  _GEN_10364;
  wire  _GEN_10366;
  wire [5:0] _GEN_10367;
  wire [1:0] _GEN_10372;
  wire  _GEN_10376;
  wire [6:0] _GEN_10436;
  wire [6:0] _GEN_10443;
  wire  _GEN_10450;
  wire  _GEN_10451;
  wire  _GEN_10453;
  wire  _GEN_10454;
  wire  _GEN_10456;
  wire [5:0] _GEN_10457;
  wire [1:0] _GEN_10462;
  wire  _GEN_10466;
  wire [6:0] _GEN_10526;
  wire [6:0] _GEN_10533;
  wire  _GEN_10540;
  wire  _GEN_10541;
  wire  _GEN_10543;
  wire  _GEN_10544;
  wire  _GEN_10546;
  wire [5:0] _GEN_10547;
  wire [1:0] _GEN_10552;
  wire  _GEN_10556;
  wire [6:0] _GEN_10616;
  wire [6:0] _GEN_10623;
  wire  _GEN_10630;
  wire  _GEN_10631;
  wire  _GEN_10633;
  wire  _GEN_10634;
  wire  _GEN_10636;
  wire [5:0] _GEN_10637;
  wire [1:0] _GEN_10642;
  wire  _GEN_10646;
  wire [6:0] _GEN_10706;
  wire [6:0] _GEN_10713;
  wire  _GEN_10720;
  wire  _GEN_10721;
  wire  _GEN_10723;
  wire  _GEN_10724;
  wire  _GEN_10726;
  wire [5:0] _GEN_10727;
  wire [1:0] _GEN_10732;
  wire  _GEN_10736;
  wire [6:0] _GEN_10796;
  wire [6:0] _GEN_10803;
  wire  _GEN_10810;
  wire  _GEN_10811;
  wire  _GEN_10813;
  wire  _GEN_10814;
  wire  _GEN_10816;
  wire [5:0] _GEN_10817;
  wire [1:0] _GEN_10822;
  wire  _GEN_10826;
  wire [6:0] _GEN_10886;
  wire [6:0] _GEN_10893;
  wire  _GEN_10900;
  wire  _GEN_10901;
  wire  _GEN_10903;
  wire  _GEN_10904;
  wire  _GEN_10906;
  wire [5:0] _GEN_10907;
  wire [1:0] _GEN_10912;
  wire  _GEN_10916;
  wire [6:0] _GEN_10976;
  wire [6:0] _GEN_10983;
  wire  _GEN_10990;
  wire  _GEN_10991;
  wire  _GEN_10993;
  wire  _GEN_10994;
  wire  _GEN_10996;
  wire [5:0] _GEN_10997;
  wire [1:0] _GEN_11002;
  wire  _GEN_11006;
  wire [6:0] _GEN_11066;
  wire [6:0] _GEN_11073;
  wire  _GEN_11080;
  wire  _GEN_11081;
  wire  _GEN_11083;
  wire  _GEN_11084;
  wire  _GEN_11086;
  wire [5:0] _GEN_11087;
  wire [1:0] _GEN_11092;
  wire  _GEN_11096;
  wire [6:0] _GEN_11156;
  wire [6:0] _GEN_11163;
  wire  _GEN_11170;
  wire  _GEN_11171;
  wire  _GEN_11173;
  wire  _GEN_11174;
  wire  _GEN_11176;
  wire [5:0] _GEN_11177;
  wire [1:0] _GEN_11182;
  wire  _GEN_11186;
  wire [6:0] _GEN_11246;
  wire [6:0] _GEN_11253;
  wire  _GEN_11260;
  wire  _GEN_11261;
  wire  _GEN_11263;
  wire  _GEN_11264;
  wire  _GEN_11266;
  wire [5:0] _GEN_11267;
  wire [1:0] _GEN_11272;
  wire  _GEN_11276;
  wire [6:0] _GEN_11336;
  wire [6:0] _GEN_11343;
  wire  _GEN_11350;
  wire  _GEN_11351;
  wire  _GEN_11353;
  wire  _GEN_11354;
  wire  _GEN_11356;
  wire [5:0] _GEN_11357;
  wire [1:0] _GEN_11362;
  wire  _GEN_11366;
  wire [6:0] _GEN_11426;
  wire [6:0] _GEN_11433;
  wire  _GEN_11440;
  wire  _GEN_11441;
  wire  _GEN_11443;
  wire  _GEN_11444;
  wire  _GEN_11446;
  wire [5:0] _GEN_11447;
  wire [1:0] _GEN_11452;
  wire  _GEN_11456;
  wire [6:0] _GEN_11516;
  wire [6:0] _GEN_11523;
  wire  _GEN_11530;
  wire  _GEN_11531;
  wire  _GEN_11533;
  wire  _GEN_11534;
  wire  _GEN_11536;
  wire [5:0] _GEN_11537;
  wire [1:0] _GEN_11542;
  wire  _GEN_11546;
  wire [6:0] _GEN_11606;
  wire [6:0] _GEN_11613;
  wire  _GEN_11620;
  wire  _GEN_11621;
  wire  _GEN_11623;
  wire  _GEN_11624;
  wire  _GEN_11626;
  wire [5:0] _GEN_11627;
  wire [1:0] _GEN_11632;
  wire  _GEN_11636;
  wire [6:0] _GEN_11696;
  wire [6:0] _GEN_11703;
  wire  _GEN_11710;
  wire  _GEN_11711;
  wire  _GEN_11713;
  wire  _GEN_11714;
  wire  _GEN_11716;
  wire [5:0] _GEN_11717;
  wire [1:0] _GEN_11722;
  wire  _GEN_11726;
  wire [6:0] _GEN_11786;
  wire [6:0] _GEN_11793;
  wire  _GEN_11800;
  wire  _GEN_11801;
  wire  _GEN_11803;
  wire  _GEN_11804;
  wire  _GEN_11806;
  wire [5:0] _GEN_11807;
  wire [1:0] _GEN_11812;
  wire  _GEN_11816;
  wire [6:0] _GEN_11876;
  wire [6:0] _GEN_11883;
  wire  _GEN_11890;
  wire  _GEN_11891;
  wire  _GEN_11893;
  wire  _GEN_11894;
  wire  _GEN_11896;
  wire [5:0] _GEN_11897;
  wire [1:0] _GEN_11902;
  wire  _GEN_11906;
  wire [6:0] _GEN_11966;
  wire [6:0] _GEN_11973;
  wire  _GEN_11980;
  wire  _GEN_11981;
  wire  _GEN_11983;
  wire  _GEN_11984;
  wire  _GEN_11986;
  wire [5:0] _GEN_11987;
  wire [1:0] _GEN_11992;
  wire  _GEN_11996;
  wire [6:0] _GEN_12056;
  wire [6:0] _GEN_12063;
  wire  _GEN_12070;
  wire  _GEN_12071;
  wire  _GEN_12073;
  wire  _GEN_12074;
  wire  _GEN_12076;
  wire [5:0] _GEN_12077;
  wire [1:0] _GEN_12082;
  wire  _GEN_12086;
  wire [6:0] _GEN_157_pdst;
  wire [6:0] _GEN_164_stale_pdst;
  wire  _GEN_171_is_fencei;
  wire  _GEN_172_is_store;
  wire  _GEN_174_is_load;
  wire  _GEN_175_is_sys_pc2epc;
  wire  _GEN_177_flush_on_commit;
  wire [5:0] _GEN_178_ldst;
  wire [1:0] _GEN_183_dst_rtype;
  wire  _GEN_187_fp_val;
  wire  _GEN_195;
  wire  _GEN_12094;
  wire  _GEN_12095;
  wire  _GEN_12096;
  wire  _GEN_12097;
  wire  _GEN_12098;
  wire  _GEN_12099;
  wire  _GEN_12100;
  wire  _GEN_12101;
  wire  _GEN_12102;
  wire  _GEN_12103;
  wire  _GEN_12104;
  wire  _GEN_12105;
  wire  _GEN_12106;
  wire  _GEN_12107;
  wire  _GEN_12108;
  wire  _GEN_12109;
  wire  _GEN_12110;
  wire  _GEN_12111;
  wire  _GEN_12112;
  wire  _GEN_12113;
  wire  _GEN_12114;
  wire  _GEN_12115;
  wire  _GEN_12116;
  wire  _GEN_12117;
  wire  _GEN_12118;
  wire  _GEN_12119;
  wire  _GEN_12120;
  wire  _GEN_12121;
  wire  _GEN_12122;
  wire  _GEN_12123;
  wire  _GEN_12124;
  wire  _GEN_12125;
  wire  _GEN_12126;
  wire  _GEN_12127;
  wire  _GEN_12128;
  wire  _GEN_12129;
  wire  _GEN_12130;
  wire  _GEN_12131;
  wire  _GEN_12132;
  wire  _T_4046;
  wire [1:0] _GEN_196_dst_rtype;
  wire  _T_4059;
  wire [1:0] _GEN_197_dst_rtype;
  wire  _T_4072;
  wire  _T_4073;
  wire  _T_4074;
  wire  _T_4077;
  wire  _GEN_19153;
  wire  _GEN_19154;
  wire  _GEN_19155;
  wire  _GEN_19156;
  wire  _GEN_19157;
  wire  _GEN_19158;
  wire  _GEN_19159;
  wire  _GEN_19160;
  wire  _GEN_19161;
  wire  _GEN_19162;
  wire  _GEN_19163;
  wire  _GEN_19164;
  wire  _GEN_19165;
  wire  _GEN_19166;
  wire  _GEN_19167;
  wire  _GEN_19168;
  wire  _GEN_19169;
  wire  _GEN_19170;
  wire  _GEN_19171;
  wire  _GEN_19172;
  wire  _GEN_19173;
  wire  _GEN_19174;
  wire  _GEN_19175;
  wire  _GEN_19176;
  wire  _GEN_19177;
  wire  _GEN_19178;
  wire  _GEN_19179;
  wire  _GEN_19180;
  wire  _GEN_19181;
  wire  _GEN_19182;
  wire  _GEN_19183;
  wire  _GEN_19184;
  wire  _GEN_19185;
  wire  _GEN_19186;
  wire  _GEN_19187;
  wire  _GEN_19188;
  wire  _GEN_19189;
  wire  _GEN_19190;
  wire  _GEN_19191;
  wire  _GEN_19192;
  wire  _GEN_19193;
  wire  _GEN_19194;
  wire  _GEN_19195;
  wire  _GEN_19196;
  wire  _GEN_19197;
  wire  _GEN_19198;
  wire  _GEN_19199;
  wire  _GEN_19200;
  wire  _GEN_19201;
  wire  _GEN_19202;
  wire  _GEN_19203;
  wire  _GEN_19204;
  wire  _GEN_19205;
  wire  _GEN_19206;
  wire  _GEN_19207;
  wire  _GEN_19208;
  wire  _GEN_19209;
  wire  _GEN_19210;
  wire  _GEN_19211;
  wire  _GEN_19212;
  wire  _GEN_19213;
  wire  _GEN_19214;
  wire  _GEN_19215;
  wire  _GEN_19216;
  wire  _GEN_19217;
  wire  _GEN_19218;
  wire  _GEN_19219;
  wire  _GEN_19220;
  wire  _GEN_19221;
  wire  _GEN_19222;
  wire  _GEN_19223;
  wire  _GEN_19224;
  wire  _GEN_19225;
  wire  _GEN_19226;
  wire  _GEN_19227;
  wire  _GEN_19228;
  wire  _GEN_19229;
  wire  _GEN_19230;
  wire  _GEN_19231;
  wire  _GEN_19232;
  wire [7:0] _T_4090;
  wire  _T_4092;
  wire  _T_4093;
  wire  _T_4094;
  wire  _T_4095;
  wire  _T_4108;
  wire  _T_4109;
  wire  _T_4110;
  wire [7:0] _T_4111;
  wire [7:0] _T_4112;
  wire [7:0] _GEN_19237;
  wire  _GEN_19238;
  wire [7:0] _GEN_19240;
  wire [7:0] _T_4113;
  wire  _T_4115;
  wire  _T_4116;
  wire  _T_4118;
  wire  _T_4133;
  wire [7:0] _T_4135;
  wire [7:0] _GEN_19241;
  wire  _GEN_19242;
  wire [7:0] _GEN_19244;
  wire [7:0] _T_4136;
  wire  _T_4138;
  wire  _T_4139;
  wire  _T_4141;
  wire  _T_4156;
  wire [7:0] _T_4158;
  wire [7:0] _GEN_19245;
  wire  _GEN_19246;
  wire [7:0] _GEN_19248;
  wire [7:0] _T_4159;
  wire  _T_4161;
  wire  _T_4162;
  wire  _T_4164;
  wire  _T_4179;
  wire [7:0] _T_4181;
  wire [7:0] _GEN_19249;
  wire  _GEN_19250;
  wire [7:0] _GEN_19252;
  wire [7:0] _T_4182;
  wire  _T_4184;
  wire  _T_4185;
  wire  _T_4187;
  wire  _T_4202;
  wire [7:0] _T_4204;
  wire [7:0] _GEN_19253;
  wire  _GEN_19254;
  wire [7:0] _GEN_19256;
  wire [7:0] _T_4205;
  wire  _T_4207;
  wire  _T_4208;
  wire  _T_4210;
  wire  _T_4225;
  wire [7:0] _T_4227;
  wire [7:0] _GEN_19257;
  wire  _GEN_19258;
  wire [7:0] _GEN_19260;
  wire [7:0] _T_4228;
  wire  _T_4230;
  wire  _T_4231;
  wire  _T_4233;
  wire  _T_4248;
  wire [7:0] _T_4250;
  wire [7:0] _GEN_19261;
  wire  _GEN_19262;
  wire [7:0] _GEN_19264;
  wire [7:0] _T_4251;
  wire  _T_4253;
  wire  _T_4254;
  wire  _T_4256;
  wire  _T_4271;
  wire [7:0] _T_4273;
  wire [7:0] _GEN_19265;
  wire  _GEN_19266;
  wire [7:0] _GEN_19268;
  wire [7:0] _T_4274;
  wire  _T_4276;
  wire  _T_4277;
  wire  _T_4279;
  wire  _T_4294;
  wire [7:0] _T_4296;
  wire [7:0] _GEN_19269;
  wire  _GEN_19270;
  wire [7:0] _GEN_19272;
  wire [7:0] _T_4297;
  wire  _T_4299;
  wire  _T_4300;
  wire  _T_4302;
  wire  _T_4317;
  wire [7:0] _T_4319;
  wire [7:0] _GEN_19273;
  wire  _GEN_19274;
  wire [7:0] _GEN_19276;
  wire [7:0] _T_4320;
  wire  _T_4322;
  wire  _T_4323;
  wire  _T_4325;
  wire  _T_4340;
  wire [7:0] _T_4342;
  wire [7:0] _GEN_19277;
  wire  _GEN_19278;
  wire [7:0] _GEN_19280;
  wire [7:0] _T_4343;
  wire  _T_4345;
  wire  _T_4346;
  wire  _T_4348;
  wire  _T_4363;
  wire [7:0] _T_4365;
  wire [7:0] _GEN_19281;
  wire  _GEN_19282;
  wire [7:0] _GEN_19284;
  wire [7:0] _T_4366;
  wire  _T_4368;
  wire  _T_4369;
  wire  _T_4371;
  wire  _T_4386;
  wire [7:0] _T_4388;
  wire [7:0] _GEN_19285;
  wire  _GEN_19286;
  wire [7:0] _GEN_19288;
  wire [7:0] _T_4389;
  wire  _T_4391;
  wire  _T_4392;
  wire  _T_4394;
  wire  _T_4409;
  wire [7:0] _T_4411;
  wire [7:0] _GEN_19289;
  wire  _GEN_19290;
  wire [7:0] _GEN_19292;
  wire [7:0] _T_4412;
  wire  _T_4414;
  wire  _T_4415;
  wire  _T_4417;
  wire  _T_4432;
  wire [7:0] _T_4434;
  wire [7:0] _GEN_19293;
  wire  _GEN_19294;
  wire [7:0] _GEN_19296;
  wire [7:0] _T_4435;
  wire  _T_4437;
  wire  _T_4438;
  wire  _T_4440;
  wire  _T_4455;
  wire [7:0] _T_4457;
  wire [7:0] _GEN_19297;
  wire  _GEN_19298;
  wire [7:0] _GEN_19300;
  wire [7:0] _T_4458;
  wire  _T_4460;
  wire  _T_4461;
  wire  _T_4463;
  wire  _T_4478;
  wire [7:0] _T_4480;
  wire [7:0] _GEN_19301;
  wire  _GEN_19302;
  wire [7:0] _GEN_19304;
  wire [7:0] _T_4481;
  wire  _T_4483;
  wire  _T_4484;
  wire  _T_4486;
  wire  _T_4501;
  wire [7:0] _T_4503;
  wire [7:0] _GEN_19305;
  wire  _GEN_19306;
  wire [7:0] _GEN_19308;
  wire [7:0] _T_4504;
  wire  _T_4506;
  wire  _T_4507;
  wire  _T_4509;
  wire  _T_4524;
  wire [7:0] _T_4526;
  wire [7:0] _GEN_19309;
  wire  _GEN_19310;
  wire [7:0] _GEN_19312;
  wire [7:0] _T_4527;
  wire  _T_4529;
  wire  _T_4530;
  wire  _T_4532;
  wire  _T_4547;
  wire [7:0] _T_4549;
  wire [7:0] _GEN_19313;
  wire  _GEN_19314;
  wire [7:0] _GEN_19316;
  wire [7:0] _T_4550;
  wire  _T_4552;
  wire  _T_4553;
  wire  _T_4555;
  wire  _T_4570;
  wire [7:0] _T_4572;
  wire [7:0] _GEN_19317;
  wire  _GEN_19318;
  wire [7:0] _GEN_19320;
  wire [7:0] _T_4573;
  wire  _T_4575;
  wire  _T_4576;
  wire  _T_4578;
  wire  _T_4593;
  wire [7:0] _T_4595;
  wire [7:0] _GEN_19321;
  wire  _GEN_19322;
  wire [7:0] _GEN_19324;
  wire [7:0] _T_4596;
  wire  _T_4598;
  wire  _T_4599;
  wire  _T_4601;
  wire  _T_4616;
  wire [7:0] _T_4618;
  wire [7:0] _GEN_19325;
  wire  _GEN_19326;
  wire [7:0] _GEN_19328;
  wire [7:0] _T_4619;
  wire  _T_4621;
  wire  _T_4622;
  wire  _T_4624;
  wire  _T_4639;
  wire [7:0] _T_4641;
  wire [7:0] _GEN_19329;
  wire  _GEN_19330;
  wire [7:0] _GEN_19332;
  wire [7:0] _T_4642;
  wire  _T_4644;
  wire  _T_4645;
  wire  _T_4647;
  wire  _T_4662;
  wire [7:0] _T_4664;
  wire [7:0] _GEN_19333;
  wire  _GEN_19334;
  wire [7:0] _GEN_19336;
  wire [7:0] _T_4665;
  wire  _T_4667;
  wire  _T_4668;
  wire  _T_4670;
  wire  _T_4685;
  wire [7:0] _T_4687;
  wire [7:0] _GEN_19337;
  wire  _GEN_19338;
  wire [7:0] _GEN_19340;
  wire [7:0] _T_4688;
  wire  _T_4690;
  wire  _T_4691;
  wire  _T_4693;
  wire  _T_4708;
  wire [7:0] _T_4710;
  wire [7:0] _GEN_19341;
  wire  _GEN_19342;
  wire [7:0] _GEN_19344;
  wire [7:0] _T_4711;
  wire  _T_4713;
  wire  _T_4714;
  wire  _T_4716;
  wire  _T_4731;
  wire [7:0] _T_4733;
  wire [7:0] _GEN_19345;
  wire  _GEN_19346;
  wire [7:0] _GEN_19348;
  wire [7:0] _T_4734;
  wire  _T_4736;
  wire  _T_4737;
  wire  _T_4739;
  wire  _T_4754;
  wire [7:0] _T_4756;
  wire [7:0] _GEN_19349;
  wire  _GEN_19350;
  wire [7:0] _GEN_19352;
  wire [7:0] _T_4757;
  wire  _T_4759;
  wire  _T_4760;
  wire  _T_4762;
  wire  _T_4777;
  wire [7:0] _T_4779;
  wire [7:0] _GEN_19353;
  wire  _GEN_19354;
  wire [7:0] _GEN_19356;
  wire [7:0] _T_4780;
  wire  _T_4782;
  wire  _T_4783;
  wire  _T_4785;
  wire  _T_4800;
  wire [7:0] _T_4802;
  wire [7:0] _GEN_19357;
  wire  _GEN_19358;
  wire [7:0] _GEN_19360;
  wire [7:0] _T_4803;
  wire  _T_4805;
  wire  _T_4806;
  wire  _T_4808;
  wire  _T_4823;
  wire [7:0] _T_4825;
  wire [7:0] _GEN_19361;
  wire  _GEN_19362;
  wire [7:0] _GEN_19364;
  wire [7:0] _T_4826;
  wire  _T_4828;
  wire  _T_4829;
  wire  _T_4831;
  wire  _T_4846;
  wire [7:0] _T_4848;
  wire [7:0] _GEN_19365;
  wire  _GEN_19366;
  wire [7:0] _GEN_19368;
  wire [7:0] _T_4849;
  wire  _T_4851;
  wire  _T_4852;
  wire  _T_4854;
  wire  _T_4869;
  wire [7:0] _T_4871;
  wire [7:0] _GEN_19369;
  wire  _GEN_19370;
  wire [7:0] _GEN_19372;
  wire [7:0] _T_4872;
  wire  _T_4874;
  wire  _T_4875;
  wire  _T_4877;
  wire  _T_4892;
  wire [7:0] _T_4894;
  wire [7:0] _GEN_19373;
  wire  _GEN_19374;
  wire [7:0] _GEN_19376;
  wire [7:0] _T_4895;
  wire  _T_4897;
  wire  _T_4898;
  wire  _T_4900;
  wire  _T_4915;
  wire [7:0] _T_4917;
  wire [7:0] _GEN_19377;
  wire  _GEN_19378;
  wire [7:0] _GEN_19380;
  wire [7:0] _T_4918;
  wire  _T_4920;
  wire  _T_4921;
  wire  _T_4923;
  wire  _T_4938;
  wire [7:0] _T_4940;
  wire [7:0] _GEN_19381;
  wire  _GEN_19382;
  wire [7:0] _GEN_19384;
  wire [7:0] _T_4941;
  wire  _T_4943;
  wire  _T_4944;
  wire  _T_4946;
  wire  _T_4961;
  wire [7:0] _T_4963;
  wire [7:0] _GEN_19385;
  wire  _GEN_19386;
  wire [7:0] _GEN_19388;
  wire [7:0] _T_4964;
  wire  _T_4966;
  wire  _T_4967;
  wire  _T_4969;
  wire  _T_4984;
  wire [7:0] _T_4986;
  wire [7:0] _GEN_19389;
  wire  _GEN_19390;
  wire [7:0] _GEN_19392;
  wire [7:0] _T_4987;
  wire  _T_4989;
  wire  _T_4990;
  wire  _T_4992;
  wire  _T_5007;
  wire [7:0] _T_5009;
  wire [7:0] _GEN_19393;
  wire  _GEN_19394;
  wire [7:0] _GEN_19396;
  wire  _GEN_19397;
  wire  _GEN_19398;
  wire  _GEN_19399;
  wire  _GEN_19400;
  wire  _GEN_19401;
  wire  _GEN_19402;
  wire  _GEN_19403;
  wire  _GEN_19404;
  wire  _GEN_19405;
  wire  _GEN_19406;
  wire  _GEN_19407;
  wire  _GEN_19408;
  wire  _GEN_19409;
  wire  _GEN_19410;
  wire  _GEN_19411;
  wire  _GEN_19412;
  wire  _GEN_19413;
  wire  _GEN_19414;
  wire  _GEN_19415;
  wire  _GEN_19416;
  wire  _GEN_19417;
  wire  _GEN_19418;
  wire  _GEN_19419;
  wire  _GEN_19420;
  wire  _GEN_19421;
  wire  _GEN_19422;
  wire  _GEN_19423;
  wire  _GEN_19424;
  wire  _GEN_19425;
  wire  _GEN_19426;
  wire  _GEN_19427;
  wire  _GEN_19428;
  wire  _GEN_19429;
  wire  _GEN_19430;
  wire  _GEN_19431;
  wire  _GEN_19432;
  wire  _GEN_19433;
  wire  _GEN_19434;
  wire  _GEN_19435;
  wire  _GEN_19436;
  wire  _GEN_19437;
  wire  _GEN_19438;
  wire  _GEN_19439;
  wire  _GEN_19440;
  wire  _GEN_19441;
  wire  _GEN_19442;
  wire  _GEN_19443;
  wire  _GEN_19444;
  wire  _GEN_19445;
  wire  _GEN_19446;
  wire  _GEN_19447;
  wire  _GEN_19448;
  wire  _GEN_19449;
  wire  _GEN_19450;
  wire  _GEN_19451;
  wire  _GEN_19452;
  wire  _GEN_19453;
  wire  _GEN_19454;
  wire  _GEN_19455;
  wire  _GEN_19456;
  wire  _GEN_19457;
  wire  _GEN_19458;
  wire  _GEN_19459;
  wire  _GEN_19460;
  wire  _GEN_19461;
  wire  _GEN_19462;
  wire  _GEN_19463;
  wire  _GEN_19464;
  wire  _GEN_19465;
  wire  _GEN_19466;
  wire  _GEN_19467;
  wire  _GEN_19468;
  wire  _GEN_19469;
  wire  _GEN_19470;
  wire  _GEN_19471;
  wire  _GEN_19472;
  wire  _GEN_19473;
  wire  _GEN_19474;
  wire  _GEN_19475;
  wire  _GEN_19476;
  wire  _GEN_200;
  wire  _GEN_201_is_store;
  wire  _GEN_19544;
  wire  _GEN_19546;
  wire  _GEN_19634;
  wire  _GEN_19636;
  wire  _GEN_19724;
  wire  _GEN_19726;
  wire  _GEN_19814;
  wire  _GEN_19816;
  wire  _GEN_19904;
  wire  _GEN_19906;
  wire  _GEN_19994;
  wire  _GEN_19996;
  wire  _GEN_20084;
  wire  _GEN_20086;
  wire  _GEN_20174;
  wire  _GEN_20176;
  wire  _GEN_20264;
  wire  _GEN_20266;
  wire  _GEN_20354;
  wire  _GEN_20356;
  wire  _GEN_20444;
  wire  _GEN_20446;
  wire  _GEN_20534;
  wire  _GEN_20536;
  wire  _GEN_20624;
  wire  _GEN_20626;
  wire  _GEN_20714;
  wire  _GEN_20716;
  wire  _GEN_20804;
  wire  _GEN_20806;
  wire  _GEN_20894;
  wire  _GEN_20896;
  wire  _GEN_20984;
  wire  _GEN_20986;
  wire  _GEN_21074;
  wire  _GEN_21076;
  wire  _GEN_21164;
  wire  _GEN_21166;
  wire  _GEN_21254;
  wire  _GEN_21256;
  wire  _GEN_21344;
  wire  _GEN_21346;
  wire  _GEN_21434;
  wire  _GEN_21436;
  wire  _GEN_21524;
  wire  _GEN_21526;
  wire  _GEN_21614;
  wire  _GEN_21616;
  wire  _GEN_21704;
  wire  _GEN_21706;
  wire  _GEN_21794;
  wire  _GEN_21796;
  wire  _GEN_21884;
  wire  _GEN_21886;
  wire  _GEN_21974;
  wire  _GEN_21976;
  wire  _GEN_22064;
  wire  _GEN_22066;
  wire  _GEN_22154;
  wire  _GEN_22156;
  wire  _GEN_22244;
  wire  _GEN_22246;
  wire  _GEN_22334;
  wire  _GEN_22336;
  wire  _GEN_22424;
  wire  _GEN_22426;
  wire  _GEN_22514;
  wire  _GEN_22516;
  wire  _GEN_22604;
  wire  _GEN_22606;
  wire  _GEN_22694;
  wire  _GEN_22696;
  wire  _GEN_22784;
  wire  _GEN_22786;
  wire  _GEN_22874;
  wire  _GEN_22876;
  wire  _GEN_22964;
  wire  _GEN_22966;
  wire  _GEN_202_is_load;
  wire  _GEN_203;
  wire  _GEN_22987;
  wire  _GEN_22988;
  wire  _GEN_22989;
  wire  _GEN_22990;
  wire  _GEN_22991;
  wire  _GEN_22992;
  wire  _GEN_22993;
  wire  _GEN_22994;
  wire  _GEN_22995;
  wire  _GEN_22996;
  wire  _GEN_22997;
  wire  _GEN_22998;
  wire  _GEN_22999;
  wire  _GEN_23000;
  wire  _GEN_23001;
  wire  _GEN_23002;
  wire  _GEN_23003;
  wire  _GEN_23004;
  wire  _GEN_23005;
  wire  _GEN_23006;
  wire  _GEN_23007;
  wire  _GEN_23008;
  wire  _GEN_23009;
  wire  _GEN_23010;
  wire  _GEN_23011;
  wire  _GEN_23012;
  wire  _GEN_23013;
  wire  _GEN_23014;
  wire  _GEN_23015;
  wire  _GEN_23016;
  wire  _GEN_23017;
  wire  _GEN_23018;
  wire  _GEN_23019;
  wire  _GEN_23020;
  wire  _GEN_23021;
  wire  _GEN_23022;
  wire  _GEN_23023;
  wire  _GEN_23024;
  wire  _GEN_23025;
  wire  _T_5045;
  wire [7:0] _T_5048;
  wire [6:0] _T_5049;
  wire [6:0] _T_5050;
  wire [5:0] _T_5054;
  wire  _GEN_204;
  wire  _GEN_23026;
  wire  _GEN_23027;
  wire  _GEN_23028;
  wire  _GEN_23029;
  wire  _GEN_23030;
  wire  _GEN_23031;
  wire  _GEN_23032;
  wire  _GEN_23033;
  wire  _GEN_23034;
  wire  _GEN_23035;
  wire  _GEN_23036;
  wire  _GEN_23037;
  wire  _GEN_23038;
  wire  _GEN_23039;
  wire  _GEN_23040;
  wire  _GEN_23041;
  wire  _GEN_23042;
  wire  _GEN_23043;
  wire  _GEN_23044;
  wire  _GEN_23045;
  wire  _GEN_23046;
  wire  _GEN_23047;
  wire  _GEN_23048;
  wire  _GEN_23049;
  wire  _GEN_23050;
  wire  _GEN_23051;
  wire  _GEN_23052;
  wire  _GEN_23053;
  wire  _GEN_23054;
  wire  _GEN_23055;
  wire  _GEN_23056;
  wire  _GEN_23057;
  wire  _GEN_23058;
  wire  _GEN_23059;
  wire  _GEN_23060;
  wire  _GEN_23061;
  wire  _GEN_23062;
  wire  _GEN_23063;
  wire  _GEN_23064;
  wire  _GEN_208;
  wire  _GEN_23305;
  wire  _GEN_23306;
  wire  _GEN_23307;
  wire  _GEN_23308;
  wire  _GEN_23309;
  wire  _GEN_23310;
  wire  _GEN_23311;
  wire  _GEN_23312;
  wire  _GEN_23313;
  wire  _GEN_23314;
  wire  _GEN_23315;
  wire  _GEN_23316;
  wire  _GEN_23317;
  wire  _GEN_23318;
  wire  _GEN_23319;
  wire  _GEN_23320;
  wire  _GEN_23321;
  wire  _GEN_23322;
  wire  _GEN_23323;
  wire  _GEN_23324;
  wire  _GEN_23325;
  wire  _GEN_23326;
  wire  _GEN_23327;
  wire  _GEN_23328;
  wire  _GEN_23329;
  wire  _GEN_23330;
  wire  _GEN_23331;
  wire  _GEN_23332;
  wire  _GEN_23333;
  wire  _GEN_23334;
  wire  _GEN_23335;
  wire  _GEN_23336;
  wire  _GEN_23337;
  wire  _GEN_23338;
  wire  _GEN_23339;
  wire  _GEN_23340;
  wire  _GEN_23341;
  wire  _GEN_23342;
  wire  _GEN_23343;
  wire  _T_5113;
  wire  _T_5114;
  wire  _T_5116;
  wire  _T_5118;
  wire  _T_5120;
  wire [5:0] _T_5127;
  wire  _T_5130;
  wire  _T_5131;
  wire  _T_5133;
  wire  _T_5135;
  wire  _T_5137;
  wire  _GEN_209_ldst_val;
  wire [6:0] _GEN_23396;
  wire  _GEN_23421;
  wire [6:0] _GEN_23486;
  wire  _GEN_23511;
  wire [6:0] _GEN_23576;
  wire  _GEN_23601;
  wire [6:0] _GEN_23666;
  wire  _GEN_23691;
  wire [6:0] _GEN_23756;
  wire  _GEN_23781;
  wire [6:0] _GEN_23846;
  wire  _GEN_23871;
  wire [6:0] _GEN_23936;
  wire  _GEN_23961;
  wire [6:0] _GEN_24026;
  wire  _GEN_24051;
  wire [6:0] _GEN_24116;
  wire  _GEN_24141;
  wire [6:0] _GEN_24206;
  wire  _GEN_24231;
  wire [6:0] _GEN_24296;
  wire  _GEN_24321;
  wire [6:0] _GEN_24386;
  wire  _GEN_24411;
  wire [6:0] _GEN_24476;
  wire  _GEN_24501;
  wire [6:0] _GEN_24566;
  wire  _GEN_24591;
  wire [6:0] _GEN_24656;
  wire  _GEN_24681;
  wire [6:0] _GEN_24746;
  wire  _GEN_24771;
  wire [6:0] _GEN_24836;
  wire  _GEN_24861;
  wire [6:0] _GEN_24926;
  wire  _GEN_24951;
  wire [6:0] _GEN_25016;
  wire  _GEN_25041;
  wire [6:0] _GEN_25106;
  wire  _GEN_25131;
  wire [6:0] _GEN_25196;
  wire  _GEN_25221;
  wire [6:0] _GEN_25286;
  wire  _GEN_25311;
  wire [6:0] _GEN_25376;
  wire  _GEN_25401;
  wire [6:0] _GEN_25466;
  wire  _GEN_25491;
  wire [6:0] _GEN_25556;
  wire  _GEN_25581;
  wire [6:0] _GEN_25646;
  wire  _GEN_25671;
  wire [6:0] _GEN_25736;
  wire  _GEN_25761;
  wire [6:0] _GEN_25826;
  wire  _GEN_25851;
  wire [6:0] _GEN_25916;
  wire  _GEN_25941;
  wire [6:0] _GEN_26006;
  wire  _GEN_26031;
  wire [6:0] _GEN_26096;
  wire  _GEN_26121;
  wire [6:0] _GEN_26186;
  wire  _GEN_26211;
  wire [6:0] _GEN_26276;
  wire  _GEN_26301;
  wire [6:0] _GEN_26366;
  wire  _GEN_26391;
  wire [6:0] _GEN_26456;
  wire  _GEN_26481;
  wire [6:0] _GEN_26546;
  wire  _GEN_26571;
  wire [6:0] _GEN_26636;
  wire  _GEN_26661;
  wire [6:0] _GEN_26726;
  wire  _GEN_26751;
  wire [6:0] _GEN_26816;
  wire  _GEN_26841;
  wire  _T_5142;
  wire [6:0] _GEN_210_pdst;
  wire  _T_5143;
  wire  _T_5144;
  wire  _T_5146;
  wire  _T_5148;
  wire  _T_5150;
  wire  _GEN_212;
  wire  _GEN_26934;
  wire  _GEN_26935;
  wire  _GEN_26936;
  wire  _GEN_26937;
  wire  _GEN_26938;
  wire  _GEN_26939;
  wire  _GEN_26940;
  wire  _GEN_26941;
  wire  _GEN_26942;
  wire  _GEN_26943;
  wire  _GEN_26944;
  wire  _GEN_26945;
  wire  _GEN_26946;
  wire  _GEN_26947;
  wire  _GEN_26948;
  wire  _GEN_26949;
  wire  _GEN_26950;
  wire  _GEN_26951;
  wire  _GEN_26952;
  wire  _GEN_26953;
  wire  _GEN_26954;
  wire  _GEN_26955;
  wire  _GEN_26956;
  wire  _GEN_26957;
  wire  _GEN_26958;
  wire  _GEN_26959;
  wire  _GEN_26960;
  wire  _GEN_26961;
  wire  _GEN_26962;
  wire  _GEN_26963;
  wire  _GEN_26964;
  wire  _GEN_26965;
  wire  _GEN_26966;
  wire  _GEN_26967;
  wire  _GEN_26968;
  wire  _GEN_26969;
  wire  _GEN_26970;
  wire  _GEN_26971;
  wire  _GEN_26972;
  wire  _T_5190;
  wire  _T_5191;
  wire  _T_5193;
  wire  _T_5195;
  wire  _T_5197;
  wire [5:0] _T_5204;
  wire  _T_5207;
  wire  _T_5208;
  wire  _T_5210;
  wire  _T_5212;
  wire  _T_5214;
  wire  _GEN_213_ldst_val;
  wire [6:0] _GEN_27025;
  wire  _GEN_27050;
  wire [6:0] _GEN_27115;
  wire  _GEN_27140;
  wire [6:0] _GEN_27205;
  wire  _GEN_27230;
  wire [6:0] _GEN_27295;
  wire  _GEN_27320;
  wire [6:0] _GEN_27385;
  wire  _GEN_27410;
  wire [6:0] _GEN_27475;
  wire  _GEN_27500;
  wire [6:0] _GEN_27565;
  wire  _GEN_27590;
  wire [6:0] _GEN_27655;
  wire  _GEN_27680;
  wire [6:0] _GEN_27745;
  wire  _GEN_27770;
  wire [6:0] _GEN_27835;
  wire  _GEN_27860;
  wire [6:0] _GEN_27925;
  wire  _GEN_27950;
  wire [6:0] _GEN_28015;
  wire  _GEN_28040;
  wire [6:0] _GEN_28105;
  wire  _GEN_28130;
  wire [6:0] _GEN_28195;
  wire  _GEN_28220;
  wire [6:0] _GEN_28285;
  wire  _GEN_28310;
  wire [6:0] _GEN_28375;
  wire  _GEN_28400;
  wire [6:0] _GEN_28465;
  wire  _GEN_28490;
  wire [6:0] _GEN_28555;
  wire  _GEN_28580;
  wire [6:0] _GEN_28645;
  wire  _GEN_28670;
  wire [6:0] _GEN_28735;
  wire  _GEN_28760;
  wire [6:0] _GEN_28825;
  wire  _GEN_28850;
  wire [6:0] _GEN_28915;
  wire  _GEN_28940;
  wire [6:0] _GEN_29005;
  wire  _GEN_29030;
  wire [6:0] _GEN_29095;
  wire  _GEN_29120;
  wire [6:0] _GEN_29185;
  wire  _GEN_29210;
  wire [6:0] _GEN_29275;
  wire  _GEN_29300;
  wire [6:0] _GEN_29365;
  wire  _GEN_29390;
  wire [6:0] _GEN_29455;
  wire  _GEN_29480;
  wire [6:0] _GEN_29545;
  wire  _GEN_29570;
  wire [6:0] _GEN_29635;
  wire  _GEN_29660;
  wire [6:0] _GEN_29725;
  wire  _GEN_29750;
  wire [6:0] _GEN_29815;
  wire  _GEN_29840;
  wire [6:0] _GEN_29905;
  wire  _GEN_29930;
  wire [6:0] _GEN_29995;
  wire  _GEN_30020;
  wire [6:0] _GEN_30085;
  wire  _GEN_30110;
  wire [6:0] _GEN_30175;
  wire  _GEN_30200;
  wire [6:0] _GEN_30265;
  wire  _GEN_30290;
  wire [6:0] _GEN_30355;
  wire  _GEN_30380;
  wire [6:0] _GEN_30445;
  wire  _GEN_30470;
  wire  _T_5219;
  wire [6:0] _GEN_214_pdst;
  wire  _T_5220;
  wire  _T_5221;
  wire  _T_5223;
  wire  _T_5225;
  wire  _T_5227;
  wire  _GEN_216;
  wire  _GEN_30563;
  wire  _GEN_30564;
  wire  _GEN_30565;
  wire  _GEN_30566;
  wire  _GEN_30567;
  wire  _GEN_30568;
  wire  _GEN_30569;
  wire  _GEN_30570;
  wire  _GEN_30571;
  wire  _GEN_30572;
  wire  _GEN_30573;
  wire  _GEN_30574;
  wire  _GEN_30575;
  wire  _GEN_30576;
  wire  _GEN_30577;
  wire  _GEN_30578;
  wire  _GEN_30579;
  wire  _GEN_30580;
  wire  _GEN_30581;
  wire  _GEN_30582;
  wire  _GEN_30583;
  wire  _GEN_30584;
  wire  _GEN_30585;
  wire  _GEN_30586;
  wire  _GEN_30587;
  wire  _GEN_30588;
  wire  _GEN_30589;
  wire  _GEN_30590;
  wire  _GEN_30591;
  wire  _GEN_30592;
  wire  _GEN_30593;
  wire  _GEN_30594;
  wire  _GEN_30595;
  wire  _GEN_30596;
  wire  _GEN_30597;
  wire  _GEN_30598;
  wire  _GEN_30599;
  wire  _GEN_30600;
  wire  _GEN_30601;
  wire  _T_5267;
  wire  _T_5268;
  wire  _T_5270;
  wire  _T_5272;
  wire  _T_5274;
  wire [5:0] _T_5281;
  wire  _T_5284;
  wire  _T_5285;
  wire  _T_5287;
  wire  _T_5289;
  wire  _T_5291;
  wire  _GEN_217_ldst_val;
  wire [6:0] _GEN_30654;
  wire  _GEN_30679;
  wire [6:0] _GEN_30744;
  wire  _GEN_30769;
  wire [6:0] _GEN_30834;
  wire  _GEN_30859;
  wire [6:0] _GEN_30924;
  wire  _GEN_30949;
  wire [6:0] _GEN_31014;
  wire  _GEN_31039;
  wire [6:0] _GEN_31104;
  wire  _GEN_31129;
  wire [6:0] _GEN_31194;
  wire  _GEN_31219;
  wire [6:0] _GEN_31284;
  wire  _GEN_31309;
  wire [6:0] _GEN_31374;
  wire  _GEN_31399;
  wire [6:0] _GEN_31464;
  wire  _GEN_31489;
  wire [6:0] _GEN_31554;
  wire  _GEN_31579;
  wire [6:0] _GEN_31644;
  wire  _GEN_31669;
  wire [6:0] _GEN_31734;
  wire  _GEN_31759;
  wire [6:0] _GEN_31824;
  wire  _GEN_31849;
  wire [6:0] _GEN_31914;
  wire  _GEN_31939;
  wire [6:0] _GEN_32004;
  wire  _GEN_32029;
  wire [6:0] _GEN_32094;
  wire  _GEN_32119;
  wire [6:0] _GEN_32184;
  wire  _GEN_32209;
  wire [6:0] _GEN_32274;
  wire  _GEN_32299;
  wire [6:0] _GEN_32364;
  wire  _GEN_32389;
  wire [6:0] _GEN_32454;
  wire  _GEN_32479;
  wire [6:0] _GEN_32544;
  wire  _GEN_32569;
  wire [6:0] _GEN_32634;
  wire  _GEN_32659;
  wire [6:0] _GEN_32724;
  wire  _GEN_32749;
  wire [6:0] _GEN_32814;
  wire  _GEN_32839;
  wire [6:0] _GEN_32904;
  wire  _GEN_32929;
  wire [6:0] _GEN_32994;
  wire  _GEN_33019;
  wire [6:0] _GEN_33084;
  wire  _GEN_33109;
  wire [6:0] _GEN_33174;
  wire  _GEN_33199;
  wire [6:0] _GEN_33264;
  wire  _GEN_33289;
  wire [6:0] _GEN_33354;
  wire  _GEN_33379;
  wire [6:0] _GEN_33444;
  wire  _GEN_33469;
  wire [6:0] _GEN_33534;
  wire  _GEN_33559;
  wire [6:0] _GEN_33624;
  wire  _GEN_33649;
  wire [6:0] _GEN_33714;
  wire  _GEN_33739;
  wire [6:0] _GEN_33804;
  wire  _GEN_33829;
  wire [6:0] _GEN_33894;
  wire  _GEN_33919;
  wire [6:0] _GEN_33984;
  wire  _GEN_34009;
  wire [6:0] _GEN_34074;
  wire  _GEN_34099;
  wire  _T_5296;
  wire [6:0] _GEN_218_pdst;
  wire  _T_5297;
  wire  _T_5298;
  wire  _T_5300;
  wire  _T_5302;
  wire  _T_5304;
  wire  _GEN_220;
  wire  _GEN_34192;
  wire  _GEN_34193;
  wire  _GEN_34194;
  wire  _GEN_34195;
  wire  _GEN_34196;
  wire  _GEN_34197;
  wire  _GEN_34198;
  wire  _GEN_34199;
  wire  _GEN_34200;
  wire  _GEN_34201;
  wire  _GEN_34202;
  wire  _GEN_34203;
  wire  _GEN_34204;
  wire  _GEN_34205;
  wire  _GEN_34206;
  wire  _GEN_34207;
  wire  _GEN_34208;
  wire  _GEN_34209;
  wire  _GEN_34210;
  wire  _GEN_34211;
  wire  _GEN_34212;
  wire  _GEN_34213;
  wire  _GEN_34214;
  wire  _GEN_34215;
  wire  _GEN_34216;
  wire  _GEN_34217;
  wire  _GEN_34218;
  wire  _GEN_34219;
  wire  _GEN_34220;
  wire  _GEN_34221;
  wire  _GEN_34222;
  wire  _GEN_34223;
  wire  _GEN_34224;
  wire  _GEN_34225;
  wire  _GEN_34226;
  wire  _GEN_34227;
  wire  _GEN_34228;
  wire  _GEN_34229;
  wire  _GEN_34230;
  wire  _T_5344;
  wire  _T_5345;
  wire  _T_5347;
  wire  _T_5349;
  wire  _T_5351;
  wire [5:0] _T_5358;
  wire  _T_5361;
  wire  _T_5362;
  wire  _T_5364;
  wire  _T_5366;
  wire  _T_5368;
  wire  _GEN_221_ldst_val;
  wire [6:0] _GEN_34283;
  wire  _GEN_34308;
  wire [6:0] _GEN_34373;
  wire  _GEN_34398;
  wire [6:0] _GEN_34463;
  wire  _GEN_34488;
  wire [6:0] _GEN_34553;
  wire  _GEN_34578;
  wire [6:0] _GEN_34643;
  wire  _GEN_34668;
  wire [6:0] _GEN_34733;
  wire  _GEN_34758;
  wire [6:0] _GEN_34823;
  wire  _GEN_34848;
  wire [6:0] _GEN_34913;
  wire  _GEN_34938;
  wire [6:0] _GEN_35003;
  wire  _GEN_35028;
  wire [6:0] _GEN_35093;
  wire  _GEN_35118;
  wire [6:0] _GEN_35183;
  wire  _GEN_35208;
  wire [6:0] _GEN_35273;
  wire  _GEN_35298;
  wire [6:0] _GEN_35363;
  wire  _GEN_35388;
  wire [6:0] _GEN_35453;
  wire  _GEN_35478;
  wire [6:0] _GEN_35543;
  wire  _GEN_35568;
  wire [6:0] _GEN_35633;
  wire  _GEN_35658;
  wire [6:0] _GEN_35723;
  wire  _GEN_35748;
  wire [6:0] _GEN_35813;
  wire  _GEN_35838;
  wire [6:0] _GEN_35903;
  wire  _GEN_35928;
  wire [6:0] _GEN_35993;
  wire  _GEN_36018;
  wire [6:0] _GEN_36083;
  wire  _GEN_36108;
  wire [6:0] _GEN_36173;
  wire  _GEN_36198;
  wire [6:0] _GEN_36263;
  wire  _GEN_36288;
  wire [6:0] _GEN_36353;
  wire  _GEN_36378;
  wire [6:0] _GEN_36443;
  wire  _GEN_36468;
  wire [6:0] _GEN_36533;
  wire  _GEN_36558;
  wire [6:0] _GEN_36623;
  wire  _GEN_36648;
  wire [6:0] _GEN_36713;
  wire  _GEN_36738;
  wire [6:0] _GEN_36803;
  wire  _GEN_36828;
  wire [6:0] _GEN_36893;
  wire  _GEN_36918;
  wire [6:0] _GEN_36983;
  wire  _GEN_37008;
  wire [6:0] _GEN_37073;
  wire  _GEN_37098;
  wire [6:0] _GEN_37163;
  wire  _GEN_37188;
  wire [6:0] _GEN_37253;
  wire  _GEN_37278;
  wire [6:0] _GEN_37343;
  wire  _GEN_37368;
  wire [6:0] _GEN_37433;
  wire  _GEN_37458;
  wire [6:0] _GEN_37523;
  wire  _GEN_37548;
  wire [6:0] _GEN_37613;
  wire  _GEN_37638;
  wire [6:0] _GEN_37703;
  wire  _GEN_37728;
  wire  _T_5373;
  wire [6:0] _GEN_222_pdst;
  wire  _T_5374;
  wire  _T_5375;
  wire  _T_5377;
  wire  _T_5379;
  wire  _T_5381;
  wire  _GEN_224;
  wire  _GEN_37821;
  wire  _GEN_37822;
  wire  _GEN_37823;
  wire  _GEN_37824;
  wire  _GEN_37825;
  wire  _GEN_37826;
  wire  _GEN_37827;
  wire  _GEN_37828;
  wire  _GEN_37829;
  wire  _GEN_37830;
  wire  _GEN_37831;
  wire  _GEN_37832;
  wire  _GEN_37833;
  wire  _GEN_37834;
  wire  _GEN_37835;
  wire  _GEN_37836;
  wire  _GEN_37837;
  wire  _GEN_37838;
  wire  _GEN_37839;
  wire  _GEN_37840;
  wire  _GEN_37841;
  wire  _GEN_37842;
  wire  _GEN_37843;
  wire  _GEN_37844;
  wire  _GEN_37845;
  wire  _GEN_37846;
  wire  _GEN_37847;
  wire  _GEN_37848;
  wire  _GEN_37849;
  wire  _GEN_37850;
  wire  _GEN_37851;
  wire  _GEN_37852;
  wire  _GEN_37853;
  wire  _GEN_37854;
  wire  _GEN_37855;
  wire  _GEN_37856;
  wire  _GEN_37857;
  wire  _GEN_37858;
  wire  _GEN_37859;
  wire  _T_5421;
  wire  _T_5422;
  wire  _T_5424;
  wire  _T_5426;
  wire  _T_5428;
  wire [5:0] _T_5435;
  wire  _T_5438;
  wire  _T_5439;
  wire  _T_5441;
  wire  _T_5443;
  wire  _T_5445;
  wire  _GEN_225_ldst_val;
  wire [6:0] _GEN_37912;
  wire  _GEN_37937;
  wire [6:0] _GEN_38002;
  wire  _GEN_38027;
  wire [6:0] _GEN_38092;
  wire  _GEN_38117;
  wire [6:0] _GEN_38182;
  wire  _GEN_38207;
  wire [6:0] _GEN_38272;
  wire  _GEN_38297;
  wire [6:0] _GEN_38362;
  wire  _GEN_38387;
  wire [6:0] _GEN_38452;
  wire  _GEN_38477;
  wire [6:0] _GEN_38542;
  wire  _GEN_38567;
  wire [6:0] _GEN_38632;
  wire  _GEN_38657;
  wire [6:0] _GEN_38722;
  wire  _GEN_38747;
  wire [6:0] _GEN_38812;
  wire  _GEN_38837;
  wire [6:0] _GEN_38902;
  wire  _GEN_38927;
  wire [6:0] _GEN_38992;
  wire  _GEN_39017;
  wire [6:0] _GEN_39082;
  wire  _GEN_39107;
  wire [6:0] _GEN_39172;
  wire  _GEN_39197;
  wire [6:0] _GEN_39262;
  wire  _GEN_39287;
  wire [6:0] _GEN_39352;
  wire  _GEN_39377;
  wire [6:0] _GEN_39442;
  wire  _GEN_39467;
  wire [6:0] _GEN_39532;
  wire  _GEN_39557;
  wire [6:0] _GEN_39622;
  wire  _GEN_39647;
  wire [6:0] _GEN_39712;
  wire  _GEN_39737;
  wire [6:0] _GEN_39802;
  wire  _GEN_39827;
  wire [6:0] _GEN_39892;
  wire  _GEN_39917;
  wire [6:0] _GEN_39982;
  wire  _GEN_40007;
  wire [6:0] _GEN_40072;
  wire  _GEN_40097;
  wire [6:0] _GEN_40162;
  wire  _GEN_40187;
  wire [6:0] _GEN_40252;
  wire  _GEN_40277;
  wire [6:0] _GEN_40342;
  wire  _GEN_40367;
  wire [6:0] _GEN_40432;
  wire  _GEN_40457;
  wire [6:0] _GEN_40522;
  wire  _GEN_40547;
  wire [6:0] _GEN_40612;
  wire  _GEN_40637;
  wire [6:0] _GEN_40702;
  wire  _GEN_40727;
  wire [6:0] _GEN_40792;
  wire  _GEN_40817;
  wire [6:0] _GEN_40882;
  wire  _GEN_40907;
  wire [6:0] _GEN_40972;
  wire  _GEN_40997;
  wire [6:0] _GEN_41062;
  wire  _GEN_41087;
  wire [6:0] _GEN_41152;
  wire  _GEN_41177;
  wire [6:0] _GEN_41242;
  wire  _GEN_41267;
  wire [6:0] _GEN_41332;
  wire  _GEN_41357;
  wire  _T_5450;
  wire [6:0] _GEN_226_pdst;
  wire  _T_5451;
  wire  _T_5452;
  wire  _T_5454;
  wire  _T_5456;
  wire  _T_5458;
  reg  _T_5637_0;
  reg [31:0] _RAND_553;
  reg  _T_5637_1;
  reg [31:0] _RAND_554;
  reg  _T_5637_2;
  reg [31:0] _RAND_555;
  reg  _T_5637_3;
  reg [31:0] _RAND_556;
  reg  _T_5637_4;
  reg [31:0] _RAND_557;
  reg  _T_5637_5;
  reg [31:0] _RAND_558;
  reg  _T_5637_6;
  reg [31:0] _RAND_559;
  reg  _T_5637_7;
  reg [31:0] _RAND_560;
  reg  _T_5637_8;
  reg [31:0] _RAND_561;
  reg  _T_5637_9;
  reg [31:0] _RAND_562;
  reg  _T_5637_10;
  reg [31:0] _RAND_563;
  reg  _T_5637_11;
  reg [31:0] _RAND_564;
  reg  _T_5637_12;
  reg [31:0] _RAND_565;
  reg  _T_5637_13;
  reg [31:0] _RAND_566;
  reg  _T_5637_14;
  reg [31:0] _RAND_567;
  reg  _T_5637_15;
  reg [31:0] _RAND_568;
  reg  _T_5637_16;
  reg [31:0] _RAND_569;
  reg  _T_5637_17;
  reg [31:0] _RAND_570;
  reg  _T_5637_18;
  reg [31:0] _RAND_571;
  reg  _T_5637_19;
  reg [31:0] _RAND_572;
  reg  _T_5637_20;
  reg [31:0] _RAND_573;
  reg  _T_5637_21;
  reg [31:0] _RAND_574;
  reg  _T_5637_22;
  reg [31:0] _RAND_575;
  reg  _T_5637_23;
  reg [31:0] _RAND_576;
  reg  _T_5637_24;
  reg [31:0] _RAND_577;
  reg  _T_5637_25;
  reg [31:0] _RAND_578;
  reg  _T_5637_26;
  reg [31:0] _RAND_579;
  reg  _T_5637_27;
  reg [31:0] _RAND_580;
  reg  _T_5637_28;
  reg [31:0] _RAND_581;
  reg  _T_5637_29;
  reg [31:0] _RAND_582;
  reg  _T_5637_30;
  reg [31:0] _RAND_583;
  reg  _T_5637_31;
  reg [31:0] _RAND_584;
  reg  _T_5637_32;
  reg [31:0] _RAND_585;
  reg  _T_5637_33;
  reg [31:0] _RAND_586;
  reg  _T_5637_34;
  reg [31:0] _RAND_587;
  reg  _T_5637_35;
  reg [31:0] _RAND_588;
  reg  _T_5637_36;
  reg [31:0] _RAND_589;
  reg  _T_5637_37;
  reg [31:0] _RAND_590;
  reg  _T_5637_38;
  reg [31:0] _RAND_591;
  reg  _T_5637_39;
  reg [31:0] _RAND_592;
  reg  _T_5764 [0:39];
  reg [31:0] _RAND_593;
  wire  _T_5764__T_6441_data;
  wire [5:0] _T_5764__T_6441_addr;
  reg [31:0] _RAND_594;
  wire  _T_5764__T_6468_data;
  wire [5:0] _T_5764__T_6468_addr;
  reg [31:0] _RAND_595;
  wire  _T_5764__T_6581_data;
  wire [5:0] _T_5764__T_6581_addr;
  reg [31:0] _RAND_596;
  wire  _T_5764__T_7692_data;
  wire [5:0] _T_5764__T_7692_addr;
  reg [31:0] _RAND_597;
  wire  _T_5764__T_7769_data;
  wire [5:0] _T_5764__T_7769_addr;
  reg [31:0] _RAND_598;
  wire  _T_5764__T_7846_data;
  wire [5:0] _T_5764__T_7846_addr;
  reg [31:0] _RAND_599;
  wire  _T_5764__T_7923_data;
  wire [5:0] _T_5764__T_7923_addr;
  reg [31:0] _RAND_600;
  wire  _T_5764__T_8000_data;
  wire [5:0] _T_5764__T_8000_addr;
  reg [31:0] _RAND_601;
  wire  _T_5764__T_6317_data;
  wire [5:0] _T_5764__T_6317_addr;
  wire  _T_5764__T_6317_mask;
  wire  _T_5764__T_6317_en;
  wire  _T_5764__T_6383_data;
  wire [5:0] _T_5764__T_6383_addr;
  wire  _T_5764__T_6383_mask;
  wire  _T_5764__T_6383_en;
  wire  _T_5764__T_6392_data;
  wire [5:0] _T_5764__T_6392_addr;
  wire  _T_5764__T_6392_mask;
  wire  _T_5764__T_6392_en;
  wire  _T_5764__T_6401_data;
  wire [5:0] _T_5764__T_6401_addr;
  wire  _T_5764__T_6401_mask;
  wire  _T_5764__T_6401_en;
  wire  _T_5764__T_6410_data;
  wire [5:0] _T_5764__T_6410_addr;
  wire  _T_5764__T_6410_mask;
  wire  _T_5764__T_6410_en;
  wire  _T_5764__T_6419_data;
  wire [5:0] _T_5764__T_6419_addr;
  wire  _T_5764__T_6419_mask;
  wire  _T_5764__T_6419_en;
  wire  _T_5764__T_6428_data;
  wire [5:0] _T_5764__T_6428_addr;
  wire  _T_5764__T_6428_mask;
  wire  _T_5764__T_6428_en;
  wire  _T_5764__T_6455_data;
  wire [5:0] _T_5764__T_6455_addr;
  wire  _T_5764__T_6455_mask;
  wire  _T_5764__T_6455_en;
  reg [7:0] _T_5936_0_br_mask;
  reg [31:0] _RAND_602;
  reg [6:0] _T_5936_0_pdst;
  reg [31:0] _RAND_603;
  reg [6:0] _T_5936_0_stale_pdst;
  reg [31:0] _RAND_604;
  reg  _T_5936_0_is_fencei;
  reg [31:0] _RAND_605;
  reg  _T_5936_0_is_store;
  reg [31:0] _RAND_606;
  reg  _T_5936_0_is_load;
  reg [31:0] _RAND_607;
  reg  _T_5936_0_is_sys_pc2epc;
  reg [31:0] _RAND_608;
  reg  _T_5936_0_flush_on_commit;
  reg [31:0] _RAND_609;
  reg [5:0] _T_5936_0_ldst;
  reg [31:0] _RAND_610;
  reg  _T_5936_0_ldst_val;
  reg [31:0] _RAND_611;
  reg [1:0] _T_5936_0_dst_rtype;
  reg [31:0] _RAND_612;
  reg  _T_5936_0_fp_val;
  reg [31:0] _RAND_613;
  reg [7:0] _T_5936_1_br_mask;
  reg [31:0] _RAND_614;
  reg [6:0] _T_5936_1_pdst;
  reg [31:0] _RAND_615;
  reg [6:0] _T_5936_1_stale_pdst;
  reg [31:0] _RAND_616;
  reg  _T_5936_1_is_fencei;
  reg [31:0] _RAND_617;
  reg  _T_5936_1_is_store;
  reg [31:0] _RAND_618;
  reg  _T_5936_1_is_load;
  reg [31:0] _RAND_619;
  reg  _T_5936_1_is_sys_pc2epc;
  reg [31:0] _RAND_620;
  reg  _T_5936_1_flush_on_commit;
  reg [31:0] _RAND_621;
  reg [5:0] _T_5936_1_ldst;
  reg [31:0] _RAND_622;
  reg  _T_5936_1_ldst_val;
  reg [31:0] _RAND_623;
  reg [1:0] _T_5936_1_dst_rtype;
  reg [31:0] _RAND_624;
  reg  _T_5936_1_fp_val;
  reg [31:0] _RAND_625;
  reg [7:0] _T_5936_2_br_mask;
  reg [31:0] _RAND_626;
  reg [6:0] _T_5936_2_pdst;
  reg [31:0] _RAND_627;
  reg [6:0] _T_5936_2_stale_pdst;
  reg [31:0] _RAND_628;
  reg  _T_5936_2_is_fencei;
  reg [31:0] _RAND_629;
  reg  _T_5936_2_is_store;
  reg [31:0] _RAND_630;
  reg  _T_5936_2_is_load;
  reg [31:0] _RAND_631;
  reg  _T_5936_2_is_sys_pc2epc;
  reg [31:0] _RAND_632;
  reg  _T_5936_2_flush_on_commit;
  reg [31:0] _RAND_633;
  reg [5:0] _T_5936_2_ldst;
  reg [31:0] _RAND_634;
  reg  _T_5936_2_ldst_val;
  reg [31:0] _RAND_635;
  reg [1:0] _T_5936_2_dst_rtype;
  reg [31:0] _RAND_636;
  reg  _T_5936_2_fp_val;
  reg [31:0] _RAND_637;
  reg [7:0] _T_5936_3_br_mask;
  reg [31:0] _RAND_638;
  reg [6:0] _T_5936_3_pdst;
  reg [31:0] _RAND_639;
  reg [6:0] _T_5936_3_stale_pdst;
  reg [31:0] _RAND_640;
  reg  _T_5936_3_is_fencei;
  reg [31:0] _RAND_641;
  reg  _T_5936_3_is_store;
  reg [31:0] _RAND_642;
  reg  _T_5936_3_is_load;
  reg [31:0] _RAND_643;
  reg  _T_5936_3_is_sys_pc2epc;
  reg [31:0] _RAND_644;
  reg  _T_5936_3_flush_on_commit;
  reg [31:0] _RAND_645;
  reg [5:0] _T_5936_3_ldst;
  reg [31:0] _RAND_646;
  reg  _T_5936_3_ldst_val;
  reg [31:0] _RAND_647;
  reg [1:0] _T_5936_3_dst_rtype;
  reg [31:0] _RAND_648;
  reg  _T_5936_3_fp_val;
  reg [31:0] _RAND_649;
  reg [7:0] _T_5936_4_br_mask;
  reg [31:0] _RAND_650;
  reg [6:0] _T_5936_4_pdst;
  reg [31:0] _RAND_651;
  reg [6:0] _T_5936_4_stale_pdst;
  reg [31:0] _RAND_652;
  reg  _T_5936_4_is_fencei;
  reg [31:0] _RAND_653;
  reg  _T_5936_4_is_store;
  reg [31:0] _RAND_654;
  reg  _T_5936_4_is_load;
  reg [31:0] _RAND_655;
  reg  _T_5936_4_is_sys_pc2epc;
  reg [31:0] _RAND_656;
  reg  _T_5936_4_flush_on_commit;
  reg [31:0] _RAND_657;
  reg [5:0] _T_5936_4_ldst;
  reg [31:0] _RAND_658;
  reg  _T_5936_4_ldst_val;
  reg [31:0] _RAND_659;
  reg [1:0] _T_5936_4_dst_rtype;
  reg [31:0] _RAND_660;
  reg  _T_5936_4_fp_val;
  reg [31:0] _RAND_661;
  reg [7:0] _T_5936_5_br_mask;
  reg [31:0] _RAND_662;
  reg [6:0] _T_5936_5_pdst;
  reg [31:0] _RAND_663;
  reg [6:0] _T_5936_5_stale_pdst;
  reg [31:0] _RAND_664;
  reg  _T_5936_5_is_fencei;
  reg [31:0] _RAND_665;
  reg  _T_5936_5_is_store;
  reg [31:0] _RAND_666;
  reg  _T_5936_5_is_load;
  reg [31:0] _RAND_667;
  reg  _T_5936_5_is_sys_pc2epc;
  reg [31:0] _RAND_668;
  reg  _T_5936_5_flush_on_commit;
  reg [31:0] _RAND_669;
  reg [5:0] _T_5936_5_ldst;
  reg [31:0] _RAND_670;
  reg  _T_5936_5_ldst_val;
  reg [31:0] _RAND_671;
  reg [1:0] _T_5936_5_dst_rtype;
  reg [31:0] _RAND_672;
  reg  _T_5936_5_fp_val;
  reg [31:0] _RAND_673;
  reg [7:0] _T_5936_6_br_mask;
  reg [31:0] _RAND_674;
  reg [6:0] _T_5936_6_pdst;
  reg [31:0] _RAND_675;
  reg [6:0] _T_5936_6_stale_pdst;
  reg [31:0] _RAND_676;
  reg  _T_5936_6_is_fencei;
  reg [31:0] _RAND_677;
  reg  _T_5936_6_is_store;
  reg [31:0] _RAND_678;
  reg  _T_5936_6_is_load;
  reg [31:0] _RAND_679;
  reg  _T_5936_6_is_sys_pc2epc;
  reg [31:0] _RAND_680;
  reg  _T_5936_6_flush_on_commit;
  reg [31:0] _RAND_681;
  reg [5:0] _T_5936_6_ldst;
  reg [31:0] _RAND_682;
  reg  _T_5936_6_ldst_val;
  reg [31:0] _RAND_683;
  reg [1:0] _T_5936_6_dst_rtype;
  reg [31:0] _RAND_684;
  reg  _T_5936_6_fp_val;
  reg [31:0] _RAND_685;
  reg [7:0] _T_5936_7_br_mask;
  reg [31:0] _RAND_686;
  reg [6:0] _T_5936_7_pdst;
  reg [31:0] _RAND_687;
  reg [6:0] _T_5936_7_stale_pdst;
  reg [31:0] _RAND_688;
  reg  _T_5936_7_is_fencei;
  reg [31:0] _RAND_689;
  reg  _T_5936_7_is_store;
  reg [31:0] _RAND_690;
  reg  _T_5936_7_is_load;
  reg [31:0] _RAND_691;
  reg  _T_5936_7_is_sys_pc2epc;
  reg [31:0] _RAND_692;
  reg  _T_5936_7_flush_on_commit;
  reg [31:0] _RAND_693;
  reg [5:0] _T_5936_7_ldst;
  reg [31:0] _RAND_694;
  reg  _T_5936_7_ldst_val;
  reg [31:0] _RAND_695;
  reg [1:0] _T_5936_7_dst_rtype;
  reg [31:0] _RAND_696;
  reg  _T_5936_7_fp_val;
  reg [31:0] _RAND_697;
  reg [7:0] _T_5936_8_br_mask;
  reg [31:0] _RAND_698;
  reg [6:0] _T_5936_8_pdst;
  reg [31:0] _RAND_699;
  reg [6:0] _T_5936_8_stale_pdst;
  reg [31:0] _RAND_700;
  reg  _T_5936_8_is_fencei;
  reg [31:0] _RAND_701;
  reg  _T_5936_8_is_store;
  reg [31:0] _RAND_702;
  reg  _T_5936_8_is_load;
  reg [31:0] _RAND_703;
  reg  _T_5936_8_is_sys_pc2epc;
  reg [31:0] _RAND_704;
  reg  _T_5936_8_flush_on_commit;
  reg [31:0] _RAND_705;
  reg [5:0] _T_5936_8_ldst;
  reg [31:0] _RAND_706;
  reg  _T_5936_8_ldst_val;
  reg [31:0] _RAND_707;
  reg [1:0] _T_5936_8_dst_rtype;
  reg [31:0] _RAND_708;
  reg  _T_5936_8_fp_val;
  reg [31:0] _RAND_709;
  reg [7:0] _T_5936_9_br_mask;
  reg [31:0] _RAND_710;
  reg [6:0] _T_5936_9_pdst;
  reg [31:0] _RAND_711;
  reg [6:0] _T_5936_9_stale_pdst;
  reg [31:0] _RAND_712;
  reg  _T_5936_9_is_fencei;
  reg [31:0] _RAND_713;
  reg  _T_5936_9_is_store;
  reg [31:0] _RAND_714;
  reg  _T_5936_9_is_load;
  reg [31:0] _RAND_715;
  reg  _T_5936_9_is_sys_pc2epc;
  reg [31:0] _RAND_716;
  reg  _T_5936_9_flush_on_commit;
  reg [31:0] _RAND_717;
  reg [5:0] _T_5936_9_ldst;
  reg [31:0] _RAND_718;
  reg  _T_5936_9_ldst_val;
  reg [31:0] _RAND_719;
  reg [1:0] _T_5936_9_dst_rtype;
  reg [31:0] _RAND_720;
  reg  _T_5936_9_fp_val;
  reg [31:0] _RAND_721;
  reg [7:0] _T_5936_10_br_mask;
  reg [31:0] _RAND_722;
  reg [6:0] _T_5936_10_pdst;
  reg [31:0] _RAND_723;
  reg [6:0] _T_5936_10_stale_pdst;
  reg [31:0] _RAND_724;
  reg  _T_5936_10_is_fencei;
  reg [31:0] _RAND_725;
  reg  _T_5936_10_is_store;
  reg [31:0] _RAND_726;
  reg  _T_5936_10_is_load;
  reg [31:0] _RAND_727;
  reg  _T_5936_10_is_sys_pc2epc;
  reg [31:0] _RAND_728;
  reg  _T_5936_10_flush_on_commit;
  reg [31:0] _RAND_729;
  reg [5:0] _T_5936_10_ldst;
  reg [31:0] _RAND_730;
  reg  _T_5936_10_ldst_val;
  reg [31:0] _RAND_731;
  reg [1:0] _T_5936_10_dst_rtype;
  reg [31:0] _RAND_732;
  reg  _T_5936_10_fp_val;
  reg [31:0] _RAND_733;
  reg [7:0] _T_5936_11_br_mask;
  reg [31:0] _RAND_734;
  reg [6:0] _T_5936_11_pdst;
  reg [31:0] _RAND_735;
  reg [6:0] _T_5936_11_stale_pdst;
  reg [31:0] _RAND_736;
  reg  _T_5936_11_is_fencei;
  reg [31:0] _RAND_737;
  reg  _T_5936_11_is_store;
  reg [31:0] _RAND_738;
  reg  _T_5936_11_is_load;
  reg [31:0] _RAND_739;
  reg  _T_5936_11_is_sys_pc2epc;
  reg [31:0] _RAND_740;
  reg  _T_5936_11_flush_on_commit;
  reg [31:0] _RAND_741;
  reg [5:0] _T_5936_11_ldst;
  reg [31:0] _RAND_742;
  reg  _T_5936_11_ldst_val;
  reg [31:0] _RAND_743;
  reg [1:0] _T_5936_11_dst_rtype;
  reg [31:0] _RAND_744;
  reg  _T_5936_11_fp_val;
  reg [31:0] _RAND_745;
  reg [7:0] _T_5936_12_br_mask;
  reg [31:0] _RAND_746;
  reg [6:0] _T_5936_12_pdst;
  reg [31:0] _RAND_747;
  reg [6:0] _T_5936_12_stale_pdst;
  reg [31:0] _RAND_748;
  reg  _T_5936_12_is_fencei;
  reg [31:0] _RAND_749;
  reg  _T_5936_12_is_store;
  reg [31:0] _RAND_750;
  reg  _T_5936_12_is_load;
  reg [31:0] _RAND_751;
  reg  _T_5936_12_is_sys_pc2epc;
  reg [31:0] _RAND_752;
  reg  _T_5936_12_flush_on_commit;
  reg [31:0] _RAND_753;
  reg [5:0] _T_5936_12_ldst;
  reg [31:0] _RAND_754;
  reg  _T_5936_12_ldst_val;
  reg [31:0] _RAND_755;
  reg [1:0] _T_5936_12_dst_rtype;
  reg [31:0] _RAND_756;
  reg  _T_5936_12_fp_val;
  reg [31:0] _RAND_757;
  reg [7:0] _T_5936_13_br_mask;
  reg [31:0] _RAND_758;
  reg [6:0] _T_5936_13_pdst;
  reg [31:0] _RAND_759;
  reg [6:0] _T_5936_13_stale_pdst;
  reg [31:0] _RAND_760;
  reg  _T_5936_13_is_fencei;
  reg [31:0] _RAND_761;
  reg  _T_5936_13_is_store;
  reg [31:0] _RAND_762;
  reg  _T_5936_13_is_load;
  reg [31:0] _RAND_763;
  reg  _T_5936_13_is_sys_pc2epc;
  reg [31:0] _RAND_764;
  reg  _T_5936_13_flush_on_commit;
  reg [31:0] _RAND_765;
  reg [5:0] _T_5936_13_ldst;
  reg [31:0] _RAND_766;
  reg  _T_5936_13_ldst_val;
  reg [31:0] _RAND_767;
  reg [1:0] _T_5936_13_dst_rtype;
  reg [31:0] _RAND_768;
  reg  _T_5936_13_fp_val;
  reg [31:0] _RAND_769;
  reg [7:0] _T_5936_14_br_mask;
  reg [31:0] _RAND_770;
  reg [6:0] _T_5936_14_pdst;
  reg [31:0] _RAND_771;
  reg [6:0] _T_5936_14_stale_pdst;
  reg [31:0] _RAND_772;
  reg  _T_5936_14_is_fencei;
  reg [31:0] _RAND_773;
  reg  _T_5936_14_is_store;
  reg [31:0] _RAND_774;
  reg  _T_5936_14_is_load;
  reg [31:0] _RAND_775;
  reg  _T_5936_14_is_sys_pc2epc;
  reg [31:0] _RAND_776;
  reg  _T_5936_14_flush_on_commit;
  reg [31:0] _RAND_777;
  reg [5:0] _T_5936_14_ldst;
  reg [31:0] _RAND_778;
  reg  _T_5936_14_ldst_val;
  reg [31:0] _RAND_779;
  reg [1:0] _T_5936_14_dst_rtype;
  reg [31:0] _RAND_780;
  reg  _T_5936_14_fp_val;
  reg [31:0] _RAND_781;
  reg [7:0] _T_5936_15_br_mask;
  reg [31:0] _RAND_782;
  reg [6:0] _T_5936_15_pdst;
  reg [31:0] _RAND_783;
  reg [6:0] _T_5936_15_stale_pdst;
  reg [31:0] _RAND_784;
  reg  _T_5936_15_is_fencei;
  reg [31:0] _RAND_785;
  reg  _T_5936_15_is_store;
  reg [31:0] _RAND_786;
  reg  _T_5936_15_is_load;
  reg [31:0] _RAND_787;
  reg  _T_5936_15_is_sys_pc2epc;
  reg [31:0] _RAND_788;
  reg  _T_5936_15_flush_on_commit;
  reg [31:0] _RAND_789;
  reg [5:0] _T_5936_15_ldst;
  reg [31:0] _RAND_790;
  reg  _T_5936_15_ldst_val;
  reg [31:0] _RAND_791;
  reg [1:0] _T_5936_15_dst_rtype;
  reg [31:0] _RAND_792;
  reg  _T_5936_15_fp_val;
  reg [31:0] _RAND_793;
  reg [7:0] _T_5936_16_br_mask;
  reg [31:0] _RAND_794;
  reg [6:0] _T_5936_16_pdst;
  reg [31:0] _RAND_795;
  reg [6:0] _T_5936_16_stale_pdst;
  reg [31:0] _RAND_796;
  reg  _T_5936_16_is_fencei;
  reg [31:0] _RAND_797;
  reg  _T_5936_16_is_store;
  reg [31:0] _RAND_798;
  reg  _T_5936_16_is_load;
  reg [31:0] _RAND_799;
  reg  _T_5936_16_is_sys_pc2epc;
  reg [31:0] _RAND_800;
  reg  _T_5936_16_flush_on_commit;
  reg [31:0] _RAND_801;
  reg [5:0] _T_5936_16_ldst;
  reg [31:0] _RAND_802;
  reg  _T_5936_16_ldst_val;
  reg [31:0] _RAND_803;
  reg [1:0] _T_5936_16_dst_rtype;
  reg [31:0] _RAND_804;
  reg  _T_5936_16_fp_val;
  reg [31:0] _RAND_805;
  reg [7:0] _T_5936_17_br_mask;
  reg [31:0] _RAND_806;
  reg [6:0] _T_5936_17_pdst;
  reg [31:0] _RAND_807;
  reg [6:0] _T_5936_17_stale_pdst;
  reg [31:0] _RAND_808;
  reg  _T_5936_17_is_fencei;
  reg [31:0] _RAND_809;
  reg  _T_5936_17_is_store;
  reg [31:0] _RAND_810;
  reg  _T_5936_17_is_load;
  reg [31:0] _RAND_811;
  reg  _T_5936_17_is_sys_pc2epc;
  reg [31:0] _RAND_812;
  reg  _T_5936_17_flush_on_commit;
  reg [31:0] _RAND_813;
  reg [5:0] _T_5936_17_ldst;
  reg [31:0] _RAND_814;
  reg  _T_5936_17_ldst_val;
  reg [31:0] _RAND_815;
  reg [1:0] _T_5936_17_dst_rtype;
  reg [31:0] _RAND_816;
  reg  _T_5936_17_fp_val;
  reg [31:0] _RAND_817;
  reg [7:0] _T_5936_18_br_mask;
  reg [31:0] _RAND_818;
  reg [6:0] _T_5936_18_pdst;
  reg [31:0] _RAND_819;
  reg [6:0] _T_5936_18_stale_pdst;
  reg [31:0] _RAND_820;
  reg  _T_5936_18_is_fencei;
  reg [31:0] _RAND_821;
  reg  _T_5936_18_is_store;
  reg [31:0] _RAND_822;
  reg  _T_5936_18_is_load;
  reg [31:0] _RAND_823;
  reg  _T_5936_18_is_sys_pc2epc;
  reg [31:0] _RAND_824;
  reg  _T_5936_18_flush_on_commit;
  reg [31:0] _RAND_825;
  reg [5:0] _T_5936_18_ldst;
  reg [31:0] _RAND_826;
  reg  _T_5936_18_ldst_val;
  reg [31:0] _RAND_827;
  reg [1:0] _T_5936_18_dst_rtype;
  reg [31:0] _RAND_828;
  reg  _T_5936_18_fp_val;
  reg [31:0] _RAND_829;
  reg [7:0] _T_5936_19_br_mask;
  reg [31:0] _RAND_830;
  reg [6:0] _T_5936_19_pdst;
  reg [31:0] _RAND_831;
  reg [6:0] _T_5936_19_stale_pdst;
  reg [31:0] _RAND_832;
  reg  _T_5936_19_is_fencei;
  reg [31:0] _RAND_833;
  reg  _T_5936_19_is_store;
  reg [31:0] _RAND_834;
  reg  _T_5936_19_is_load;
  reg [31:0] _RAND_835;
  reg  _T_5936_19_is_sys_pc2epc;
  reg [31:0] _RAND_836;
  reg  _T_5936_19_flush_on_commit;
  reg [31:0] _RAND_837;
  reg [5:0] _T_5936_19_ldst;
  reg [31:0] _RAND_838;
  reg  _T_5936_19_ldst_val;
  reg [31:0] _RAND_839;
  reg [1:0] _T_5936_19_dst_rtype;
  reg [31:0] _RAND_840;
  reg  _T_5936_19_fp_val;
  reg [31:0] _RAND_841;
  reg [7:0] _T_5936_20_br_mask;
  reg [31:0] _RAND_842;
  reg [6:0] _T_5936_20_pdst;
  reg [31:0] _RAND_843;
  reg [6:0] _T_5936_20_stale_pdst;
  reg [31:0] _RAND_844;
  reg  _T_5936_20_is_fencei;
  reg [31:0] _RAND_845;
  reg  _T_5936_20_is_store;
  reg [31:0] _RAND_846;
  reg  _T_5936_20_is_load;
  reg [31:0] _RAND_847;
  reg  _T_5936_20_is_sys_pc2epc;
  reg [31:0] _RAND_848;
  reg  _T_5936_20_flush_on_commit;
  reg [31:0] _RAND_849;
  reg [5:0] _T_5936_20_ldst;
  reg [31:0] _RAND_850;
  reg  _T_5936_20_ldst_val;
  reg [31:0] _RAND_851;
  reg [1:0] _T_5936_20_dst_rtype;
  reg [31:0] _RAND_852;
  reg  _T_5936_20_fp_val;
  reg [31:0] _RAND_853;
  reg [7:0] _T_5936_21_br_mask;
  reg [31:0] _RAND_854;
  reg [6:0] _T_5936_21_pdst;
  reg [31:0] _RAND_855;
  reg [6:0] _T_5936_21_stale_pdst;
  reg [31:0] _RAND_856;
  reg  _T_5936_21_is_fencei;
  reg [31:0] _RAND_857;
  reg  _T_5936_21_is_store;
  reg [31:0] _RAND_858;
  reg  _T_5936_21_is_load;
  reg [31:0] _RAND_859;
  reg  _T_5936_21_is_sys_pc2epc;
  reg [31:0] _RAND_860;
  reg  _T_5936_21_flush_on_commit;
  reg [31:0] _RAND_861;
  reg [5:0] _T_5936_21_ldst;
  reg [31:0] _RAND_862;
  reg  _T_5936_21_ldst_val;
  reg [31:0] _RAND_863;
  reg [1:0] _T_5936_21_dst_rtype;
  reg [31:0] _RAND_864;
  reg  _T_5936_21_fp_val;
  reg [31:0] _RAND_865;
  reg [7:0] _T_5936_22_br_mask;
  reg [31:0] _RAND_866;
  reg [6:0] _T_5936_22_pdst;
  reg [31:0] _RAND_867;
  reg [6:0] _T_5936_22_stale_pdst;
  reg [31:0] _RAND_868;
  reg  _T_5936_22_is_fencei;
  reg [31:0] _RAND_869;
  reg  _T_5936_22_is_store;
  reg [31:0] _RAND_870;
  reg  _T_5936_22_is_load;
  reg [31:0] _RAND_871;
  reg  _T_5936_22_is_sys_pc2epc;
  reg [31:0] _RAND_872;
  reg  _T_5936_22_flush_on_commit;
  reg [31:0] _RAND_873;
  reg [5:0] _T_5936_22_ldst;
  reg [31:0] _RAND_874;
  reg  _T_5936_22_ldst_val;
  reg [31:0] _RAND_875;
  reg [1:0] _T_5936_22_dst_rtype;
  reg [31:0] _RAND_876;
  reg  _T_5936_22_fp_val;
  reg [31:0] _RAND_877;
  reg [7:0] _T_5936_23_br_mask;
  reg [31:0] _RAND_878;
  reg [6:0] _T_5936_23_pdst;
  reg [31:0] _RAND_879;
  reg [6:0] _T_5936_23_stale_pdst;
  reg [31:0] _RAND_880;
  reg  _T_5936_23_is_fencei;
  reg [31:0] _RAND_881;
  reg  _T_5936_23_is_store;
  reg [31:0] _RAND_882;
  reg  _T_5936_23_is_load;
  reg [31:0] _RAND_883;
  reg  _T_5936_23_is_sys_pc2epc;
  reg [31:0] _RAND_884;
  reg  _T_5936_23_flush_on_commit;
  reg [31:0] _RAND_885;
  reg [5:0] _T_5936_23_ldst;
  reg [31:0] _RAND_886;
  reg  _T_5936_23_ldst_val;
  reg [31:0] _RAND_887;
  reg [1:0] _T_5936_23_dst_rtype;
  reg [31:0] _RAND_888;
  reg  _T_5936_23_fp_val;
  reg [31:0] _RAND_889;
  reg [7:0] _T_5936_24_br_mask;
  reg [31:0] _RAND_890;
  reg [6:0] _T_5936_24_pdst;
  reg [31:0] _RAND_891;
  reg [6:0] _T_5936_24_stale_pdst;
  reg [31:0] _RAND_892;
  reg  _T_5936_24_is_fencei;
  reg [31:0] _RAND_893;
  reg  _T_5936_24_is_store;
  reg [31:0] _RAND_894;
  reg  _T_5936_24_is_load;
  reg [31:0] _RAND_895;
  reg  _T_5936_24_is_sys_pc2epc;
  reg [31:0] _RAND_896;
  reg  _T_5936_24_flush_on_commit;
  reg [31:0] _RAND_897;
  reg [5:0] _T_5936_24_ldst;
  reg [31:0] _RAND_898;
  reg  _T_5936_24_ldst_val;
  reg [31:0] _RAND_899;
  reg [1:0] _T_5936_24_dst_rtype;
  reg [31:0] _RAND_900;
  reg  _T_5936_24_fp_val;
  reg [31:0] _RAND_901;
  reg [7:0] _T_5936_25_br_mask;
  reg [31:0] _RAND_902;
  reg [6:0] _T_5936_25_pdst;
  reg [31:0] _RAND_903;
  reg [6:0] _T_5936_25_stale_pdst;
  reg [31:0] _RAND_904;
  reg  _T_5936_25_is_fencei;
  reg [31:0] _RAND_905;
  reg  _T_5936_25_is_store;
  reg [31:0] _RAND_906;
  reg  _T_5936_25_is_load;
  reg [31:0] _RAND_907;
  reg  _T_5936_25_is_sys_pc2epc;
  reg [31:0] _RAND_908;
  reg  _T_5936_25_flush_on_commit;
  reg [31:0] _RAND_909;
  reg [5:0] _T_5936_25_ldst;
  reg [31:0] _RAND_910;
  reg  _T_5936_25_ldst_val;
  reg [31:0] _RAND_911;
  reg [1:0] _T_5936_25_dst_rtype;
  reg [31:0] _RAND_912;
  reg  _T_5936_25_fp_val;
  reg [31:0] _RAND_913;
  reg [7:0] _T_5936_26_br_mask;
  reg [31:0] _RAND_914;
  reg [6:0] _T_5936_26_pdst;
  reg [31:0] _RAND_915;
  reg [6:0] _T_5936_26_stale_pdst;
  reg [31:0] _RAND_916;
  reg  _T_5936_26_is_fencei;
  reg [31:0] _RAND_917;
  reg  _T_5936_26_is_store;
  reg [31:0] _RAND_918;
  reg  _T_5936_26_is_load;
  reg [31:0] _RAND_919;
  reg  _T_5936_26_is_sys_pc2epc;
  reg [31:0] _RAND_920;
  reg  _T_5936_26_flush_on_commit;
  reg [31:0] _RAND_921;
  reg [5:0] _T_5936_26_ldst;
  reg [31:0] _RAND_922;
  reg  _T_5936_26_ldst_val;
  reg [31:0] _RAND_923;
  reg [1:0] _T_5936_26_dst_rtype;
  reg [31:0] _RAND_924;
  reg  _T_5936_26_fp_val;
  reg [31:0] _RAND_925;
  reg [7:0] _T_5936_27_br_mask;
  reg [31:0] _RAND_926;
  reg [6:0] _T_5936_27_pdst;
  reg [31:0] _RAND_927;
  reg [6:0] _T_5936_27_stale_pdst;
  reg [31:0] _RAND_928;
  reg  _T_5936_27_is_fencei;
  reg [31:0] _RAND_929;
  reg  _T_5936_27_is_store;
  reg [31:0] _RAND_930;
  reg  _T_5936_27_is_load;
  reg [31:0] _RAND_931;
  reg  _T_5936_27_is_sys_pc2epc;
  reg [31:0] _RAND_932;
  reg  _T_5936_27_flush_on_commit;
  reg [31:0] _RAND_933;
  reg [5:0] _T_5936_27_ldst;
  reg [31:0] _RAND_934;
  reg  _T_5936_27_ldst_val;
  reg [31:0] _RAND_935;
  reg [1:0] _T_5936_27_dst_rtype;
  reg [31:0] _RAND_936;
  reg  _T_5936_27_fp_val;
  reg [31:0] _RAND_937;
  reg [7:0] _T_5936_28_br_mask;
  reg [31:0] _RAND_938;
  reg [6:0] _T_5936_28_pdst;
  reg [31:0] _RAND_939;
  reg [6:0] _T_5936_28_stale_pdst;
  reg [31:0] _RAND_940;
  reg  _T_5936_28_is_fencei;
  reg [31:0] _RAND_941;
  reg  _T_5936_28_is_store;
  reg [31:0] _RAND_942;
  reg  _T_5936_28_is_load;
  reg [31:0] _RAND_943;
  reg  _T_5936_28_is_sys_pc2epc;
  reg [31:0] _RAND_944;
  reg  _T_5936_28_flush_on_commit;
  reg [31:0] _RAND_945;
  reg [5:0] _T_5936_28_ldst;
  reg [31:0] _RAND_946;
  reg  _T_5936_28_ldst_val;
  reg [31:0] _RAND_947;
  reg [1:0] _T_5936_28_dst_rtype;
  reg [31:0] _RAND_948;
  reg  _T_5936_28_fp_val;
  reg [31:0] _RAND_949;
  reg [7:0] _T_5936_29_br_mask;
  reg [31:0] _RAND_950;
  reg [6:0] _T_5936_29_pdst;
  reg [31:0] _RAND_951;
  reg [6:0] _T_5936_29_stale_pdst;
  reg [31:0] _RAND_952;
  reg  _T_5936_29_is_fencei;
  reg [31:0] _RAND_953;
  reg  _T_5936_29_is_store;
  reg [31:0] _RAND_954;
  reg  _T_5936_29_is_load;
  reg [31:0] _RAND_955;
  reg  _T_5936_29_is_sys_pc2epc;
  reg [31:0] _RAND_956;
  reg  _T_5936_29_flush_on_commit;
  reg [31:0] _RAND_957;
  reg [5:0] _T_5936_29_ldst;
  reg [31:0] _RAND_958;
  reg  _T_5936_29_ldst_val;
  reg [31:0] _RAND_959;
  reg [1:0] _T_5936_29_dst_rtype;
  reg [31:0] _RAND_960;
  reg  _T_5936_29_fp_val;
  reg [31:0] _RAND_961;
  reg [7:0] _T_5936_30_br_mask;
  reg [31:0] _RAND_962;
  reg [6:0] _T_5936_30_pdst;
  reg [31:0] _RAND_963;
  reg [6:0] _T_5936_30_stale_pdst;
  reg [31:0] _RAND_964;
  reg  _T_5936_30_is_fencei;
  reg [31:0] _RAND_965;
  reg  _T_5936_30_is_store;
  reg [31:0] _RAND_966;
  reg  _T_5936_30_is_load;
  reg [31:0] _RAND_967;
  reg  _T_5936_30_is_sys_pc2epc;
  reg [31:0] _RAND_968;
  reg  _T_5936_30_flush_on_commit;
  reg [31:0] _RAND_969;
  reg [5:0] _T_5936_30_ldst;
  reg [31:0] _RAND_970;
  reg  _T_5936_30_ldst_val;
  reg [31:0] _RAND_971;
  reg [1:0] _T_5936_30_dst_rtype;
  reg [31:0] _RAND_972;
  reg  _T_5936_30_fp_val;
  reg [31:0] _RAND_973;
  reg [7:0] _T_5936_31_br_mask;
  reg [31:0] _RAND_974;
  reg [6:0] _T_5936_31_pdst;
  reg [31:0] _RAND_975;
  reg [6:0] _T_5936_31_stale_pdst;
  reg [31:0] _RAND_976;
  reg  _T_5936_31_is_fencei;
  reg [31:0] _RAND_977;
  reg  _T_5936_31_is_store;
  reg [31:0] _RAND_978;
  reg  _T_5936_31_is_load;
  reg [31:0] _RAND_979;
  reg  _T_5936_31_is_sys_pc2epc;
  reg [31:0] _RAND_980;
  reg  _T_5936_31_flush_on_commit;
  reg [31:0] _RAND_981;
  reg [5:0] _T_5936_31_ldst;
  reg [31:0] _RAND_982;
  reg  _T_5936_31_ldst_val;
  reg [31:0] _RAND_983;
  reg [1:0] _T_5936_31_dst_rtype;
  reg [31:0] _RAND_984;
  reg  _T_5936_31_fp_val;
  reg [31:0] _RAND_985;
  reg [7:0] _T_5936_32_br_mask;
  reg [31:0] _RAND_986;
  reg [6:0] _T_5936_32_pdst;
  reg [31:0] _RAND_987;
  reg [6:0] _T_5936_32_stale_pdst;
  reg [31:0] _RAND_988;
  reg  _T_5936_32_is_fencei;
  reg [31:0] _RAND_989;
  reg  _T_5936_32_is_store;
  reg [31:0] _RAND_990;
  reg  _T_5936_32_is_load;
  reg [31:0] _RAND_991;
  reg  _T_5936_32_is_sys_pc2epc;
  reg [31:0] _RAND_992;
  reg  _T_5936_32_flush_on_commit;
  reg [31:0] _RAND_993;
  reg [5:0] _T_5936_32_ldst;
  reg [31:0] _RAND_994;
  reg  _T_5936_32_ldst_val;
  reg [31:0] _RAND_995;
  reg [1:0] _T_5936_32_dst_rtype;
  reg [31:0] _RAND_996;
  reg  _T_5936_32_fp_val;
  reg [31:0] _RAND_997;
  reg [7:0] _T_5936_33_br_mask;
  reg [31:0] _RAND_998;
  reg [6:0] _T_5936_33_pdst;
  reg [31:0] _RAND_999;
  reg [6:0] _T_5936_33_stale_pdst;
  reg [31:0] _RAND_1000;
  reg  _T_5936_33_is_fencei;
  reg [31:0] _RAND_1001;
  reg  _T_5936_33_is_store;
  reg [31:0] _RAND_1002;
  reg  _T_5936_33_is_load;
  reg [31:0] _RAND_1003;
  reg  _T_5936_33_is_sys_pc2epc;
  reg [31:0] _RAND_1004;
  reg  _T_5936_33_flush_on_commit;
  reg [31:0] _RAND_1005;
  reg [5:0] _T_5936_33_ldst;
  reg [31:0] _RAND_1006;
  reg  _T_5936_33_ldst_val;
  reg [31:0] _RAND_1007;
  reg [1:0] _T_5936_33_dst_rtype;
  reg [31:0] _RAND_1008;
  reg  _T_5936_33_fp_val;
  reg [31:0] _RAND_1009;
  reg [7:0] _T_5936_34_br_mask;
  reg [31:0] _RAND_1010;
  reg [6:0] _T_5936_34_pdst;
  reg [31:0] _RAND_1011;
  reg [6:0] _T_5936_34_stale_pdst;
  reg [31:0] _RAND_1012;
  reg  _T_5936_34_is_fencei;
  reg [31:0] _RAND_1013;
  reg  _T_5936_34_is_store;
  reg [31:0] _RAND_1014;
  reg  _T_5936_34_is_load;
  reg [31:0] _RAND_1015;
  reg  _T_5936_34_is_sys_pc2epc;
  reg [31:0] _RAND_1016;
  reg  _T_5936_34_flush_on_commit;
  reg [31:0] _RAND_1017;
  reg [5:0] _T_5936_34_ldst;
  reg [31:0] _RAND_1018;
  reg  _T_5936_34_ldst_val;
  reg [31:0] _RAND_1019;
  reg [1:0] _T_5936_34_dst_rtype;
  reg [31:0] _RAND_1020;
  reg  _T_5936_34_fp_val;
  reg [31:0] _RAND_1021;
  reg [7:0] _T_5936_35_br_mask;
  reg [31:0] _RAND_1022;
  reg [6:0] _T_5936_35_pdst;
  reg [31:0] _RAND_1023;
  reg [6:0] _T_5936_35_stale_pdst;
  reg [31:0] _RAND_1024;
  reg  _T_5936_35_is_fencei;
  reg [31:0] _RAND_1025;
  reg  _T_5936_35_is_store;
  reg [31:0] _RAND_1026;
  reg  _T_5936_35_is_load;
  reg [31:0] _RAND_1027;
  reg  _T_5936_35_is_sys_pc2epc;
  reg [31:0] _RAND_1028;
  reg  _T_5936_35_flush_on_commit;
  reg [31:0] _RAND_1029;
  reg [5:0] _T_5936_35_ldst;
  reg [31:0] _RAND_1030;
  reg  _T_5936_35_ldst_val;
  reg [31:0] _RAND_1031;
  reg [1:0] _T_5936_35_dst_rtype;
  reg [31:0] _RAND_1032;
  reg  _T_5936_35_fp_val;
  reg [31:0] _RAND_1033;
  reg [7:0] _T_5936_36_br_mask;
  reg [31:0] _RAND_1034;
  reg [6:0] _T_5936_36_pdst;
  reg [31:0] _RAND_1035;
  reg [6:0] _T_5936_36_stale_pdst;
  reg [31:0] _RAND_1036;
  reg  _T_5936_36_is_fencei;
  reg [31:0] _RAND_1037;
  reg  _T_5936_36_is_store;
  reg [31:0] _RAND_1038;
  reg  _T_5936_36_is_load;
  reg [31:0] _RAND_1039;
  reg  _T_5936_36_is_sys_pc2epc;
  reg [31:0] _RAND_1040;
  reg  _T_5936_36_flush_on_commit;
  reg [31:0] _RAND_1041;
  reg [5:0] _T_5936_36_ldst;
  reg [31:0] _RAND_1042;
  reg  _T_5936_36_ldst_val;
  reg [31:0] _RAND_1043;
  reg [1:0] _T_5936_36_dst_rtype;
  reg [31:0] _RAND_1044;
  reg  _T_5936_36_fp_val;
  reg [31:0] _RAND_1045;
  reg [7:0] _T_5936_37_br_mask;
  reg [31:0] _RAND_1046;
  reg [6:0] _T_5936_37_pdst;
  reg [31:0] _RAND_1047;
  reg [6:0] _T_5936_37_stale_pdst;
  reg [31:0] _RAND_1048;
  reg  _T_5936_37_is_fencei;
  reg [31:0] _RAND_1049;
  reg  _T_5936_37_is_store;
  reg [31:0] _RAND_1050;
  reg  _T_5936_37_is_load;
  reg [31:0] _RAND_1051;
  reg  _T_5936_37_is_sys_pc2epc;
  reg [31:0] _RAND_1052;
  reg  _T_5936_37_flush_on_commit;
  reg [31:0] _RAND_1053;
  reg [5:0] _T_5936_37_ldst;
  reg [31:0] _RAND_1054;
  reg  _T_5936_37_ldst_val;
  reg [31:0] _RAND_1055;
  reg [1:0] _T_5936_37_dst_rtype;
  reg [31:0] _RAND_1056;
  reg  _T_5936_37_fp_val;
  reg [31:0] _RAND_1057;
  reg [7:0] _T_5936_38_br_mask;
  reg [31:0] _RAND_1058;
  reg [6:0] _T_5936_38_pdst;
  reg [31:0] _RAND_1059;
  reg [6:0] _T_5936_38_stale_pdst;
  reg [31:0] _RAND_1060;
  reg  _T_5936_38_is_fencei;
  reg [31:0] _RAND_1061;
  reg  _T_5936_38_is_store;
  reg [31:0] _RAND_1062;
  reg  _T_5936_38_is_load;
  reg [31:0] _RAND_1063;
  reg  _T_5936_38_is_sys_pc2epc;
  reg [31:0] _RAND_1064;
  reg  _T_5936_38_flush_on_commit;
  reg [31:0] _RAND_1065;
  reg [5:0] _T_5936_38_ldst;
  reg [31:0] _RAND_1066;
  reg  _T_5936_38_ldst_val;
  reg [31:0] _RAND_1067;
  reg [1:0] _T_5936_38_dst_rtype;
  reg [31:0] _RAND_1068;
  reg  _T_5936_38_fp_val;
  reg [31:0] _RAND_1069;
  reg [7:0] _T_5936_39_br_mask;
  reg [31:0] _RAND_1070;
  reg [6:0] _T_5936_39_pdst;
  reg [31:0] _RAND_1071;
  reg [6:0] _T_5936_39_stale_pdst;
  reg [31:0] _RAND_1072;
  reg  _T_5936_39_is_fencei;
  reg [31:0] _RAND_1073;
  reg  _T_5936_39_is_store;
  reg [31:0] _RAND_1074;
  reg  _T_5936_39_is_load;
  reg [31:0] _RAND_1075;
  reg  _T_5936_39_is_sys_pc2epc;
  reg [31:0] _RAND_1076;
  reg  _T_5936_39_flush_on_commit;
  reg [31:0] _RAND_1077;
  reg [5:0] _T_5936_39_ldst;
  reg [31:0] _RAND_1078;
  reg  _T_5936_39_ldst_val;
  reg [31:0] _RAND_1079;
  reg [1:0] _T_5936_39_dst_rtype;
  reg [31:0] _RAND_1080;
  reg  _T_5936_39_fp_val;
  reg [31:0] _RAND_1081;
  reg  _T_6309 [0:39];
  reg [31:0] _RAND_1082;
  wire  _T_6309__T_6576_data;
  wire [5:0] _T_6309__T_6576_addr;
  reg [31:0] _RAND_1083;
  wire  _T_6309__T_6332_data;
  wire [5:0] _T_6309__T_6332_addr;
  wire  _T_6309__T_6332_mask;
  wire  _T_6309__T_6332_en;
  wire  _T_6309__T_6562_data;
  wire [5:0] _T_6309__T_6562_addr;
  wire  _T_6309__T_6562_mask;
  wire  _T_6309__T_6562_en;
  wire  _T_6309__T_6571_data;
  wire [5:0] _T_6309__T_6571_addr;
  wire  _T_6309__T_6571_mask;
  wire  _T_6309__T_6571_en;
  wire  _T_6309__T_6652_data;
  wire [5:0] _T_6309__T_6652_addr;
  wire  _T_6309__T_6652_mask;
  wire  _T_6309__T_6652_en;
  reg [4:0] _T_6312 [0:39];
  reg [31:0] _RAND_1084;
  wire [4:0] _T_6312__T_7581_data;
  wire [5:0] _T_6312__T_7581_addr;
  reg [31:0] _RAND_1085;
  wire [4:0] _T_6312__T_6333_data;
  wire [5:0] _T_6312__T_6333_addr;
  wire  _T_6312__T_6333_mask;
  wire  _T_6312__T_6333_en;
  wire [4:0] _T_6312__T_6546_data;
  wire [5:0] _T_6312__T_6546_addr;
  wire  _T_6312__T_6546_mask;
  wire  _T_6312__T_6546_en;
  wire [4:0] _T_6312__T_6554_data;
  wire [5:0] _T_6312__T_6554_addr;
  wire  _T_6312__T_6554_mask;
  wire  _T_6312__T_6554_en;
  wire  _GEN_41370;
  wire  _GEN_41371;
  wire  _GEN_41372;
  wire  _GEN_41373;
  wire  _GEN_41374;
  wire  _GEN_41375;
  wire  _GEN_41376;
  wire  _GEN_41377;
  wire  _GEN_41378;
  wire  _GEN_41379;
  wire  _GEN_41380;
  wire  _GEN_41381;
  wire  _GEN_41382;
  wire  _GEN_41383;
  wire  _GEN_41384;
  wire  _GEN_41385;
  wire  _GEN_41386;
  wire  _GEN_41387;
  wire  _GEN_41388;
  wire  _GEN_41389;
  wire  _GEN_41390;
  wire  _GEN_41391;
  wire  _GEN_41392;
  wire  _GEN_41393;
  wire  _GEN_41394;
  wire  _GEN_41395;
  wire  _GEN_41396;
  wire  _GEN_41397;
  wire  _GEN_41398;
  wire  _GEN_41399;
  wire  _GEN_41400;
  wire  _GEN_41401;
  wire  _GEN_41402;
  wire  _GEN_41403;
  wire  _GEN_41404;
  wire  _GEN_41405;
  wire  _GEN_41406;
  wire  _GEN_41407;
  wire  _GEN_41408;
  wire  _GEN_41409;
  wire  _T_6319;
  wire  _T_6321;
  wire  _T_6322;
  wire [7:0] _GEN_253;
  wire [7:0] _GEN_42370;
  wire [7:0] _GEN_42371;
  wire [7:0] _GEN_42372;
  wire [7:0] _GEN_42373;
  wire [7:0] _GEN_42374;
  wire [7:0] _GEN_42375;
  wire [7:0] _GEN_42376;
  wire [7:0] _GEN_42377;
  wire [7:0] _GEN_42378;
  wire [7:0] _GEN_42379;
  wire [7:0] _GEN_42380;
  wire [7:0] _GEN_42381;
  wire [7:0] _GEN_42382;
  wire [7:0] _GEN_42383;
  wire [7:0] _GEN_42384;
  wire [7:0] _GEN_42385;
  wire [7:0] _GEN_42386;
  wire [7:0] _GEN_42387;
  wire [7:0] _GEN_42388;
  wire [7:0] _GEN_42389;
  wire [7:0] _GEN_42390;
  wire [7:0] _GEN_42391;
  wire [7:0] _GEN_42392;
  wire [7:0] _GEN_42393;
  wire [7:0] _GEN_42394;
  wire [7:0] _GEN_42395;
  wire [7:0] _GEN_42396;
  wire [7:0] _GEN_42397;
  wire [7:0] _GEN_42398;
  wire [7:0] _GEN_42399;
  wire [7:0] _GEN_42400;
  wire [7:0] _GEN_42401;
  wire [7:0] _GEN_42402;
  wire [7:0] _GEN_42403;
  wire [7:0] _GEN_42404;
  wire [7:0] _GEN_42405;
  wire [7:0] _GEN_42406;
  wire [7:0] _GEN_42407;
  wire [7:0] _GEN_42408;
  wire [7:0] _GEN_42409;
  wire [6:0] _GEN_281;
  wire [6:0] _GEN_43490;
  wire [6:0] _GEN_43491;
  wire [6:0] _GEN_43492;
  wire [6:0] _GEN_43493;
  wire [6:0] _GEN_43494;
  wire [6:0] _GEN_43495;
  wire [6:0] _GEN_43496;
  wire [6:0] _GEN_43497;
  wire [6:0] _GEN_43498;
  wire [6:0] _GEN_43499;
  wire [6:0] _GEN_43500;
  wire [6:0] _GEN_43501;
  wire [6:0] _GEN_43502;
  wire [6:0] _GEN_43503;
  wire [6:0] _GEN_43504;
  wire [6:0] _GEN_43505;
  wire [6:0] _GEN_43506;
  wire [6:0] _GEN_43507;
  wire [6:0] _GEN_43508;
  wire [6:0] _GEN_43509;
  wire [6:0] _GEN_43510;
  wire [6:0] _GEN_43511;
  wire [6:0] _GEN_43512;
  wire [6:0] _GEN_43513;
  wire [6:0] _GEN_43514;
  wire [6:0] _GEN_43515;
  wire [6:0] _GEN_43516;
  wire [6:0] _GEN_43517;
  wire [6:0] _GEN_43518;
  wire [6:0] _GEN_43519;
  wire [6:0] _GEN_43520;
  wire [6:0] _GEN_43521;
  wire [6:0] _GEN_43522;
  wire [6:0] _GEN_43523;
  wire [6:0] _GEN_43524;
  wire [6:0] _GEN_43525;
  wire [6:0] _GEN_43526;
  wire [6:0] _GEN_43527;
  wire [6:0] _GEN_43528;
  wire [6:0] _GEN_43529;
  wire [6:0] _GEN_288;
  wire [6:0] _GEN_43770;
  wire [6:0] _GEN_43771;
  wire [6:0] _GEN_43772;
  wire [6:0] _GEN_43773;
  wire [6:0] _GEN_43774;
  wire [6:0] _GEN_43775;
  wire [6:0] _GEN_43776;
  wire [6:0] _GEN_43777;
  wire [6:0] _GEN_43778;
  wire [6:0] _GEN_43779;
  wire [6:0] _GEN_43780;
  wire [6:0] _GEN_43781;
  wire [6:0] _GEN_43782;
  wire [6:0] _GEN_43783;
  wire [6:0] _GEN_43784;
  wire [6:0] _GEN_43785;
  wire [6:0] _GEN_43786;
  wire [6:0] _GEN_43787;
  wire [6:0] _GEN_43788;
  wire [6:0] _GEN_43789;
  wire [6:0] _GEN_43790;
  wire [6:0] _GEN_43791;
  wire [6:0] _GEN_43792;
  wire [6:0] _GEN_43793;
  wire [6:0] _GEN_43794;
  wire [6:0] _GEN_43795;
  wire [6:0] _GEN_43796;
  wire [6:0] _GEN_43797;
  wire [6:0] _GEN_43798;
  wire [6:0] _GEN_43799;
  wire [6:0] _GEN_43800;
  wire [6:0] _GEN_43801;
  wire [6:0] _GEN_43802;
  wire [6:0] _GEN_43803;
  wire [6:0] _GEN_43804;
  wire [6:0] _GEN_43805;
  wire [6:0] _GEN_43806;
  wire [6:0] _GEN_43807;
  wire [6:0] _GEN_43808;
  wire [6:0] _GEN_43809;
  wire  _GEN_295;
  wire  _GEN_44050;
  wire  _GEN_44051;
  wire  _GEN_44052;
  wire  _GEN_44053;
  wire  _GEN_44054;
  wire  _GEN_44055;
  wire  _GEN_44056;
  wire  _GEN_44057;
  wire  _GEN_44058;
  wire  _GEN_44059;
  wire  _GEN_44060;
  wire  _GEN_44061;
  wire  _GEN_44062;
  wire  _GEN_44063;
  wire  _GEN_44064;
  wire  _GEN_44065;
  wire  _GEN_44066;
  wire  _GEN_44067;
  wire  _GEN_44068;
  wire  _GEN_44069;
  wire  _GEN_44070;
  wire  _GEN_44071;
  wire  _GEN_44072;
  wire  _GEN_44073;
  wire  _GEN_44074;
  wire  _GEN_44075;
  wire  _GEN_44076;
  wire  _GEN_44077;
  wire  _GEN_44078;
  wire  _GEN_44079;
  wire  _GEN_44080;
  wire  _GEN_44081;
  wire  _GEN_44082;
  wire  _GEN_44083;
  wire  _GEN_44084;
  wire  _GEN_44085;
  wire  _GEN_44086;
  wire  _GEN_44087;
  wire  _GEN_44088;
  wire  _GEN_44089;
  wire  _GEN_296;
  wire  _GEN_44090;
  wire  _GEN_44091;
  wire  _GEN_44092;
  wire  _GEN_44093;
  wire  _GEN_44094;
  wire  _GEN_44095;
  wire  _GEN_44096;
  wire  _GEN_44097;
  wire  _GEN_44098;
  wire  _GEN_44099;
  wire  _GEN_44100;
  wire  _GEN_44101;
  wire  _GEN_44102;
  wire  _GEN_44103;
  wire  _GEN_44104;
  wire  _GEN_44105;
  wire  _GEN_44106;
  wire  _GEN_44107;
  wire  _GEN_44108;
  wire  _GEN_44109;
  wire  _GEN_44110;
  wire  _GEN_44111;
  wire  _GEN_44112;
  wire  _GEN_44113;
  wire  _GEN_44114;
  wire  _GEN_44115;
  wire  _GEN_44116;
  wire  _GEN_44117;
  wire  _GEN_44118;
  wire  _GEN_44119;
  wire  _GEN_44120;
  wire  _GEN_44121;
  wire  _GEN_44122;
  wire  _GEN_44123;
  wire  _GEN_44124;
  wire  _GEN_44125;
  wire  _GEN_44126;
  wire  _GEN_44127;
  wire  _GEN_44128;
  wire  _GEN_44129;
  wire  _GEN_298;
  wire  _GEN_44170;
  wire  _GEN_44171;
  wire  _GEN_44172;
  wire  _GEN_44173;
  wire  _GEN_44174;
  wire  _GEN_44175;
  wire  _GEN_44176;
  wire  _GEN_44177;
  wire  _GEN_44178;
  wire  _GEN_44179;
  wire  _GEN_44180;
  wire  _GEN_44181;
  wire  _GEN_44182;
  wire  _GEN_44183;
  wire  _GEN_44184;
  wire  _GEN_44185;
  wire  _GEN_44186;
  wire  _GEN_44187;
  wire  _GEN_44188;
  wire  _GEN_44189;
  wire  _GEN_44190;
  wire  _GEN_44191;
  wire  _GEN_44192;
  wire  _GEN_44193;
  wire  _GEN_44194;
  wire  _GEN_44195;
  wire  _GEN_44196;
  wire  _GEN_44197;
  wire  _GEN_44198;
  wire  _GEN_44199;
  wire  _GEN_44200;
  wire  _GEN_44201;
  wire  _GEN_44202;
  wire  _GEN_44203;
  wire  _GEN_44204;
  wire  _GEN_44205;
  wire  _GEN_44206;
  wire  _GEN_44207;
  wire  _GEN_44208;
  wire  _GEN_44209;
  wire  _GEN_299;
  wire  _GEN_44210;
  wire  _GEN_44211;
  wire  _GEN_44212;
  wire  _GEN_44213;
  wire  _GEN_44214;
  wire  _GEN_44215;
  wire  _GEN_44216;
  wire  _GEN_44217;
  wire  _GEN_44218;
  wire  _GEN_44219;
  wire  _GEN_44220;
  wire  _GEN_44221;
  wire  _GEN_44222;
  wire  _GEN_44223;
  wire  _GEN_44224;
  wire  _GEN_44225;
  wire  _GEN_44226;
  wire  _GEN_44227;
  wire  _GEN_44228;
  wire  _GEN_44229;
  wire  _GEN_44230;
  wire  _GEN_44231;
  wire  _GEN_44232;
  wire  _GEN_44233;
  wire  _GEN_44234;
  wire  _GEN_44235;
  wire  _GEN_44236;
  wire  _GEN_44237;
  wire  _GEN_44238;
  wire  _GEN_44239;
  wire  _GEN_44240;
  wire  _GEN_44241;
  wire  _GEN_44242;
  wire  _GEN_44243;
  wire  _GEN_44244;
  wire  _GEN_44245;
  wire  _GEN_44246;
  wire  _GEN_44247;
  wire  _GEN_44248;
  wire  _GEN_44249;
  wire  _GEN_301;
  wire  _GEN_44290;
  wire  _GEN_44291;
  wire  _GEN_44292;
  wire  _GEN_44293;
  wire  _GEN_44294;
  wire  _GEN_44295;
  wire  _GEN_44296;
  wire  _GEN_44297;
  wire  _GEN_44298;
  wire  _GEN_44299;
  wire  _GEN_44300;
  wire  _GEN_44301;
  wire  _GEN_44302;
  wire  _GEN_44303;
  wire  _GEN_44304;
  wire  _GEN_44305;
  wire  _GEN_44306;
  wire  _GEN_44307;
  wire  _GEN_44308;
  wire  _GEN_44309;
  wire  _GEN_44310;
  wire  _GEN_44311;
  wire  _GEN_44312;
  wire  _GEN_44313;
  wire  _GEN_44314;
  wire  _GEN_44315;
  wire  _GEN_44316;
  wire  _GEN_44317;
  wire  _GEN_44318;
  wire  _GEN_44319;
  wire  _GEN_44320;
  wire  _GEN_44321;
  wire  _GEN_44322;
  wire  _GEN_44323;
  wire  _GEN_44324;
  wire  _GEN_44325;
  wire  _GEN_44326;
  wire  _GEN_44327;
  wire  _GEN_44328;
  wire  _GEN_44329;
  wire [5:0] _GEN_302;
  wire [5:0] _GEN_44330;
  wire [5:0] _GEN_44331;
  wire [5:0] _GEN_44332;
  wire [5:0] _GEN_44333;
  wire [5:0] _GEN_44334;
  wire [5:0] _GEN_44335;
  wire [5:0] _GEN_44336;
  wire [5:0] _GEN_44337;
  wire [5:0] _GEN_44338;
  wire [5:0] _GEN_44339;
  wire [5:0] _GEN_44340;
  wire [5:0] _GEN_44341;
  wire [5:0] _GEN_44342;
  wire [5:0] _GEN_44343;
  wire [5:0] _GEN_44344;
  wire [5:0] _GEN_44345;
  wire [5:0] _GEN_44346;
  wire [5:0] _GEN_44347;
  wire [5:0] _GEN_44348;
  wire [5:0] _GEN_44349;
  wire [5:0] _GEN_44350;
  wire [5:0] _GEN_44351;
  wire [5:0] _GEN_44352;
  wire [5:0] _GEN_44353;
  wire [5:0] _GEN_44354;
  wire [5:0] _GEN_44355;
  wire [5:0] _GEN_44356;
  wire [5:0] _GEN_44357;
  wire [5:0] _GEN_44358;
  wire [5:0] _GEN_44359;
  wire [5:0] _GEN_44360;
  wire [5:0] _GEN_44361;
  wire [5:0] _GEN_44362;
  wire [5:0] _GEN_44363;
  wire [5:0] _GEN_44364;
  wire [5:0] _GEN_44365;
  wire [5:0] _GEN_44366;
  wire [5:0] _GEN_44367;
  wire [5:0] _GEN_44368;
  wire [5:0] _GEN_44369;
  wire  _GEN_306;
  wire  _GEN_44490;
  wire  _GEN_44491;
  wire  _GEN_44492;
  wire  _GEN_44493;
  wire  _GEN_44494;
  wire  _GEN_44495;
  wire  _GEN_44496;
  wire  _GEN_44497;
  wire  _GEN_44498;
  wire  _GEN_44499;
  wire  _GEN_44500;
  wire  _GEN_44501;
  wire  _GEN_44502;
  wire  _GEN_44503;
  wire  _GEN_44504;
  wire  _GEN_44505;
  wire  _GEN_44506;
  wire  _GEN_44507;
  wire  _GEN_44508;
  wire  _GEN_44509;
  wire  _GEN_44510;
  wire  _GEN_44511;
  wire  _GEN_44512;
  wire  _GEN_44513;
  wire  _GEN_44514;
  wire  _GEN_44515;
  wire  _GEN_44516;
  wire  _GEN_44517;
  wire  _GEN_44518;
  wire  _GEN_44519;
  wire  _GEN_44520;
  wire  _GEN_44521;
  wire  _GEN_44522;
  wire  _GEN_44523;
  wire  _GEN_44524;
  wire  _GEN_44525;
  wire  _GEN_44526;
  wire  _GEN_44527;
  wire  _GEN_44528;
  wire  _GEN_44529;
  wire [1:0] _GEN_307;
  wire [1:0] _GEN_44530;
  wire [1:0] _GEN_44531;
  wire [1:0] _GEN_44532;
  wire [1:0] _GEN_44533;
  wire [1:0] _GEN_44534;
  wire [1:0] _GEN_44535;
  wire [1:0] _GEN_44536;
  wire [1:0] _GEN_44537;
  wire [1:0] _GEN_44538;
  wire [1:0] _GEN_44539;
  wire [1:0] _GEN_44540;
  wire [1:0] _GEN_44541;
  wire [1:0] _GEN_44542;
  wire [1:0] _GEN_44543;
  wire [1:0] _GEN_44544;
  wire [1:0] _GEN_44545;
  wire [1:0] _GEN_44546;
  wire [1:0] _GEN_44547;
  wire [1:0] _GEN_44548;
  wire [1:0] _GEN_44549;
  wire [1:0] _GEN_44550;
  wire [1:0] _GEN_44551;
  wire [1:0] _GEN_44552;
  wire [1:0] _GEN_44553;
  wire [1:0] _GEN_44554;
  wire [1:0] _GEN_44555;
  wire [1:0] _GEN_44556;
  wire [1:0] _GEN_44557;
  wire [1:0] _GEN_44558;
  wire [1:0] _GEN_44559;
  wire [1:0] _GEN_44560;
  wire [1:0] _GEN_44561;
  wire [1:0] _GEN_44562;
  wire [1:0] _GEN_44563;
  wire [1:0] _GEN_44564;
  wire [1:0] _GEN_44565;
  wire [1:0] _GEN_44566;
  wire [1:0] _GEN_44567;
  wire [1:0] _GEN_44568;
  wire [1:0] _GEN_44569;
  wire  _GEN_311;
  wire  _GEN_44690;
  wire  _GEN_44691;
  wire  _GEN_44692;
  wire  _GEN_44693;
  wire  _GEN_44694;
  wire  _GEN_44695;
  wire  _GEN_44696;
  wire  _GEN_44697;
  wire  _GEN_44698;
  wire  _GEN_44699;
  wire  _GEN_44700;
  wire  _GEN_44701;
  wire  _GEN_44702;
  wire  _GEN_44703;
  wire  _GEN_44704;
  wire  _GEN_44705;
  wire  _GEN_44706;
  wire  _GEN_44707;
  wire  _GEN_44708;
  wire  _GEN_44709;
  wire  _GEN_44710;
  wire  _GEN_44711;
  wire  _GEN_44712;
  wire  _GEN_44713;
  wire  _GEN_44714;
  wire  _GEN_44715;
  wire  _GEN_44716;
  wire  _GEN_44717;
  wire  _GEN_44718;
  wire  _GEN_44719;
  wire  _GEN_44720;
  wire  _GEN_44721;
  wire  _GEN_44722;
  wire  _GEN_44723;
  wire  _GEN_44724;
  wire  _GEN_44725;
  wire  _GEN_44726;
  wire  _GEN_44727;
  wire  _GEN_44728;
  wire  _GEN_44729;
  wire  _GEN_320;
  wire  _GEN_45050;
  wire  _GEN_45051;
  wire  _GEN_45052;
  wire  _GEN_45053;
  wire  _GEN_45054;
  wire  _GEN_45055;
  wire  _GEN_45056;
  wire  _GEN_45057;
  wire  _GEN_45058;
  wire  _GEN_45059;
  wire  _GEN_45060;
  wire  _GEN_45061;
  wire  _GEN_45062;
  wire  _GEN_45063;
  wire  _GEN_45064;
  wire  _GEN_45065;
  wire  _GEN_45066;
  wire  _GEN_45067;
  wire  _GEN_45068;
  wire  _GEN_45069;
  wire  _GEN_45070;
  wire  _GEN_45071;
  wire  _GEN_45072;
  wire  _GEN_45073;
  wire  _GEN_45074;
  wire  _GEN_45075;
  wire  _GEN_45076;
  wire  _GEN_45077;
  wire  _GEN_45078;
  wire  _GEN_45079;
  wire  _GEN_45080;
  wire  _GEN_45081;
  wire  _GEN_45082;
  wire  _GEN_45083;
  wire  _GEN_45084;
  wire  _GEN_45085;
  wire  _GEN_45086;
  wire  _GEN_45087;
  wire  _GEN_45088;
  wire  _T_6349;
  wire  _T_6351;
  wire  _T_6353;
  wire [5:0] _T_6354;
  wire  _T_6355;
  wire  _T_6357;
  wire  _T_6359;
  wire  _GEN_45169;
  wire  _GEN_45170;
  wire  _GEN_45171;
  wire  _GEN_45172;
  wire  _GEN_45173;
  wire  _GEN_45174;
  wire  _GEN_45175;
  wire  _GEN_45176;
  wire  _GEN_45177;
  wire  _GEN_45178;
  wire  _GEN_45179;
  wire  _GEN_45180;
  wire  _GEN_45181;
  wire  _GEN_45182;
  wire  _GEN_45183;
  wire  _GEN_45184;
  wire  _GEN_45185;
  wire  _GEN_45186;
  wire  _GEN_45187;
  wire  _GEN_45188;
  wire  _GEN_45189;
  wire  _GEN_45190;
  wire  _GEN_45191;
  wire  _GEN_45192;
  wire  _GEN_45193;
  wire  _GEN_45194;
  wire  _GEN_45195;
  wire  _GEN_45196;
  wire  _GEN_45197;
  wire  _GEN_45198;
  wire  _GEN_45199;
  wire  _GEN_45200;
  wire  _GEN_45201;
  wire  _GEN_45202;
  wire  _GEN_45203;
  wire  _GEN_45204;
  wire  _GEN_45205;
  wire  _GEN_45206;
  wire  _GEN_45207;
  wire  _GEN_45208;
  wire [7:0] _GEN_46173;
  wire [7:0] _GEN_46174;
  wire [7:0] _GEN_46175;
  wire [7:0] _GEN_46176;
  wire [7:0] _GEN_46177;
  wire [7:0] _GEN_46178;
  wire [7:0] _GEN_46179;
  wire [7:0] _GEN_46180;
  wire [7:0] _GEN_46181;
  wire [7:0] _GEN_46182;
  wire [7:0] _GEN_46183;
  wire [7:0] _GEN_46184;
  wire [7:0] _GEN_46185;
  wire [7:0] _GEN_46186;
  wire [7:0] _GEN_46187;
  wire [7:0] _GEN_46188;
  wire [7:0] _GEN_46189;
  wire [7:0] _GEN_46190;
  wire [7:0] _GEN_46191;
  wire [7:0] _GEN_46192;
  wire [7:0] _GEN_46193;
  wire [7:0] _GEN_46194;
  wire [7:0] _GEN_46195;
  wire [7:0] _GEN_46196;
  wire [7:0] _GEN_46197;
  wire [7:0] _GEN_46198;
  wire [7:0] _GEN_46199;
  wire [7:0] _GEN_46200;
  wire [7:0] _GEN_46201;
  wire [7:0] _GEN_46202;
  wire [7:0] _GEN_46203;
  wire [7:0] _GEN_46204;
  wire [7:0] _GEN_46205;
  wire [7:0] _GEN_46206;
  wire [7:0] _GEN_46207;
  wire [7:0] _GEN_46208;
  wire [7:0] _GEN_46209;
  wire [7:0] _GEN_46210;
  wire [7:0] _GEN_46211;
  wire [7:0] _GEN_46212;
  wire [6:0] _GEN_47293;
  wire [6:0] _GEN_47294;
  wire [6:0] _GEN_47295;
  wire [6:0] _GEN_47296;
  wire [6:0] _GEN_47297;
  wire [6:0] _GEN_47298;
  wire [6:0] _GEN_47299;
  wire [6:0] _GEN_47300;
  wire [6:0] _GEN_47301;
  wire [6:0] _GEN_47302;
  wire [6:0] _GEN_47303;
  wire [6:0] _GEN_47304;
  wire [6:0] _GEN_47305;
  wire [6:0] _GEN_47306;
  wire [6:0] _GEN_47307;
  wire [6:0] _GEN_47308;
  wire [6:0] _GEN_47309;
  wire [6:0] _GEN_47310;
  wire [6:0] _GEN_47311;
  wire [6:0] _GEN_47312;
  wire [6:0] _GEN_47313;
  wire [6:0] _GEN_47314;
  wire [6:0] _GEN_47315;
  wire [6:0] _GEN_47316;
  wire [6:0] _GEN_47317;
  wire [6:0] _GEN_47318;
  wire [6:0] _GEN_47319;
  wire [6:0] _GEN_47320;
  wire [6:0] _GEN_47321;
  wire [6:0] _GEN_47322;
  wire [6:0] _GEN_47323;
  wire [6:0] _GEN_47324;
  wire [6:0] _GEN_47325;
  wire [6:0] _GEN_47326;
  wire [6:0] _GEN_47327;
  wire [6:0] _GEN_47328;
  wire [6:0] _GEN_47329;
  wire [6:0] _GEN_47330;
  wire [6:0] _GEN_47331;
  wire [6:0] _GEN_47332;
  wire [6:0] _GEN_47573;
  wire [6:0] _GEN_47574;
  wire [6:0] _GEN_47575;
  wire [6:0] _GEN_47576;
  wire [6:0] _GEN_47577;
  wire [6:0] _GEN_47578;
  wire [6:0] _GEN_47579;
  wire [6:0] _GEN_47580;
  wire [6:0] _GEN_47581;
  wire [6:0] _GEN_47582;
  wire [6:0] _GEN_47583;
  wire [6:0] _GEN_47584;
  wire [6:0] _GEN_47585;
  wire [6:0] _GEN_47586;
  wire [6:0] _GEN_47587;
  wire [6:0] _GEN_47588;
  wire [6:0] _GEN_47589;
  wire [6:0] _GEN_47590;
  wire [6:0] _GEN_47591;
  wire [6:0] _GEN_47592;
  wire [6:0] _GEN_47593;
  wire [6:0] _GEN_47594;
  wire [6:0] _GEN_47595;
  wire [6:0] _GEN_47596;
  wire [6:0] _GEN_47597;
  wire [6:0] _GEN_47598;
  wire [6:0] _GEN_47599;
  wire [6:0] _GEN_47600;
  wire [6:0] _GEN_47601;
  wire [6:0] _GEN_47602;
  wire [6:0] _GEN_47603;
  wire [6:0] _GEN_47604;
  wire [6:0] _GEN_47605;
  wire [6:0] _GEN_47606;
  wire [6:0] _GEN_47607;
  wire [6:0] _GEN_47608;
  wire [6:0] _GEN_47609;
  wire [6:0] _GEN_47610;
  wire [6:0] _GEN_47611;
  wire [6:0] _GEN_47612;
  wire  _GEN_47853;
  wire  _GEN_47854;
  wire  _GEN_47855;
  wire  _GEN_47856;
  wire  _GEN_47857;
  wire  _GEN_47858;
  wire  _GEN_47859;
  wire  _GEN_47860;
  wire  _GEN_47861;
  wire  _GEN_47862;
  wire  _GEN_47863;
  wire  _GEN_47864;
  wire  _GEN_47865;
  wire  _GEN_47866;
  wire  _GEN_47867;
  wire  _GEN_47868;
  wire  _GEN_47869;
  wire  _GEN_47870;
  wire  _GEN_47871;
  wire  _GEN_47872;
  wire  _GEN_47873;
  wire  _GEN_47874;
  wire  _GEN_47875;
  wire  _GEN_47876;
  wire  _GEN_47877;
  wire  _GEN_47878;
  wire  _GEN_47879;
  wire  _GEN_47880;
  wire  _GEN_47881;
  wire  _GEN_47882;
  wire  _GEN_47883;
  wire  _GEN_47884;
  wire  _GEN_47885;
  wire  _GEN_47886;
  wire  _GEN_47887;
  wire  _GEN_47888;
  wire  _GEN_47889;
  wire  _GEN_47890;
  wire  _GEN_47891;
  wire  _GEN_47892;
  wire  _GEN_47893;
  wire  _GEN_47894;
  wire  _GEN_47895;
  wire  _GEN_47896;
  wire  _GEN_47897;
  wire  _GEN_47898;
  wire  _GEN_47899;
  wire  _GEN_47900;
  wire  _GEN_47901;
  wire  _GEN_47902;
  wire  _GEN_47903;
  wire  _GEN_47904;
  wire  _GEN_47905;
  wire  _GEN_47906;
  wire  _GEN_47907;
  wire  _GEN_47908;
  wire  _GEN_47909;
  wire  _GEN_47910;
  wire  _GEN_47911;
  wire  _GEN_47912;
  wire  _GEN_47913;
  wire  _GEN_47914;
  wire  _GEN_47915;
  wire  _GEN_47916;
  wire  _GEN_47917;
  wire  _GEN_47918;
  wire  _GEN_47919;
  wire  _GEN_47920;
  wire  _GEN_47921;
  wire  _GEN_47922;
  wire  _GEN_47923;
  wire  _GEN_47924;
  wire  _GEN_47925;
  wire  _GEN_47926;
  wire  _GEN_47927;
  wire  _GEN_47928;
  wire  _GEN_47929;
  wire  _GEN_47930;
  wire  _GEN_47931;
  wire  _GEN_47932;
  wire  _GEN_47973;
  wire  _GEN_47974;
  wire  _GEN_47975;
  wire  _GEN_47976;
  wire  _GEN_47977;
  wire  _GEN_47978;
  wire  _GEN_47979;
  wire  _GEN_47980;
  wire  _GEN_47981;
  wire  _GEN_47982;
  wire  _GEN_47983;
  wire  _GEN_47984;
  wire  _GEN_47985;
  wire  _GEN_47986;
  wire  _GEN_47987;
  wire  _GEN_47988;
  wire  _GEN_47989;
  wire  _GEN_47990;
  wire  _GEN_47991;
  wire  _GEN_47992;
  wire  _GEN_47993;
  wire  _GEN_47994;
  wire  _GEN_47995;
  wire  _GEN_47996;
  wire  _GEN_47997;
  wire  _GEN_47998;
  wire  _GEN_47999;
  wire  _GEN_48000;
  wire  _GEN_48001;
  wire  _GEN_48002;
  wire  _GEN_48003;
  wire  _GEN_48004;
  wire  _GEN_48005;
  wire  _GEN_48006;
  wire  _GEN_48007;
  wire  _GEN_48008;
  wire  _GEN_48009;
  wire  _GEN_48010;
  wire  _GEN_48011;
  wire  _GEN_48012;
  wire  _GEN_48013;
  wire  _GEN_48014;
  wire  _GEN_48015;
  wire  _GEN_48016;
  wire  _GEN_48017;
  wire  _GEN_48018;
  wire  _GEN_48019;
  wire  _GEN_48020;
  wire  _GEN_48021;
  wire  _GEN_48022;
  wire  _GEN_48023;
  wire  _GEN_48024;
  wire  _GEN_48025;
  wire  _GEN_48026;
  wire  _GEN_48027;
  wire  _GEN_48028;
  wire  _GEN_48029;
  wire  _GEN_48030;
  wire  _GEN_48031;
  wire  _GEN_48032;
  wire  _GEN_48033;
  wire  _GEN_48034;
  wire  _GEN_48035;
  wire  _GEN_48036;
  wire  _GEN_48037;
  wire  _GEN_48038;
  wire  _GEN_48039;
  wire  _GEN_48040;
  wire  _GEN_48041;
  wire  _GEN_48042;
  wire  _GEN_48043;
  wire  _GEN_48044;
  wire  _GEN_48045;
  wire  _GEN_48046;
  wire  _GEN_48047;
  wire  _GEN_48048;
  wire  _GEN_48049;
  wire  _GEN_48050;
  wire  _GEN_48051;
  wire  _GEN_48052;
  wire  _GEN_48093;
  wire  _GEN_48094;
  wire  _GEN_48095;
  wire  _GEN_48096;
  wire  _GEN_48097;
  wire  _GEN_48098;
  wire  _GEN_48099;
  wire  _GEN_48100;
  wire  _GEN_48101;
  wire  _GEN_48102;
  wire  _GEN_48103;
  wire  _GEN_48104;
  wire  _GEN_48105;
  wire  _GEN_48106;
  wire  _GEN_48107;
  wire  _GEN_48108;
  wire  _GEN_48109;
  wire  _GEN_48110;
  wire  _GEN_48111;
  wire  _GEN_48112;
  wire  _GEN_48113;
  wire  _GEN_48114;
  wire  _GEN_48115;
  wire  _GEN_48116;
  wire  _GEN_48117;
  wire  _GEN_48118;
  wire  _GEN_48119;
  wire  _GEN_48120;
  wire  _GEN_48121;
  wire  _GEN_48122;
  wire  _GEN_48123;
  wire  _GEN_48124;
  wire  _GEN_48125;
  wire  _GEN_48126;
  wire  _GEN_48127;
  wire  _GEN_48128;
  wire  _GEN_48129;
  wire  _GEN_48130;
  wire  _GEN_48131;
  wire  _GEN_48132;
  wire [5:0] _GEN_48133;
  wire [5:0] _GEN_48134;
  wire [5:0] _GEN_48135;
  wire [5:0] _GEN_48136;
  wire [5:0] _GEN_48137;
  wire [5:0] _GEN_48138;
  wire [5:0] _GEN_48139;
  wire [5:0] _GEN_48140;
  wire [5:0] _GEN_48141;
  wire [5:0] _GEN_48142;
  wire [5:0] _GEN_48143;
  wire [5:0] _GEN_48144;
  wire [5:0] _GEN_48145;
  wire [5:0] _GEN_48146;
  wire [5:0] _GEN_48147;
  wire [5:0] _GEN_48148;
  wire [5:0] _GEN_48149;
  wire [5:0] _GEN_48150;
  wire [5:0] _GEN_48151;
  wire [5:0] _GEN_48152;
  wire [5:0] _GEN_48153;
  wire [5:0] _GEN_48154;
  wire [5:0] _GEN_48155;
  wire [5:0] _GEN_48156;
  wire [5:0] _GEN_48157;
  wire [5:0] _GEN_48158;
  wire [5:0] _GEN_48159;
  wire [5:0] _GEN_48160;
  wire [5:0] _GEN_48161;
  wire [5:0] _GEN_48162;
  wire [5:0] _GEN_48163;
  wire [5:0] _GEN_48164;
  wire [5:0] _GEN_48165;
  wire [5:0] _GEN_48166;
  wire [5:0] _GEN_48167;
  wire [5:0] _GEN_48168;
  wire [5:0] _GEN_48169;
  wire [5:0] _GEN_48170;
  wire [5:0] _GEN_48171;
  wire [5:0] _GEN_48172;
  wire  _GEN_48293;
  wire  _GEN_48294;
  wire  _GEN_48295;
  wire  _GEN_48296;
  wire  _GEN_48297;
  wire  _GEN_48298;
  wire  _GEN_48299;
  wire  _GEN_48300;
  wire  _GEN_48301;
  wire  _GEN_48302;
  wire  _GEN_48303;
  wire  _GEN_48304;
  wire  _GEN_48305;
  wire  _GEN_48306;
  wire  _GEN_48307;
  wire  _GEN_48308;
  wire  _GEN_48309;
  wire  _GEN_48310;
  wire  _GEN_48311;
  wire  _GEN_48312;
  wire  _GEN_48313;
  wire  _GEN_48314;
  wire  _GEN_48315;
  wire  _GEN_48316;
  wire  _GEN_48317;
  wire  _GEN_48318;
  wire  _GEN_48319;
  wire  _GEN_48320;
  wire  _GEN_48321;
  wire  _GEN_48322;
  wire  _GEN_48323;
  wire  _GEN_48324;
  wire  _GEN_48325;
  wire  _GEN_48326;
  wire  _GEN_48327;
  wire  _GEN_48328;
  wire  _GEN_48329;
  wire  _GEN_48330;
  wire  _GEN_48331;
  wire  _GEN_48332;
  wire [1:0] _GEN_48333;
  wire [1:0] _GEN_48334;
  wire [1:0] _GEN_48335;
  wire [1:0] _GEN_48336;
  wire [1:0] _GEN_48337;
  wire [1:0] _GEN_48338;
  wire [1:0] _GEN_48339;
  wire [1:0] _GEN_48340;
  wire [1:0] _GEN_48341;
  wire [1:0] _GEN_48342;
  wire [1:0] _GEN_48343;
  wire [1:0] _GEN_48344;
  wire [1:0] _GEN_48345;
  wire [1:0] _GEN_48346;
  wire [1:0] _GEN_48347;
  wire [1:0] _GEN_48348;
  wire [1:0] _GEN_48349;
  wire [1:0] _GEN_48350;
  wire [1:0] _GEN_48351;
  wire [1:0] _GEN_48352;
  wire [1:0] _GEN_48353;
  wire [1:0] _GEN_48354;
  wire [1:0] _GEN_48355;
  wire [1:0] _GEN_48356;
  wire [1:0] _GEN_48357;
  wire [1:0] _GEN_48358;
  wire [1:0] _GEN_48359;
  wire [1:0] _GEN_48360;
  wire [1:0] _GEN_48361;
  wire [1:0] _GEN_48362;
  wire [1:0] _GEN_48363;
  wire [1:0] _GEN_48364;
  wire [1:0] _GEN_48365;
  wire [1:0] _GEN_48366;
  wire [1:0] _GEN_48367;
  wire [1:0] _GEN_48368;
  wire [1:0] _GEN_48369;
  wire [1:0] _GEN_48370;
  wire [1:0] _GEN_48371;
  wire [1:0] _GEN_48372;
  wire  _GEN_48493;
  wire  _GEN_48494;
  wire  _GEN_48495;
  wire  _GEN_48496;
  wire  _GEN_48497;
  wire  _GEN_48498;
  wire  _GEN_48499;
  wire  _GEN_48500;
  wire  _GEN_48501;
  wire  _GEN_48502;
  wire  _GEN_48503;
  wire  _GEN_48504;
  wire  _GEN_48505;
  wire  _GEN_48506;
  wire  _GEN_48507;
  wire  _GEN_48508;
  wire  _GEN_48509;
  wire  _GEN_48510;
  wire  _GEN_48511;
  wire  _GEN_48512;
  wire  _GEN_48513;
  wire  _GEN_48514;
  wire  _GEN_48515;
  wire  _GEN_48516;
  wire  _GEN_48517;
  wire  _GEN_48518;
  wire  _GEN_48519;
  wire  _GEN_48520;
  wire  _GEN_48521;
  wire  _GEN_48522;
  wire  _GEN_48523;
  wire  _GEN_48524;
  wire  _GEN_48525;
  wire  _GEN_48526;
  wire  _GEN_48527;
  wire  _GEN_48528;
  wire  _GEN_48529;
  wire  _GEN_48530;
  wire  _GEN_48531;
  wire  _GEN_48532;
  wire  _T_6381;
  wire [5:0] _T_6382;
  wire  _T_6390;
  wire [5:0] _T_6391;
  wire  _T_6399;
  wire [5:0] _T_6400;
  wire  _T_6408;
  wire [5:0] _T_6409;
  wire  _T_6417;
  wire [5:0] _T_6418;
  wire  _T_6424;
  wire [5:0] _T_6427;
  wire  _GEN_323;
  wire  _GEN_48835;
  wire  _GEN_48836;
  wire  _GEN_48837;
  wire  _GEN_48838;
  wire  _GEN_48839;
  wire  _GEN_48840;
  wire  _GEN_48841;
  wire  _GEN_48842;
  wire  _GEN_48843;
  wire  _GEN_48844;
  wire  _GEN_48845;
  wire  _GEN_48846;
  wire  _GEN_48847;
  wire  _GEN_48848;
  wire  _GEN_48849;
  wire  _GEN_48850;
  wire  _GEN_48851;
  wire  _GEN_48852;
  wire  _GEN_48853;
  wire  _GEN_48854;
  wire  _GEN_48855;
  wire  _GEN_48856;
  wire  _GEN_48857;
  wire  _GEN_48858;
  wire  _GEN_48859;
  wire  _GEN_48860;
  wire  _GEN_48861;
  wire  _GEN_48862;
  wire  _GEN_48863;
  wire  _GEN_48864;
  wire  _GEN_48865;
  wire  _GEN_48866;
  wire  _GEN_48867;
  wire  _GEN_48868;
  wire  _GEN_48869;
  wire  _GEN_48870;
  wire  _GEN_48871;
  wire  _GEN_48872;
  wire  _GEN_48873;
  wire  _T_6437;
  wire  _T_6439;
  wire [5:0] _T_6440;
  wire  _T_6443;
  wire  _T_6445;
  wire  _T_6447;
  wire  _T_6451;
  wire [5:0] _T_6454;
  wire  _GEN_324;
  wire  _GEN_48879;
  wire  _GEN_48880;
  wire  _GEN_48881;
  wire  _GEN_48882;
  wire  _GEN_48883;
  wire  _GEN_48884;
  wire  _GEN_48885;
  wire  _GEN_48886;
  wire  _GEN_48887;
  wire  _GEN_48888;
  wire  _GEN_48889;
  wire  _GEN_48890;
  wire  _GEN_48891;
  wire  _GEN_48892;
  wire  _GEN_48893;
  wire  _GEN_48894;
  wire  _GEN_48895;
  wire  _GEN_48896;
  wire  _GEN_48897;
  wire  _GEN_48898;
  wire  _GEN_48899;
  wire  _GEN_48900;
  wire  _GEN_48901;
  wire  _GEN_48902;
  wire  _GEN_48903;
  wire  _GEN_48904;
  wire  _GEN_48905;
  wire  _GEN_48906;
  wire  _GEN_48907;
  wire  _GEN_48908;
  wire  _GEN_48909;
  wire  _GEN_48910;
  wire  _GEN_48911;
  wire  _GEN_48912;
  wire  _GEN_48913;
  wire  _GEN_48914;
  wire  _GEN_48915;
  wire  _GEN_48916;
  wire  _GEN_48917;
  wire  _T_6464;
  wire  _T_6466;
  wire [5:0] _T_6467;
  wire  _T_6470;
  wire  _T_6472;
  wire  _T_6474;
  wire  _T_6542;
  wire [5:0] _T_6545;
  wire  _T_6550;
  wire [5:0] _T_6553;
  wire  _T_6558;
  wire [5:0] _T_6561;
  wire  _T_6567;
  wire [5:0] _T_6570;
  wire  _GEN_330;
  wire  _GEN_49339;
  wire  _GEN_49340;
  wire  _GEN_49341;
  wire  _GEN_49342;
  wire  _GEN_49343;
  wire  _GEN_49344;
  wire  _GEN_49345;
  wire  _GEN_49346;
  wire  _GEN_49347;
  wire  _GEN_49348;
  wire  _GEN_49349;
  wire  _GEN_49350;
  wire  _GEN_49351;
  wire  _GEN_49352;
  wire  _GEN_49353;
  wire  _GEN_49354;
  wire  _GEN_49355;
  wire  _GEN_49356;
  wire  _GEN_49357;
  wire  _GEN_49358;
  wire  _GEN_49359;
  wire  _GEN_49360;
  wire  _GEN_49361;
  wire  _GEN_49362;
  wire  _GEN_49363;
  wire  _GEN_49364;
  wire  _GEN_49365;
  wire  _GEN_49366;
  wire  _GEN_49367;
  wire  _GEN_49368;
  wire  _GEN_49369;
  wire  _GEN_49370;
  wire  _GEN_49371;
  wire  _GEN_49372;
  wire  _GEN_49373;
  wire  _GEN_49374;
  wire  _GEN_49375;
  wire  _GEN_49376;
  wire  _GEN_49377;
  wire  _T_6577;
  wire  _T_6583;
  wire  _GEN_331;
  wire  _T_6584;
  wire  _T_6587;
  wire [5:0] _T_6589;
  wire [6:0] _GEN_49431;
  wire [6:0] _GEN_49438;
  wire  _GEN_49445;
  wire  _GEN_49446;
  wire  _GEN_49448;
  wire  _GEN_49449;
  wire  _GEN_49451;
  wire [5:0] _GEN_49452;
  wire [1:0] _GEN_49457;
  wire  _GEN_49461;
  wire [6:0] _GEN_49521;
  wire [6:0] _GEN_49528;
  wire  _GEN_49535;
  wire  _GEN_49536;
  wire  _GEN_49538;
  wire  _GEN_49539;
  wire  _GEN_49541;
  wire [5:0] _GEN_49542;
  wire [1:0] _GEN_49547;
  wire  _GEN_49551;
  wire [6:0] _GEN_49611;
  wire [6:0] _GEN_49618;
  wire  _GEN_49625;
  wire  _GEN_49626;
  wire  _GEN_49628;
  wire  _GEN_49629;
  wire  _GEN_49631;
  wire [5:0] _GEN_49632;
  wire [1:0] _GEN_49637;
  wire  _GEN_49641;
  wire [6:0] _GEN_49701;
  wire [6:0] _GEN_49708;
  wire  _GEN_49715;
  wire  _GEN_49716;
  wire  _GEN_49718;
  wire  _GEN_49719;
  wire  _GEN_49721;
  wire [5:0] _GEN_49722;
  wire [1:0] _GEN_49727;
  wire  _GEN_49731;
  wire [6:0] _GEN_49791;
  wire [6:0] _GEN_49798;
  wire  _GEN_49805;
  wire  _GEN_49806;
  wire  _GEN_49808;
  wire  _GEN_49809;
  wire  _GEN_49811;
  wire [5:0] _GEN_49812;
  wire [1:0] _GEN_49817;
  wire  _GEN_49821;
  wire [6:0] _GEN_49881;
  wire [6:0] _GEN_49888;
  wire  _GEN_49895;
  wire  _GEN_49896;
  wire  _GEN_49898;
  wire  _GEN_49899;
  wire  _GEN_49901;
  wire [5:0] _GEN_49902;
  wire [1:0] _GEN_49907;
  wire  _GEN_49911;
  wire [6:0] _GEN_49971;
  wire [6:0] _GEN_49978;
  wire  _GEN_49985;
  wire  _GEN_49986;
  wire  _GEN_49988;
  wire  _GEN_49989;
  wire  _GEN_49991;
  wire [5:0] _GEN_49992;
  wire [1:0] _GEN_49997;
  wire  _GEN_50001;
  wire [6:0] _GEN_50061;
  wire [6:0] _GEN_50068;
  wire  _GEN_50075;
  wire  _GEN_50076;
  wire  _GEN_50078;
  wire  _GEN_50079;
  wire  _GEN_50081;
  wire [5:0] _GEN_50082;
  wire [1:0] _GEN_50087;
  wire  _GEN_50091;
  wire [6:0] _GEN_50151;
  wire [6:0] _GEN_50158;
  wire  _GEN_50165;
  wire  _GEN_50166;
  wire  _GEN_50168;
  wire  _GEN_50169;
  wire  _GEN_50171;
  wire [5:0] _GEN_50172;
  wire [1:0] _GEN_50177;
  wire  _GEN_50181;
  wire [6:0] _GEN_50241;
  wire [6:0] _GEN_50248;
  wire  _GEN_50255;
  wire  _GEN_50256;
  wire  _GEN_50258;
  wire  _GEN_50259;
  wire  _GEN_50261;
  wire [5:0] _GEN_50262;
  wire [1:0] _GEN_50267;
  wire  _GEN_50271;
  wire [6:0] _GEN_50331;
  wire [6:0] _GEN_50338;
  wire  _GEN_50345;
  wire  _GEN_50346;
  wire  _GEN_50348;
  wire  _GEN_50349;
  wire  _GEN_50351;
  wire [5:0] _GEN_50352;
  wire [1:0] _GEN_50357;
  wire  _GEN_50361;
  wire [6:0] _GEN_50421;
  wire [6:0] _GEN_50428;
  wire  _GEN_50435;
  wire  _GEN_50436;
  wire  _GEN_50438;
  wire  _GEN_50439;
  wire  _GEN_50441;
  wire [5:0] _GEN_50442;
  wire [1:0] _GEN_50447;
  wire  _GEN_50451;
  wire [6:0] _GEN_50511;
  wire [6:0] _GEN_50518;
  wire  _GEN_50525;
  wire  _GEN_50526;
  wire  _GEN_50528;
  wire  _GEN_50529;
  wire  _GEN_50531;
  wire [5:0] _GEN_50532;
  wire [1:0] _GEN_50537;
  wire  _GEN_50541;
  wire [6:0] _GEN_50601;
  wire [6:0] _GEN_50608;
  wire  _GEN_50615;
  wire  _GEN_50616;
  wire  _GEN_50618;
  wire  _GEN_50619;
  wire  _GEN_50621;
  wire [5:0] _GEN_50622;
  wire [1:0] _GEN_50627;
  wire  _GEN_50631;
  wire [6:0] _GEN_50691;
  wire [6:0] _GEN_50698;
  wire  _GEN_50705;
  wire  _GEN_50706;
  wire  _GEN_50708;
  wire  _GEN_50709;
  wire  _GEN_50711;
  wire [5:0] _GEN_50712;
  wire [1:0] _GEN_50717;
  wire  _GEN_50721;
  wire [6:0] _GEN_50781;
  wire [6:0] _GEN_50788;
  wire  _GEN_50795;
  wire  _GEN_50796;
  wire  _GEN_50798;
  wire  _GEN_50799;
  wire  _GEN_50801;
  wire [5:0] _GEN_50802;
  wire [1:0] _GEN_50807;
  wire  _GEN_50811;
  wire [6:0] _GEN_50871;
  wire [6:0] _GEN_50878;
  wire  _GEN_50885;
  wire  _GEN_50886;
  wire  _GEN_50888;
  wire  _GEN_50889;
  wire  _GEN_50891;
  wire [5:0] _GEN_50892;
  wire [1:0] _GEN_50897;
  wire  _GEN_50901;
  wire [6:0] _GEN_50961;
  wire [6:0] _GEN_50968;
  wire  _GEN_50975;
  wire  _GEN_50976;
  wire  _GEN_50978;
  wire  _GEN_50979;
  wire  _GEN_50981;
  wire [5:0] _GEN_50982;
  wire [1:0] _GEN_50987;
  wire  _GEN_50991;
  wire [6:0] _GEN_51051;
  wire [6:0] _GEN_51058;
  wire  _GEN_51065;
  wire  _GEN_51066;
  wire  _GEN_51068;
  wire  _GEN_51069;
  wire  _GEN_51071;
  wire [5:0] _GEN_51072;
  wire [1:0] _GEN_51077;
  wire  _GEN_51081;
  wire [6:0] _GEN_51141;
  wire [6:0] _GEN_51148;
  wire  _GEN_51155;
  wire  _GEN_51156;
  wire  _GEN_51158;
  wire  _GEN_51159;
  wire  _GEN_51161;
  wire [5:0] _GEN_51162;
  wire [1:0] _GEN_51167;
  wire  _GEN_51171;
  wire [6:0] _GEN_51231;
  wire [6:0] _GEN_51238;
  wire  _GEN_51245;
  wire  _GEN_51246;
  wire  _GEN_51248;
  wire  _GEN_51249;
  wire  _GEN_51251;
  wire [5:0] _GEN_51252;
  wire [1:0] _GEN_51257;
  wire  _GEN_51261;
  wire [6:0] _GEN_51321;
  wire [6:0] _GEN_51328;
  wire  _GEN_51335;
  wire  _GEN_51336;
  wire  _GEN_51338;
  wire  _GEN_51339;
  wire  _GEN_51341;
  wire [5:0] _GEN_51342;
  wire [1:0] _GEN_51347;
  wire  _GEN_51351;
  wire [6:0] _GEN_51411;
  wire [6:0] _GEN_51418;
  wire  _GEN_51425;
  wire  _GEN_51426;
  wire  _GEN_51428;
  wire  _GEN_51429;
  wire  _GEN_51431;
  wire [5:0] _GEN_51432;
  wire [1:0] _GEN_51437;
  wire  _GEN_51441;
  wire [6:0] _GEN_51501;
  wire [6:0] _GEN_51508;
  wire  _GEN_51515;
  wire  _GEN_51516;
  wire  _GEN_51518;
  wire  _GEN_51519;
  wire  _GEN_51521;
  wire [5:0] _GEN_51522;
  wire [1:0] _GEN_51527;
  wire  _GEN_51531;
  wire [6:0] _GEN_51591;
  wire [6:0] _GEN_51598;
  wire  _GEN_51605;
  wire  _GEN_51606;
  wire  _GEN_51608;
  wire  _GEN_51609;
  wire  _GEN_51611;
  wire [5:0] _GEN_51612;
  wire [1:0] _GEN_51617;
  wire  _GEN_51621;
  wire [6:0] _GEN_51681;
  wire [6:0] _GEN_51688;
  wire  _GEN_51695;
  wire  _GEN_51696;
  wire  _GEN_51698;
  wire  _GEN_51699;
  wire  _GEN_51701;
  wire [5:0] _GEN_51702;
  wire [1:0] _GEN_51707;
  wire  _GEN_51711;
  wire [6:0] _GEN_51771;
  wire [6:0] _GEN_51778;
  wire  _GEN_51785;
  wire  _GEN_51786;
  wire  _GEN_51788;
  wire  _GEN_51789;
  wire  _GEN_51791;
  wire [5:0] _GEN_51792;
  wire [1:0] _GEN_51797;
  wire  _GEN_51801;
  wire [6:0] _GEN_51861;
  wire [6:0] _GEN_51868;
  wire  _GEN_51875;
  wire  _GEN_51876;
  wire  _GEN_51878;
  wire  _GEN_51879;
  wire  _GEN_51881;
  wire [5:0] _GEN_51882;
  wire [1:0] _GEN_51887;
  wire  _GEN_51891;
  wire [6:0] _GEN_51951;
  wire [6:0] _GEN_51958;
  wire  _GEN_51965;
  wire  _GEN_51966;
  wire  _GEN_51968;
  wire  _GEN_51969;
  wire  _GEN_51971;
  wire [5:0] _GEN_51972;
  wire [1:0] _GEN_51977;
  wire  _GEN_51981;
  wire [6:0] _GEN_52041;
  wire [6:0] _GEN_52048;
  wire  _GEN_52055;
  wire  _GEN_52056;
  wire  _GEN_52058;
  wire  _GEN_52059;
  wire  _GEN_52061;
  wire [5:0] _GEN_52062;
  wire [1:0] _GEN_52067;
  wire  _GEN_52071;
  wire [6:0] _GEN_52131;
  wire [6:0] _GEN_52138;
  wire  _GEN_52145;
  wire  _GEN_52146;
  wire  _GEN_52148;
  wire  _GEN_52149;
  wire  _GEN_52151;
  wire [5:0] _GEN_52152;
  wire [1:0] _GEN_52157;
  wire  _GEN_52161;
  wire [6:0] _GEN_52221;
  wire [6:0] _GEN_52228;
  wire  _GEN_52235;
  wire  _GEN_52236;
  wire  _GEN_52238;
  wire  _GEN_52239;
  wire  _GEN_52241;
  wire [5:0] _GEN_52242;
  wire [1:0] _GEN_52247;
  wire  _GEN_52251;
  wire [6:0] _GEN_52311;
  wire [6:0] _GEN_52318;
  wire  _GEN_52325;
  wire  _GEN_52326;
  wire  _GEN_52328;
  wire  _GEN_52329;
  wire  _GEN_52331;
  wire [5:0] _GEN_52332;
  wire [1:0] _GEN_52337;
  wire  _GEN_52341;
  wire [6:0] _GEN_52401;
  wire [6:0] _GEN_52408;
  wire  _GEN_52415;
  wire  _GEN_52416;
  wire  _GEN_52418;
  wire  _GEN_52419;
  wire  _GEN_52421;
  wire [5:0] _GEN_52422;
  wire [1:0] _GEN_52427;
  wire  _GEN_52431;
  wire [6:0] _GEN_52491;
  wire [6:0] _GEN_52498;
  wire  _GEN_52505;
  wire  _GEN_52506;
  wire  _GEN_52508;
  wire  _GEN_52509;
  wire  _GEN_52511;
  wire [5:0] _GEN_52512;
  wire [1:0] _GEN_52517;
  wire  _GEN_52521;
  wire [6:0] _GEN_52581;
  wire [6:0] _GEN_52588;
  wire  _GEN_52595;
  wire  _GEN_52596;
  wire  _GEN_52598;
  wire  _GEN_52599;
  wire  _GEN_52601;
  wire [5:0] _GEN_52602;
  wire [1:0] _GEN_52607;
  wire  _GEN_52611;
  wire [6:0] _GEN_52671;
  wire [6:0] _GEN_52678;
  wire  _GEN_52685;
  wire  _GEN_52686;
  wire  _GEN_52688;
  wire  _GEN_52689;
  wire  _GEN_52691;
  wire [5:0] _GEN_52692;
  wire [1:0] _GEN_52697;
  wire  _GEN_52701;
  wire [6:0] _GEN_52761;
  wire [6:0] _GEN_52768;
  wire  _GEN_52775;
  wire  _GEN_52776;
  wire  _GEN_52778;
  wire  _GEN_52779;
  wire  _GEN_52781;
  wire [5:0] _GEN_52782;
  wire [1:0] _GEN_52787;
  wire  _GEN_52791;
  wire [6:0] _GEN_52851;
  wire [6:0] _GEN_52858;
  wire  _GEN_52865;
  wire  _GEN_52866;
  wire  _GEN_52868;
  wire  _GEN_52869;
  wire  _GEN_52871;
  wire [5:0] _GEN_52872;
  wire [1:0] _GEN_52877;
  wire  _GEN_52881;
  wire [6:0] _GEN_384_pdst;
  wire [6:0] _GEN_391_stale_pdst;
  wire  _GEN_398_is_fencei;
  wire  _GEN_399_is_store;
  wire  _GEN_401_is_load;
  wire  _GEN_402_is_sys_pc2epc;
  wire  _GEN_404_flush_on_commit;
  wire [5:0] _GEN_405_ldst;
  wire [1:0] _GEN_410_dst_rtype;
  wire  _GEN_414_fp_val;
  wire  _GEN_422;
  wire  _GEN_52889;
  wire  _GEN_52890;
  wire  _GEN_52891;
  wire  _GEN_52892;
  wire  _GEN_52893;
  wire  _GEN_52894;
  wire  _GEN_52895;
  wire  _GEN_52896;
  wire  _GEN_52897;
  wire  _GEN_52898;
  wire  _GEN_52899;
  wire  _GEN_52900;
  wire  _GEN_52901;
  wire  _GEN_52902;
  wire  _GEN_52903;
  wire  _GEN_52904;
  wire  _GEN_52905;
  wire  _GEN_52906;
  wire  _GEN_52907;
  wire  _GEN_52908;
  wire  _GEN_52909;
  wire  _GEN_52910;
  wire  _GEN_52911;
  wire  _GEN_52912;
  wire  _GEN_52913;
  wire  _GEN_52914;
  wire  _GEN_52915;
  wire  _GEN_52916;
  wire  _GEN_52917;
  wire  _GEN_52918;
  wire  _GEN_52919;
  wire  _GEN_52920;
  wire  _GEN_52921;
  wire  _GEN_52922;
  wire  _GEN_52923;
  wire  _GEN_52924;
  wire  _GEN_52925;
  wire  _GEN_52926;
  wire  _GEN_52927;
  wire  _T_6610;
  wire [1:0] _GEN_423_dst_rtype;
  wire  _T_6623;
  wire [1:0] _GEN_424_dst_rtype;
  wire  _T_6636;
  wire  _T_6637;
  wire  _T_6638;
  wire  _T_6641;
  wire  _GEN_59948;
  wire  _GEN_59949;
  wire  _GEN_59950;
  wire  _GEN_59951;
  wire  _GEN_59952;
  wire  _GEN_59953;
  wire  _GEN_59954;
  wire  _GEN_59955;
  wire  _GEN_59956;
  wire  _GEN_59957;
  wire  _GEN_59958;
  wire  _GEN_59959;
  wire  _GEN_59960;
  wire  _GEN_59961;
  wire  _GEN_59962;
  wire  _GEN_59963;
  wire  _GEN_59964;
  wire  _GEN_59965;
  wire  _GEN_59966;
  wire  _GEN_59967;
  wire  _GEN_59968;
  wire  _GEN_59969;
  wire  _GEN_59970;
  wire  _GEN_59971;
  wire  _GEN_59972;
  wire  _GEN_59973;
  wire  _GEN_59974;
  wire  _GEN_59975;
  wire  _GEN_59976;
  wire  _GEN_59977;
  wire  _GEN_59978;
  wire  _GEN_59979;
  wire  _GEN_59980;
  wire  _GEN_59981;
  wire  _GEN_59982;
  wire  _GEN_59983;
  wire  _GEN_59984;
  wire  _GEN_59985;
  wire  _GEN_59986;
  wire  _GEN_59987;
  wire  _GEN_59988;
  wire  _GEN_59989;
  wire  _GEN_59990;
  wire  _GEN_59991;
  wire  _GEN_59992;
  wire  _GEN_59993;
  wire  _GEN_59994;
  wire  _GEN_59995;
  wire  _GEN_59996;
  wire  _GEN_59997;
  wire  _GEN_59998;
  wire  _GEN_59999;
  wire  _GEN_60000;
  wire  _GEN_60001;
  wire  _GEN_60002;
  wire  _GEN_60003;
  wire  _GEN_60004;
  wire  _GEN_60005;
  wire  _GEN_60006;
  wire  _GEN_60007;
  wire  _GEN_60008;
  wire  _GEN_60009;
  wire  _GEN_60010;
  wire  _GEN_60011;
  wire  _GEN_60012;
  wire  _GEN_60013;
  wire  _GEN_60014;
  wire  _GEN_60015;
  wire  _GEN_60016;
  wire  _GEN_60017;
  wire  _GEN_60018;
  wire  _GEN_60019;
  wire  _GEN_60020;
  wire  _GEN_60021;
  wire  _GEN_60022;
  wire  _GEN_60023;
  wire  _GEN_60024;
  wire  _GEN_60025;
  wire  _GEN_60026;
  wire  _GEN_60027;
  wire [7:0] _T_6654;
  wire  _T_6656;
  wire  _T_6657;
  wire  _T_6659;
  wire  _T_6674;
  wire [7:0] _T_6676;
  wire [7:0] _GEN_60032;
  wire  _GEN_60033;
  wire [7:0] _GEN_60035;
  wire [7:0] _T_6677;
  wire  _T_6679;
  wire  _T_6680;
  wire  _T_6682;
  wire  _T_6697;
  wire [7:0] _T_6699;
  wire [7:0] _GEN_60036;
  wire  _GEN_60037;
  wire [7:0] _GEN_60039;
  wire [7:0] _T_6700;
  wire  _T_6702;
  wire  _T_6703;
  wire  _T_6705;
  wire  _T_6720;
  wire [7:0] _T_6722;
  wire [7:0] _GEN_60040;
  wire  _GEN_60041;
  wire [7:0] _GEN_60043;
  wire [7:0] _T_6723;
  wire  _T_6725;
  wire  _T_6726;
  wire  _T_6728;
  wire  _T_6743;
  wire [7:0] _T_6745;
  wire [7:0] _GEN_60044;
  wire  _GEN_60045;
  wire [7:0] _GEN_60047;
  wire [7:0] _T_6746;
  wire  _T_6748;
  wire  _T_6749;
  wire  _T_6751;
  wire  _T_6766;
  wire [7:0] _T_6768;
  wire [7:0] _GEN_60048;
  wire  _GEN_60049;
  wire [7:0] _GEN_60051;
  wire [7:0] _T_6769;
  wire  _T_6771;
  wire  _T_6772;
  wire  _T_6774;
  wire  _T_6789;
  wire [7:0] _T_6791;
  wire [7:0] _GEN_60052;
  wire  _GEN_60053;
  wire [7:0] _GEN_60055;
  wire [7:0] _T_6792;
  wire  _T_6794;
  wire  _T_6795;
  wire  _T_6797;
  wire  _T_6812;
  wire [7:0] _T_6814;
  wire [7:0] _GEN_60056;
  wire  _GEN_60057;
  wire [7:0] _GEN_60059;
  wire [7:0] _T_6815;
  wire  _T_6817;
  wire  _T_6818;
  wire  _T_6820;
  wire  _T_6835;
  wire [7:0] _T_6837;
  wire [7:0] _GEN_60060;
  wire  _GEN_60061;
  wire [7:0] _GEN_60063;
  wire [7:0] _T_6838;
  wire  _T_6840;
  wire  _T_6841;
  wire  _T_6843;
  wire  _T_6858;
  wire [7:0] _T_6860;
  wire [7:0] _GEN_60064;
  wire  _GEN_60065;
  wire [7:0] _GEN_60067;
  wire [7:0] _T_6861;
  wire  _T_6863;
  wire  _T_6864;
  wire  _T_6866;
  wire  _T_6881;
  wire [7:0] _T_6883;
  wire [7:0] _GEN_60068;
  wire  _GEN_60069;
  wire [7:0] _GEN_60071;
  wire [7:0] _T_6884;
  wire  _T_6886;
  wire  _T_6887;
  wire  _T_6889;
  wire  _T_6904;
  wire [7:0] _T_6906;
  wire [7:0] _GEN_60072;
  wire  _GEN_60073;
  wire [7:0] _GEN_60075;
  wire [7:0] _T_6907;
  wire  _T_6909;
  wire  _T_6910;
  wire  _T_6912;
  wire  _T_6927;
  wire [7:0] _T_6929;
  wire [7:0] _GEN_60076;
  wire  _GEN_60077;
  wire [7:0] _GEN_60079;
  wire [7:0] _T_6930;
  wire  _T_6932;
  wire  _T_6933;
  wire  _T_6935;
  wire  _T_6950;
  wire [7:0] _T_6952;
  wire [7:0] _GEN_60080;
  wire  _GEN_60081;
  wire [7:0] _GEN_60083;
  wire [7:0] _T_6953;
  wire  _T_6955;
  wire  _T_6956;
  wire  _T_6958;
  wire  _T_6973;
  wire [7:0] _T_6975;
  wire [7:0] _GEN_60084;
  wire  _GEN_60085;
  wire [7:0] _GEN_60087;
  wire [7:0] _T_6976;
  wire  _T_6978;
  wire  _T_6979;
  wire  _T_6981;
  wire  _T_6996;
  wire [7:0] _T_6998;
  wire [7:0] _GEN_60088;
  wire  _GEN_60089;
  wire [7:0] _GEN_60091;
  wire [7:0] _T_6999;
  wire  _T_7001;
  wire  _T_7002;
  wire  _T_7004;
  wire  _T_7019;
  wire [7:0] _T_7021;
  wire [7:0] _GEN_60092;
  wire  _GEN_60093;
  wire [7:0] _GEN_60095;
  wire [7:0] _T_7022;
  wire  _T_7024;
  wire  _T_7025;
  wire  _T_7027;
  wire  _T_7042;
  wire [7:0] _T_7044;
  wire [7:0] _GEN_60096;
  wire  _GEN_60097;
  wire [7:0] _GEN_60099;
  wire [7:0] _T_7045;
  wire  _T_7047;
  wire  _T_7048;
  wire  _T_7050;
  wire  _T_7065;
  wire [7:0] _T_7067;
  wire [7:0] _GEN_60100;
  wire  _GEN_60101;
  wire [7:0] _GEN_60103;
  wire [7:0] _T_7068;
  wire  _T_7070;
  wire  _T_7071;
  wire  _T_7073;
  wire  _T_7088;
  wire [7:0] _T_7090;
  wire [7:0] _GEN_60104;
  wire  _GEN_60105;
  wire [7:0] _GEN_60107;
  wire [7:0] _T_7091;
  wire  _T_7093;
  wire  _T_7094;
  wire  _T_7096;
  wire  _T_7111;
  wire [7:0] _T_7113;
  wire [7:0] _GEN_60108;
  wire  _GEN_60109;
  wire [7:0] _GEN_60111;
  wire [7:0] _T_7114;
  wire  _T_7116;
  wire  _T_7117;
  wire  _T_7119;
  wire  _T_7134;
  wire [7:0] _T_7136;
  wire [7:0] _GEN_60112;
  wire  _GEN_60113;
  wire [7:0] _GEN_60115;
  wire [7:0] _T_7137;
  wire  _T_7139;
  wire  _T_7140;
  wire  _T_7142;
  wire  _T_7157;
  wire [7:0] _T_7159;
  wire [7:0] _GEN_60116;
  wire  _GEN_60117;
  wire [7:0] _GEN_60119;
  wire [7:0] _T_7160;
  wire  _T_7162;
  wire  _T_7163;
  wire  _T_7165;
  wire  _T_7180;
  wire [7:0] _T_7182;
  wire [7:0] _GEN_60120;
  wire  _GEN_60121;
  wire [7:0] _GEN_60123;
  wire [7:0] _T_7183;
  wire  _T_7185;
  wire  _T_7186;
  wire  _T_7188;
  wire  _T_7203;
  wire [7:0] _T_7205;
  wire [7:0] _GEN_60124;
  wire  _GEN_60125;
  wire [7:0] _GEN_60127;
  wire [7:0] _T_7206;
  wire  _T_7208;
  wire  _T_7209;
  wire  _T_7211;
  wire  _T_7226;
  wire [7:0] _T_7228;
  wire [7:0] _GEN_60128;
  wire  _GEN_60129;
  wire [7:0] _GEN_60131;
  wire [7:0] _T_7229;
  wire  _T_7231;
  wire  _T_7232;
  wire  _T_7234;
  wire  _T_7249;
  wire [7:0] _T_7251;
  wire [7:0] _GEN_60132;
  wire  _GEN_60133;
  wire [7:0] _GEN_60135;
  wire [7:0] _T_7252;
  wire  _T_7254;
  wire  _T_7255;
  wire  _T_7257;
  wire  _T_7272;
  wire [7:0] _T_7274;
  wire [7:0] _GEN_60136;
  wire  _GEN_60137;
  wire [7:0] _GEN_60139;
  wire [7:0] _T_7275;
  wire  _T_7277;
  wire  _T_7278;
  wire  _T_7280;
  wire  _T_7295;
  wire [7:0] _T_7297;
  wire [7:0] _GEN_60140;
  wire  _GEN_60141;
  wire [7:0] _GEN_60143;
  wire [7:0] _T_7298;
  wire  _T_7300;
  wire  _T_7301;
  wire  _T_7303;
  wire  _T_7318;
  wire [7:0] _T_7320;
  wire [7:0] _GEN_60144;
  wire  _GEN_60145;
  wire [7:0] _GEN_60147;
  wire [7:0] _T_7321;
  wire  _T_7323;
  wire  _T_7324;
  wire  _T_7326;
  wire  _T_7341;
  wire [7:0] _T_7343;
  wire [7:0] _GEN_60148;
  wire  _GEN_60149;
  wire [7:0] _GEN_60151;
  wire [7:0] _T_7344;
  wire  _T_7346;
  wire  _T_7347;
  wire  _T_7349;
  wire  _T_7364;
  wire [7:0] _T_7366;
  wire [7:0] _GEN_60152;
  wire  _GEN_60153;
  wire [7:0] _GEN_60155;
  wire [7:0] _T_7367;
  wire  _T_7369;
  wire  _T_7370;
  wire  _T_7372;
  wire  _T_7387;
  wire [7:0] _T_7389;
  wire [7:0] _GEN_60156;
  wire  _GEN_60157;
  wire [7:0] _GEN_60159;
  wire [7:0] _T_7390;
  wire  _T_7392;
  wire  _T_7393;
  wire  _T_7395;
  wire  _T_7410;
  wire [7:0] _T_7412;
  wire [7:0] _GEN_60160;
  wire  _GEN_60161;
  wire [7:0] _GEN_60163;
  wire [7:0] _T_7413;
  wire  _T_7415;
  wire  _T_7416;
  wire  _T_7418;
  wire  _T_7433;
  wire [7:0] _T_7435;
  wire [7:0] _GEN_60164;
  wire  _GEN_60165;
  wire [7:0] _GEN_60167;
  wire [7:0] _T_7436;
  wire  _T_7438;
  wire  _T_7439;
  wire  _T_7441;
  wire  _T_7456;
  wire [7:0] _T_7458;
  wire [7:0] _GEN_60168;
  wire  _GEN_60169;
  wire [7:0] _GEN_60171;
  wire [7:0] _T_7459;
  wire  _T_7461;
  wire  _T_7462;
  wire  _T_7464;
  wire  _T_7479;
  wire [7:0] _T_7481;
  wire [7:0] _GEN_60172;
  wire  _GEN_60173;
  wire [7:0] _GEN_60175;
  wire [7:0] _T_7482;
  wire  _T_7484;
  wire  _T_7485;
  wire  _T_7487;
  wire  _T_7502;
  wire [7:0] _T_7504;
  wire [7:0] _GEN_60176;
  wire  _GEN_60177;
  wire [7:0] _GEN_60179;
  wire [7:0] _T_7505;
  wire  _T_7507;
  wire  _T_7508;
  wire  _T_7510;
  wire  _T_7525;
  wire [7:0] _T_7527;
  wire [7:0] _GEN_60180;
  wire  _GEN_60181;
  wire [7:0] _GEN_60183;
  wire [7:0] _T_7528;
  wire  _T_7530;
  wire  _T_7531;
  wire  _T_7533;
  wire  _T_7548;
  wire [7:0] _T_7550;
  wire [7:0] _GEN_60184;
  wire  _GEN_60185;
  wire [7:0] _GEN_60187;
  wire [7:0] _T_7551;
  wire  _T_7553;
  wire  _T_7554;
  wire  _T_7556;
  wire  _T_7571;
  wire [7:0] _T_7573;
  wire [7:0] _GEN_60188;
  wire  _GEN_60189;
  wire [7:0] _GEN_60191;
  wire  _GEN_60192;
  wire  _GEN_60193;
  wire  _GEN_60194;
  wire  _GEN_60195;
  wire  _GEN_60196;
  wire  _GEN_60197;
  wire  _GEN_60198;
  wire  _GEN_60199;
  wire  _GEN_60200;
  wire  _GEN_60201;
  wire  _GEN_60202;
  wire  _GEN_60203;
  wire  _GEN_60204;
  wire  _GEN_60205;
  wire  _GEN_60206;
  wire  _GEN_60207;
  wire  _GEN_60208;
  wire  _GEN_60209;
  wire  _GEN_60210;
  wire  _GEN_60211;
  wire  _GEN_60212;
  wire  _GEN_60213;
  wire  _GEN_60214;
  wire  _GEN_60215;
  wire  _GEN_60216;
  wire  _GEN_60217;
  wire  _GEN_60218;
  wire  _GEN_60219;
  wire  _GEN_60220;
  wire  _GEN_60221;
  wire  _GEN_60222;
  wire  _GEN_60223;
  wire  _GEN_60224;
  wire  _GEN_60225;
  wire  _GEN_60226;
  wire  _GEN_60227;
  wire  _GEN_60228;
  wire  _GEN_60229;
  wire  _GEN_60230;
  wire  _GEN_60231;
  wire  _GEN_60232;
  wire  _GEN_60233;
  wire  _GEN_60234;
  wire  _GEN_60235;
  wire  _GEN_60236;
  wire  _GEN_60237;
  wire  _GEN_60238;
  wire  _GEN_60239;
  wire  _GEN_60240;
  wire  _GEN_60241;
  wire  _GEN_60242;
  wire  _GEN_60243;
  wire  _GEN_60244;
  wire  _GEN_60245;
  wire  _GEN_60246;
  wire  _GEN_60247;
  wire  _GEN_60248;
  wire  _GEN_60249;
  wire  _GEN_60250;
  wire  _GEN_60251;
  wire  _GEN_60252;
  wire  _GEN_60253;
  wire  _GEN_60254;
  wire  _GEN_60255;
  wire  _GEN_60256;
  wire  _GEN_60257;
  wire  _GEN_60258;
  wire  _GEN_60259;
  wire  _GEN_60260;
  wire  _GEN_60261;
  wire  _GEN_60262;
  wire  _GEN_60263;
  wire  _GEN_60264;
  wire  _GEN_60265;
  wire  _GEN_60266;
  wire  _GEN_60267;
  wire  _GEN_60268;
  wire  _GEN_60269;
  wire  _GEN_60270;
  wire  _GEN_60271;
  wire  _GEN_427;
  wire  _GEN_428_is_store;
  wire  _GEN_60339;
  wire  _GEN_60341;
  wire  _GEN_60429;
  wire  _GEN_60431;
  wire  _GEN_60519;
  wire  _GEN_60521;
  wire  _GEN_60609;
  wire  _GEN_60611;
  wire  _GEN_60699;
  wire  _GEN_60701;
  wire  _GEN_60789;
  wire  _GEN_60791;
  wire  _GEN_60879;
  wire  _GEN_60881;
  wire  _GEN_60969;
  wire  _GEN_60971;
  wire  _GEN_61059;
  wire  _GEN_61061;
  wire  _GEN_61149;
  wire  _GEN_61151;
  wire  _GEN_61239;
  wire  _GEN_61241;
  wire  _GEN_61329;
  wire  _GEN_61331;
  wire  _GEN_61419;
  wire  _GEN_61421;
  wire  _GEN_61509;
  wire  _GEN_61511;
  wire  _GEN_61599;
  wire  _GEN_61601;
  wire  _GEN_61689;
  wire  _GEN_61691;
  wire  _GEN_61779;
  wire  _GEN_61781;
  wire  _GEN_61869;
  wire  _GEN_61871;
  wire  _GEN_61959;
  wire  _GEN_61961;
  wire  _GEN_62049;
  wire  _GEN_62051;
  wire  _GEN_62139;
  wire  _GEN_62141;
  wire  _GEN_62229;
  wire  _GEN_62231;
  wire  _GEN_62319;
  wire  _GEN_62321;
  wire  _GEN_62409;
  wire  _GEN_62411;
  wire  _GEN_62499;
  wire  _GEN_62501;
  wire  _GEN_62589;
  wire  _GEN_62591;
  wire  _GEN_62679;
  wire  _GEN_62681;
  wire  _GEN_62769;
  wire  _GEN_62771;
  wire  _GEN_62859;
  wire  _GEN_62861;
  wire  _GEN_62949;
  wire  _GEN_62951;
  wire  _GEN_63039;
  wire  _GEN_63041;
  wire  _GEN_63129;
  wire  _GEN_63131;
  wire  _GEN_63219;
  wire  _GEN_63221;
  wire  _GEN_63309;
  wire  _GEN_63311;
  wire  _GEN_63399;
  wire  _GEN_63401;
  wire  _GEN_63489;
  wire  _GEN_63491;
  wire  _GEN_63579;
  wire  _GEN_63581;
  wire  _GEN_63669;
  wire  _GEN_63671;
  wire  _GEN_63759;
  wire  _GEN_63761;
  wire  _GEN_429_is_load;
  wire  _GEN_430;
  wire  _GEN_63782;
  wire  _GEN_63783;
  wire  _GEN_63784;
  wire  _GEN_63785;
  wire  _GEN_63786;
  wire  _GEN_63787;
  wire  _GEN_63788;
  wire  _GEN_63789;
  wire  _GEN_63790;
  wire  _GEN_63791;
  wire  _GEN_63792;
  wire  _GEN_63793;
  wire  _GEN_63794;
  wire  _GEN_63795;
  wire  _GEN_63796;
  wire  _GEN_63797;
  wire  _GEN_63798;
  wire  _GEN_63799;
  wire  _GEN_63800;
  wire  _GEN_63801;
  wire  _GEN_63802;
  wire  _GEN_63803;
  wire  _GEN_63804;
  wire  _GEN_63805;
  wire  _GEN_63806;
  wire  _GEN_63807;
  wire  _GEN_63808;
  wire  _GEN_63809;
  wire  _GEN_63810;
  wire  _GEN_63811;
  wire  _GEN_63812;
  wire  _GEN_63813;
  wire  _GEN_63814;
  wire  _GEN_63815;
  wire  _GEN_63816;
  wire  _GEN_63817;
  wire  _GEN_63818;
  wire  _GEN_63819;
  wire  _GEN_63820;
  wire  _GEN_431;
  wire  _GEN_63821;
  wire  _GEN_63822;
  wire  _GEN_63823;
  wire  _GEN_63824;
  wire  _GEN_63825;
  wire  _GEN_63826;
  wire  _GEN_63827;
  wire  _GEN_63828;
  wire  _GEN_63829;
  wire  _GEN_63830;
  wire  _GEN_63831;
  wire  _GEN_63832;
  wire  _GEN_63833;
  wire  _GEN_63834;
  wire  _GEN_63835;
  wire  _GEN_63836;
  wire  _GEN_63837;
  wire  _GEN_63838;
  wire  _GEN_63839;
  wire  _GEN_63840;
  wire  _GEN_63841;
  wire  _GEN_63842;
  wire  _GEN_63843;
  wire  _GEN_63844;
  wire  _GEN_63845;
  wire  _GEN_63846;
  wire  _GEN_63847;
  wire  _GEN_63848;
  wire  _GEN_63849;
  wire  _GEN_63850;
  wire  _GEN_63851;
  wire  _GEN_63852;
  wire  _GEN_63853;
  wire  _GEN_63854;
  wire  _GEN_63855;
  wire  _GEN_63856;
  wire  _GEN_63857;
  wire  _GEN_63858;
  wire  _GEN_63859;
  wire  _GEN_435;
  wire  _GEN_64100;
  wire  _GEN_64101;
  wire  _GEN_64102;
  wire  _GEN_64103;
  wire  _GEN_64104;
  wire  _GEN_64105;
  wire  _GEN_64106;
  wire  _GEN_64107;
  wire  _GEN_64108;
  wire  _GEN_64109;
  wire  _GEN_64110;
  wire  _GEN_64111;
  wire  _GEN_64112;
  wire  _GEN_64113;
  wire  _GEN_64114;
  wire  _GEN_64115;
  wire  _GEN_64116;
  wire  _GEN_64117;
  wire  _GEN_64118;
  wire  _GEN_64119;
  wire  _GEN_64120;
  wire  _GEN_64121;
  wire  _GEN_64122;
  wire  _GEN_64123;
  wire  _GEN_64124;
  wire  _GEN_64125;
  wire  _GEN_64126;
  wire  _GEN_64127;
  wire  _GEN_64128;
  wire  _GEN_64129;
  wire  _GEN_64130;
  wire  _GEN_64131;
  wire  _GEN_64132;
  wire  _GEN_64133;
  wire  _GEN_64134;
  wire  _GEN_64135;
  wire  _GEN_64136;
  wire  _GEN_64137;
  wire  _GEN_64138;
  wire  _T_7677;
  wire  _T_7678;
  wire  _T_7680;
  wire  _T_7682;
  wire  _T_7684;
  wire [5:0] _T_7691;
  wire  _T_7694;
  wire  _T_7695;
  wire  _T_7697;
  wire  _T_7699;
  wire  _T_7701;
  wire  _GEN_436_ldst_val;
  wire [6:0] _GEN_64191;
  wire  _GEN_64216;
  wire [6:0] _GEN_64281;
  wire  _GEN_64306;
  wire [6:0] _GEN_64371;
  wire  _GEN_64396;
  wire [6:0] _GEN_64461;
  wire  _GEN_64486;
  wire [6:0] _GEN_64551;
  wire  _GEN_64576;
  wire [6:0] _GEN_64641;
  wire  _GEN_64666;
  wire [6:0] _GEN_64731;
  wire  _GEN_64756;
  wire [6:0] _GEN_64821;
  wire  _GEN_64846;
  wire [6:0] _GEN_64911;
  wire  _GEN_64936;
  wire [6:0] _GEN_65001;
  wire  _GEN_65026;
  wire [6:0] _GEN_65091;
  wire  _GEN_65116;
  wire [6:0] _GEN_65181;
  wire  _GEN_65206;
  wire [6:0] _GEN_65271;
  wire  _GEN_65296;
  wire [6:0] _GEN_65361;
  wire  _GEN_65386;
  wire [6:0] _GEN_65451;
  wire  _GEN_65476;
  wire [6:0] _GEN_65541;
  wire  _GEN_65566;
  wire [6:0] _GEN_65631;
  wire  _GEN_65656;
  wire [6:0] _GEN_65721;
  wire  _GEN_65746;
  wire [6:0] _GEN_65811;
  wire  _GEN_65836;
  wire [6:0] _GEN_65901;
  wire  _GEN_65926;
  wire [6:0] _GEN_65991;
  wire  _GEN_66016;
  wire [6:0] _GEN_66081;
  wire  _GEN_66106;
  wire [6:0] _GEN_66171;
  wire  _GEN_66196;
  wire [6:0] _GEN_66261;
  wire  _GEN_66286;
  wire [6:0] _GEN_66351;
  wire  _GEN_66376;
  wire [6:0] _GEN_66441;
  wire  _GEN_66466;
  wire [6:0] _GEN_66531;
  wire  _GEN_66556;
  wire [6:0] _GEN_66621;
  wire  _GEN_66646;
  wire [6:0] _GEN_66711;
  wire  _GEN_66736;
  wire [6:0] _GEN_66801;
  wire  _GEN_66826;
  wire [6:0] _GEN_66891;
  wire  _GEN_66916;
  wire [6:0] _GEN_66981;
  wire  _GEN_67006;
  wire [6:0] _GEN_67071;
  wire  _GEN_67096;
  wire [6:0] _GEN_67161;
  wire  _GEN_67186;
  wire [6:0] _GEN_67251;
  wire  _GEN_67276;
  wire [6:0] _GEN_67341;
  wire  _GEN_67366;
  wire [6:0] _GEN_67431;
  wire  _GEN_67456;
  wire [6:0] _GEN_67521;
  wire  _GEN_67546;
  wire [6:0] _GEN_67611;
  wire  _GEN_67636;
  wire  _T_7706;
  wire [6:0] _GEN_437_pdst;
  wire  _T_7707;
  wire  _T_7708;
  wire  _T_7710;
  wire  _T_7712;
  wire  _T_7714;
  wire  _GEN_439;
  wire  _GEN_67729;
  wire  _GEN_67730;
  wire  _GEN_67731;
  wire  _GEN_67732;
  wire  _GEN_67733;
  wire  _GEN_67734;
  wire  _GEN_67735;
  wire  _GEN_67736;
  wire  _GEN_67737;
  wire  _GEN_67738;
  wire  _GEN_67739;
  wire  _GEN_67740;
  wire  _GEN_67741;
  wire  _GEN_67742;
  wire  _GEN_67743;
  wire  _GEN_67744;
  wire  _GEN_67745;
  wire  _GEN_67746;
  wire  _GEN_67747;
  wire  _GEN_67748;
  wire  _GEN_67749;
  wire  _GEN_67750;
  wire  _GEN_67751;
  wire  _GEN_67752;
  wire  _GEN_67753;
  wire  _GEN_67754;
  wire  _GEN_67755;
  wire  _GEN_67756;
  wire  _GEN_67757;
  wire  _GEN_67758;
  wire  _GEN_67759;
  wire  _GEN_67760;
  wire  _GEN_67761;
  wire  _GEN_67762;
  wire  _GEN_67763;
  wire  _GEN_67764;
  wire  _GEN_67765;
  wire  _GEN_67766;
  wire  _GEN_67767;
  wire  _T_7754;
  wire  _T_7755;
  wire  _T_7757;
  wire  _T_7759;
  wire  _T_7761;
  wire [5:0] _T_7768;
  wire  _T_7771;
  wire  _T_7772;
  wire  _T_7774;
  wire  _T_7776;
  wire  _T_7778;
  wire  _GEN_440_ldst_val;
  wire [6:0] _GEN_67820;
  wire  _GEN_67845;
  wire [6:0] _GEN_67910;
  wire  _GEN_67935;
  wire [6:0] _GEN_68000;
  wire  _GEN_68025;
  wire [6:0] _GEN_68090;
  wire  _GEN_68115;
  wire [6:0] _GEN_68180;
  wire  _GEN_68205;
  wire [6:0] _GEN_68270;
  wire  _GEN_68295;
  wire [6:0] _GEN_68360;
  wire  _GEN_68385;
  wire [6:0] _GEN_68450;
  wire  _GEN_68475;
  wire [6:0] _GEN_68540;
  wire  _GEN_68565;
  wire [6:0] _GEN_68630;
  wire  _GEN_68655;
  wire [6:0] _GEN_68720;
  wire  _GEN_68745;
  wire [6:0] _GEN_68810;
  wire  _GEN_68835;
  wire [6:0] _GEN_68900;
  wire  _GEN_68925;
  wire [6:0] _GEN_68990;
  wire  _GEN_69015;
  wire [6:0] _GEN_69080;
  wire  _GEN_69105;
  wire [6:0] _GEN_69170;
  wire  _GEN_69195;
  wire [6:0] _GEN_69260;
  wire  _GEN_69285;
  wire [6:0] _GEN_69350;
  wire  _GEN_69375;
  wire [6:0] _GEN_69440;
  wire  _GEN_69465;
  wire [6:0] _GEN_69530;
  wire  _GEN_69555;
  wire [6:0] _GEN_69620;
  wire  _GEN_69645;
  wire [6:0] _GEN_69710;
  wire  _GEN_69735;
  wire [6:0] _GEN_69800;
  wire  _GEN_69825;
  wire [6:0] _GEN_69890;
  wire  _GEN_69915;
  wire [6:0] _GEN_69980;
  wire  _GEN_70005;
  wire [6:0] _GEN_70070;
  wire  _GEN_70095;
  wire [6:0] _GEN_70160;
  wire  _GEN_70185;
  wire [6:0] _GEN_70250;
  wire  _GEN_70275;
  wire [6:0] _GEN_70340;
  wire  _GEN_70365;
  wire [6:0] _GEN_70430;
  wire  _GEN_70455;
  wire [6:0] _GEN_70520;
  wire  _GEN_70545;
  wire [6:0] _GEN_70610;
  wire  _GEN_70635;
  wire [6:0] _GEN_70700;
  wire  _GEN_70725;
  wire [6:0] _GEN_70790;
  wire  _GEN_70815;
  wire [6:0] _GEN_70880;
  wire  _GEN_70905;
  wire [6:0] _GEN_70970;
  wire  _GEN_70995;
  wire [6:0] _GEN_71060;
  wire  _GEN_71085;
  wire [6:0] _GEN_71150;
  wire  _GEN_71175;
  wire [6:0] _GEN_71240;
  wire  _GEN_71265;
  wire  _T_7783;
  wire [6:0] _GEN_441_pdst;
  wire  _T_7784;
  wire  _T_7785;
  wire  _T_7787;
  wire  _T_7789;
  wire  _T_7791;
  wire  _GEN_443;
  wire  _GEN_71358;
  wire  _GEN_71359;
  wire  _GEN_71360;
  wire  _GEN_71361;
  wire  _GEN_71362;
  wire  _GEN_71363;
  wire  _GEN_71364;
  wire  _GEN_71365;
  wire  _GEN_71366;
  wire  _GEN_71367;
  wire  _GEN_71368;
  wire  _GEN_71369;
  wire  _GEN_71370;
  wire  _GEN_71371;
  wire  _GEN_71372;
  wire  _GEN_71373;
  wire  _GEN_71374;
  wire  _GEN_71375;
  wire  _GEN_71376;
  wire  _GEN_71377;
  wire  _GEN_71378;
  wire  _GEN_71379;
  wire  _GEN_71380;
  wire  _GEN_71381;
  wire  _GEN_71382;
  wire  _GEN_71383;
  wire  _GEN_71384;
  wire  _GEN_71385;
  wire  _GEN_71386;
  wire  _GEN_71387;
  wire  _GEN_71388;
  wire  _GEN_71389;
  wire  _GEN_71390;
  wire  _GEN_71391;
  wire  _GEN_71392;
  wire  _GEN_71393;
  wire  _GEN_71394;
  wire  _GEN_71395;
  wire  _GEN_71396;
  wire  _T_7831;
  wire  _T_7832;
  wire  _T_7834;
  wire  _T_7836;
  wire  _T_7838;
  wire [5:0] _T_7845;
  wire  _T_7848;
  wire  _T_7849;
  wire  _T_7851;
  wire  _T_7853;
  wire  _T_7855;
  wire  _GEN_444_ldst_val;
  wire [6:0] _GEN_71449;
  wire  _GEN_71474;
  wire [6:0] _GEN_71539;
  wire  _GEN_71564;
  wire [6:0] _GEN_71629;
  wire  _GEN_71654;
  wire [6:0] _GEN_71719;
  wire  _GEN_71744;
  wire [6:0] _GEN_71809;
  wire  _GEN_71834;
  wire [6:0] _GEN_71899;
  wire  _GEN_71924;
  wire [6:0] _GEN_71989;
  wire  _GEN_72014;
  wire [6:0] _GEN_72079;
  wire  _GEN_72104;
  wire [6:0] _GEN_72169;
  wire  _GEN_72194;
  wire [6:0] _GEN_72259;
  wire  _GEN_72284;
  wire [6:0] _GEN_72349;
  wire  _GEN_72374;
  wire [6:0] _GEN_72439;
  wire  _GEN_72464;
  wire [6:0] _GEN_72529;
  wire  _GEN_72554;
  wire [6:0] _GEN_72619;
  wire  _GEN_72644;
  wire [6:0] _GEN_72709;
  wire  _GEN_72734;
  wire [6:0] _GEN_72799;
  wire  _GEN_72824;
  wire [6:0] _GEN_72889;
  wire  _GEN_72914;
  wire [6:0] _GEN_72979;
  wire  _GEN_73004;
  wire [6:0] _GEN_73069;
  wire  _GEN_73094;
  wire [6:0] _GEN_73159;
  wire  _GEN_73184;
  wire [6:0] _GEN_73249;
  wire  _GEN_73274;
  wire [6:0] _GEN_73339;
  wire  _GEN_73364;
  wire [6:0] _GEN_73429;
  wire  _GEN_73454;
  wire [6:0] _GEN_73519;
  wire  _GEN_73544;
  wire [6:0] _GEN_73609;
  wire  _GEN_73634;
  wire [6:0] _GEN_73699;
  wire  _GEN_73724;
  wire [6:0] _GEN_73789;
  wire  _GEN_73814;
  wire [6:0] _GEN_73879;
  wire  _GEN_73904;
  wire [6:0] _GEN_73969;
  wire  _GEN_73994;
  wire [6:0] _GEN_74059;
  wire  _GEN_74084;
  wire [6:0] _GEN_74149;
  wire  _GEN_74174;
  wire [6:0] _GEN_74239;
  wire  _GEN_74264;
  wire [6:0] _GEN_74329;
  wire  _GEN_74354;
  wire [6:0] _GEN_74419;
  wire  _GEN_74444;
  wire [6:0] _GEN_74509;
  wire  _GEN_74534;
  wire [6:0] _GEN_74599;
  wire  _GEN_74624;
  wire [6:0] _GEN_74689;
  wire  _GEN_74714;
  wire [6:0] _GEN_74779;
  wire  _GEN_74804;
  wire [6:0] _GEN_74869;
  wire  _GEN_74894;
  wire  _T_7860;
  wire [6:0] _GEN_445_pdst;
  wire  _T_7861;
  wire  _T_7862;
  wire  _T_7864;
  wire  _T_7866;
  wire  _T_7868;
  wire  _GEN_447;
  wire  _GEN_74987;
  wire  _GEN_74988;
  wire  _GEN_74989;
  wire  _GEN_74990;
  wire  _GEN_74991;
  wire  _GEN_74992;
  wire  _GEN_74993;
  wire  _GEN_74994;
  wire  _GEN_74995;
  wire  _GEN_74996;
  wire  _GEN_74997;
  wire  _GEN_74998;
  wire  _GEN_74999;
  wire  _GEN_75000;
  wire  _GEN_75001;
  wire  _GEN_75002;
  wire  _GEN_75003;
  wire  _GEN_75004;
  wire  _GEN_75005;
  wire  _GEN_75006;
  wire  _GEN_75007;
  wire  _GEN_75008;
  wire  _GEN_75009;
  wire  _GEN_75010;
  wire  _GEN_75011;
  wire  _GEN_75012;
  wire  _GEN_75013;
  wire  _GEN_75014;
  wire  _GEN_75015;
  wire  _GEN_75016;
  wire  _GEN_75017;
  wire  _GEN_75018;
  wire  _GEN_75019;
  wire  _GEN_75020;
  wire  _GEN_75021;
  wire  _GEN_75022;
  wire  _GEN_75023;
  wire  _GEN_75024;
  wire  _GEN_75025;
  wire  _T_7908;
  wire  _T_7909;
  wire  _T_7911;
  wire  _T_7913;
  wire  _T_7915;
  wire [5:0] _T_7922;
  wire  _T_7925;
  wire  _T_7926;
  wire  _T_7928;
  wire  _T_7930;
  wire  _T_7932;
  wire  _GEN_448_ldst_val;
  wire [6:0] _GEN_75078;
  wire  _GEN_75103;
  wire [6:0] _GEN_75168;
  wire  _GEN_75193;
  wire [6:0] _GEN_75258;
  wire  _GEN_75283;
  wire [6:0] _GEN_75348;
  wire  _GEN_75373;
  wire [6:0] _GEN_75438;
  wire  _GEN_75463;
  wire [6:0] _GEN_75528;
  wire  _GEN_75553;
  wire [6:0] _GEN_75618;
  wire  _GEN_75643;
  wire [6:0] _GEN_75708;
  wire  _GEN_75733;
  wire [6:0] _GEN_75798;
  wire  _GEN_75823;
  wire [6:0] _GEN_75888;
  wire  _GEN_75913;
  wire [6:0] _GEN_75978;
  wire  _GEN_76003;
  wire [6:0] _GEN_76068;
  wire  _GEN_76093;
  wire [6:0] _GEN_76158;
  wire  _GEN_76183;
  wire [6:0] _GEN_76248;
  wire  _GEN_76273;
  wire [6:0] _GEN_76338;
  wire  _GEN_76363;
  wire [6:0] _GEN_76428;
  wire  _GEN_76453;
  wire [6:0] _GEN_76518;
  wire  _GEN_76543;
  wire [6:0] _GEN_76608;
  wire  _GEN_76633;
  wire [6:0] _GEN_76698;
  wire  _GEN_76723;
  wire [6:0] _GEN_76788;
  wire  _GEN_76813;
  wire [6:0] _GEN_76878;
  wire  _GEN_76903;
  wire [6:0] _GEN_76968;
  wire  _GEN_76993;
  wire [6:0] _GEN_77058;
  wire  _GEN_77083;
  wire [6:0] _GEN_77148;
  wire  _GEN_77173;
  wire [6:0] _GEN_77238;
  wire  _GEN_77263;
  wire [6:0] _GEN_77328;
  wire  _GEN_77353;
  wire [6:0] _GEN_77418;
  wire  _GEN_77443;
  wire [6:0] _GEN_77508;
  wire  _GEN_77533;
  wire [6:0] _GEN_77598;
  wire  _GEN_77623;
  wire [6:0] _GEN_77688;
  wire  _GEN_77713;
  wire [6:0] _GEN_77778;
  wire  _GEN_77803;
  wire [6:0] _GEN_77868;
  wire  _GEN_77893;
  wire [6:0] _GEN_77958;
  wire  _GEN_77983;
  wire [6:0] _GEN_78048;
  wire  _GEN_78073;
  wire [6:0] _GEN_78138;
  wire  _GEN_78163;
  wire [6:0] _GEN_78228;
  wire  _GEN_78253;
  wire [6:0] _GEN_78318;
  wire  _GEN_78343;
  wire [6:0] _GEN_78408;
  wire  _GEN_78433;
  wire [6:0] _GEN_78498;
  wire  _GEN_78523;
  wire  _T_7937;
  wire [6:0] _GEN_449_pdst;
  wire  _T_7938;
  wire  _T_7939;
  wire  _T_7941;
  wire  _T_7943;
  wire  _T_7945;
  wire  _GEN_451;
  wire  _GEN_78616;
  wire  _GEN_78617;
  wire  _GEN_78618;
  wire  _GEN_78619;
  wire  _GEN_78620;
  wire  _GEN_78621;
  wire  _GEN_78622;
  wire  _GEN_78623;
  wire  _GEN_78624;
  wire  _GEN_78625;
  wire  _GEN_78626;
  wire  _GEN_78627;
  wire  _GEN_78628;
  wire  _GEN_78629;
  wire  _GEN_78630;
  wire  _GEN_78631;
  wire  _GEN_78632;
  wire  _GEN_78633;
  wire  _GEN_78634;
  wire  _GEN_78635;
  wire  _GEN_78636;
  wire  _GEN_78637;
  wire  _GEN_78638;
  wire  _GEN_78639;
  wire  _GEN_78640;
  wire  _GEN_78641;
  wire  _GEN_78642;
  wire  _GEN_78643;
  wire  _GEN_78644;
  wire  _GEN_78645;
  wire  _GEN_78646;
  wire  _GEN_78647;
  wire  _GEN_78648;
  wire  _GEN_78649;
  wire  _GEN_78650;
  wire  _GEN_78651;
  wire  _GEN_78652;
  wire  _GEN_78653;
  wire  _GEN_78654;
  wire  _T_7985;
  wire  _T_7986;
  wire  _T_7988;
  wire  _T_7990;
  wire  _T_7992;
  wire [5:0] _T_7999;
  wire  _T_8002;
  wire  _T_8003;
  wire  _T_8005;
  wire  _T_8007;
  wire  _T_8009;
  wire  _GEN_452_ldst_val;
  wire [6:0] _GEN_78707;
  wire  _GEN_78732;
  wire [6:0] _GEN_78797;
  wire  _GEN_78822;
  wire [6:0] _GEN_78887;
  wire  _GEN_78912;
  wire [6:0] _GEN_78977;
  wire  _GEN_79002;
  wire [6:0] _GEN_79067;
  wire  _GEN_79092;
  wire [6:0] _GEN_79157;
  wire  _GEN_79182;
  wire [6:0] _GEN_79247;
  wire  _GEN_79272;
  wire [6:0] _GEN_79337;
  wire  _GEN_79362;
  wire [6:0] _GEN_79427;
  wire  _GEN_79452;
  wire [6:0] _GEN_79517;
  wire  _GEN_79542;
  wire [6:0] _GEN_79607;
  wire  _GEN_79632;
  wire [6:0] _GEN_79697;
  wire  _GEN_79722;
  wire [6:0] _GEN_79787;
  wire  _GEN_79812;
  wire [6:0] _GEN_79877;
  wire  _GEN_79902;
  wire [6:0] _GEN_79967;
  wire  _GEN_79992;
  wire [6:0] _GEN_80057;
  wire  _GEN_80082;
  wire [6:0] _GEN_80147;
  wire  _GEN_80172;
  wire [6:0] _GEN_80237;
  wire  _GEN_80262;
  wire [6:0] _GEN_80327;
  wire  _GEN_80352;
  wire [6:0] _GEN_80417;
  wire  _GEN_80442;
  wire [6:0] _GEN_80507;
  wire  _GEN_80532;
  wire [6:0] _GEN_80597;
  wire  _GEN_80622;
  wire [6:0] _GEN_80687;
  wire  _GEN_80712;
  wire [6:0] _GEN_80777;
  wire  _GEN_80802;
  wire [6:0] _GEN_80867;
  wire  _GEN_80892;
  wire [6:0] _GEN_80957;
  wire  _GEN_80982;
  wire [6:0] _GEN_81047;
  wire  _GEN_81072;
  wire [6:0] _GEN_81137;
  wire  _GEN_81162;
  wire [6:0] _GEN_81227;
  wire  _GEN_81252;
  wire [6:0] _GEN_81317;
  wire  _GEN_81342;
  wire [6:0] _GEN_81407;
  wire  _GEN_81432;
  wire [6:0] _GEN_81497;
  wire  _GEN_81522;
  wire [6:0] _GEN_81587;
  wire  _GEN_81612;
  wire [6:0] _GEN_81677;
  wire  _GEN_81702;
  wire [6:0] _GEN_81767;
  wire  _GEN_81792;
  wire [6:0] _GEN_81857;
  wire  _GEN_81882;
  wire [6:0] _GEN_81947;
  wire  _GEN_81972;
  wire [6:0] _GEN_82037;
  wire  _GEN_82062;
  wire [6:0] _GEN_82127;
  wire  _GEN_82152;
  wire  _T_8014;
  wire [6:0] _GEN_453_pdst;
  wire  _T_8015;
  wire  _T_8016;
  wire  _T_8018;
  wire  _T_8020;
  wire  _T_8022;
  wire  _T_8032;
  wire  _T_8033;
  wire  _T_8034;
  wire  _T_8038;
  wire  _T_8039;
  wire  _T_8045;
  wire  _T_8046;
  wire  _T_8049;
  wire  _T_8051;
  wire  _T_8052;
  wire  _T_8053;
  wire  _T_8054;
  wire  _T_8056;
  wire  _T_8057;
  wire  _T_8059;
  wire  _T_8060;
  wire  will_throw_exception;
  wire  _T_8062;
  wire  _T_8063;
  wire  _T_8066;
  wire  _T_8072;
  wire  _T_8073;
  wire  is_mini_exception;
  wire  _T_8075;
  wire  _T_8076;
  wire  _T_8077;
  wire  _T_8078;
  wire  insn_sys_pc2epc;
  wire  refetch_inst;
  wire [63:0] _T_8080;
  wire [5:0] _T_8082;
  wire [4:0] _T_8083;
  wire [39:0] _GEN_440;
  wire [39:0] _T_8086;
  wire  _T_8087;
  wire [4:0] _T_8090;
  wire [39:0] _GEN_441;
  wire [39:0] _T_8093;
  wire [39:0] _GEN_82168;
  wire [39:0] _T_8094;
  wire  _T_8095;
  wire [23:0] _T_8099;
  wire [63:0] _T_8100;
  wire [2:0] _T_8103;
  wire [63:0] _GEN_444;
  wire [64:0] _T_8104;
  wire [63:0] _T_8105;
  wire [2:0] _T_8108;
  wire [63:0] _GEN_445;
  wire [64:0] _T_8109;
  wire [63:0] flush_pc;
  wire  _T_8110;
  wire  _T_8111;
  wire  _T_8112;
  wire  _T_8113;
  wire  flush_val;
  reg  _T_8115;
  reg [31:0] _RAND_1086;
  wire  _T_8117;
  wire [63:0] _T_8118;
  reg [63:0] _T_8120;
  reg [63:0] _RAND_1087;
  wire  _T_8122;
  reg  com_lsu_misspec;
  reg [31:0] _RAND_1088;
  wire  _T_8125;
  wire  _T_8126;
  wire  _T_8128;
  wire  _T_8130;
  wire  _T_8132;
  wire  fflags_val_0;
  wire  fflags_val_1;
  wire [4:0] fflags_0;
  wire [4:0] fflags_1;
  wire  _T_8147;
  wire  _T_8148;
  wire  _T_8150;
  wire  _T_8151;
  wire [4:0] _T_8153;
  wire  _T_8155;
  wire  _T_8156;
  wire  _T_8158;
  wire  _T_8159;
  wire  _T_8161;
  wire  _T_8163;
  wire  _T_8165;
  wire  _T_8168;
  wire  _T_8171;
  wire  _T_8173;
  wire  _T_8175;
  wire  _T_8177;
  wire  _T_8178;
  wire  _T_8179;
  wire  _T_8181;
  wire  _T_8182;
  wire [4:0] _T_8184;
  wire  _T_8186;
  wire  _T_8187;
  wire  _T_8189;
  wire  _T_8190;
  wire  _T_8192;
  wire  _T_8194;
  wire  _T_8196;
  wire  _T_8199;
  wire  _T_8202;
  wire  _T_8204;
  wire  _T_8206;
  wire  _T_8208;
  wire  _T_8209;
  wire [4:0] _T_8210;
  wire [7:0] next_xcpt_uop_br_mask;
  wire [6:0] next_xcpt_uop_rob_idx;
  wire [63:0] next_xcpt_uop_exc_cause;
  wire  enq_xcpts_0;
  wire  enq_xcpts_1;
  wire  _T_8227;
  wire  _T_8228;
  wire  _T_8229;
  wire  _T_8231;
  wire  _T_8232;
  wire  _T_8233;
  wire  _T_8234;
  wire  _T_8236;
  wire  _T_8237;
  wire  _T_8238;
  wire  _T_8239;
  wire [7:0] _T_8240;
  wire  _T_8241;
  wire [7:0] _T_8242;
  wire  _T_8243;
  wire  _T_8244;
  wire  _T_8245;
  wire [7:0] _T_8246_br_mask;
  wire [6:0] _T_8246_rob_idx;
  wire  _T_8252;
  wire  _T_8253;
  wire [7:0] _T_8254;
  wire  _T_8255;
  wire [7:0] _T_8256;
  wire  _T_8257;
  wire  _T_8258;
  wire [4:0] _T_8260;
  wire [39:0] _T_8261;
  wire  _GEN_82169;
  wire [7:0] _GEN_82194;
  wire [6:0] _GEN_82218;
  wire [63:0] _GEN_82231;
  wire [63:0] _GEN_82260;
  wire  _T_8264;
  wire  _T_8265;
  wire  _T_8268;
  wire [7:0] _GEN_82285;
  wire [6:0] _GEN_82309;
  wire [63:0] _GEN_82322;
  wire [7:0] _GEN_479_br_mask;
  wire [6:0] _GEN_503_rob_idx;
  wire [63:0] _GEN_516_exc_cause;
  wire [63:0] _GEN_545_exc_cause;
  wire  _T_8289;
  wire [3:0] _GEN_448;
  wire [3:0] _T_8292;
  wire [39:0] _GEN_449;
  wire [40:0] _T_8293;
  wire [39:0] _T_8294;
  wire [39:0] _T_8295;
  wire  _GEN_82351;
  wire [7:0] _GEN_82376;
  wire [6:0] _GEN_82400;
  wire [63:0] _GEN_82413;
  wire [63:0] _GEN_82442;
  wire  _GEN_82443;
  wire [7:0] _GEN_82468;
  wire [6:0] _GEN_82492;
  wire [63:0] _GEN_82505;
  wire [63:0] _GEN_82534;
  wire  _GEN_82535;
  wire [7:0] _GEN_82560;
  wire [6:0] _GEN_82584;
  wire [63:0] _GEN_82597;
  wire [63:0] _GEN_82626;
  wire [7:0] _T_8297;
  wire [7:0] _T_8298;
  wire [7:0] _T_8300;
  wire  _T_8302;
  wire  _T_8303;
  wire  _T_8304;
  wire  _GEN_82627;
  wire  _T_8311;
  wire  _T_8313;
  wire  _T_8315;
  wire  _T_8317;
  wire  _T_8318;
  wire  _T_8320;
  wire  _T_8322;
  wire  _T_8324;
  wire [6:0] _T_8326;
  wire [6:0] _GEN_452;
  wire  _T_8327;
  wire  _T_8328;
  wire  _T_8330;
  wire  _T_8332;
  wire  _T_8334;
  wire [1:0] _T_8335;
  wire  _T_8337;
  wire [1:0] _T_8338;
  wire [1:0] _T_8339;
  wire [1:0] _T_8340;
  wire  _T_8342;
  wire  _T_8343;
  wire  _T_8344;
  wire  _T_8345;
  wire  _T_8347;
  wire  _T_8348;
  wire  _T_8350;
  wire [6:0] _T_8353;
  wire [5:0] _T_8354;
  wire [5:0] _T_8355;
  wire [5:0] _GEN_82628;
  wire  _T_8357;
  wire  _T_8358;
  wire  _T_8360;
  wire [6:0] _T_8363;
  wire [6:0] _T_8364;
  wire [5:0] _T_8365;
  wire [5:0] _T_8366;
  wire  _T_8371;
  wire [7:0] _T_8374;
  wire [6:0] _T_8375;
  wire [6:0] _T_8376;
  wire  _T_8379;
  wire  _T_8381;
  wire  _T_8382;
  wire  _T_8384;
  wire [6:0] _T_8387;
  wire [5:0] _T_8388;
  wire [5:0] _T_8389;
  wire [5:0] _GEN_82629;
  wire [6:0] _GEN_82630;
  wire [6:0] _GEN_82631;
  wire  full;
  wire  _T_8400;
  wire  _T_8401;
  wire  _T_8402;
  wire  _T_8404;
  wire  _T_8405;
  wire  _T_8406;
  wire [1:0] _GEN_82632;
  wire  _T_8407;
  wire [1:0] _GEN_82633;
  wire [1:0] _GEN_82634;
  wire [1:0] _GEN_82635;
  wire [1:0] _GEN_82636;
  wire  _T_8410;
  wire [1:0] _GEN_82637;
  wire [1:0] _GEN_82638;
  wire  _T_8411;
  wire [1:0] _GEN_82639;
  wire [1:0] _GEN_82640;
  wire [1:0] _GEN_82641;
  wire  _T_8412;
  wire  _T_8413;
  wire  _T_8414;
  wire  _T_8415;
  wire  _T_8417;
  wire  _T_8421;
  wire  _GEN_546;
  wire  _GEN_82642;
  assign _GEN_421 = {{1'd0}, rob_tail};
  assign rob_tail_idx = _GEN_421 << 1'h1;
  assign _T_2772__T_2805_addr = _T_2804;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2772__T_2805_data = _T_2772[_T_2772__T_2805_addr];
  `else
  assign _T_2772__T_2805_data = _T_2772__T_2805_addr >= 5'h14 ? _RAND_9[36:0] : _T_2772[_T_2772__T_2805_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2772__T_8084_addr = _T_8083;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2772__T_8084_data = _T_2772[_T_2772__T_8084_addr];
  `else
  assign _T_2772__T_8084_data = _T_2772__T_8084_addr >= 5'h14 ? _RAND_10[36:0] : _T_2772[_T_2772__T_8084_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2772__T_2788_data = _GEN_112;
  assign _T_2772__T_2788_addr = _T_2787;
  assign _T_2772__T_2788_mask = _GEN_561;
  assign _T_2772__T_2788_en = _GEN_561;
  assign _GEN_112 = _T_2779[36:0];
  assign _T_2775__T_2811_addr = _T_2810;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2775__T_2811_data = _T_2775[_T_2775__T_2811_addr];
  `else
  assign _T_2775__T_2811_data = _T_2775__T_2811_addr >= 5'h14 ? _RAND_12[36:0] : _T_2775[_T_2775__T_2811_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2775__T_8091_addr = _T_8090;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2775__T_8091_data = _T_2775[_T_2775__T_8091_addr];
  `else
  assign _T_2775__T_8091_data = _T_2775__T_8091_addr >= 5'h14 ? _RAND_13[36:0] : _T_2775[_T_2775__T_8091_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2775__T_2784_data = _GEN_112;
  assign _T_2775__T_2784_addr = _T_2783;
  assign _T_2775__T_2784_mask = _GEN_557;
  assign _T_2775__T_2784_en = _GEN_557;
  assign _T_2776 = io_enq_valids_0 | io_enq_valids_1;
  assign _T_2779 = io_enq_uops_0_pc >> 2'h3;
  assign _T_2780 = rob_tail[0];
  assign _T_2782 = rob_tail >> 1'h1;
  assign _T_2783 = _T_2782[4:0];
  assign _T_2787 = _T_2782[4:0];
  assign _GEN_553 = _T_2780 ? 1'h0 : 1'h1;
  assign _GEN_557 = _T_2776 ? _T_2780 : 1'h0;
  assign _GEN_561 = _T_2776 ? _GEN_553 : 1'h0;
  assign _T_2790 = io_get_pc_rob_idx >> 1'h1;
  assign _T_2791 = _T_2790[0];
  assign _T_2793 = _T_2790 >> 1'h1;
  assign _T_2795 = _T_2793 == 7'h13;
  assign _T_2798 = _T_2793 + 7'h1;
  assign _T_2799 = _T_2798[6:0];
  assign _T_2800 = _T_2795 ? 7'h0 : _T_2799;
  assign _T_2803 = _T_2791 ? _T_2800 : _T_2793;
  assign _T_2804 = _T_2803[4:0];
  assign _GEN_423 = {{3'd0}, _T_2772__T_2805_data};
  assign _T_2807 = _GEN_423 << 2'h3;
  assign _T_2810 = _T_2793[4:0];
  assign _GEN_424 = {{3'd0}, _T_2775__T_2811_data};
  assign _T_2813 = _GEN_424 << 2'h3;
  assign _T_2819 = _T_2791 ? _T_2813 : _T_2807;
  assign _T_2821 = _T_2791 ? _T_2807 : _T_2813;
  assign _T_2822 = _T_2815[39:0];
  assign _T_2823 = _T_2822[39];
  assign _T_2827 = _T_2823 ? 24'hffffff : 24'h0;
  assign curr_row_pc = {_T_2827,_T_2822};
  assign _T_2828 = _T_2817[39:0];
  assign _T_2829 = _T_2828[39];
  assign _T_2833 = _T_2829 ? 24'hffffff : 24'h0;
  assign next_row_pc = {_T_2833,_T_2828};
  assign _T_2834 = io_get_pc_rob_idx[0];
  assign _T_2836 = {_T_2834,2'h0};
  assign _GEN_428 = {{61'd0}, _T_2836};
  assign _T_2837 = curr_row_pc + _GEN_428;
  assign _T_2838 = _T_2837[63:0];
  assign _T_2841 = _T_2834 + 1'h1;
  assign curr_idx = _T_2841[0:0];
  assign _GEN_563 = curr_idx ? rob_getpc_curr_vals_1 : rob_getpc_curr_vals_0;
  assign _T_2846 = _GEN_0 & curr_idx;
  assign _T_2848 = {curr_idx,2'h0};
  assign _GEN_429 = {{61'd0}, _T_2848};
  assign _T_2849 = curr_row_pc + _GEN_429;
  assign curr_row_next_pc = _T_2849[63:0];
  assign _T_2850 = {rob_getpc_next_vals_1,rob_getpc_next_vals_0};
  assign _T_2851 = _T_2850[0];
  assign next_bank_idx = _T_2851 ? 1'h0 : 1'h1;
  assign rob_pc_hob_next_val = rob_getpc_next_vals_0 | rob_getpc_next_vals_1;
  assign _T_2855 = {io_enq_valids_1,io_enq_valids_0};
  assign _T_2856 = _T_2855[0];
  assign bypass_next_bank_idx = _T_2856 ? 1'h0 : 1'h1;
  assign _T_2860 = $signed(io_enq_uops_0_pc);
  assign _T_2862 = $signed(_T_2860) & $signed(-40'sh8);
  assign _T_2863 = $signed(_T_2862);
  assign _T_2864 = $unsigned(_T_2863);
  assign _T_2866 = {bypass_next_bank_idx,2'h0};
  assign _GEN_436 = {{37'd0}, _T_2866};
  assign _T_2867 = _T_2864 + _GEN_436;
  assign bypass_next_pc = _T_2867[39:0];
  assign _T_2869 = rob_pc_hob_next_val | _T_2776;
  assign _T_2870 = _T_2869 | curr_row_next_pc_val;
  assign _T_2872 = {next_bank_idx,2'h0};
  assign _GEN_437 = {{61'd0}, _T_2872};
  assign _T_2873 = next_row_pc + _GEN_437;
  assign _T_2874 = _T_2873[63:0];
  assign _T_2875 = rob_pc_hob_next_val ? _T_2874 : {{24'd0}, bypass_next_pc};
  assign _T_2876 = curr_row_next_pc_val ? curr_row_next_pc : _T_2875;
  assign row_metadata_brob_idx__T_2896_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx__T_2896_data = row_metadata_brob_idx[row_metadata_brob_idx__T_2896_addr];
  `else
  assign row_metadata_brob_idx__T_2896_data = row_metadata_brob_idx__T_2896_addr >= 6'h28 ? _RAND_16[5:0] : row_metadata_brob_idx[row_metadata_brob_idx__T_2896_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx__T_2900_addr = _T_2899;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx__T_2900_data = row_metadata_brob_idx[row_metadata_brob_idx__T_2900_addr];
  `else
  assign row_metadata_brob_idx__T_2900_data = row_metadata_brob_idx__T_2900_addr >= 6'h28 ? _RAND_17[5:0] : row_metadata_brob_idx[row_metadata_brob_idx__T_2900_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_brob_idx__T_2886_data = io_enq_uops_0_brob_idx;
  assign row_metadata_brob_idx__T_2886_addr = rob_tail;
  assign row_metadata_brob_idx__T_2886_mask = _T_2885;
  assign row_metadata_brob_idx__T_2886_en = _T_2885;
  assign row_metadata_has_brorjalr__T_2894_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr__T_2894_data = row_metadata_has_brorjalr[row_metadata_has_brorjalr__T_2894_addr];
  `else
  assign row_metadata_has_brorjalr__T_2894_data = row_metadata_has_brorjalr__T_2894_addr >= 6'h28 ? _RAND_19[0:0] : row_metadata_has_brorjalr[row_metadata_has_brorjalr__T_2894_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign row_metadata_has_brorjalr__T_2887_data = io_enq_has_br_or_jalr_in_packet;
  assign row_metadata_has_brorjalr__T_2887_addr = rob_tail;
  assign row_metadata_has_brorjalr__T_2887_mask = _T_2885;
  assign row_metadata_has_brorjalr__T_2887_en = _T_2885;
  assign row_metadata_has_brorjalr__T_2892_data = 1'h0;
  assign row_metadata_has_brorjalr__T_2892_addr = rob_tail;
  assign row_metadata_has_brorjalr__T_2892_mask = io_clear_brob;
  assign row_metadata_has_brorjalr__T_2892_en = io_clear_brob;
  assign _T_2885 = _T_2776 & io_enq_new_packet;
  assign _T_2890 = io_enq_new_packet == 1'h0;
  assign _T_2891 = _T_2776 & _T_2890;
  assign _GEN_564 = _T_2891 ? io_enq_partial_stall : r_partial_row;
  assign _GEN_570 = _T_2885 ? io_enq_partial_stall : _GEN_564;
  assign _T_2895 = finished_committing_row & row_metadata_has_brorjalr__T_2894_data;
  assign _T_2899 = _T_2790[5:0];
  assign _T_2901 = io_enq_valids_0 & io_enq_uops_0_is_unique;
  assign _T_2902 = io_enq_valids_1 & io_enq_uops_1_is_unique;
  assign _T_2903 = _T_2901 | _T_2902;
  assign _T_3200__T_3877_addr = _T_3876;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_3877_data = _T_3200[_T_3200__T_3877_addr];
  `else
  assign _T_3200__T_3877_data = _T_3200__T_3877_addr >= 6'h28 ? _RAND_61[0:0] : _T_3200[_T_3200__T_3877_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_3904_addr = _T_3903;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_3904_data = _T_3200[_T_3200__T_3904_addr];
  `else
  assign _T_3200__T_3904_data = _T_3200__T_3904_addr >= 6'h28 ? _RAND_62[0:0] : _T_3200[_T_3200__T_3904_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_4017_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_4017_data = _T_3200[_T_3200__T_4017_addr];
  `else
  assign _T_3200__T_4017_data = _T_3200__T_4017_addr >= 6'h28 ? _RAND_63[0:0] : _T_3200[_T_3200__T_4017_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5128_addr = _T_5127;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5128_data = _T_3200[_T_3200__T_5128_addr];
  `else
  assign _T_3200__T_5128_data = _T_3200__T_5128_addr >= 6'h28 ? _RAND_64[0:0] : _T_3200[_T_3200__T_5128_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5205_addr = _T_5204;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5205_data = _T_3200[_T_3200__T_5205_addr];
  `else
  assign _T_3200__T_5205_data = _T_3200__T_5205_addr >= 6'h28 ? _RAND_65[0:0] : _T_3200[_T_3200__T_5205_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5282_addr = _T_5281;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5282_data = _T_3200[_T_3200__T_5282_addr];
  `else
  assign _T_3200__T_5282_data = _T_3200__T_5282_addr >= 6'h28 ? _RAND_66[0:0] : _T_3200[_T_3200__T_5282_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5359_addr = _T_5358;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5359_data = _T_3200[_T_3200__T_5359_addr];
  `else
  assign _T_3200__T_5359_data = _T_3200__T_5359_addr >= 6'h28 ? _RAND_67[0:0] : _T_3200[_T_3200__T_5359_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5436_addr = _T_5435;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_5436_data = _T_3200[_T_3200__T_5436_addr];
  `else
  assign _T_3200__T_5436_data = _T_3200__T_5436_addr >= 6'h28 ? _RAND_68[0:0] : _T_3200[_T_3200__T_5436_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3200__T_3753_data = _T_3758;
  assign _T_3200__T_3753_addr = rob_tail;
  assign _T_3200__T_3753_mask = io_enq_valids_0;
  assign _T_3200__T_3753_en = io_enq_valids_0;
  assign _T_3200__T_3819_data = 1'h0;
  assign _T_3200__T_3819_addr = _T_3818;
  assign _T_3200__T_3819_mask = _T_3817;
  assign _T_3200__T_3819_en = _T_3817;
  assign _T_3200__T_3828_data = 1'h0;
  assign _T_3200__T_3828_addr = _T_3827;
  assign _T_3200__T_3828_mask = _T_3826;
  assign _T_3200__T_3828_en = _T_3826;
  assign _T_3200__T_3837_data = 1'h0;
  assign _T_3200__T_3837_addr = _T_3836;
  assign _T_3200__T_3837_mask = _T_3835;
  assign _T_3200__T_3837_en = _T_3835;
  assign _T_3200__T_3846_data = 1'h0;
  assign _T_3200__T_3846_addr = _T_3845;
  assign _T_3200__T_3846_mask = _T_3844;
  assign _T_3200__T_3846_en = _T_3844;
  assign _T_3200__T_3855_data = 1'h0;
  assign _T_3200__T_3855_addr = _T_3854;
  assign _T_3200__T_3855_mask = _T_3853;
  assign _T_3200__T_3855_en = _T_3853;
  assign _T_3200__T_3864_data = 1'h0;
  assign _T_3200__T_3864_addr = _T_3863;
  assign _T_3200__T_3864_mask = _T_3860;
  assign _T_3200__T_3864_en = _T_3860;
  assign _T_3200__T_3891_data = 1'h0;
  assign _T_3200__T_3891_addr = _T_3890;
  assign _T_3200__T_3891_mask = _T_3887;
  assign _T_3200__T_3891_en = _T_3887;
  assign _T_3745__T_4012_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3745__T_4012_data = _T_3745[_T_3745__T_4012_addr];
  `else
  assign _T_3745__T_4012_data = _T_3745__T_4012_addr >= 6'h28 ? _RAND_550[0:0] : _T_3745[_T_3745__T_4012_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3745__T_3768_data = io_enq_uops_0_exception;
  assign _T_3745__T_3768_addr = rob_tail;
  assign _T_3745__T_3768_mask = io_enq_valids_0;
  assign _T_3745__T_3768_en = io_enq_valids_0;
  assign _T_3745__T_3998_data = 1'h1;
  assign _T_3745__T_3998_addr = _T_3997;
  assign _T_3745__T_3998_mask = _T_3994;
  assign _T_3745__T_3998_en = _T_3994;
  assign _T_3745__T_4007_data = 1'h1;
  assign _T_3745__T_4007_addr = _T_4006;
  assign _T_3745__T_4007_mask = _T_4003;
  assign _T_3745__T_4007_en = _T_4003;
  assign _T_3745__T_4088_data = 1'h0;
  assign _T_3745__T_4088_addr = _T_4025;
  assign _T_3745__T_4088_mask = _T_4077;
  assign _T_3745__T_4088_en = _T_4077;
  assign _T_3748__T_5017_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3748__T_5017_data = _T_3748[_T_3748__T_5017_addr];
  `else
  assign _T_3748__T_5017_data = _T_3748__T_5017_addr >= 6'h28 ? _RAND_552[4:0] : _T_3748[_T_3748__T_5017_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3748__T_3769_data = 5'h0;
  assign _T_3748__T_3769_addr = rob_tail;
  assign _T_3748__T_3769_mask = io_enq_valids_0;
  assign _T_3748__T_3769_en = io_enq_valids_0;
  assign _T_3748__T_3982_data = io_fflags_0_bits_flags;
  assign _T_3748__T_3982_addr = _T_3981;
  assign _T_3748__T_3982_mask = _T_3978;
  assign _T_3748__T_3982_en = _T_3978;
  assign _T_3748__T_3990_data = io_fflags_1_bits_flags;
  assign _T_3748__T_3990_addr = _T_3989;
  assign _T_3748__T_3990_mask = _T_3986;
  assign _T_3748__T_3990_en = _T_3986;
  assign _GEN_575 = 6'h0 == rob_tail ? 1'h1 : _T_3073_0;
  assign _GEN_576 = 6'h1 == rob_tail ? 1'h1 : _T_3073_1;
  assign _GEN_577 = 6'h2 == rob_tail ? 1'h1 : _T_3073_2;
  assign _GEN_578 = 6'h3 == rob_tail ? 1'h1 : _T_3073_3;
  assign _GEN_579 = 6'h4 == rob_tail ? 1'h1 : _T_3073_4;
  assign _GEN_580 = 6'h5 == rob_tail ? 1'h1 : _T_3073_5;
  assign _GEN_581 = 6'h6 == rob_tail ? 1'h1 : _T_3073_6;
  assign _GEN_582 = 6'h7 == rob_tail ? 1'h1 : _T_3073_7;
  assign _GEN_583 = 6'h8 == rob_tail ? 1'h1 : _T_3073_8;
  assign _GEN_584 = 6'h9 == rob_tail ? 1'h1 : _T_3073_9;
  assign _GEN_585 = 6'ha == rob_tail ? 1'h1 : _T_3073_10;
  assign _GEN_586 = 6'hb == rob_tail ? 1'h1 : _T_3073_11;
  assign _GEN_587 = 6'hc == rob_tail ? 1'h1 : _T_3073_12;
  assign _GEN_588 = 6'hd == rob_tail ? 1'h1 : _T_3073_13;
  assign _GEN_589 = 6'he == rob_tail ? 1'h1 : _T_3073_14;
  assign _GEN_590 = 6'hf == rob_tail ? 1'h1 : _T_3073_15;
  assign _GEN_591 = 6'h10 == rob_tail ? 1'h1 : _T_3073_16;
  assign _GEN_592 = 6'h11 == rob_tail ? 1'h1 : _T_3073_17;
  assign _GEN_593 = 6'h12 == rob_tail ? 1'h1 : _T_3073_18;
  assign _GEN_594 = 6'h13 == rob_tail ? 1'h1 : _T_3073_19;
  assign _GEN_595 = 6'h14 == rob_tail ? 1'h1 : _T_3073_20;
  assign _GEN_596 = 6'h15 == rob_tail ? 1'h1 : _T_3073_21;
  assign _GEN_597 = 6'h16 == rob_tail ? 1'h1 : _T_3073_22;
  assign _GEN_598 = 6'h17 == rob_tail ? 1'h1 : _T_3073_23;
  assign _GEN_599 = 6'h18 == rob_tail ? 1'h1 : _T_3073_24;
  assign _GEN_600 = 6'h19 == rob_tail ? 1'h1 : _T_3073_25;
  assign _GEN_601 = 6'h1a == rob_tail ? 1'h1 : _T_3073_26;
  assign _GEN_602 = 6'h1b == rob_tail ? 1'h1 : _T_3073_27;
  assign _GEN_603 = 6'h1c == rob_tail ? 1'h1 : _T_3073_28;
  assign _GEN_604 = 6'h1d == rob_tail ? 1'h1 : _T_3073_29;
  assign _GEN_605 = 6'h1e == rob_tail ? 1'h1 : _T_3073_30;
  assign _GEN_606 = 6'h1f == rob_tail ? 1'h1 : _T_3073_31;
  assign _GEN_607 = 6'h20 == rob_tail ? 1'h1 : _T_3073_32;
  assign _GEN_608 = 6'h21 == rob_tail ? 1'h1 : _T_3073_33;
  assign _GEN_609 = 6'h22 == rob_tail ? 1'h1 : _T_3073_34;
  assign _GEN_610 = 6'h23 == rob_tail ? 1'h1 : _T_3073_35;
  assign _GEN_611 = 6'h24 == rob_tail ? 1'h1 : _T_3073_36;
  assign _GEN_612 = 6'h25 == rob_tail ? 1'h1 : _T_3073_37;
  assign _GEN_613 = 6'h26 == rob_tail ? 1'h1 : _T_3073_38;
  assign _GEN_614 = 6'h27 == rob_tail ? 1'h1 : _T_3073_39;
  assign _T_3755 = io_enq_uops_0_is_fence == 1'h0;
  assign _T_3757 = io_enq_uops_0_is_fencei == 1'h0;
  assign _T_3758 = _T_3755 & _T_3757;
  assign _GEN_1575 = 6'h0 == rob_tail ? _GEN_26 : _T_3372_0_br_mask;
  assign _GEN_1576 = 6'h1 == rob_tail ? _GEN_26 : _T_3372_1_br_mask;
  assign _GEN_1577 = 6'h2 == rob_tail ? _GEN_26 : _T_3372_2_br_mask;
  assign _GEN_1578 = 6'h3 == rob_tail ? _GEN_26 : _T_3372_3_br_mask;
  assign _GEN_1579 = 6'h4 == rob_tail ? _GEN_26 : _T_3372_4_br_mask;
  assign _GEN_1580 = 6'h5 == rob_tail ? _GEN_26 : _T_3372_5_br_mask;
  assign _GEN_1581 = 6'h6 == rob_tail ? _GEN_26 : _T_3372_6_br_mask;
  assign _GEN_1582 = 6'h7 == rob_tail ? _GEN_26 : _T_3372_7_br_mask;
  assign _GEN_1583 = 6'h8 == rob_tail ? _GEN_26 : _T_3372_8_br_mask;
  assign _GEN_1584 = 6'h9 == rob_tail ? _GEN_26 : _T_3372_9_br_mask;
  assign _GEN_1585 = 6'ha == rob_tail ? _GEN_26 : _T_3372_10_br_mask;
  assign _GEN_1586 = 6'hb == rob_tail ? _GEN_26 : _T_3372_11_br_mask;
  assign _GEN_1587 = 6'hc == rob_tail ? _GEN_26 : _T_3372_12_br_mask;
  assign _GEN_1588 = 6'hd == rob_tail ? _GEN_26 : _T_3372_13_br_mask;
  assign _GEN_1589 = 6'he == rob_tail ? _GEN_26 : _T_3372_14_br_mask;
  assign _GEN_1590 = 6'hf == rob_tail ? _GEN_26 : _T_3372_15_br_mask;
  assign _GEN_1591 = 6'h10 == rob_tail ? _GEN_26 : _T_3372_16_br_mask;
  assign _GEN_1592 = 6'h11 == rob_tail ? _GEN_26 : _T_3372_17_br_mask;
  assign _GEN_1593 = 6'h12 == rob_tail ? _GEN_26 : _T_3372_18_br_mask;
  assign _GEN_1594 = 6'h13 == rob_tail ? _GEN_26 : _T_3372_19_br_mask;
  assign _GEN_1595 = 6'h14 == rob_tail ? _GEN_26 : _T_3372_20_br_mask;
  assign _GEN_1596 = 6'h15 == rob_tail ? _GEN_26 : _T_3372_21_br_mask;
  assign _GEN_1597 = 6'h16 == rob_tail ? _GEN_26 : _T_3372_22_br_mask;
  assign _GEN_1598 = 6'h17 == rob_tail ? _GEN_26 : _T_3372_23_br_mask;
  assign _GEN_1599 = 6'h18 == rob_tail ? _GEN_26 : _T_3372_24_br_mask;
  assign _GEN_1600 = 6'h19 == rob_tail ? _GEN_26 : _T_3372_25_br_mask;
  assign _GEN_1601 = 6'h1a == rob_tail ? _GEN_26 : _T_3372_26_br_mask;
  assign _GEN_1602 = 6'h1b == rob_tail ? _GEN_26 : _T_3372_27_br_mask;
  assign _GEN_1603 = 6'h1c == rob_tail ? _GEN_26 : _T_3372_28_br_mask;
  assign _GEN_1604 = 6'h1d == rob_tail ? _GEN_26 : _T_3372_29_br_mask;
  assign _GEN_1605 = 6'h1e == rob_tail ? _GEN_26 : _T_3372_30_br_mask;
  assign _GEN_1606 = 6'h1f == rob_tail ? _GEN_26 : _T_3372_31_br_mask;
  assign _GEN_1607 = 6'h20 == rob_tail ? _GEN_26 : _T_3372_32_br_mask;
  assign _GEN_1608 = 6'h21 == rob_tail ? _GEN_26 : _T_3372_33_br_mask;
  assign _GEN_1609 = 6'h22 == rob_tail ? _GEN_26 : _T_3372_34_br_mask;
  assign _GEN_1610 = 6'h23 == rob_tail ? _GEN_26 : _T_3372_35_br_mask;
  assign _GEN_1611 = 6'h24 == rob_tail ? _GEN_26 : _T_3372_36_br_mask;
  assign _GEN_1612 = 6'h25 == rob_tail ? _GEN_26 : _T_3372_37_br_mask;
  assign _GEN_1613 = 6'h26 == rob_tail ? _GEN_26 : _T_3372_38_br_mask;
  assign _GEN_1614 = 6'h27 == rob_tail ? _GEN_26 : _T_3372_39_br_mask;
  assign _GEN_2695 = 6'h0 == rob_tail ? _GEN_54 : _T_3372_0_pdst;
  assign _GEN_2696 = 6'h1 == rob_tail ? _GEN_54 : _T_3372_1_pdst;
  assign _GEN_2697 = 6'h2 == rob_tail ? _GEN_54 : _T_3372_2_pdst;
  assign _GEN_2698 = 6'h3 == rob_tail ? _GEN_54 : _T_3372_3_pdst;
  assign _GEN_2699 = 6'h4 == rob_tail ? _GEN_54 : _T_3372_4_pdst;
  assign _GEN_2700 = 6'h5 == rob_tail ? _GEN_54 : _T_3372_5_pdst;
  assign _GEN_2701 = 6'h6 == rob_tail ? _GEN_54 : _T_3372_6_pdst;
  assign _GEN_2702 = 6'h7 == rob_tail ? _GEN_54 : _T_3372_7_pdst;
  assign _GEN_2703 = 6'h8 == rob_tail ? _GEN_54 : _T_3372_8_pdst;
  assign _GEN_2704 = 6'h9 == rob_tail ? _GEN_54 : _T_3372_9_pdst;
  assign _GEN_2705 = 6'ha == rob_tail ? _GEN_54 : _T_3372_10_pdst;
  assign _GEN_2706 = 6'hb == rob_tail ? _GEN_54 : _T_3372_11_pdst;
  assign _GEN_2707 = 6'hc == rob_tail ? _GEN_54 : _T_3372_12_pdst;
  assign _GEN_2708 = 6'hd == rob_tail ? _GEN_54 : _T_3372_13_pdst;
  assign _GEN_2709 = 6'he == rob_tail ? _GEN_54 : _T_3372_14_pdst;
  assign _GEN_2710 = 6'hf == rob_tail ? _GEN_54 : _T_3372_15_pdst;
  assign _GEN_2711 = 6'h10 == rob_tail ? _GEN_54 : _T_3372_16_pdst;
  assign _GEN_2712 = 6'h11 == rob_tail ? _GEN_54 : _T_3372_17_pdst;
  assign _GEN_2713 = 6'h12 == rob_tail ? _GEN_54 : _T_3372_18_pdst;
  assign _GEN_2714 = 6'h13 == rob_tail ? _GEN_54 : _T_3372_19_pdst;
  assign _GEN_2715 = 6'h14 == rob_tail ? _GEN_54 : _T_3372_20_pdst;
  assign _GEN_2716 = 6'h15 == rob_tail ? _GEN_54 : _T_3372_21_pdst;
  assign _GEN_2717 = 6'h16 == rob_tail ? _GEN_54 : _T_3372_22_pdst;
  assign _GEN_2718 = 6'h17 == rob_tail ? _GEN_54 : _T_3372_23_pdst;
  assign _GEN_2719 = 6'h18 == rob_tail ? _GEN_54 : _T_3372_24_pdst;
  assign _GEN_2720 = 6'h19 == rob_tail ? _GEN_54 : _T_3372_25_pdst;
  assign _GEN_2721 = 6'h1a == rob_tail ? _GEN_54 : _T_3372_26_pdst;
  assign _GEN_2722 = 6'h1b == rob_tail ? _GEN_54 : _T_3372_27_pdst;
  assign _GEN_2723 = 6'h1c == rob_tail ? _GEN_54 : _T_3372_28_pdst;
  assign _GEN_2724 = 6'h1d == rob_tail ? _GEN_54 : _T_3372_29_pdst;
  assign _GEN_2725 = 6'h1e == rob_tail ? _GEN_54 : _T_3372_30_pdst;
  assign _GEN_2726 = 6'h1f == rob_tail ? _GEN_54 : _T_3372_31_pdst;
  assign _GEN_2727 = 6'h20 == rob_tail ? _GEN_54 : _T_3372_32_pdst;
  assign _GEN_2728 = 6'h21 == rob_tail ? _GEN_54 : _T_3372_33_pdst;
  assign _GEN_2729 = 6'h22 == rob_tail ? _GEN_54 : _T_3372_34_pdst;
  assign _GEN_2730 = 6'h23 == rob_tail ? _GEN_54 : _T_3372_35_pdst;
  assign _GEN_2731 = 6'h24 == rob_tail ? _GEN_54 : _T_3372_36_pdst;
  assign _GEN_2732 = 6'h25 == rob_tail ? _GEN_54 : _T_3372_37_pdst;
  assign _GEN_2733 = 6'h26 == rob_tail ? _GEN_54 : _T_3372_38_pdst;
  assign _GEN_2734 = 6'h27 == rob_tail ? _GEN_54 : _T_3372_39_pdst;
  assign _GEN_2975 = 6'h0 == rob_tail ? _GEN_61 : _T_3372_0_stale_pdst;
  assign _GEN_2976 = 6'h1 == rob_tail ? _GEN_61 : _T_3372_1_stale_pdst;
  assign _GEN_2977 = 6'h2 == rob_tail ? _GEN_61 : _T_3372_2_stale_pdst;
  assign _GEN_2978 = 6'h3 == rob_tail ? _GEN_61 : _T_3372_3_stale_pdst;
  assign _GEN_2979 = 6'h4 == rob_tail ? _GEN_61 : _T_3372_4_stale_pdst;
  assign _GEN_2980 = 6'h5 == rob_tail ? _GEN_61 : _T_3372_5_stale_pdst;
  assign _GEN_2981 = 6'h6 == rob_tail ? _GEN_61 : _T_3372_6_stale_pdst;
  assign _GEN_2982 = 6'h7 == rob_tail ? _GEN_61 : _T_3372_7_stale_pdst;
  assign _GEN_2983 = 6'h8 == rob_tail ? _GEN_61 : _T_3372_8_stale_pdst;
  assign _GEN_2984 = 6'h9 == rob_tail ? _GEN_61 : _T_3372_9_stale_pdst;
  assign _GEN_2985 = 6'ha == rob_tail ? _GEN_61 : _T_3372_10_stale_pdst;
  assign _GEN_2986 = 6'hb == rob_tail ? _GEN_61 : _T_3372_11_stale_pdst;
  assign _GEN_2987 = 6'hc == rob_tail ? _GEN_61 : _T_3372_12_stale_pdst;
  assign _GEN_2988 = 6'hd == rob_tail ? _GEN_61 : _T_3372_13_stale_pdst;
  assign _GEN_2989 = 6'he == rob_tail ? _GEN_61 : _T_3372_14_stale_pdst;
  assign _GEN_2990 = 6'hf == rob_tail ? _GEN_61 : _T_3372_15_stale_pdst;
  assign _GEN_2991 = 6'h10 == rob_tail ? _GEN_61 : _T_3372_16_stale_pdst;
  assign _GEN_2992 = 6'h11 == rob_tail ? _GEN_61 : _T_3372_17_stale_pdst;
  assign _GEN_2993 = 6'h12 == rob_tail ? _GEN_61 : _T_3372_18_stale_pdst;
  assign _GEN_2994 = 6'h13 == rob_tail ? _GEN_61 : _T_3372_19_stale_pdst;
  assign _GEN_2995 = 6'h14 == rob_tail ? _GEN_61 : _T_3372_20_stale_pdst;
  assign _GEN_2996 = 6'h15 == rob_tail ? _GEN_61 : _T_3372_21_stale_pdst;
  assign _GEN_2997 = 6'h16 == rob_tail ? _GEN_61 : _T_3372_22_stale_pdst;
  assign _GEN_2998 = 6'h17 == rob_tail ? _GEN_61 : _T_3372_23_stale_pdst;
  assign _GEN_2999 = 6'h18 == rob_tail ? _GEN_61 : _T_3372_24_stale_pdst;
  assign _GEN_3000 = 6'h19 == rob_tail ? _GEN_61 : _T_3372_25_stale_pdst;
  assign _GEN_3001 = 6'h1a == rob_tail ? _GEN_61 : _T_3372_26_stale_pdst;
  assign _GEN_3002 = 6'h1b == rob_tail ? _GEN_61 : _T_3372_27_stale_pdst;
  assign _GEN_3003 = 6'h1c == rob_tail ? _GEN_61 : _T_3372_28_stale_pdst;
  assign _GEN_3004 = 6'h1d == rob_tail ? _GEN_61 : _T_3372_29_stale_pdst;
  assign _GEN_3005 = 6'h1e == rob_tail ? _GEN_61 : _T_3372_30_stale_pdst;
  assign _GEN_3006 = 6'h1f == rob_tail ? _GEN_61 : _T_3372_31_stale_pdst;
  assign _GEN_3007 = 6'h20 == rob_tail ? _GEN_61 : _T_3372_32_stale_pdst;
  assign _GEN_3008 = 6'h21 == rob_tail ? _GEN_61 : _T_3372_33_stale_pdst;
  assign _GEN_3009 = 6'h22 == rob_tail ? _GEN_61 : _T_3372_34_stale_pdst;
  assign _GEN_3010 = 6'h23 == rob_tail ? _GEN_61 : _T_3372_35_stale_pdst;
  assign _GEN_3011 = 6'h24 == rob_tail ? _GEN_61 : _T_3372_36_stale_pdst;
  assign _GEN_3012 = 6'h25 == rob_tail ? _GEN_61 : _T_3372_37_stale_pdst;
  assign _GEN_3013 = 6'h26 == rob_tail ? _GEN_61 : _T_3372_38_stale_pdst;
  assign _GEN_3014 = 6'h27 == rob_tail ? _GEN_61 : _T_3372_39_stale_pdst;
  assign _GEN_3255 = 6'h0 == rob_tail ? _GEN_68 : _T_3372_0_is_fencei;
  assign _GEN_3256 = 6'h1 == rob_tail ? _GEN_68 : _T_3372_1_is_fencei;
  assign _GEN_3257 = 6'h2 == rob_tail ? _GEN_68 : _T_3372_2_is_fencei;
  assign _GEN_3258 = 6'h3 == rob_tail ? _GEN_68 : _T_3372_3_is_fencei;
  assign _GEN_3259 = 6'h4 == rob_tail ? _GEN_68 : _T_3372_4_is_fencei;
  assign _GEN_3260 = 6'h5 == rob_tail ? _GEN_68 : _T_3372_5_is_fencei;
  assign _GEN_3261 = 6'h6 == rob_tail ? _GEN_68 : _T_3372_6_is_fencei;
  assign _GEN_3262 = 6'h7 == rob_tail ? _GEN_68 : _T_3372_7_is_fencei;
  assign _GEN_3263 = 6'h8 == rob_tail ? _GEN_68 : _T_3372_8_is_fencei;
  assign _GEN_3264 = 6'h9 == rob_tail ? _GEN_68 : _T_3372_9_is_fencei;
  assign _GEN_3265 = 6'ha == rob_tail ? _GEN_68 : _T_3372_10_is_fencei;
  assign _GEN_3266 = 6'hb == rob_tail ? _GEN_68 : _T_3372_11_is_fencei;
  assign _GEN_3267 = 6'hc == rob_tail ? _GEN_68 : _T_3372_12_is_fencei;
  assign _GEN_3268 = 6'hd == rob_tail ? _GEN_68 : _T_3372_13_is_fencei;
  assign _GEN_3269 = 6'he == rob_tail ? _GEN_68 : _T_3372_14_is_fencei;
  assign _GEN_3270 = 6'hf == rob_tail ? _GEN_68 : _T_3372_15_is_fencei;
  assign _GEN_3271 = 6'h10 == rob_tail ? _GEN_68 : _T_3372_16_is_fencei;
  assign _GEN_3272 = 6'h11 == rob_tail ? _GEN_68 : _T_3372_17_is_fencei;
  assign _GEN_3273 = 6'h12 == rob_tail ? _GEN_68 : _T_3372_18_is_fencei;
  assign _GEN_3274 = 6'h13 == rob_tail ? _GEN_68 : _T_3372_19_is_fencei;
  assign _GEN_3275 = 6'h14 == rob_tail ? _GEN_68 : _T_3372_20_is_fencei;
  assign _GEN_3276 = 6'h15 == rob_tail ? _GEN_68 : _T_3372_21_is_fencei;
  assign _GEN_3277 = 6'h16 == rob_tail ? _GEN_68 : _T_3372_22_is_fencei;
  assign _GEN_3278 = 6'h17 == rob_tail ? _GEN_68 : _T_3372_23_is_fencei;
  assign _GEN_3279 = 6'h18 == rob_tail ? _GEN_68 : _T_3372_24_is_fencei;
  assign _GEN_3280 = 6'h19 == rob_tail ? _GEN_68 : _T_3372_25_is_fencei;
  assign _GEN_3281 = 6'h1a == rob_tail ? _GEN_68 : _T_3372_26_is_fencei;
  assign _GEN_3282 = 6'h1b == rob_tail ? _GEN_68 : _T_3372_27_is_fencei;
  assign _GEN_3283 = 6'h1c == rob_tail ? _GEN_68 : _T_3372_28_is_fencei;
  assign _GEN_3284 = 6'h1d == rob_tail ? _GEN_68 : _T_3372_29_is_fencei;
  assign _GEN_3285 = 6'h1e == rob_tail ? _GEN_68 : _T_3372_30_is_fencei;
  assign _GEN_3286 = 6'h1f == rob_tail ? _GEN_68 : _T_3372_31_is_fencei;
  assign _GEN_3287 = 6'h20 == rob_tail ? _GEN_68 : _T_3372_32_is_fencei;
  assign _GEN_3288 = 6'h21 == rob_tail ? _GEN_68 : _T_3372_33_is_fencei;
  assign _GEN_3289 = 6'h22 == rob_tail ? _GEN_68 : _T_3372_34_is_fencei;
  assign _GEN_3290 = 6'h23 == rob_tail ? _GEN_68 : _T_3372_35_is_fencei;
  assign _GEN_3291 = 6'h24 == rob_tail ? _GEN_68 : _T_3372_36_is_fencei;
  assign _GEN_3292 = 6'h25 == rob_tail ? _GEN_68 : _T_3372_37_is_fencei;
  assign _GEN_3293 = 6'h26 == rob_tail ? _GEN_68 : _T_3372_38_is_fencei;
  assign _GEN_3294 = 6'h27 == rob_tail ? _GEN_68 : _T_3372_39_is_fencei;
  assign _GEN_3295 = 6'h0 == rob_tail ? _GEN_69 : _T_3372_0_is_store;
  assign _GEN_3296 = 6'h1 == rob_tail ? _GEN_69 : _T_3372_1_is_store;
  assign _GEN_3297 = 6'h2 == rob_tail ? _GEN_69 : _T_3372_2_is_store;
  assign _GEN_3298 = 6'h3 == rob_tail ? _GEN_69 : _T_3372_3_is_store;
  assign _GEN_3299 = 6'h4 == rob_tail ? _GEN_69 : _T_3372_4_is_store;
  assign _GEN_3300 = 6'h5 == rob_tail ? _GEN_69 : _T_3372_5_is_store;
  assign _GEN_3301 = 6'h6 == rob_tail ? _GEN_69 : _T_3372_6_is_store;
  assign _GEN_3302 = 6'h7 == rob_tail ? _GEN_69 : _T_3372_7_is_store;
  assign _GEN_3303 = 6'h8 == rob_tail ? _GEN_69 : _T_3372_8_is_store;
  assign _GEN_3304 = 6'h9 == rob_tail ? _GEN_69 : _T_3372_9_is_store;
  assign _GEN_3305 = 6'ha == rob_tail ? _GEN_69 : _T_3372_10_is_store;
  assign _GEN_3306 = 6'hb == rob_tail ? _GEN_69 : _T_3372_11_is_store;
  assign _GEN_3307 = 6'hc == rob_tail ? _GEN_69 : _T_3372_12_is_store;
  assign _GEN_3308 = 6'hd == rob_tail ? _GEN_69 : _T_3372_13_is_store;
  assign _GEN_3309 = 6'he == rob_tail ? _GEN_69 : _T_3372_14_is_store;
  assign _GEN_3310 = 6'hf == rob_tail ? _GEN_69 : _T_3372_15_is_store;
  assign _GEN_3311 = 6'h10 == rob_tail ? _GEN_69 : _T_3372_16_is_store;
  assign _GEN_3312 = 6'h11 == rob_tail ? _GEN_69 : _T_3372_17_is_store;
  assign _GEN_3313 = 6'h12 == rob_tail ? _GEN_69 : _T_3372_18_is_store;
  assign _GEN_3314 = 6'h13 == rob_tail ? _GEN_69 : _T_3372_19_is_store;
  assign _GEN_3315 = 6'h14 == rob_tail ? _GEN_69 : _T_3372_20_is_store;
  assign _GEN_3316 = 6'h15 == rob_tail ? _GEN_69 : _T_3372_21_is_store;
  assign _GEN_3317 = 6'h16 == rob_tail ? _GEN_69 : _T_3372_22_is_store;
  assign _GEN_3318 = 6'h17 == rob_tail ? _GEN_69 : _T_3372_23_is_store;
  assign _GEN_3319 = 6'h18 == rob_tail ? _GEN_69 : _T_3372_24_is_store;
  assign _GEN_3320 = 6'h19 == rob_tail ? _GEN_69 : _T_3372_25_is_store;
  assign _GEN_3321 = 6'h1a == rob_tail ? _GEN_69 : _T_3372_26_is_store;
  assign _GEN_3322 = 6'h1b == rob_tail ? _GEN_69 : _T_3372_27_is_store;
  assign _GEN_3323 = 6'h1c == rob_tail ? _GEN_69 : _T_3372_28_is_store;
  assign _GEN_3324 = 6'h1d == rob_tail ? _GEN_69 : _T_3372_29_is_store;
  assign _GEN_3325 = 6'h1e == rob_tail ? _GEN_69 : _T_3372_30_is_store;
  assign _GEN_3326 = 6'h1f == rob_tail ? _GEN_69 : _T_3372_31_is_store;
  assign _GEN_3327 = 6'h20 == rob_tail ? _GEN_69 : _T_3372_32_is_store;
  assign _GEN_3328 = 6'h21 == rob_tail ? _GEN_69 : _T_3372_33_is_store;
  assign _GEN_3329 = 6'h22 == rob_tail ? _GEN_69 : _T_3372_34_is_store;
  assign _GEN_3330 = 6'h23 == rob_tail ? _GEN_69 : _T_3372_35_is_store;
  assign _GEN_3331 = 6'h24 == rob_tail ? _GEN_69 : _T_3372_36_is_store;
  assign _GEN_3332 = 6'h25 == rob_tail ? _GEN_69 : _T_3372_37_is_store;
  assign _GEN_3333 = 6'h26 == rob_tail ? _GEN_69 : _T_3372_38_is_store;
  assign _GEN_3334 = 6'h27 == rob_tail ? _GEN_69 : _T_3372_39_is_store;
  assign _GEN_3375 = 6'h0 == rob_tail ? _GEN_71 : _T_3372_0_is_load;
  assign _GEN_3376 = 6'h1 == rob_tail ? _GEN_71 : _T_3372_1_is_load;
  assign _GEN_3377 = 6'h2 == rob_tail ? _GEN_71 : _T_3372_2_is_load;
  assign _GEN_3378 = 6'h3 == rob_tail ? _GEN_71 : _T_3372_3_is_load;
  assign _GEN_3379 = 6'h4 == rob_tail ? _GEN_71 : _T_3372_4_is_load;
  assign _GEN_3380 = 6'h5 == rob_tail ? _GEN_71 : _T_3372_5_is_load;
  assign _GEN_3381 = 6'h6 == rob_tail ? _GEN_71 : _T_3372_6_is_load;
  assign _GEN_3382 = 6'h7 == rob_tail ? _GEN_71 : _T_3372_7_is_load;
  assign _GEN_3383 = 6'h8 == rob_tail ? _GEN_71 : _T_3372_8_is_load;
  assign _GEN_3384 = 6'h9 == rob_tail ? _GEN_71 : _T_3372_9_is_load;
  assign _GEN_3385 = 6'ha == rob_tail ? _GEN_71 : _T_3372_10_is_load;
  assign _GEN_3386 = 6'hb == rob_tail ? _GEN_71 : _T_3372_11_is_load;
  assign _GEN_3387 = 6'hc == rob_tail ? _GEN_71 : _T_3372_12_is_load;
  assign _GEN_3388 = 6'hd == rob_tail ? _GEN_71 : _T_3372_13_is_load;
  assign _GEN_3389 = 6'he == rob_tail ? _GEN_71 : _T_3372_14_is_load;
  assign _GEN_3390 = 6'hf == rob_tail ? _GEN_71 : _T_3372_15_is_load;
  assign _GEN_3391 = 6'h10 == rob_tail ? _GEN_71 : _T_3372_16_is_load;
  assign _GEN_3392 = 6'h11 == rob_tail ? _GEN_71 : _T_3372_17_is_load;
  assign _GEN_3393 = 6'h12 == rob_tail ? _GEN_71 : _T_3372_18_is_load;
  assign _GEN_3394 = 6'h13 == rob_tail ? _GEN_71 : _T_3372_19_is_load;
  assign _GEN_3395 = 6'h14 == rob_tail ? _GEN_71 : _T_3372_20_is_load;
  assign _GEN_3396 = 6'h15 == rob_tail ? _GEN_71 : _T_3372_21_is_load;
  assign _GEN_3397 = 6'h16 == rob_tail ? _GEN_71 : _T_3372_22_is_load;
  assign _GEN_3398 = 6'h17 == rob_tail ? _GEN_71 : _T_3372_23_is_load;
  assign _GEN_3399 = 6'h18 == rob_tail ? _GEN_71 : _T_3372_24_is_load;
  assign _GEN_3400 = 6'h19 == rob_tail ? _GEN_71 : _T_3372_25_is_load;
  assign _GEN_3401 = 6'h1a == rob_tail ? _GEN_71 : _T_3372_26_is_load;
  assign _GEN_3402 = 6'h1b == rob_tail ? _GEN_71 : _T_3372_27_is_load;
  assign _GEN_3403 = 6'h1c == rob_tail ? _GEN_71 : _T_3372_28_is_load;
  assign _GEN_3404 = 6'h1d == rob_tail ? _GEN_71 : _T_3372_29_is_load;
  assign _GEN_3405 = 6'h1e == rob_tail ? _GEN_71 : _T_3372_30_is_load;
  assign _GEN_3406 = 6'h1f == rob_tail ? _GEN_71 : _T_3372_31_is_load;
  assign _GEN_3407 = 6'h20 == rob_tail ? _GEN_71 : _T_3372_32_is_load;
  assign _GEN_3408 = 6'h21 == rob_tail ? _GEN_71 : _T_3372_33_is_load;
  assign _GEN_3409 = 6'h22 == rob_tail ? _GEN_71 : _T_3372_34_is_load;
  assign _GEN_3410 = 6'h23 == rob_tail ? _GEN_71 : _T_3372_35_is_load;
  assign _GEN_3411 = 6'h24 == rob_tail ? _GEN_71 : _T_3372_36_is_load;
  assign _GEN_3412 = 6'h25 == rob_tail ? _GEN_71 : _T_3372_37_is_load;
  assign _GEN_3413 = 6'h26 == rob_tail ? _GEN_71 : _T_3372_38_is_load;
  assign _GEN_3414 = 6'h27 == rob_tail ? _GEN_71 : _T_3372_39_is_load;
  assign _GEN_3415 = 6'h0 == rob_tail ? _GEN_72 : _T_3372_0_is_sys_pc2epc;
  assign _GEN_3416 = 6'h1 == rob_tail ? _GEN_72 : _T_3372_1_is_sys_pc2epc;
  assign _GEN_3417 = 6'h2 == rob_tail ? _GEN_72 : _T_3372_2_is_sys_pc2epc;
  assign _GEN_3418 = 6'h3 == rob_tail ? _GEN_72 : _T_3372_3_is_sys_pc2epc;
  assign _GEN_3419 = 6'h4 == rob_tail ? _GEN_72 : _T_3372_4_is_sys_pc2epc;
  assign _GEN_3420 = 6'h5 == rob_tail ? _GEN_72 : _T_3372_5_is_sys_pc2epc;
  assign _GEN_3421 = 6'h6 == rob_tail ? _GEN_72 : _T_3372_6_is_sys_pc2epc;
  assign _GEN_3422 = 6'h7 == rob_tail ? _GEN_72 : _T_3372_7_is_sys_pc2epc;
  assign _GEN_3423 = 6'h8 == rob_tail ? _GEN_72 : _T_3372_8_is_sys_pc2epc;
  assign _GEN_3424 = 6'h9 == rob_tail ? _GEN_72 : _T_3372_9_is_sys_pc2epc;
  assign _GEN_3425 = 6'ha == rob_tail ? _GEN_72 : _T_3372_10_is_sys_pc2epc;
  assign _GEN_3426 = 6'hb == rob_tail ? _GEN_72 : _T_3372_11_is_sys_pc2epc;
  assign _GEN_3427 = 6'hc == rob_tail ? _GEN_72 : _T_3372_12_is_sys_pc2epc;
  assign _GEN_3428 = 6'hd == rob_tail ? _GEN_72 : _T_3372_13_is_sys_pc2epc;
  assign _GEN_3429 = 6'he == rob_tail ? _GEN_72 : _T_3372_14_is_sys_pc2epc;
  assign _GEN_3430 = 6'hf == rob_tail ? _GEN_72 : _T_3372_15_is_sys_pc2epc;
  assign _GEN_3431 = 6'h10 == rob_tail ? _GEN_72 : _T_3372_16_is_sys_pc2epc;
  assign _GEN_3432 = 6'h11 == rob_tail ? _GEN_72 : _T_3372_17_is_sys_pc2epc;
  assign _GEN_3433 = 6'h12 == rob_tail ? _GEN_72 : _T_3372_18_is_sys_pc2epc;
  assign _GEN_3434 = 6'h13 == rob_tail ? _GEN_72 : _T_3372_19_is_sys_pc2epc;
  assign _GEN_3435 = 6'h14 == rob_tail ? _GEN_72 : _T_3372_20_is_sys_pc2epc;
  assign _GEN_3436 = 6'h15 == rob_tail ? _GEN_72 : _T_3372_21_is_sys_pc2epc;
  assign _GEN_3437 = 6'h16 == rob_tail ? _GEN_72 : _T_3372_22_is_sys_pc2epc;
  assign _GEN_3438 = 6'h17 == rob_tail ? _GEN_72 : _T_3372_23_is_sys_pc2epc;
  assign _GEN_3439 = 6'h18 == rob_tail ? _GEN_72 : _T_3372_24_is_sys_pc2epc;
  assign _GEN_3440 = 6'h19 == rob_tail ? _GEN_72 : _T_3372_25_is_sys_pc2epc;
  assign _GEN_3441 = 6'h1a == rob_tail ? _GEN_72 : _T_3372_26_is_sys_pc2epc;
  assign _GEN_3442 = 6'h1b == rob_tail ? _GEN_72 : _T_3372_27_is_sys_pc2epc;
  assign _GEN_3443 = 6'h1c == rob_tail ? _GEN_72 : _T_3372_28_is_sys_pc2epc;
  assign _GEN_3444 = 6'h1d == rob_tail ? _GEN_72 : _T_3372_29_is_sys_pc2epc;
  assign _GEN_3445 = 6'h1e == rob_tail ? _GEN_72 : _T_3372_30_is_sys_pc2epc;
  assign _GEN_3446 = 6'h1f == rob_tail ? _GEN_72 : _T_3372_31_is_sys_pc2epc;
  assign _GEN_3447 = 6'h20 == rob_tail ? _GEN_72 : _T_3372_32_is_sys_pc2epc;
  assign _GEN_3448 = 6'h21 == rob_tail ? _GEN_72 : _T_3372_33_is_sys_pc2epc;
  assign _GEN_3449 = 6'h22 == rob_tail ? _GEN_72 : _T_3372_34_is_sys_pc2epc;
  assign _GEN_3450 = 6'h23 == rob_tail ? _GEN_72 : _T_3372_35_is_sys_pc2epc;
  assign _GEN_3451 = 6'h24 == rob_tail ? _GEN_72 : _T_3372_36_is_sys_pc2epc;
  assign _GEN_3452 = 6'h25 == rob_tail ? _GEN_72 : _T_3372_37_is_sys_pc2epc;
  assign _GEN_3453 = 6'h26 == rob_tail ? _GEN_72 : _T_3372_38_is_sys_pc2epc;
  assign _GEN_3454 = 6'h27 == rob_tail ? _GEN_72 : _T_3372_39_is_sys_pc2epc;
  assign _GEN_3495 = 6'h0 == rob_tail ? _GEN_74 : _T_3372_0_flush_on_commit;
  assign _GEN_3496 = 6'h1 == rob_tail ? _GEN_74 : _T_3372_1_flush_on_commit;
  assign _GEN_3497 = 6'h2 == rob_tail ? _GEN_74 : _T_3372_2_flush_on_commit;
  assign _GEN_3498 = 6'h3 == rob_tail ? _GEN_74 : _T_3372_3_flush_on_commit;
  assign _GEN_3499 = 6'h4 == rob_tail ? _GEN_74 : _T_3372_4_flush_on_commit;
  assign _GEN_3500 = 6'h5 == rob_tail ? _GEN_74 : _T_3372_5_flush_on_commit;
  assign _GEN_3501 = 6'h6 == rob_tail ? _GEN_74 : _T_3372_6_flush_on_commit;
  assign _GEN_3502 = 6'h7 == rob_tail ? _GEN_74 : _T_3372_7_flush_on_commit;
  assign _GEN_3503 = 6'h8 == rob_tail ? _GEN_74 : _T_3372_8_flush_on_commit;
  assign _GEN_3504 = 6'h9 == rob_tail ? _GEN_74 : _T_3372_9_flush_on_commit;
  assign _GEN_3505 = 6'ha == rob_tail ? _GEN_74 : _T_3372_10_flush_on_commit;
  assign _GEN_3506 = 6'hb == rob_tail ? _GEN_74 : _T_3372_11_flush_on_commit;
  assign _GEN_3507 = 6'hc == rob_tail ? _GEN_74 : _T_3372_12_flush_on_commit;
  assign _GEN_3508 = 6'hd == rob_tail ? _GEN_74 : _T_3372_13_flush_on_commit;
  assign _GEN_3509 = 6'he == rob_tail ? _GEN_74 : _T_3372_14_flush_on_commit;
  assign _GEN_3510 = 6'hf == rob_tail ? _GEN_74 : _T_3372_15_flush_on_commit;
  assign _GEN_3511 = 6'h10 == rob_tail ? _GEN_74 : _T_3372_16_flush_on_commit;
  assign _GEN_3512 = 6'h11 == rob_tail ? _GEN_74 : _T_3372_17_flush_on_commit;
  assign _GEN_3513 = 6'h12 == rob_tail ? _GEN_74 : _T_3372_18_flush_on_commit;
  assign _GEN_3514 = 6'h13 == rob_tail ? _GEN_74 : _T_3372_19_flush_on_commit;
  assign _GEN_3515 = 6'h14 == rob_tail ? _GEN_74 : _T_3372_20_flush_on_commit;
  assign _GEN_3516 = 6'h15 == rob_tail ? _GEN_74 : _T_3372_21_flush_on_commit;
  assign _GEN_3517 = 6'h16 == rob_tail ? _GEN_74 : _T_3372_22_flush_on_commit;
  assign _GEN_3518 = 6'h17 == rob_tail ? _GEN_74 : _T_3372_23_flush_on_commit;
  assign _GEN_3519 = 6'h18 == rob_tail ? _GEN_74 : _T_3372_24_flush_on_commit;
  assign _GEN_3520 = 6'h19 == rob_tail ? _GEN_74 : _T_3372_25_flush_on_commit;
  assign _GEN_3521 = 6'h1a == rob_tail ? _GEN_74 : _T_3372_26_flush_on_commit;
  assign _GEN_3522 = 6'h1b == rob_tail ? _GEN_74 : _T_3372_27_flush_on_commit;
  assign _GEN_3523 = 6'h1c == rob_tail ? _GEN_74 : _T_3372_28_flush_on_commit;
  assign _GEN_3524 = 6'h1d == rob_tail ? _GEN_74 : _T_3372_29_flush_on_commit;
  assign _GEN_3525 = 6'h1e == rob_tail ? _GEN_74 : _T_3372_30_flush_on_commit;
  assign _GEN_3526 = 6'h1f == rob_tail ? _GEN_74 : _T_3372_31_flush_on_commit;
  assign _GEN_3527 = 6'h20 == rob_tail ? _GEN_74 : _T_3372_32_flush_on_commit;
  assign _GEN_3528 = 6'h21 == rob_tail ? _GEN_74 : _T_3372_33_flush_on_commit;
  assign _GEN_3529 = 6'h22 == rob_tail ? _GEN_74 : _T_3372_34_flush_on_commit;
  assign _GEN_3530 = 6'h23 == rob_tail ? _GEN_74 : _T_3372_35_flush_on_commit;
  assign _GEN_3531 = 6'h24 == rob_tail ? _GEN_74 : _T_3372_36_flush_on_commit;
  assign _GEN_3532 = 6'h25 == rob_tail ? _GEN_74 : _T_3372_37_flush_on_commit;
  assign _GEN_3533 = 6'h26 == rob_tail ? _GEN_74 : _T_3372_38_flush_on_commit;
  assign _GEN_3534 = 6'h27 == rob_tail ? _GEN_74 : _T_3372_39_flush_on_commit;
  assign _GEN_3535 = 6'h0 == rob_tail ? _GEN_75 : _T_3372_0_ldst;
  assign _GEN_3536 = 6'h1 == rob_tail ? _GEN_75 : _T_3372_1_ldst;
  assign _GEN_3537 = 6'h2 == rob_tail ? _GEN_75 : _T_3372_2_ldst;
  assign _GEN_3538 = 6'h3 == rob_tail ? _GEN_75 : _T_3372_3_ldst;
  assign _GEN_3539 = 6'h4 == rob_tail ? _GEN_75 : _T_3372_4_ldst;
  assign _GEN_3540 = 6'h5 == rob_tail ? _GEN_75 : _T_3372_5_ldst;
  assign _GEN_3541 = 6'h6 == rob_tail ? _GEN_75 : _T_3372_6_ldst;
  assign _GEN_3542 = 6'h7 == rob_tail ? _GEN_75 : _T_3372_7_ldst;
  assign _GEN_3543 = 6'h8 == rob_tail ? _GEN_75 : _T_3372_8_ldst;
  assign _GEN_3544 = 6'h9 == rob_tail ? _GEN_75 : _T_3372_9_ldst;
  assign _GEN_3545 = 6'ha == rob_tail ? _GEN_75 : _T_3372_10_ldst;
  assign _GEN_3546 = 6'hb == rob_tail ? _GEN_75 : _T_3372_11_ldst;
  assign _GEN_3547 = 6'hc == rob_tail ? _GEN_75 : _T_3372_12_ldst;
  assign _GEN_3548 = 6'hd == rob_tail ? _GEN_75 : _T_3372_13_ldst;
  assign _GEN_3549 = 6'he == rob_tail ? _GEN_75 : _T_3372_14_ldst;
  assign _GEN_3550 = 6'hf == rob_tail ? _GEN_75 : _T_3372_15_ldst;
  assign _GEN_3551 = 6'h10 == rob_tail ? _GEN_75 : _T_3372_16_ldst;
  assign _GEN_3552 = 6'h11 == rob_tail ? _GEN_75 : _T_3372_17_ldst;
  assign _GEN_3553 = 6'h12 == rob_tail ? _GEN_75 : _T_3372_18_ldst;
  assign _GEN_3554 = 6'h13 == rob_tail ? _GEN_75 : _T_3372_19_ldst;
  assign _GEN_3555 = 6'h14 == rob_tail ? _GEN_75 : _T_3372_20_ldst;
  assign _GEN_3556 = 6'h15 == rob_tail ? _GEN_75 : _T_3372_21_ldst;
  assign _GEN_3557 = 6'h16 == rob_tail ? _GEN_75 : _T_3372_22_ldst;
  assign _GEN_3558 = 6'h17 == rob_tail ? _GEN_75 : _T_3372_23_ldst;
  assign _GEN_3559 = 6'h18 == rob_tail ? _GEN_75 : _T_3372_24_ldst;
  assign _GEN_3560 = 6'h19 == rob_tail ? _GEN_75 : _T_3372_25_ldst;
  assign _GEN_3561 = 6'h1a == rob_tail ? _GEN_75 : _T_3372_26_ldst;
  assign _GEN_3562 = 6'h1b == rob_tail ? _GEN_75 : _T_3372_27_ldst;
  assign _GEN_3563 = 6'h1c == rob_tail ? _GEN_75 : _T_3372_28_ldst;
  assign _GEN_3564 = 6'h1d == rob_tail ? _GEN_75 : _T_3372_29_ldst;
  assign _GEN_3565 = 6'h1e == rob_tail ? _GEN_75 : _T_3372_30_ldst;
  assign _GEN_3566 = 6'h1f == rob_tail ? _GEN_75 : _T_3372_31_ldst;
  assign _GEN_3567 = 6'h20 == rob_tail ? _GEN_75 : _T_3372_32_ldst;
  assign _GEN_3568 = 6'h21 == rob_tail ? _GEN_75 : _T_3372_33_ldst;
  assign _GEN_3569 = 6'h22 == rob_tail ? _GEN_75 : _T_3372_34_ldst;
  assign _GEN_3570 = 6'h23 == rob_tail ? _GEN_75 : _T_3372_35_ldst;
  assign _GEN_3571 = 6'h24 == rob_tail ? _GEN_75 : _T_3372_36_ldst;
  assign _GEN_3572 = 6'h25 == rob_tail ? _GEN_75 : _T_3372_37_ldst;
  assign _GEN_3573 = 6'h26 == rob_tail ? _GEN_75 : _T_3372_38_ldst;
  assign _GEN_3574 = 6'h27 == rob_tail ? _GEN_75 : _T_3372_39_ldst;
  assign _GEN_3695 = 6'h0 == rob_tail ? _GEN_79 : _T_3372_0_ldst_val;
  assign _GEN_3696 = 6'h1 == rob_tail ? _GEN_79 : _T_3372_1_ldst_val;
  assign _GEN_3697 = 6'h2 == rob_tail ? _GEN_79 : _T_3372_2_ldst_val;
  assign _GEN_3698 = 6'h3 == rob_tail ? _GEN_79 : _T_3372_3_ldst_val;
  assign _GEN_3699 = 6'h4 == rob_tail ? _GEN_79 : _T_3372_4_ldst_val;
  assign _GEN_3700 = 6'h5 == rob_tail ? _GEN_79 : _T_3372_5_ldst_val;
  assign _GEN_3701 = 6'h6 == rob_tail ? _GEN_79 : _T_3372_6_ldst_val;
  assign _GEN_3702 = 6'h7 == rob_tail ? _GEN_79 : _T_3372_7_ldst_val;
  assign _GEN_3703 = 6'h8 == rob_tail ? _GEN_79 : _T_3372_8_ldst_val;
  assign _GEN_3704 = 6'h9 == rob_tail ? _GEN_79 : _T_3372_9_ldst_val;
  assign _GEN_3705 = 6'ha == rob_tail ? _GEN_79 : _T_3372_10_ldst_val;
  assign _GEN_3706 = 6'hb == rob_tail ? _GEN_79 : _T_3372_11_ldst_val;
  assign _GEN_3707 = 6'hc == rob_tail ? _GEN_79 : _T_3372_12_ldst_val;
  assign _GEN_3708 = 6'hd == rob_tail ? _GEN_79 : _T_3372_13_ldst_val;
  assign _GEN_3709 = 6'he == rob_tail ? _GEN_79 : _T_3372_14_ldst_val;
  assign _GEN_3710 = 6'hf == rob_tail ? _GEN_79 : _T_3372_15_ldst_val;
  assign _GEN_3711 = 6'h10 == rob_tail ? _GEN_79 : _T_3372_16_ldst_val;
  assign _GEN_3712 = 6'h11 == rob_tail ? _GEN_79 : _T_3372_17_ldst_val;
  assign _GEN_3713 = 6'h12 == rob_tail ? _GEN_79 : _T_3372_18_ldst_val;
  assign _GEN_3714 = 6'h13 == rob_tail ? _GEN_79 : _T_3372_19_ldst_val;
  assign _GEN_3715 = 6'h14 == rob_tail ? _GEN_79 : _T_3372_20_ldst_val;
  assign _GEN_3716 = 6'h15 == rob_tail ? _GEN_79 : _T_3372_21_ldst_val;
  assign _GEN_3717 = 6'h16 == rob_tail ? _GEN_79 : _T_3372_22_ldst_val;
  assign _GEN_3718 = 6'h17 == rob_tail ? _GEN_79 : _T_3372_23_ldst_val;
  assign _GEN_3719 = 6'h18 == rob_tail ? _GEN_79 : _T_3372_24_ldst_val;
  assign _GEN_3720 = 6'h19 == rob_tail ? _GEN_79 : _T_3372_25_ldst_val;
  assign _GEN_3721 = 6'h1a == rob_tail ? _GEN_79 : _T_3372_26_ldst_val;
  assign _GEN_3722 = 6'h1b == rob_tail ? _GEN_79 : _T_3372_27_ldst_val;
  assign _GEN_3723 = 6'h1c == rob_tail ? _GEN_79 : _T_3372_28_ldst_val;
  assign _GEN_3724 = 6'h1d == rob_tail ? _GEN_79 : _T_3372_29_ldst_val;
  assign _GEN_3725 = 6'h1e == rob_tail ? _GEN_79 : _T_3372_30_ldst_val;
  assign _GEN_3726 = 6'h1f == rob_tail ? _GEN_79 : _T_3372_31_ldst_val;
  assign _GEN_3727 = 6'h20 == rob_tail ? _GEN_79 : _T_3372_32_ldst_val;
  assign _GEN_3728 = 6'h21 == rob_tail ? _GEN_79 : _T_3372_33_ldst_val;
  assign _GEN_3729 = 6'h22 == rob_tail ? _GEN_79 : _T_3372_34_ldst_val;
  assign _GEN_3730 = 6'h23 == rob_tail ? _GEN_79 : _T_3372_35_ldst_val;
  assign _GEN_3731 = 6'h24 == rob_tail ? _GEN_79 : _T_3372_36_ldst_val;
  assign _GEN_3732 = 6'h25 == rob_tail ? _GEN_79 : _T_3372_37_ldst_val;
  assign _GEN_3733 = 6'h26 == rob_tail ? _GEN_79 : _T_3372_38_ldst_val;
  assign _GEN_3734 = 6'h27 == rob_tail ? _GEN_79 : _T_3372_39_ldst_val;
  assign _GEN_3735 = 6'h0 == rob_tail ? _GEN_80 : _T_3372_0_dst_rtype;
  assign _GEN_3736 = 6'h1 == rob_tail ? _GEN_80 : _T_3372_1_dst_rtype;
  assign _GEN_3737 = 6'h2 == rob_tail ? _GEN_80 : _T_3372_2_dst_rtype;
  assign _GEN_3738 = 6'h3 == rob_tail ? _GEN_80 : _T_3372_3_dst_rtype;
  assign _GEN_3739 = 6'h4 == rob_tail ? _GEN_80 : _T_3372_4_dst_rtype;
  assign _GEN_3740 = 6'h5 == rob_tail ? _GEN_80 : _T_3372_5_dst_rtype;
  assign _GEN_3741 = 6'h6 == rob_tail ? _GEN_80 : _T_3372_6_dst_rtype;
  assign _GEN_3742 = 6'h7 == rob_tail ? _GEN_80 : _T_3372_7_dst_rtype;
  assign _GEN_3743 = 6'h8 == rob_tail ? _GEN_80 : _T_3372_8_dst_rtype;
  assign _GEN_3744 = 6'h9 == rob_tail ? _GEN_80 : _T_3372_9_dst_rtype;
  assign _GEN_3745 = 6'ha == rob_tail ? _GEN_80 : _T_3372_10_dst_rtype;
  assign _GEN_3746 = 6'hb == rob_tail ? _GEN_80 : _T_3372_11_dst_rtype;
  assign _GEN_3747 = 6'hc == rob_tail ? _GEN_80 : _T_3372_12_dst_rtype;
  assign _GEN_3748 = 6'hd == rob_tail ? _GEN_80 : _T_3372_13_dst_rtype;
  assign _GEN_3749 = 6'he == rob_tail ? _GEN_80 : _T_3372_14_dst_rtype;
  assign _GEN_3750 = 6'hf == rob_tail ? _GEN_80 : _T_3372_15_dst_rtype;
  assign _GEN_3751 = 6'h10 == rob_tail ? _GEN_80 : _T_3372_16_dst_rtype;
  assign _GEN_3752 = 6'h11 == rob_tail ? _GEN_80 : _T_3372_17_dst_rtype;
  assign _GEN_3753 = 6'h12 == rob_tail ? _GEN_80 : _T_3372_18_dst_rtype;
  assign _GEN_3754 = 6'h13 == rob_tail ? _GEN_80 : _T_3372_19_dst_rtype;
  assign _GEN_3755 = 6'h14 == rob_tail ? _GEN_80 : _T_3372_20_dst_rtype;
  assign _GEN_3756 = 6'h15 == rob_tail ? _GEN_80 : _T_3372_21_dst_rtype;
  assign _GEN_3757 = 6'h16 == rob_tail ? _GEN_80 : _T_3372_22_dst_rtype;
  assign _GEN_3758 = 6'h17 == rob_tail ? _GEN_80 : _T_3372_23_dst_rtype;
  assign _GEN_3759 = 6'h18 == rob_tail ? _GEN_80 : _T_3372_24_dst_rtype;
  assign _GEN_3760 = 6'h19 == rob_tail ? _GEN_80 : _T_3372_25_dst_rtype;
  assign _GEN_3761 = 6'h1a == rob_tail ? _GEN_80 : _T_3372_26_dst_rtype;
  assign _GEN_3762 = 6'h1b == rob_tail ? _GEN_80 : _T_3372_27_dst_rtype;
  assign _GEN_3763 = 6'h1c == rob_tail ? _GEN_80 : _T_3372_28_dst_rtype;
  assign _GEN_3764 = 6'h1d == rob_tail ? _GEN_80 : _T_3372_29_dst_rtype;
  assign _GEN_3765 = 6'h1e == rob_tail ? _GEN_80 : _T_3372_30_dst_rtype;
  assign _GEN_3766 = 6'h1f == rob_tail ? _GEN_80 : _T_3372_31_dst_rtype;
  assign _GEN_3767 = 6'h20 == rob_tail ? _GEN_80 : _T_3372_32_dst_rtype;
  assign _GEN_3768 = 6'h21 == rob_tail ? _GEN_80 : _T_3372_33_dst_rtype;
  assign _GEN_3769 = 6'h22 == rob_tail ? _GEN_80 : _T_3372_34_dst_rtype;
  assign _GEN_3770 = 6'h23 == rob_tail ? _GEN_80 : _T_3372_35_dst_rtype;
  assign _GEN_3771 = 6'h24 == rob_tail ? _GEN_80 : _T_3372_36_dst_rtype;
  assign _GEN_3772 = 6'h25 == rob_tail ? _GEN_80 : _T_3372_37_dst_rtype;
  assign _GEN_3773 = 6'h26 == rob_tail ? _GEN_80 : _T_3372_38_dst_rtype;
  assign _GEN_3774 = 6'h27 == rob_tail ? _GEN_80 : _T_3372_39_dst_rtype;
  assign _GEN_3895 = 6'h0 == rob_tail ? _GEN_84 : _T_3372_0_fp_val;
  assign _GEN_3896 = 6'h1 == rob_tail ? _GEN_84 : _T_3372_1_fp_val;
  assign _GEN_3897 = 6'h2 == rob_tail ? _GEN_84 : _T_3372_2_fp_val;
  assign _GEN_3898 = 6'h3 == rob_tail ? _GEN_84 : _T_3372_3_fp_val;
  assign _GEN_3899 = 6'h4 == rob_tail ? _GEN_84 : _T_3372_4_fp_val;
  assign _GEN_3900 = 6'h5 == rob_tail ? _GEN_84 : _T_3372_5_fp_val;
  assign _GEN_3901 = 6'h6 == rob_tail ? _GEN_84 : _T_3372_6_fp_val;
  assign _GEN_3902 = 6'h7 == rob_tail ? _GEN_84 : _T_3372_7_fp_val;
  assign _GEN_3903 = 6'h8 == rob_tail ? _GEN_84 : _T_3372_8_fp_val;
  assign _GEN_3904 = 6'h9 == rob_tail ? _GEN_84 : _T_3372_9_fp_val;
  assign _GEN_3905 = 6'ha == rob_tail ? _GEN_84 : _T_3372_10_fp_val;
  assign _GEN_3906 = 6'hb == rob_tail ? _GEN_84 : _T_3372_11_fp_val;
  assign _GEN_3907 = 6'hc == rob_tail ? _GEN_84 : _T_3372_12_fp_val;
  assign _GEN_3908 = 6'hd == rob_tail ? _GEN_84 : _T_3372_13_fp_val;
  assign _GEN_3909 = 6'he == rob_tail ? _GEN_84 : _T_3372_14_fp_val;
  assign _GEN_3910 = 6'hf == rob_tail ? _GEN_84 : _T_3372_15_fp_val;
  assign _GEN_3911 = 6'h10 == rob_tail ? _GEN_84 : _T_3372_16_fp_val;
  assign _GEN_3912 = 6'h11 == rob_tail ? _GEN_84 : _T_3372_17_fp_val;
  assign _GEN_3913 = 6'h12 == rob_tail ? _GEN_84 : _T_3372_18_fp_val;
  assign _GEN_3914 = 6'h13 == rob_tail ? _GEN_84 : _T_3372_19_fp_val;
  assign _GEN_3915 = 6'h14 == rob_tail ? _GEN_84 : _T_3372_20_fp_val;
  assign _GEN_3916 = 6'h15 == rob_tail ? _GEN_84 : _T_3372_21_fp_val;
  assign _GEN_3917 = 6'h16 == rob_tail ? _GEN_84 : _T_3372_22_fp_val;
  assign _GEN_3918 = 6'h17 == rob_tail ? _GEN_84 : _T_3372_23_fp_val;
  assign _GEN_3919 = 6'h18 == rob_tail ? _GEN_84 : _T_3372_24_fp_val;
  assign _GEN_3920 = 6'h19 == rob_tail ? _GEN_84 : _T_3372_25_fp_val;
  assign _GEN_3921 = 6'h1a == rob_tail ? _GEN_84 : _T_3372_26_fp_val;
  assign _GEN_3922 = 6'h1b == rob_tail ? _GEN_84 : _T_3372_27_fp_val;
  assign _GEN_3923 = 6'h1c == rob_tail ? _GEN_84 : _T_3372_28_fp_val;
  assign _GEN_3924 = 6'h1d == rob_tail ? _GEN_84 : _T_3372_29_fp_val;
  assign _GEN_3925 = 6'h1e == rob_tail ? _GEN_84 : _T_3372_30_fp_val;
  assign _GEN_3926 = 6'h1f == rob_tail ? _GEN_84 : _T_3372_31_fp_val;
  assign _GEN_3927 = 6'h20 == rob_tail ? _GEN_84 : _T_3372_32_fp_val;
  assign _GEN_3928 = 6'h21 == rob_tail ? _GEN_84 : _T_3372_33_fp_val;
  assign _GEN_3929 = 6'h22 == rob_tail ? _GEN_84 : _T_3372_34_fp_val;
  assign _GEN_3930 = 6'h23 == rob_tail ? _GEN_84 : _T_3372_35_fp_val;
  assign _GEN_3931 = 6'h24 == rob_tail ? _GEN_84 : _T_3372_36_fp_val;
  assign _GEN_3932 = 6'h25 == rob_tail ? _GEN_84 : _T_3372_37_fp_val;
  assign _GEN_3933 = 6'h26 == rob_tail ? _GEN_84 : _T_3372_38_fp_val;
  assign _GEN_3934 = 6'h27 == rob_tail ? _GEN_84 : _T_3372_39_fp_val;
  assign _GEN_4255 = 6'h1 == rob_tail ? _T_3073_1 : _T_3073_0;
  assign _GEN_4256 = 6'h2 == rob_tail ? _T_3073_2 : _GEN_4255;
  assign _GEN_4257 = 6'h3 == rob_tail ? _T_3073_3 : _GEN_4256;
  assign _GEN_4258 = 6'h4 == rob_tail ? _T_3073_4 : _GEN_4257;
  assign _GEN_4259 = 6'h5 == rob_tail ? _T_3073_5 : _GEN_4258;
  assign _GEN_4260 = 6'h6 == rob_tail ? _T_3073_6 : _GEN_4259;
  assign _GEN_4261 = 6'h7 == rob_tail ? _T_3073_7 : _GEN_4260;
  assign _GEN_4262 = 6'h8 == rob_tail ? _T_3073_8 : _GEN_4261;
  assign _GEN_4263 = 6'h9 == rob_tail ? _T_3073_9 : _GEN_4262;
  assign _GEN_4264 = 6'ha == rob_tail ? _T_3073_10 : _GEN_4263;
  assign _GEN_4265 = 6'hb == rob_tail ? _T_3073_11 : _GEN_4264;
  assign _GEN_4266 = 6'hc == rob_tail ? _T_3073_12 : _GEN_4265;
  assign _GEN_4267 = 6'hd == rob_tail ? _T_3073_13 : _GEN_4266;
  assign _GEN_4268 = 6'he == rob_tail ? _T_3073_14 : _GEN_4267;
  assign _GEN_4269 = 6'hf == rob_tail ? _T_3073_15 : _GEN_4268;
  assign _GEN_4270 = 6'h10 == rob_tail ? _T_3073_16 : _GEN_4269;
  assign _GEN_4271 = 6'h11 == rob_tail ? _T_3073_17 : _GEN_4270;
  assign _GEN_4272 = 6'h12 == rob_tail ? _T_3073_18 : _GEN_4271;
  assign _GEN_4273 = 6'h13 == rob_tail ? _T_3073_19 : _GEN_4272;
  assign _GEN_4274 = 6'h14 == rob_tail ? _T_3073_20 : _GEN_4273;
  assign _GEN_4275 = 6'h15 == rob_tail ? _T_3073_21 : _GEN_4274;
  assign _GEN_4276 = 6'h16 == rob_tail ? _T_3073_22 : _GEN_4275;
  assign _GEN_4277 = 6'h17 == rob_tail ? _T_3073_23 : _GEN_4276;
  assign _GEN_4278 = 6'h18 == rob_tail ? _T_3073_24 : _GEN_4277;
  assign _GEN_4279 = 6'h19 == rob_tail ? _T_3073_25 : _GEN_4278;
  assign _GEN_4280 = 6'h1a == rob_tail ? _T_3073_26 : _GEN_4279;
  assign _GEN_4281 = 6'h1b == rob_tail ? _T_3073_27 : _GEN_4280;
  assign _GEN_4282 = 6'h1c == rob_tail ? _T_3073_28 : _GEN_4281;
  assign _GEN_4283 = 6'h1d == rob_tail ? _T_3073_29 : _GEN_4282;
  assign _GEN_4284 = 6'h1e == rob_tail ? _T_3073_30 : _GEN_4283;
  assign _GEN_4285 = 6'h1f == rob_tail ? _T_3073_31 : _GEN_4284;
  assign _GEN_4286 = 6'h20 == rob_tail ? _T_3073_32 : _GEN_4285;
  assign _GEN_4287 = 6'h21 == rob_tail ? _T_3073_33 : _GEN_4286;
  assign _GEN_4288 = 6'h22 == rob_tail ? _T_3073_34 : _GEN_4287;
  assign _GEN_4289 = 6'h23 == rob_tail ? _T_3073_35 : _GEN_4288;
  assign _GEN_4290 = 6'h24 == rob_tail ? _T_3073_36 : _GEN_4289;
  assign _GEN_4291 = 6'h25 == rob_tail ? _T_3073_37 : _GEN_4290;
  assign _GEN_4292 = 6'h26 == rob_tail ? _T_3073_38 : _GEN_4291;
  assign _GEN_4293 = 6'h27 == rob_tail ? _T_3073_39 : _GEN_4292;
  assign _T_3785 = _GEN_93 == 1'h0;
  assign _T_3787 = _T_3785 | reset;
  assign _T_3789 = _T_3787 == 1'h0;
  assign _T_3790 = io_enq_uops_0_rob_idx[6:1];
  assign _T_3791 = _T_3790 == rob_tail;
  assign _T_3793 = _T_3791 | reset;
  assign _T_3795 = _T_3793 == 1'h0;
  assign _GEN_4374 = io_enq_valids_0 ? _GEN_575 : _T_3073_0;
  assign _GEN_4375 = io_enq_valids_0 ? _GEN_576 : _T_3073_1;
  assign _GEN_4376 = io_enq_valids_0 ? _GEN_577 : _T_3073_2;
  assign _GEN_4377 = io_enq_valids_0 ? _GEN_578 : _T_3073_3;
  assign _GEN_4378 = io_enq_valids_0 ? _GEN_579 : _T_3073_4;
  assign _GEN_4379 = io_enq_valids_0 ? _GEN_580 : _T_3073_5;
  assign _GEN_4380 = io_enq_valids_0 ? _GEN_581 : _T_3073_6;
  assign _GEN_4381 = io_enq_valids_0 ? _GEN_582 : _T_3073_7;
  assign _GEN_4382 = io_enq_valids_0 ? _GEN_583 : _T_3073_8;
  assign _GEN_4383 = io_enq_valids_0 ? _GEN_584 : _T_3073_9;
  assign _GEN_4384 = io_enq_valids_0 ? _GEN_585 : _T_3073_10;
  assign _GEN_4385 = io_enq_valids_0 ? _GEN_586 : _T_3073_11;
  assign _GEN_4386 = io_enq_valids_0 ? _GEN_587 : _T_3073_12;
  assign _GEN_4387 = io_enq_valids_0 ? _GEN_588 : _T_3073_13;
  assign _GEN_4388 = io_enq_valids_0 ? _GEN_589 : _T_3073_14;
  assign _GEN_4389 = io_enq_valids_0 ? _GEN_590 : _T_3073_15;
  assign _GEN_4390 = io_enq_valids_0 ? _GEN_591 : _T_3073_16;
  assign _GEN_4391 = io_enq_valids_0 ? _GEN_592 : _T_3073_17;
  assign _GEN_4392 = io_enq_valids_0 ? _GEN_593 : _T_3073_18;
  assign _GEN_4393 = io_enq_valids_0 ? _GEN_594 : _T_3073_19;
  assign _GEN_4394 = io_enq_valids_0 ? _GEN_595 : _T_3073_20;
  assign _GEN_4395 = io_enq_valids_0 ? _GEN_596 : _T_3073_21;
  assign _GEN_4396 = io_enq_valids_0 ? _GEN_597 : _T_3073_22;
  assign _GEN_4397 = io_enq_valids_0 ? _GEN_598 : _T_3073_23;
  assign _GEN_4398 = io_enq_valids_0 ? _GEN_599 : _T_3073_24;
  assign _GEN_4399 = io_enq_valids_0 ? _GEN_600 : _T_3073_25;
  assign _GEN_4400 = io_enq_valids_0 ? _GEN_601 : _T_3073_26;
  assign _GEN_4401 = io_enq_valids_0 ? _GEN_602 : _T_3073_27;
  assign _GEN_4402 = io_enq_valids_0 ? _GEN_603 : _T_3073_28;
  assign _GEN_4403 = io_enq_valids_0 ? _GEN_604 : _T_3073_29;
  assign _GEN_4404 = io_enq_valids_0 ? _GEN_605 : _T_3073_30;
  assign _GEN_4405 = io_enq_valids_0 ? _GEN_606 : _T_3073_31;
  assign _GEN_4406 = io_enq_valids_0 ? _GEN_607 : _T_3073_32;
  assign _GEN_4407 = io_enq_valids_0 ? _GEN_608 : _T_3073_33;
  assign _GEN_4408 = io_enq_valids_0 ? _GEN_609 : _T_3073_34;
  assign _GEN_4409 = io_enq_valids_0 ? _GEN_610 : _T_3073_35;
  assign _GEN_4410 = io_enq_valids_0 ? _GEN_611 : _T_3073_36;
  assign _GEN_4411 = io_enq_valids_0 ? _GEN_612 : _T_3073_37;
  assign _GEN_4412 = io_enq_valids_0 ? _GEN_613 : _T_3073_38;
  assign _GEN_4413 = io_enq_valids_0 ? _GEN_614 : _T_3073_39;
  assign _GEN_5378 = io_enq_valids_0 ? _GEN_1575 : _T_3372_0_br_mask;
  assign _GEN_5379 = io_enq_valids_0 ? _GEN_1576 : _T_3372_1_br_mask;
  assign _GEN_5380 = io_enq_valids_0 ? _GEN_1577 : _T_3372_2_br_mask;
  assign _GEN_5381 = io_enq_valids_0 ? _GEN_1578 : _T_3372_3_br_mask;
  assign _GEN_5382 = io_enq_valids_0 ? _GEN_1579 : _T_3372_4_br_mask;
  assign _GEN_5383 = io_enq_valids_0 ? _GEN_1580 : _T_3372_5_br_mask;
  assign _GEN_5384 = io_enq_valids_0 ? _GEN_1581 : _T_3372_6_br_mask;
  assign _GEN_5385 = io_enq_valids_0 ? _GEN_1582 : _T_3372_7_br_mask;
  assign _GEN_5386 = io_enq_valids_0 ? _GEN_1583 : _T_3372_8_br_mask;
  assign _GEN_5387 = io_enq_valids_0 ? _GEN_1584 : _T_3372_9_br_mask;
  assign _GEN_5388 = io_enq_valids_0 ? _GEN_1585 : _T_3372_10_br_mask;
  assign _GEN_5389 = io_enq_valids_0 ? _GEN_1586 : _T_3372_11_br_mask;
  assign _GEN_5390 = io_enq_valids_0 ? _GEN_1587 : _T_3372_12_br_mask;
  assign _GEN_5391 = io_enq_valids_0 ? _GEN_1588 : _T_3372_13_br_mask;
  assign _GEN_5392 = io_enq_valids_0 ? _GEN_1589 : _T_3372_14_br_mask;
  assign _GEN_5393 = io_enq_valids_0 ? _GEN_1590 : _T_3372_15_br_mask;
  assign _GEN_5394 = io_enq_valids_0 ? _GEN_1591 : _T_3372_16_br_mask;
  assign _GEN_5395 = io_enq_valids_0 ? _GEN_1592 : _T_3372_17_br_mask;
  assign _GEN_5396 = io_enq_valids_0 ? _GEN_1593 : _T_3372_18_br_mask;
  assign _GEN_5397 = io_enq_valids_0 ? _GEN_1594 : _T_3372_19_br_mask;
  assign _GEN_5398 = io_enq_valids_0 ? _GEN_1595 : _T_3372_20_br_mask;
  assign _GEN_5399 = io_enq_valids_0 ? _GEN_1596 : _T_3372_21_br_mask;
  assign _GEN_5400 = io_enq_valids_0 ? _GEN_1597 : _T_3372_22_br_mask;
  assign _GEN_5401 = io_enq_valids_0 ? _GEN_1598 : _T_3372_23_br_mask;
  assign _GEN_5402 = io_enq_valids_0 ? _GEN_1599 : _T_3372_24_br_mask;
  assign _GEN_5403 = io_enq_valids_0 ? _GEN_1600 : _T_3372_25_br_mask;
  assign _GEN_5404 = io_enq_valids_0 ? _GEN_1601 : _T_3372_26_br_mask;
  assign _GEN_5405 = io_enq_valids_0 ? _GEN_1602 : _T_3372_27_br_mask;
  assign _GEN_5406 = io_enq_valids_0 ? _GEN_1603 : _T_3372_28_br_mask;
  assign _GEN_5407 = io_enq_valids_0 ? _GEN_1604 : _T_3372_29_br_mask;
  assign _GEN_5408 = io_enq_valids_0 ? _GEN_1605 : _T_3372_30_br_mask;
  assign _GEN_5409 = io_enq_valids_0 ? _GEN_1606 : _T_3372_31_br_mask;
  assign _GEN_5410 = io_enq_valids_0 ? _GEN_1607 : _T_3372_32_br_mask;
  assign _GEN_5411 = io_enq_valids_0 ? _GEN_1608 : _T_3372_33_br_mask;
  assign _GEN_5412 = io_enq_valids_0 ? _GEN_1609 : _T_3372_34_br_mask;
  assign _GEN_5413 = io_enq_valids_0 ? _GEN_1610 : _T_3372_35_br_mask;
  assign _GEN_5414 = io_enq_valids_0 ? _GEN_1611 : _T_3372_36_br_mask;
  assign _GEN_5415 = io_enq_valids_0 ? _GEN_1612 : _T_3372_37_br_mask;
  assign _GEN_5416 = io_enq_valids_0 ? _GEN_1613 : _T_3372_38_br_mask;
  assign _GEN_5417 = io_enq_valids_0 ? _GEN_1614 : _T_3372_39_br_mask;
  assign _GEN_6498 = io_enq_valids_0 ? _GEN_2695 : _T_3372_0_pdst;
  assign _GEN_6499 = io_enq_valids_0 ? _GEN_2696 : _T_3372_1_pdst;
  assign _GEN_6500 = io_enq_valids_0 ? _GEN_2697 : _T_3372_2_pdst;
  assign _GEN_6501 = io_enq_valids_0 ? _GEN_2698 : _T_3372_3_pdst;
  assign _GEN_6502 = io_enq_valids_0 ? _GEN_2699 : _T_3372_4_pdst;
  assign _GEN_6503 = io_enq_valids_0 ? _GEN_2700 : _T_3372_5_pdst;
  assign _GEN_6504 = io_enq_valids_0 ? _GEN_2701 : _T_3372_6_pdst;
  assign _GEN_6505 = io_enq_valids_0 ? _GEN_2702 : _T_3372_7_pdst;
  assign _GEN_6506 = io_enq_valids_0 ? _GEN_2703 : _T_3372_8_pdst;
  assign _GEN_6507 = io_enq_valids_0 ? _GEN_2704 : _T_3372_9_pdst;
  assign _GEN_6508 = io_enq_valids_0 ? _GEN_2705 : _T_3372_10_pdst;
  assign _GEN_6509 = io_enq_valids_0 ? _GEN_2706 : _T_3372_11_pdst;
  assign _GEN_6510 = io_enq_valids_0 ? _GEN_2707 : _T_3372_12_pdst;
  assign _GEN_6511 = io_enq_valids_0 ? _GEN_2708 : _T_3372_13_pdst;
  assign _GEN_6512 = io_enq_valids_0 ? _GEN_2709 : _T_3372_14_pdst;
  assign _GEN_6513 = io_enq_valids_0 ? _GEN_2710 : _T_3372_15_pdst;
  assign _GEN_6514 = io_enq_valids_0 ? _GEN_2711 : _T_3372_16_pdst;
  assign _GEN_6515 = io_enq_valids_0 ? _GEN_2712 : _T_3372_17_pdst;
  assign _GEN_6516 = io_enq_valids_0 ? _GEN_2713 : _T_3372_18_pdst;
  assign _GEN_6517 = io_enq_valids_0 ? _GEN_2714 : _T_3372_19_pdst;
  assign _GEN_6518 = io_enq_valids_0 ? _GEN_2715 : _T_3372_20_pdst;
  assign _GEN_6519 = io_enq_valids_0 ? _GEN_2716 : _T_3372_21_pdst;
  assign _GEN_6520 = io_enq_valids_0 ? _GEN_2717 : _T_3372_22_pdst;
  assign _GEN_6521 = io_enq_valids_0 ? _GEN_2718 : _T_3372_23_pdst;
  assign _GEN_6522 = io_enq_valids_0 ? _GEN_2719 : _T_3372_24_pdst;
  assign _GEN_6523 = io_enq_valids_0 ? _GEN_2720 : _T_3372_25_pdst;
  assign _GEN_6524 = io_enq_valids_0 ? _GEN_2721 : _T_3372_26_pdst;
  assign _GEN_6525 = io_enq_valids_0 ? _GEN_2722 : _T_3372_27_pdst;
  assign _GEN_6526 = io_enq_valids_0 ? _GEN_2723 : _T_3372_28_pdst;
  assign _GEN_6527 = io_enq_valids_0 ? _GEN_2724 : _T_3372_29_pdst;
  assign _GEN_6528 = io_enq_valids_0 ? _GEN_2725 : _T_3372_30_pdst;
  assign _GEN_6529 = io_enq_valids_0 ? _GEN_2726 : _T_3372_31_pdst;
  assign _GEN_6530 = io_enq_valids_0 ? _GEN_2727 : _T_3372_32_pdst;
  assign _GEN_6531 = io_enq_valids_0 ? _GEN_2728 : _T_3372_33_pdst;
  assign _GEN_6532 = io_enq_valids_0 ? _GEN_2729 : _T_3372_34_pdst;
  assign _GEN_6533 = io_enq_valids_0 ? _GEN_2730 : _T_3372_35_pdst;
  assign _GEN_6534 = io_enq_valids_0 ? _GEN_2731 : _T_3372_36_pdst;
  assign _GEN_6535 = io_enq_valids_0 ? _GEN_2732 : _T_3372_37_pdst;
  assign _GEN_6536 = io_enq_valids_0 ? _GEN_2733 : _T_3372_38_pdst;
  assign _GEN_6537 = io_enq_valids_0 ? _GEN_2734 : _T_3372_39_pdst;
  assign _GEN_6778 = io_enq_valids_0 ? _GEN_2975 : _T_3372_0_stale_pdst;
  assign _GEN_6779 = io_enq_valids_0 ? _GEN_2976 : _T_3372_1_stale_pdst;
  assign _GEN_6780 = io_enq_valids_0 ? _GEN_2977 : _T_3372_2_stale_pdst;
  assign _GEN_6781 = io_enq_valids_0 ? _GEN_2978 : _T_3372_3_stale_pdst;
  assign _GEN_6782 = io_enq_valids_0 ? _GEN_2979 : _T_3372_4_stale_pdst;
  assign _GEN_6783 = io_enq_valids_0 ? _GEN_2980 : _T_3372_5_stale_pdst;
  assign _GEN_6784 = io_enq_valids_0 ? _GEN_2981 : _T_3372_6_stale_pdst;
  assign _GEN_6785 = io_enq_valids_0 ? _GEN_2982 : _T_3372_7_stale_pdst;
  assign _GEN_6786 = io_enq_valids_0 ? _GEN_2983 : _T_3372_8_stale_pdst;
  assign _GEN_6787 = io_enq_valids_0 ? _GEN_2984 : _T_3372_9_stale_pdst;
  assign _GEN_6788 = io_enq_valids_0 ? _GEN_2985 : _T_3372_10_stale_pdst;
  assign _GEN_6789 = io_enq_valids_0 ? _GEN_2986 : _T_3372_11_stale_pdst;
  assign _GEN_6790 = io_enq_valids_0 ? _GEN_2987 : _T_3372_12_stale_pdst;
  assign _GEN_6791 = io_enq_valids_0 ? _GEN_2988 : _T_3372_13_stale_pdst;
  assign _GEN_6792 = io_enq_valids_0 ? _GEN_2989 : _T_3372_14_stale_pdst;
  assign _GEN_6793 = io_enq_valids_0 ? _GEN_2990 : _T_3372_15_stale_pdst;
  assign _GEN_6794 = io_enq_valids_0 ? _GEN_2991 : _T_3372_16_stale_pdst;
  assign _GEN_6795 = io_enq_valids_0 ? _GEN_2992 : _T_3372_17_stale_pdst;
  assign _GEN_6796 = io_enq_valids_0 ? _GEN_2993 : _T_3372_18_stale_pdst;
  assign _GEN_6797 = io_enq_valids_0 ? _GEN_2994 : _T_3372_19_stale_pdst;
  assign _GEN_6798 = io_enq_valids_0 ? _GEN_2995 : _T_3372_20_stale_pdst;
  assign _GEN_6799 = io_enq_valids_0 ? _GEN_2996 : _T_3372_21_stale_pdst;
  assign _GEN_6800 = io_enq_valids_0 ? _GEN_2997 : _T_3372_22_stale_pdst;
  assign _GEN_6801 = io_enq_valids_0 ? _GEN_2998 : _T_3372_23_stale_pdst;
  assign _GEN_6802 = io_enq_valids_0 ? _GEN_2999 : _T_3372_24_stale_pdst;
  assign _GEN_6803 = io_enq_valids_0 ? _GEN_3000 : _T_3372_25_stale_pdst;
  assign _GEN_6804 = io_enq_valids_0 ? _GEN_3001 : _T_3372_26_stale_pdst;
  assign _GEN_6805 = io_enq_valids_0 ? _GEN_3002 : _T_3372_27_stale_pdst;
  assign _GEN_6806 = io_enq_valids_0 ? _GEN_3003 : _T_3372_28_stale_pdst;
  assign _GEN_6807 = io_enq_valids_0 ? _GEN_3004 : _T_3372_29_stale_pdst;
  assign _GEN_6808 = io_enq_valids_0 ? _GEN_3005 : _T_3372_30_stale_pdst;
  assign _GEN_6809 = io_enq_valids_0 ? _GEN_3006 : _T_3372_31_stale_pdst;
  assign _GEN_6810 = io_enq_valids_0 ? _GEN_3007 : _T_3372_32_stale_pdst;
  assign _GEN_6811 = io_enq_valids_0 ? _GEN_3008 : _T_3372_33_stale_pdst;
  assign _GEN_6812 = io_enq_valids_0 ? _GEN_3009 : _T_3372_34_stale_pdst;
  assign _GEN_6813 = io_enq_valids_0 ? _GEN_3010 : _T_3372_35_stale_pdst;
  assign _GEN_6814 = io_enq_valids_0 ? _GEN_3011 : _T_3372_36_stale_pdst;
  assign _GEN_6815 = io_enq_valids_0 ? _GEN_3012 : _T_3372_37_stale_pdst;
  assign _GEN_6816 = io_enq_valids_0 ? _GEN_3013 : _T_3372_38_stale_pdst;
  assign _GEN_6817 = io_enq_valids_0 ? _GEN_3014 : _T_3372_39_stale_pdst;
  assign _GEN_7058 = io_enq_valids_0 ? _GEN_3255 : _T_3372_0_is_fencei;
  assign _GEN_7059 = io_enq_valids_0 ? _GEN_3256 : _T_3372_1_is_fencei;
  assign _GEN_7060 = io_enq_valids_0 ? _GEN_3257 : _T_3372_2_is_fencei;
  assign _GEN_7061 = io_enq_valids_0 ? _GEN_3258 : _T_3372_3_is_fencei;
  assign _GEN_7062 = io_enq_valids_0 ? _GEN_3259 : _T_3372_4_is_fencei;
  assign _GEN_7063 = io_enq_valids_0 ? _GEN_3260 : _T_3372_5_is_fencei;
  assign _GEN_7064 = io_enq_valids_0 ? _GEN_3261 : _T_3372_6_is_fencei;
  assign _GEN_7065 = io_enq_valids_0 ? _GEN_3262 : _T_3372_7_is_fencei;
  assign _GEN_7066 = io_enq_valids_0 ? _GEN_3263 : _T_3372_8_is_fencei;
  assign _GEN_7067 = io_enq_valids_0 ? _GEN_3264 : _T_3372_9_is_fencei;
  assign _GEN_7068 = io_enq_valids_0 ? _GEN_3265 : _T_3372_10_is_fencei;
  assign _GEN_7069 = io_enq_valids_0 ? _GEN_3266 : _T_3372_11_is_fencei;
  assign _GEN_7070 = io_enq_valids_0 ? _GEN_3267 : _T_3372_12_is_fencei;
  assign _GEN_7071 = io_enq_valids_0 ? _GEN_3268 : _T_3372_13_is_fencei;
  assign _GEN_7072 = io_enq_valids_0 ? _GEN_3269 : _T_3372_14_is_fencei;
  assign _GEN_7073 = io_enq_valids_0 ? _GEN_3270 : _T_3372_15_is_fencei;
  assign _GEN_7074 = io_enq_valids_0 ? _GEN_3271 : _T_3372_16_is_fencei;
  assign _GEN_7075 = io_enq_valids_0 ? _GEN_3272 : _T_3372_17_is_fencei;
  assign _GEN_7076 = io_enq_valids_0 ? _GEN_3273 : _T_3372_18_is_fencei;
  assign _GEN_7077 = io_enq_valids_0 ? _GEN_3274 : _T_3372_19_is_fencei;
  assign _GEN_7078 = io_enq_valids_0 ? _GEN_3275 : _T_3372_20_is_fencei;
  assign _GEN_7079 = io_enq_valids_0 ? _GEN_3276 : _T_3372_21_is_fencei;
  assign _GEN_7080 = io_enq_valids_0 ? _GEN_3277 : _T_3372_22_is_fencei;
  assign _GEN_7081 = io_enq_valids_0 ? _GEN_3278 : _T_3372_23_is_fencei;
  assign _GEN_7082 = io_enq_valids_0 ? _GEN_3279 : _T_3372_24_is_fencei;
  assign _GEN_7083 = io_enq_valids_0 ? _GEN_3280 : _T_3372_25_is_fencei;
  assign _GEN_7084 = io_enq_valids_0 ? _GEN_3281 : _T_3372_26_is_fencei;
  assign _GEN_7085 = io_enq_valids_0 ? _GEN_3282 : _T_3372_27_is_fencei;
  assign _GEN_7086 = io_enq_valids_0 ? _GEN_3283 : _T_3372_28_is_fencei;
  assign _GEN_7087 = io_enq_valids_0 ? _GEN_3284 : _T_3372_29_is_fencei;
  assign _GEN_7088 = io_enq_valids_0 ? _GEN_3285 : _T_3372_30_is_fencei;
  assign _GEN_7089 = io_enq_valids_0 ? _GEN_3286 : _T_3372_31_is_fencei;
  assign _GEN_7090 = io_enq_valids_0 ? _GEN_3287 : _T_3372_32_is_fencei;
  assign _GEN_7091 = io_enq_valids_0 ? _GEN_3288 : _T_3372_33_is_fencei;
  assign _GEN_7092 = io_enq_valids_0 ? _GEN_3289 : _T_3372_34_is_fencei;
  assign _GEN_7093 = io_enq_valids_0 ? _GEN_3290 : _T_3372_35_is_fencei;
  assign _GEN_7094 = io_enq_valids_0 ? _GEN_3291 : _T_3372_36_is_fencei;
  assign _GEN_7095 = io_enq_valids_0 ? _GEN_3292 : _T_3372_37_is_fencei;
  assign _GEN_7096 = io_enq_valids_0 ? _GEN_3293 : _T_3372_38_is_fencei;
  assign _GEN_7097 = io_enq_valids_0 ? _GEN_3294 : _T_3372_39_is_fencei;
  assign _GEN_7098 = io_enq_valids_0 ? _GEN_3295 : _T_3372_0_is_store;
  assign _GEN_7099 = io_enq_valids_0 ? _GEN_3296 : _T_3372_1_is_store;
  assign _GEN_7100 = io_enq_valids_0 ? _GEN_3297 : _T_3372_2_is_store;
  assign _GEN_7101 = io_enq_valids_0 ? _GEN_3298 : _T_3372_3_is_store;
  assign _GEN_7102 = io_enq_valids_0 ? _GEN_3299 : _T_3372_4_is_store;
  assign _GEN_7103 = io_enq_valids_0 ? _GEN_3300 : _T_3372_5_is_store;
  assign _GEN_7104 = io_enq_valids_0 ? _GEN_3301 : _T_3372_6_is_store;
  assign _GEN_7105 = io_enq_valids_0 ? _GEN_3302 : _T_3372_7_is_store;
  assign _GEN_7106 = io_enq_valids_0 ? _GEN_3303 : _T_3372_8_is_store;
  assign _GEN_7107 = io_enq_valids_0 ? _GEN_3304 : _T_3372_9_is_store;
  assign _GEN_7108 = io_enq_valids_0 ? _GEN_3305 : _T_3372_10_is_store;
  assign _GEN_7109 = io_enq_valids_0 ? _GEN_3306 : _T_3372_11_is_store;
  assign _GEN_7110 = io_enq_valids_0 ? _GEN_3307 : _T_3372_12_is_store;
  assign _GEN_7111 = io_enq_valids_0 ? _GEN_3308 : _T_3372_13_is_store;
  assign _GEN_7112 = io_enq_valids_0 ? _GEN_3309 : _T_3372_14_is_store;
  assign _GEN_7113 = io_enq_valids_0 ? _GEN_3310 : _T_3372_15_is_store;
  assign _GEN_7114 = io_enq_valids_0 ? _GEN_3311 : _T_3372_16_is_store;
  assign _GEN_7115 = io_enq_valids_0 ? _GEN_3312 : _T_3372_17_is_store;
  assign _GEN_7116 = io_enq_valids_0 ? _GEN_3313 : _T_3372_18_is_store;
  assign _GEN_7117 = io_enq_valids_0 ? _GEN_3314 : _T_3372_19_is_store;
  assign _GEN_7118 = io_enq_valids_0 ? _GEN_3315 : _T_3372_20_is_store;
  assign _GEN_7119 = io_enq_valids_0 ? _GEN_3316 : _T_3372_21_is_store;
  assign _GEN_7120 = io_enq_valids_0 ? _GEN_3317 : _T_3372_22_is_store;
  assign _GEN_7121 = io_enq_valids_0 ? _GEN_3318 : _T_3372_23_is_store;
  assign _GEN_7122 = io_enq_valids_0 ? _GEN_3319 : _T_3372_24_is_store;
  assign _GEN_7123 = io_enq_valids_0 ? _GEN_3320 : _T_3372_25_is_store;
  assign _GEN_7124 = io_enq_valids_0 ? _GEN_3321 : _T_3372_26_is_store;
  assign _GEN_7125 = io_enq_valids_0 ? _GEN_3322 : _T_3372_27_is_store;
  assign _GEN_7126 = io_enq_valids_0 ? _GEN_3323 : _T_3372_28_is_store;
  assign _GEN_7127 = io_enq_valids_0 ? _GEN_3324 : _T_3372_29_is_store;
  assign _GEN_7128 = io_enq_valids_0 ? _GEN_3325 : _T_3372_30_is_store;
  assign _GEN_7129 = io_enq_valids_0 ? _GEN_3326 : _T_3372_31_is_store;
  assign _GEN_7130 = io_enq_valids_0 ? _GEN_3327 : _T_3372_32_is_store;
  assign _GEN_7131 = io_enq_valids_0 ? _GEN_3328 : _T_3372_33_is_store;
  assign _GEN_7132 = io_enq_valids_0 ? _GEN_3329 : _T_3372_34_is_store;
  assign _GEN_7133 = io_enq_valids_0 ? _GEN_3330 : _T_3372_35_is_store;
  assign _GEN_7134 = io_enq_valids_0 ? _GEN_3331 : _T_3372_36_is_store;
  assign _GEN_7135 = io_enq_valids_0 ? _GEN_3332 : _T_3372_37_is_store;
  assign _GEN_7136 = io_enq_valids_0 ? _GEN_3333 : _T_3372_38_is_store;
  assign _GEN_7137 = io_enq_valids_0 ? _GEN_3334 : _T_3372_39_is_store;
  assign _GEN_7178 = io_enq_valids_0 ? _GEN_3375 : _T_3372_0_is_load;
  assign _GEN_7179 = io_enq_valids_0 ? _GEN_3376 : _T_3372_1_is_load;
  assign _GEN_7180 = io_enq_valids_0 ? _GEN_3377 : _T_3372_2_is_load;
  assign _GEN_7181 = io_enq_valids_0 ? _GEN_3378 : _T_3372_3_is_load;
  assign _GEN_7182 = io_enq_valids_0 ? _GEN_3379 : _T_3372_4_is_load;
  assign _GEN_7183 = io_enq_valids_0 ? _GEN_3380 : _T_3372_5_is_load;
  assign _GEN_7184 = io_enq_valids_0 ? _GEN_3381 : _T_3372_6_is_load;
  assign _GEN_7185 = io_enq_valids_0 ? _GEN_3382 : _T_3372_7_is_load;
  assign _GEN_7186 = io_enq_valids_0 ? _GEN_3383 : _T_3372_8_is_load;
  assign _GEN_7187 = io_enq_valids_0 ? _GEN_3384 : _T_3372_9_is_load;
  assign _GEN_7188 = io_enq_valids_0 ? _GEN_3385 : _T_3372_10_is_load;
  assign _GEN_7189 = io_enq_valids_0 ? _GEN_3386 : _T_3372_11_is_load;
  assign _GEN_7190 = io_enq_valids_0 ? _GEN_3387 : _T_3372_12_is_load;
  assign _GEN_7191 = io_enq_valids_0 ? _GEN_3388 : _T_3372_13_is_load;
  assign _GEN_7192 = io_enq_valids_0 ? _GEN_3389 : _T_3372_14_is_load;
  assign _GEN_7193 = io_enq_valids_0 ? _GEN_3390 : _T_3372_15_is_load;
  assign _GEN_7194 = io_enq_valids_0 ? _GEN_3391 : _T_3372_16_is_load;
  assign _GEN_7195 = io_enq_valids_0 ? _GEN_3392 : _T_3372_17_is_load;
  assign _GEN_7196 = io_enq_valids_0 ? _GEN_3393 : _T_3372_18_is_load;
  assign _GEN_7197 = io_enq_valids_0 ? _GEN_3394 : _T_3372_19_is_load;
  assign _GEN_7198 = io_enq_valids_0 ? _GEN_3395 : _T_3372_20_is_load;
  assign _GEN_7199 = io_enq_valids_0 ? _GEN_3396 : _T_3372_21_is_load;
  assign _GEN_7200 = io_enq_valids_0 ? _GEN_3397 : _T_3372_22_is_load;
  assign _GEN_7201 = io_enq_valids_0 ? _GEN_3398 : _T_3372_23_is_load;
  assign _GEN_7202 = io_enq_valids_0 ? _GEN_3399 : _T_3372_24_is_load;
  assign _GEN_7203 = io_enq_valids_0 ? _GEN_3400 : _T_3372_25_is_load;
  assign _GEN_7204 = io_enq_valids_0 ? _GEN_3401 : _T_3372_26_is_load;
  assign _GEN_7205 = io_enq_valids_0 ? _GEN_3402 : _T_3372_27_is_load;
  assign _GEN_7206 = io_enq_valids_0 ? _GEN_3403 : _T_3372_28_is_load;
  assign _GEN_7207 = io_enq_valids_0 ? _GEN_3404 : _T_3372_29_is_load;
  assign _GEN_7208 = io_enq_valids_0 ? _GEN_3405 : _T_3372_30_is_load;
  assign _GEN_7209 = io_enq_valids_0 ? _GEN_3406 : _T_3372_31_is_load;
  assign _GEN_7210 = io_enq_valids_0 ? _GEN_3407 : _T_3372_32_is_load;
  assign _GEN_7211 = io_enq_valids_0 ? _GEN_3408 : _T_3372_33_is_load;
  assign _GEN_7212 = io_enq_valids_0 ? _GEN_3409 : _T_3372_34_is_load;
  assign _GEN_7213 = io_enq_valids_0 ? _GEN_3410 : _T_3372_35_is_load;
  assign _GEN_7214 = io_enq_valids_0 ? _GEN_3411 : _T_3372_36_is_load;
  assign _GEN_7215 = io_enq_valids_0 ? _GEN_3412 : _T_3372_37_is_load;
  assign _GEN_7216 = io_enq_valids_0 ? _GEN_3413 : _T_3372_38_is_load;
  assign _GEN_7217 = io_enq_valids_0 ? _GEN_3414 : _T_3372_39_is_load;
  assign _GEN_7218 = io_enq_valids_0 ? _GEN_3415 : _T_3372_0_is_sys_pc2epc;
  assign _GEN_7219 = io_enq_valids_0 ? _GEN_3416 : _T_3372_1_is_sys_pc2epc;
  assign _GEN_7220 = io_enq_valids_0 ? _GEN_3417 : _T_3372_2_is_sys_pc2epc;
  assign _GEN_7221 = io_enq_valids_0 ? _GEN_3418 : _T_3372_3_is_sys_pc2epc;
  assign _GEN_7222 = io_enq_valids_0 ? _GEN_3419 : _T_3372_4_is_sys_pc2epc;
  assign _GEN_7223 = io_enq_valids_0 ? _GEN_3420 : _T_3372_5_is_sys_pc2epc;
  assign _GEN_7224 = io_enq_valids_0 ? _GEN_3421 : _T_3372_6_is_sys_pc2epc;
  assign _GEN_7225 = io_enq_valids_0 ? _GEN_3422 : _T_3372_7_is_sys_pc2epc;
  assign _GEN_7226 = io_enq_valids_0 ? _GEN_3423 : _T_3372_8_is_sys_pc2epc;
  assign _GEN_7227 = io_enq_valids_0 ? _GEN_3424 : _T_3372_9_is_sys_pc2epc;
  assign _GEN_7228 = io_enq_valids_0 ? _GEN_3425 : _T_3372_10_is_sys_pc2epc;
  assign _GEN_7229 = io_enq_valids_0 ? _GEN_3426 : _T_3372_11_is_sys_pc2epc;
  assign _GEN_7230 = io_enq_valids_0 ? _GEN_3427 : _T_3372_12_is_sys_pc2epc;
  assign _GEN_7231 = io_enq_valids_0 ? _GEN_3428 : _T_3372_13_is_sys_pc2epc;
  assign _GEN_7232 = io_enq_valids_0 ? _GEN_3429 : _T_3372_14_is_sys_pc2epc;
  assign _GEN_7233 = io_enq_valids_0 ? _GEN_3430 : _T_3372_15_is_sys_pc2epc;
  assign _GEN_7234 = io_enq_valids_0 ? _GEN_3431 : _T_3372_16_is_sys_pc2epc;
  assign _GEN_7235 = io_enq_valids_0 ? _GEN_3432 : _T_3372_17_is_sys_pc2epc;
  assign _GEN_7236 = io_enq_valids_0 ? _GEN_3433 : _T_3372_18_is_sys_pc2epc;
  assign _GEN_7237 = io_enq_valids_0 ? _GEN_3434 : _T_3372_19_is_sys_pc2epc;
  assign _GEN_7238 = io_enq_valids_0 ? _GEN_3435 : _T_3372_20_is_sys_pc2epc;
  assign _GEN_7239 = io_enq_valids_0 ? _GEN_3436 : _T_3372_21_is_sys_pc2epc;
  assign _GEN_7240 = io_enq_valids_0 ? _GEN_3437 : _T_3372_22_is_sys_pc2epc;
  assign _GEN_7241 = io_enq_valids_0 ? _GEN_3438 : _T_3372_23_is_sys_pc2epc;
  assign _GEN_7242 = io_enq_valids_0 ? _GEN_3439 : _T_3372_24_is_sys_pc2epc;
  assign _GEN_7243 = io_enq_valids_0 ? _GEN_3440 : _T_3372_25_is_sys_pc2epc;
  assign _GEN_7244 = io_enq_valids_0 ? _GEN_3441 : _T_3372_26_is_sys_pc2epc;
  assign _GEN_7245 = io_enq_valids_0 ? _GEN_3442 : _T_3372_27_is_sys_pc2epc;
  assign _GEN_7246 = io_enq_valids_0 ? _GEN_3443 : _T_3372_28_is_sys_pc2epc;
  assign _GEN_7247 = io_enq_valids_0 ? _GEN_3444 : _T_3372_29_is_sys_pc2epc;
  assign _GEN_7248 = io_enq_valids_0 ? _GEN_3445 : _T_3372_30_is_sys_pc2epc;
  assign _GEN_7249 = io_enq_valids_0 ? _GEN_3446 : _T_3372_31_is_sys_pc2epc;
  assign _GEN_7250 = io_enq_valids_0 ? _GEN_3447 : _T_3372_32_is_sys_pc2epc;
  assign _GEN_7251 = io_enq_valids_0 ? _GEN_3448 : _T_3372_33_is_sys_pc2epc;
  assign _GEN_7252 = io_enq_valids_0 ? _GEN_3449 : _T_3372_34_is_sys_pc2epc;
  assign _GEN_7253 = io_enq_valids_0 ? _GEN_3450 : _T_3372_35_is_sys_pc2epc;
  assign _GEN_7254 = io_enq_valids_0 ? _GEN_3451 : _T_3372_36_is_sys_pc2epc;
  assign _GEN_7255 = io_enq_valids_0 ? _GEN_3452 : _T_3372_37_is_sys_pc2epc;
  assign _GEN_7256 = io_enq_valids_0 ? _GEN_3453 : _T_3372_38_is_sys_pc2epc;
  assign _GEN_7257 = io_enq_valids_0 ? _GEN_3454 : _T_3372_39_is_sys_pc2epc;
  assign _GEN_7298 = io_enq_valids_0 ? _GEN_3495 : _T_3372_0_flush_on_commit;
  assign _GEN_7299 = io_enq_valids_0 ? _GEN_3496 : _T_3372_1_flush_on_commit;
  assign _GEN_7300 = io_enq_valids_0 ? _GEN_3497 : _T_3372_2_flush_on_commit;
  assign _GEN_7301 = io_enq_valids_0 ? _GEN_3498 : _T_3372_3_flush_on_commit;
  assign _GEN_7302 = io_enq_valids_0 ? _GEN_3499 : _T_3372_4_flush_on_commit;
  assign _GEN_7303 = io_enq_valids_0 ? _GEN_3500 : _T_3372_5_flush_on_commit;
  assign _GEN_7304 = io_enq_valids_0 ? _GEN_3501 : _T_3372_6_flush_on_commit;
  assign _GEN_7305 = io_enq_valids_0 ? _GEN_3502 : _T_3372_7_flush_on_commit;
  assign _GEN_7306 = io_enq_valids_0 ? _GEN_3503 : _T_3372_8_flush_on_commit;
  assign _GEN_7307 = io_enq_valids_0 ? _GEN_3504 : _T_3372_9_flush_on_commit;
  assign _GEN_7308 = io_enq_valids_0 ? _GEN_3505 : _T_3372_10_flush_on_commit;
  assign _GEN_7309 = io_enq_valids_0 ? _GEN_3506 : _T_3372_11_flush_on_commit;
  assign _GEN_7310 = io_enq_valids_0 ? _GEN_3507 : _T_3372_12_flush_on_commit;
  assign _GEN_7311 = io_enq_valids_0 ? _GEN_3508 : _T_3372_13_flush_on_commit;
  assign _GEN_7312 = io_enq_valids_0 ? _GEN_3509 : _T_3372_14_flush_on_commit;
  assign _GEN_7313 = io_enq_valids_0 ? _GEN_3510 : _T_3372_15_flush_on_commit;
  assign _GEN_7314 = io_enq_valids_0 ? _GEN_3511 : _T_3372_16_flush_on_commit;
  assign _GEN_7315 = io_enq_valids_0 ? _GEN_3512 : _T_3372_17_flush_on_commit;
  assign _GEN_7316 = io_enq_valids_0 ? _GEN_3513 : _T_3372_18_flush_on_commit;
  assign _GEN_7317 = io_enq_valids_0 ? _GEN_3514 : _T_3372_19_flush_on_commit;
  assign _GEN_7318 = io_enq_valids_0 ? _GEN_3515 : _T_3372_20_flush_on_commit;
  assign _GEN_7319 = io_enq_valids_0 ? _GEN_3516 : _T_3372_21_flush_on_commit;
  assign _GEN_7320 = io_enq_valids_0 ? _GEN_3517 : _T_3372_22_flush_on_commit;
  assign _GEN_7321 = io_enq_valids_0 ? _GEN_3518 : _T_3372_23_flush_on_commit;
  assign _GEN_7322 = io_enq_valids_0 ? _GEN_3519 : _T_3372_24_flush_on_commit;
  assign _GEN_7323 = io_enq_valids_0 ? _GEN_3520 : _T_3372_25_flush_on_commit;
  assign _GEN_7324 = io_enq_valids_0 ? _GEN_3521 : _T_3372_26_flush_on_commit;
  assign _GEN_7325 = io_enq_valids_0 ? _GEN_3522 : _T_3372_27_flush_on_commit;
  assign _GEN_7326 = io_enq_valids_0 ? _GEN_3523 : _T_3372_28_flush_on_commit;
  assign _GEN_7327 = io_enq_valids_0 ? _GEN_3524 : _T_3372_29_flush_on_commit;
  assign _GEN_7328 = io_enq_valids_0 ? _GEN_3525 : _T_3372_30_flush_on_commit;
  assign _GEN_7329 = io_enq_valids_0 ? _GEN_3526 : _T_3372_31_flush_on_commit;
  assign _GEN_7330 = io_enq_valids_0 ? _GEN_3527 : _T_3372_32_flush_on_commit;
  assign _GEN_7331 = io_enq_valids_0 ? _GEN_3528 : _T_3372_33_flush_on_commit;
  assign _GEN_7332 = io_enq_valids_0 ? _GEN_3529 : _T_3372_34_flush_on_commit;
  assign _GEN_7333 = io_enq_valids_0 ? _GEN_3530 : _T_3372_35_flush_on_commit;
  assign _GEN_7334 = io_enq_valids_0 ? _GEN_3531 : _T_3372_36_flush_on_commit;
  assign _GEN_7335 = io_enq_valids_0 ? _GEN_3532 : _T_3372_37_flush_on_commit;
  assign _GEN_7336 = io_enq_valids_0 ? _GEN_3533 : _T_3372_38_flush_on_commit;
  assign _GEN_7337 = io_enq_valids_0 ? _GEN_3534 : _T_3372_39_flush_on_commit;
  assign _GEN_7338 = io_enq_valids_0 ? _GEN_3535 : _T_3372_0_ldst;
  assign _GEN_7339 = io_enq_valids_0 ? _GEN_3536 : _T_3372_1_ldst;
  assign _GEN_7340 = io_enq_valids_0 ? _GEN_3537 : _T_3372_2_ldst;
  assign _GEN_7341 = io_enq_valids_0 ? _GEN_3538 : _T_3372_3_ldst;
  assign _GEN_7342 = io_enq_valids_0 ? _GEN_3539 : _T_3372_4_ldst;
  assign _GEN_7343 = io_enq_valids_0 ? _GEN_3540 : _T_3372_5_ldst;
  assign _GEN_7344 = io_enq_valids_0 ? _GEN_3541 : _T_3372_6_ldst;
  assign _GEN_7345 = io_enq_valids_0 ? _GEN_3542 : _T_3372_7_ldst;
  assign _GEN_7346 = io_enq_valids_0 ? _GEN_3543 : _T_3372_8_ldst;
  assign _GEN_7347 = io_enq_valids_0 ? _GEN_3544 : _T_3372_9_ldst;
  assign _GEN_7348 = io_enq_valids_0 ? _GEN_3545 : _T_3372_10_ldst;
  assign _GEN_7349 = io_enq_valids_0 ? _GEN_3546 : _T_3372_11_ldst;
  assign _GEN_7350 = io_enq_valids_0 ? _GEN_3547 : _T_3372_12_ldst;
  assign _GEN_7351 = io_enq_valids_0 ? _GEN_3548 : _T_3372_13_ldst;
  assign _GEN_7352 = io_enq_valids_0 ? _GEN_3549 : _T_3372_14_ldst;
  assign _GEN_7353 = io_enq_valids_0 ? _GEN_3550 : _T_3372_15_ldst;
  assign _GEN_7354 = io_enq_valids_0 ? _GEN_3551 : _T_3372_16_ldst;
  assign _GEN_7355 = io_enq_valids_0 ? _GEN_3552 : _T_3372_17_ldst;
  assign _GEN_7356 = io_enq_valids_0 ? _GEN_3553 : _T_3372_18_ldst;
  assign _GEN_7357 = io_enq_valids_0 ? _GEN_3554 : _T_3372_19_ldst;
  assign _GEN_7358 = io_enq_valids_0 ? _GEN_3555 : _T_3372_20_ldst;
  assign _GEN_7359 = io_enq_valids_0 ? _GEN_3556 : _T_3372_21_ldst;
  assign _GEN_7360 = io_enq_valids_0 ? _GEN_3557 : _T_3372_22_ldst;
  assign _GEN_7361 = io_enq_valids_0 ? _GEN_3558 : _T_3372_23_ldst;
  assign _GEN_7362 = io_enq_valids_0 ? _GEN_3559 : _T_3372_24_ldst;
  assign _GEN_7363 = io_enq_valids_0 ? _GEN_3560 : _T_3372_25_ldst;
  assign _GEN_7364 = io_enq_valids_0 ? _GEN_3561 : _T_3372_26_ldst;
  assign _GEN_7365 = io_enq_valids_0 ? _GEN_3562 : _T_3372_27_ldst;
  assign _GEN_7366 = io_enq_valids_0 ? _GEN_3563 : _T_3372_28_ldst;
  assign _GEN_7367 = io_enq_valids_0 ? _GEN_3564 : _T_3372_29_ldst;
  assign _GEN_7368 = io_enq_valids_0 ? _GEN_3565 : _T_3372_30_ldst;
  assign _GEN_7369 = io_enq_valids_0 ? _GEN_3566 : _T_3372_31_ldst;
  assign _GEN_7370 = io_enq_valids_0 ? _GEN_3567 : _T_3372_32_ldst;
  assign _GEN_7371 = io_enq_valids_0 ? _GEN_3568 : _T_3372_33_ldst;
  assign _GEN_7372 = io_enq_valids_0 ? _GEN_3569 : _T_3372_34_ldst;
  assign _GEN_7373 = io_enq_valids_0 ? _GEN_3570 : _T_3372_35_ldst;
  assign _GEN_7374 = io_enq_valids_0 ? _GEN_3571 : _T_3372_36_ldst;
  assign _GEN_7375 = io_enq_valids_0 ? _GEN_3572 : _T_3372_37_ldst;
  assign _GEN_7376 = io_enq_valids_0 ? _GEN_3573 : _T_3372_38_ldst;
  assign _GEN_7377 = io_enq_valids_0 ? _GEN_3574 : _T_3372_39_ldst;
  assign _GEN_7498 = io_enq_valids_0 ? _GEN_3695 : _T_3372_0_ldst_val;
  assign _GEN_7499 = io_enq_valids_0 ? _GEN_3696 : _T_3372_1_ldst_val;
  assign _GEN_7500 = io_enq_valids_0 ? _GEN_3697 : _T_3372_2_ldst_val;
  assign _GEN_7501 = io_enq_valids_0 ? _GEN_3698 : _T_3372_3_ldst_val;
  assign _GEN_7502 = io_enq_valids_0 ? _GEN_3699 : _T_3372_4_ldst_val;
  assign _GEN_7503 = io_enq_valids_0 ? _GEN_3700 : _T_3372_5_ldst_val;
  assign _GEN_7504 = io_enq_valids_0 ? _GEN_3701 : _T_3372_6_ldst_val;
  assign _GEN_7505 = io_enq_valids_0 ? _GEN_3702 : _T_3372_7_ldst_val;
  assign _GEN_7506 = io_enq_valids_0 ? _GEN_3703 : _T_3372_8_ldst_val;
  assign _GEN_7507 = io_enq_valids_0 ? _GEN_3704 : _T_3372_9_ldst_val;
  assign _GEN_7508 = io_enq_valids_0 ? _GEN_3705 : _T_3372_10_ldst_val;
  assign _GEN_7509 = io_enq_valids_0 ? _GEN_3706 : _T_3372_11_ldst_val;
  assign _GEN_7510 = io_enq_valids_0 ? _GEN_3707 : _T_3372_12_ldst_val;
  assign _GEN_7511 = io_enq_valids_0 ? _GEN_3708 : _T_3372_13_ldst_val;
  assign _GEN_7512 = io_enq_valids_0 ? _GEN_3709 : _T_3372_14_ldst_val;
  assign _GEN_7513 = io_enq_valids_0 ? _GEN_3710 : _T_3372_15_ldst_val;
  assign _GEN_7514 = io_enq_valids_0 ? _GEN_3711 : _T_3372_16_ldst_val;
  assign _GEN_7515 = io_enq_valids_0 ? _GEN_3712 : _T_3372_17_ldst_val;
  assign _GEN_7516 = io_enq_valids_0 ? _GEN_3713 : _T_3372_18_ldst_val;
  assign _GEN_7517 = io_enq_valids_0 ? _GEN_3714 : _T_3372_19_ldst_val;
  assign _GEN_7518 = io_enq_valids_0 ? _GEN_3715 : _T_3372_20_ldst_val;
  assign _GEN_7519 = io_enq_valids_0 ? _GEN_3716 : _T_3372_21_ldst_val;
  assign _GEN_7520 = io_enq_valids_0 ? _GEN_3717 : _T_3372_22_ldst_val;
  assign _GEN_7521 = io_enq_valids_0 ? _GEN_3718 : _T_3372_23_ldst_val;
  assign _GEN_7522 = io_enq_valids_0 ? _GEN_3719 : _T_3372_24_ldst_val;
  assign _GEN_7523 = io_enq_valids_0 ? _GEN_3720 : _T_3372_25_ldst_val;
  assign _GEN_7524 = io_enq_valids_0 ? _GEN_3721 : _T_3372_26_ldst_val;
  assign _GEN_7525 = io_enq_valids_0 ? _GEN_3722 : _T_3372_27_ldst_val;
  assign _GEN_7526 = io_enq_valids_0 ? _GEN_3723 : _T_3372_28_ldst_val;
  assign _GEN_7527 = io_enq_valids_0 ? _GEN_3724 : _T_3372_29_ldst_val;
  assign _GEN_7528 = io_enq_valids_0 ? _GEN_3725 : _T_3372_30_ldst_val;
  assign _GEN_7529 = io_enq_valids_0 ? _GEN_3726 : _T_3372_31_ldst_val;
  assign _GEN_7530 = io_enq_valids_0 ? _GEN_3727 : _T_3372_32_ldst_val;
  assign _GEN_7531 = io_enq_valids_0 ? _GEN_3728 : _T_3372_33_ldst_val;
  assign _GEN_7532 = io_enq_valids_0 ? _GEN_3729 : _T_3372_34_ldst_val;
  assign _GEN_7533 = io_enq_valids_0 ? _GEN_3730 : _T_3372_35_ldst_val;
  assign _GEN_7534 = io_enq_valids_0 ? _GEN_3731 : _T_3372_36_ldst_val;
  assign _GEN_7535 = io_enq_valids_0 ? _GEN_3732 : _T_3372_37_ldst_val;
  assign _GEN_7536 = io_enq_valids_0 ? _GEN_3733 : _T_3372_38_ldst_val;
  assign _GEN_7537 = io_enq_valids_0 ? _GEN_3734 : _T_3372_39_ldst_val;
  assign _GEN_7538 = io_enq_valids_0 ? _GEN_3735 : _T_3372_0_dst_rtype;
  assign _GEN_7539 = io_enq_valids_0 ? _GEN_3736 : _T_3372_1_dst_rtype;
  assign _GEN_7540 = io_enq_valids_0 ? _GEN_3737 : _T_3372_2_dst_rtype;
  assign _GEN_7541 = io_enq_valids_0 ? _GEN_3738 : _T_3372_3_dst_rtype;
  assign _GEN_7542 = io_enq_valids_0 ? _GEN_3739 : _T_3372_4_dst_rtype;
  assign _GEN_7543 = io_enq_valids_0 ? _GEN_3740 : _T_3372_5_dst_rtype;
  assign _GEN_7544 = io_enq_valids_0 ? _GEN_3741 : _T_3372_6_dst_rtype;
  assign _GEN_7545 = io_enq_valids_0 ? _GEN_3742 : _T_3372_7_dst_rtype;
  assign _GEN_7546 = io_enq_valids_0 ? _GEN_3743 : _T_3372_8_dst_rtype;
  assign _GEN_7547 = io_enq_valids_0 ? _GEN_3744 : _T_3372_9_dst_rtype;
  assign _GEN_7548 = io_enq_valids_0 ? _GEN_3745 : _T_3372_10_dst_rtype;
  assign _GEN_7549 = io_enq_valids_0 ? _GEN_3746 : _T_3372_11_dst_rtype;
  assign _GEN_7550 = io_enq_valids_0 ? _GEN_3747 : _T_3372_12_dst_rtype;
  assign _GEN_7551 = io_enq_valids_0 ? _GEN_3748 : _T_3372_13_dst_rtype;
  assign _GEN_7552 = io_enq_valids_0 ? _GEN_3749 : _T_3372_14_dst_rtype;
  assign _GEN_7553 = io_enq_valids_0 ? _GEN_3750 : _T_3372_15_dst_rtype;
  assign _GEN_7554 = io_enq_valids_0 ? _GEN_3751 : _T_3372_16_dst_rtype;
  assign _GEN_7555 = io_enq_valids_0 ? _GEN_3752 : _T_3372_17_dst_rtype;
  assign _GEN_7556 = io_enq_valids_0 ? _GEN_3753 : _T_3372_18_dst_rtype;
  assign _GEN_7557 = io_enq_valids_0 ? _GEN_3754 : _T_3372_19_dst_rtype;
  assign _GEN_7558 = io_enq_valids_0 ? _GEN_3755 : _T_3372_20_dst_rtype;
  assign _GEN_7559 = io_enq_valids_0 ? _GEN_3756 : _T_3372_21_dst_rtype;
  assign _GEN_7560 = io_enq_valids_0 ? _GEN_3757 : _T_3372_22_dst_rtype;
  assign _GEN_7561 = io_enq_valids_0 ? _GEN_3758 : _T_3372_23_dst_rtype;
  assign _GEN_7562 = io_enq_valids_0 ? _GEN_3759 : _T_3372_24_dst_rtype;
  assign _GEN_7563 = io_enq_valids_0 ? _GEN_3760 : _T_3372_25_dst_rtype;
  assign _GEN_7564 = io_enq_valids_0 ? _GEN_3761 : _T_3372_26_dst_rtype;
  assign _GEN_7565 = io_enq_valids_0 ? _GEN_3762 : _T_3372_27_dst_rtype;
  assign _GEN_7566 = io_enq_valids_0 ? _GEN_3763 : _T_3372_28_dst_rtype;
  assign _GEN_7567 = io_enq_valids_0 ? _GEN_3764 : _T_3372_29_dst_rtype;
  assign _GEN_7568 = io_enq_valids_0 ? _GEN_3765 : _T_3372_30_dst_rtype;
  assign _GEN_7569 = io_enq_valids_0 ? _GEN_3766 : _T_3372_31_dst_rtype;
  assign _GEN_7570 = io_enq_valids_0 ? _GEN_3767 : _T_3372_32_dst_rtype;
  assign _GEN_7571 = io_enq_valids_0 ? _GEN_3768 : _T_3372_33_dst_rtype;
  assign _GEN_7572 = io_enq_valids_0 ? _GEN_3769 : _T_3372_34_dst_rtype;
  assign _GEN_7573 = io_enq_valids_0 ? _GEN_3770 : _T_3372_35_dst_rtype;
  assign _GEN_7574 = io_enq_valids_0 ? _GEN_3771 : _T_3372_36_dst_rtype;
  assign _GEN_7575 = io_enq_valids_0 ? _GEN_3772 : _T_3372_37_dst_rtype;
  assign _GEN_7576 = io_enq_valids_0 ? _GEN_3773 : _T_3372_38_dst_rtype;
  assign _GEN_7577 = io_enq_valids_0 ? _GEN_3774 : _T_3372_39_dst_rtype;
  assign _GEN_7698 = io_enq_valids_0 ? _GEN_3895 : _T_3372_0_fp_val;
  assign _GEN_7699 = io_enq_valids_0 ? _GEN_3896 : _T_3372_1_fp_val;
  assign _GEN_7700 = io_enq_valids_0 ? _GEN_3897 : _T_3372_2_fp_val;
  assign _GEN_7701 = io_enq_valids_0 ? _GEN_3898 : _T_3372_3_fp_val;
  assign _GEN_7702 = io_enq_valids_0 ? _GEN_3899 : _T_3372_4_fp_val;
  assign _GEN_7703 = io_enq_valids_0 ? _GEN_3900 : _T_3372_5_fp_val;
  assign _GEN_7704 = io_enq_valids_0 ? _GEN_3901 : _T_3372_6_fp_val;
  assign _GEN_7705 = io_enq_valids_0 ? _GEN_3902 : _T_3372_7_fp_val;
  assign _GEN_7706 = io_enq_valids_0 ? _GEN_3903 : _T_3372_8_fp_val;
  assign _GEN_7707 = io_enq_valids_0 ? _GEN_3904 : _T_3372_9_fp_val;
  assign _GEN_7708 = io_enq_valids_0 ? _GEN_3905 : _T_3372_10_fp_val;
  assign _GEN_7709 = io_enq_valids_0 ? _GEN_3906 : _T_3372_11_fp_val;
  assign _GEN_7710 = io_enq_valids_0 ? _GEN_3907 : _T_3372_12_fp_val;
  assign _GEN_7711 = io_enq_valids_0 ? _GEN_3908 : _T_3372_13_fp_val;
  assign _GEN_7712 = io_enq_valids_0 ? _GEN_3909 : _T_3372_14_fp_val;
  assign _GEN_7713 = io_enq_valids_0 ? _GEN_3910 : _T_3372_15_fp_val;
  assign _GEN_7714 = io_enq_valids_0 ? _GEN_3911 : _T_3372_16_fp_val;
  assign _GEN_7715 = io_enq_valids_0 ? _GEN_3912 : _T_3372_17_fp_val;
  assign _GEN_7716 = io_enq_valids_0 ? _GEN_3913 : _T_3372_18_fp_val;
  assign _GEN_7717 = io_enq_valids_0 ? _GEN_3914 : _T_3372_19_fp_val;
  assign _GEN_7718 = io_enq_valids_0 ? _GEN_3915 : _T_3372_20_fp_val;
  assign _GEN_7719 = io_enq_valids_0 ? _GEN_3916 : _T_3372_21_fp_val;
  assign _GEN_7720 = io_enq_valids_0 ? _GEN_3917 : _T_3372_22_fp_val;
  assign _GEN_7721 = io_enq_valids_0 ? _GEN_3918 : _T_3372_23_fp_val;
  assign _GEN_7722 = io_enq_valids_0 ? _GEN_3919 : _T_3372_24_fp_val;
  assign _GEN_7723 = io_enq_valids_0 ? _GEN_3920 : _T_3372_25_fp_val;
  assign _GEN_7724 = io_enq_valids_0 ? _GEN_3921 : _T_3372_26_fp_val;
  assign _GEN_7725 = io_enq_valids_0 ? _GEN_3922 : _T_3372_27_fp_val;
  assign _GEN_7726 = io_enq_valids_0 ? _GEN_3923 : _T_3372_28_fp_val;
  assign _GEN_7727 = io_enq_valids_0 ? _GEN_3924 : _T_3372_29_fp_val;
  assign _GEN_7728 = io_enq_valids_0 ? _GEN_3925 : _T_3372_30_fp_val;
  assign _GEN_7729 = io_enq_valids_0 ? _GEN_3926 : _T_3372_31_fp_val;
  assign _GEN_7730 = io_enq_valids_0 ? _GEN_3927 : _T_3372_32_fp_val;
  assign _GEN_7731 = io_enq_valids_0 ? _GEN_3928 : _T_3372_33_fp_val;
  assign _GEN_7732 = io_enq_valids_0 ? _GEN_3929 : _T_3372_34_fp_val;
  assign _GEN_7733 = io_enq_valids_0 ? _GEN_3930 : _T_3372_35_fp_val;
  assign _GEN_7734 = io_enq_valids_0 ? _GEN_3931 : _T_3372_36_fp_val;
  assign _GEN_7735 = io_enq_valids_0 ? _GEN_3932 : _T_3372_37_fp_val;
  assign _GEN_7736 = io_enq_valids_0 ? _GEN_3933 : _T_3372_38_fp_val;
  assign _GEN_7737 = io_enq_valids_0 ? _GEN_3934 : _T_3372_39_fp_val;
  assign _T_3813 = io_wb_resps_0_bits_uop_rob_idx >> 1'h1;
  assign _T_3814 = io_wb_resps_0_bits_uop_rob_idx[0];
  assign _T_3816 = _T_3814 == 1'h0;
  assign _T_3817 = io_wb_resps_0_valid & _T_3816;
  assign _T_3818 = _T_3813[5:0];
  assign _T_3822 = io_wb_resps_1_bits_uop_rob_idx >> 1'h1;
  assign _T_3823 = io_wb_resps_1_bits_uop_rob_idx[0];
  assign _T_3825 = _T_3823 == 1'h0;
  assign _T_3826 = io_wb_resps_1_valid & _T_3825;
  assign _T_3827 = _T_3822[5:0];
  assign _T_3831 = io_wb_resps_2_bits_uop_rob_idx >> 1'h1;
  assign _T_3832 = io_wb_resps_2_bits_uop_rob_idx[0];
  assign _T_3834 = _T_3832 == 1'h0;
  assign _T_3835 = io_wb_resps_2_valid & _T_3834;
  assign _T_3836 = _T_3831[5:0];
  assign _T_3840 = io_wb_resps_3_bits_uop_rob_idx >> 1'h1;
  assign _T_3841 = io_wb_resps_3_bits_uop_rob_idx[0];
  assign _T_3843 = _T_3841 == 1'h0;
  assign _T_3844 = io_wb_resps_3_valid & _T_3843;
  assign _T_3845 = _T_3840[5:0];
  assign _T_3849 = io_wb_resps_4_bits_uop_rob_idx >> 1'h1;
  assign _T_3850 = io_wb_resps_4_bits_uop_rob_idx[0];
  assign _T_3852 = _T_3850 == 1'h0;
  assign _T_3853 = io_wb_resps_4_valid & _T_3852;
  assign _T_3854 = _T_3849[5:0];
  assign _T_3857 = io_lsu_clr_bsy_rob_idx_0[0];
  assign _T_3859 = _T_3857 == 1'h0;
  assign _T_3860 = io_lsu_clr_bsy_valid_0 & _T_3859;
  assign _T_3862 = io_lsu_clr_bsy_rob_idx_0 >> 1'h1;
  assign _T_3863 = _T_3862[5:0];
  assign _GEN_8040 = 6'h1 == _T_3863 ? _T_3073_1 : _T_3073_0;
  assign _GEN_8041 = 6'h2 == _T_3863 ? _T_3073_2 : _GEN_8040;
  assign _GEN_8042 = 6'h3 == _T_3863 ? _T_3073_3 : _GEN_8041;
  assign _GEN_8043 = 6'h4 == _T_3863 ? _T_3073_4 : _GEN_8042;
  assign _GEN_8044 = 6'h5 == _T_3863 ? _T_3073_5 : _GEN_8043;
  assign _GEN_8045 = 6'h6 == _T_3863 ? _T_3073_6 : _GEN_8044;
  assign _GEN_8046 = 6'h7 == _T_3863 ? _T_3073_7 : _GEN_8045;
  assign _GEN_8047 = 6'h8 == _T_3863 ? _T_3073_8 : _GEN_8046;
  assign _GEN_8048 = 6'h9 == _T_3863 ? _T_3073_9 : _GEN_8047;
  assign _GEN_8049 = 6'ha == _T_3863 ? _T_3073_10 : _GEN_8048;
  assign _GEN_8050 = 6'hb == _T_3863 ? _T_3073_11 : _GEN_8049;
  assign _GEN_8051 = 6'hc == _T_3863 ? _T_3073_12 : _GEN_8050;
  assign _GEN_8052 = 6'hd == _T_3863 ? _T_3073_13 : _GEN_8051;
  assign _GEN_8053 = 6'he == _T_3863 ? _T_3073_14 : _GEN_8052;
  assign _GEN_8054 = 6'hf == _T_3863 ? _T_3073_15 : _GEN_8053;
  assign _GEN_8055 = 6'h10 == _T_3863 ? _T_3073_16 : _GEN_8054;
  assign _GEN_8056 = 6'h11 == _T_3863 ? _T_3073_17 : _GEN_8055;
  assign _GEN_8057 = 6'h12 == _T_3863 ? _T_3073_18 : _GEN_8056;
  assign _GEN_8058 = 6'h13 == _T_3863 ? _T_3073_19 : _GEN_8057;
  assign _GEN_8059 = 6'h14 == _T_3863 ? _T_3073_20 : _GEN_8058;
  assign _GEN_8060 = 6'h15 == _T_3863 ? _T_3073_21 : _GEN_8059;
  assign _GEN_8061 = 6'h16 == _T_3863 ? _T_3073_22 : _GEN_8060;
  assign _GEN_8062 = 6'h17 == _T_3863 ? _T_3073_23 : _GEN_8061;
  assign _GEN_8063 = 6'h18 == _T_3863 ? _T_3073_24 : _GEN_8062;
  assign _GEN_8064 = 6'h19 == _T_3863 ? _T_3073_25 : _GEN_8063;
  assign _GEN_8065 = 6'h1a == _T_3863 ? _T_3073_26 : _GEN_8064;
  assign _GEN_8066 = 6'h1b == _T_3863 ? _T_3073_27 : _GEN_8065;
  assign _GEN_8067 = 6'h1c == _T_3863 ? _T_3073_28 : _GEN_8066;
  assign _GEN_8068 = 6'h1d == _T_3863 ? _T_3073_29 : _GEN_8067;
  assign _GEN_8069 = 6'h1e == _T_3863 ? _T_3073_30 : _GEN_8068;
  assign _GEN_8070 = 6'h1f == _T_3863 ? _T_3073_31 : _GEN_8069;
  assign _GEN_8071 = 6'h20 == _T_3863 ? _T_3073_32 : _GEN_8070;
  assign _GEN_8072 = 6'h21 == _T_3863 ? _T_3073_33 : _GEN_8071;
  assign _GEN_8073 = 6'h22 == _T_3863 ? _T_3073_34 : _GEN_8072;
  assign _GEN_8074 = 6'h23 == _T_3863 ? _T_3073_35 : _GEN_8073;
  assign _GEN_8075 = 6'h24 == _T_3863 ? _T_3073_36 : _GEN_8074;
  assign _GEN_8076 = 6'h25 == _T_3863 ? _T_3073_37 : _GEN_8075;
  assign _GEN_8077 = 6'h26 == _T_3863 ? _T_3073_38 : _GEN_8076;
  assign _GEN_8078 = 6'h27 == _T_3863 ? _T_3073_39 : _GEN_8077;
  assign _T_3873 = _GEN_96 | reset;
  assign _T_3875 = _T_3873 == 1'h0;
  assign _T_3876 = _T_3862[5:0];
  assign _T_3879 = _T_3200__T_3877_data;
  assign _T_3881 = _T_3879 | reset;
  assign _T_3883 = _T_3881 == 1'h0;
  assign _T_3884 = io_lsu_clr_bsy_rob_idx_1[0];
  assign _T_3886 = _T_3884 == 1'h0;
  assign _T_3887 = io_lsu_clr_bsy_valid_1 & _T_3886;
  assign _T_3889 = io_lsu_clr_bsy_rob_idx_1 >> 1'h1;
  assign _T_3890 = _T_3889[5:0];
  assign _GEN_8084 = 6'h1 == _T_3890 ? _T_3073_1 : _T_3073_0;
  assign _GEN_8085 = 6'h2 == _T_3890 ? _T_3073_2 : _GEN_8084;
  assign _GEN_8086 = 6'h3 == _T_3890 ? _T_3073_3 : _GEN_8085;
  assign _GEN_8087 = 6'h4 == _T_3890 ? _T_3073_4 : _GEN_8086;
  assign _GEN_8088 = 6'h5 == _T_3890 ? _T_3073_5 : _GEN_8087;
  assign _GEN_8089 = 6'h6 == _T_3890 ? _T_3073_6 : _GEN_8088;
  assign _GEN_8090 = 6'h7 == _T_3890 ? _T_3073_7 : _GEN_8089;
  assign _GEN_8091 = 6'h8 == _T_3890 ? _T_3073_8 : _GEN_8090;
  assign _GEN_8092 = 6'h9 == _T_3890 ? _T_3073_9 : _GEN_8091;
  assign _GEN_8093 = 6'ha == _T_3890 ? _T_3073_10 : _GEN_8092;
  assign _GEN_8094 = 6'hb == _T_3890 ? _T_3073_11 : _GEN_8093;
  assign _GEN_8095 = 6'hc == _T_3890 ? _T_3073_12 : _GEN_8094;
  assign _GEN_8096 = 6'hd == _T_3890 ? _T_3073_13 : _GEN_8095;
  assign _GEN_8097 = 6'he == _T_3890 ? _T_3073_14 : _GEN_8096;
  assign _GEN_8098 = 6'hf == _T_3890 ? _T_3073_15 : _GEN_8097;
  assign _GEN_8099 = 6'h10 == _T_3890 ? _T_3073_16 : _GEN_8098;
  assign _GEN_8100 = 6'h11 == _T_3890 ? _T_3073_17 : _GEN_8099;
  assign _GEN_8101 = 6'h12 == _T_3890 ? _T_3073_18 : _GEN_8100;
  assign _GEN_8102 = 6'h13 == _T_3890 ? _T_3073_19 : _GEN_8101;
  assign _GEN_8103 = 6'h14 == _T_3890 ? _T_3073_20 : _GEN_8102;
  assign _GEN_8104 = 6'h15 == _T_3890 ? _T_3073_21 : _GEN_8103;
  assign _GEN_8105 = 6'h16 == _T_3890 ? _T_3073_22 : _GEN_8104;
  assign _GEN_8106 = 6'h17 == _T_3890 ? _T_3073_23 : _GEN_8105;
  assign _GEN_8107 = 6'h18 == _T_3890 ? _T_3073_24 : _GEN_8106;
  assign _GEN_8108 = 6'h19 == _T_3890 ? _T_3073_25 : _GEN_8107;
  assign _GEN_8109 = 6'h1a == _T_3890 ? _T_3073_26 : _GEN_8108;
  assign _GEN_8110 = 6'h1b == _T_3890 ? _T_3073_27 : _GEN_8109;
  assign _GEN_8111 = 6'h1c == _T_3890 ? _T_3073_28 : _GEN_8110;
  assign _GEN_8112 = 6'h1d == _T_3890 ? _T_3073_29 : _GEN_8111;
  assign _GEN_8113 = 6'h1e == _T_3890 ? _T_3073_30 : _GEN_8112;
  assign _GEN_8114 = 6'h1f == _T_3890 ? _T_3073_31 : _GEN_8113;
  assign _GEN_8115 = 6'h20 == _T_3890 ? _T_3073_32 : _GEN_8114;
  assign _GEN_8116 = 6'h21 == _T_3890 ? _T_3073_33 : _GEN_8115;
  assign _GEN_8117 = 6'h22 == _T_3890 ? _T_3073_34 : _GEN_8116;
  assign _GEN_8118 = 6'h23 == _T_3890 ? _T_3073_35 : _GEN_8117;
  assign _GEN_8119 = 6'h24 == _T_3890 ? _T_3073_36 : _GEN_8118;
  assign _GEN_8120 = 6'h25 == _T_3890 ? _T_3073_37 : _GEN_8119;
  assign _GEN_8121 = 6'h26 == _T_3890 ? _T_3073_38 : _GEN_8120;
  assign _GEN_8122 = 6'h27 == _T_3890 ? _T_3073_39 : _GEN_8121;
  assign _T_3900 = _GEN_97 | reset;
  assign _T_3902 = _T_3900 == 1'h0;
  assign _T_3903 = _T_3889[5:0];
  assign _T_3906 = _T_3200__T_3904_data;
  assign _T_3908 = _T_3906 | reset;
  assign _T_3910 = _T_3908 == 1'h0;
  assign _T_3916 = io_brinfo_rob_idx >> 1'h1;
  assign _T_3975 = io_fflags_0_bits_uop_rob_idx[0];
  assign _T_3977 = _T_3975 == 1'h0;
  assign _T_3978 = io_fflags_0_valid & _T_3977;
  assign _T_3980 = io_fflags_0_bits_uop_rob_idx >> 1'h1;
  assign _T_3981 = _T_3980[5:0];
  assign _T_3983 = io_fflags_1_bits_uop_rob_idx[0];
  assign _T_3985 = _T_3983 == 1'h0;
  assign _T_3986 = io_fflags_1_valid & _T_3985;
  assign _T_3988 = io_fflags_1_bits_uop_rob_idx >> 1'h1;
  assign _T_3989 = _T_3988[5:0];
  assign _T_3991 = io_lxcpt_bits_uop_rob_idx[0];
  assign _T_3993 = _T_3991 == 1'h0;
  assign _T_3994 = io_lxcpt_valid & _T_3993;
  assign _T_3996 = io_lxcpt_bits_uop_rob_idx >> 1'h1;
  assign _T_3997 = _T_3996[5:0];
  assign _T_4000 = io_bxcpt_bits_uop_rob_idx[0];
  assign _T_4002 = _T_4000 == 1'h0;
  assign _T_4003 = io_bxcpt_valid & _T_4002;
  assign _T_4005 = io_bxcpt_bits_uop_rob_idx >> 1'h1;
  assign _T_4006 = _T_4005[5:0];
  assign _GEN_8544 = 6'h1 == rob_head ? _T_3073_1 : _T_3073_0;
  assign _GEN_8545 = 6'h2 == rob_head ? _T_3073_2 : _GEN_8544;
  assign _GEN_8546 = 6'h3 == rob_head ? _T_3073_3 : _GEN_8545;
  assign _GEN_8547 = 6'h4 == rob_head ? _T_3073_4 : _GEN_8546;
  assign _GEN_8548 = 6'h5 == rob_head ? _T_3073_5 : _GEN_8547;
  assign _GEN_8549 = 6'h6 == rob_head ? _T_3073_6 : _GEN_8548;
  assign _GEN_8550 = 6'h7 == rob_head ? _T_3073_7 : _GEN_8549;
  assign _GEN_8551 = 6'h8 == rob_head ? _T_3073_8 : _GEN_8550;
  assign _GEN_8552 = 6'h9 == rob_head ? _T_3073_9 : _GEN_8551;
  assign _GEN_8553 = 6'ha == rob_head ? _T_3073_10 : _GEN_8552;
  assign _GEN_8554 = 6'hb == rob_head ? _T_3073_11 : _GEN_8553;
  assign _GEN_8555 = 6'hc == rob_head ? _T_3073_12 : _GEN_8554;
  assign _GEN_8556 = 6'hd == rob_head ? _T_3073_13 : _GEN_8555;
  assign _GEN_8557 = 6'he == rob_head ? _T_3073_14 : _GEN_8556;
  assign _GEN_8558 = 6'hf == rob_head ? _T_3073_15 : _GEN_8557;
  assign _GEN_8559 = 6'h10 == rob_head ? _T_3073_16 : _GEN_8558;
  assign _GEN_8560 = 6'h11 == rob_head ? _T_3073_17 : _GEN_8559;
  assign _GEN_8561 = 6'h12 == rob_head ? _T_3073_18 : _GEN_8560;
  assign _GEN_8562 = 6'h13 == rob_head ? _T_3073_19 : _GEN_8561;
  assign _GEN_8563 = 6'h14 == rob_head ? _T_3073_20 : _GEN_8562;
  assign _GEN_8564 = 6'h15 == rob_head ? _T_3073_21 : _GEN_8563;
  assign _GEN_8565 = 6'h16 == rob_head ? _T_3073_22 : _GEN_8564;
  assign _GEN_8566 = 6'h17 == rob_head ? _T_3073_23 : _GEN_8565;
  assign _GEN_8567 = 6'h18 == rob_head ? _T_3073_24 : _GEN_8566;
  assign _GEN_8568 = 6'h19 == rob_head ? _T_3073_25 : _GEN_8567;
  assign _GEN_8569 = 6'h1a == rob_head ? _T_3073_26 : _GEN_8568;
  assign _GEN_8570 = 6'h1b == rob_head ? _T_3073_27 : _GEN_8569;
  assign _GEN_8571 = 6'h1c == rob_head ? _T_3073_28 : _GEN_8570;
  assign _GEN_8572 = 6'h1d == rob_head ? _T_3073_29 : _GEN_8571;
  assign _GEN_8573 = 6'h1e == rob_head ? _T_3073_30 : _GEN_8572;
  assign _GEN_8574 = 6'h1f == rob_head ? _T_3073_31 : _GEN_8573;
  assign _GEN_8575 = 6'h20 == rob_head ? _T_3073_32 : _GEN_8574;
  assign _GEN_8576 = 6'h21 == rob_head ? _T_3073_33 : _GEN_8575;
  assign _GEN_8577 = 6'h22 == rob_head ? _T_3073_34 : _GEN_8576;
  assign _GEN_8578 = 6'h23 == rob_head ? _T_3073_35 : _GEN_8577;
  assign _GEN_8579 = 6'h24 == rob_head ? _T_3073_36 : _GEN_8578;
  assign _GEN_8580 = 6'h25 == rob_head ? _T_3073_37 : _GEN_8579;
  assign _GEN_8581 = 6'h26 == rob_head ? _T_3073_38 : _GEN_8580;
  assign _GEN_8582 = 6'h27 == rob_head ? _T_3073_39 : _GEN_8581;
  assign _T_4013 = _GEN_103 & _T_3745__T_4012_data;
  assign _T_4019 = _T_3200__T_4017_data == 1'h0;
  assign _T_4020 = _GEN_104 & _T_4019;
  assign _T_4022 = io_csr_stall == 1'h0;
  assign _T_4023 = _T_4020 & _T_4022;
  assign _T_4026 = rob_state == 2'h2;
  assign _GEN_8583 = _T_4026 ? rob_tail : rob_head;
  assign _GEN_8636 = 6'h1 == _T_4025 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_8643 = 6'h1 == _T_4025 ? _T_3372_1_stale_pdst : _T_3372_0_stale_pdst;
  assign _GEN_8650 = 6'h1 == _T_4025 ? _T_3372_1_is_fencei : _T_3372_0_is_fencei;
  assign _GEN_8651 = 6'h1 == _T_4025 ? _T_3372_1_is_store : _T_3372_0_is_store;
  assign _GEN_8653 = 6'h1 == _T_4025 ? _T_3372_1_is_load : _T_3372_0_is_load;
  assign _GEN_8654 = 6'h1 == _T_4025 ? _T_3372_1_is_sys_pc2epc : _T_3372_0_is_sys_pc2epc;
  assign _GEN_8656 = 6'h1 == _T_4025 ? _T_3372_1_flush_on_commit : _T_3372_0_flush_on_commit;
  assign _GEN_8657 = 6'h1 == _T_4025 ? _T_3372_1_ldst : _T_3372_0_ldst;
  assign _GEN_8662 = 6'h1 == _T_4025 ? _T_3372_1_dst_rtype : _T_3372_0_dst_rtype;
  assign _GEN_8666 = 6'h1 == _T_4025 ? _T_3372_1_fp_val : _T_3372_0_fp_val;
  assign _GEN_8726 = 6'h2 == _T_4025 ? _T_3372_2_pdst : _GEN_8636;
  assign _GEN_8733 = 6'h2 == _T_4025 ? _T_3372_2_stale_pdst : _GEN_8643;
  assign _GEN_8740 = 6'h2 == _T_4025 ? _T_3372_2_is_fencei : _GEN_8650;
  assign _GEN_8741 = 6'h2 == _T_4025 ? _T_3372_2_is_store : _GEN_8651;
  assign _GEN_8743 = 6'h2 == _T_4025 ? _T_3372_2_is_load : _GEN_8653;
  assign _GEN_8744 = 6'h2 == _T_4025 ? _T_3372_2_is_sys_pc2epc : _GEN_8654;
  assign _GEN_8746 = 6'h2 == _T_4025 ? _T_3372_2_flush_on_commit : _GEN_8656;
  assign _GEN_8747 = 6'h2 == _T_4025 ? _T_3372_2_ldst : _GEN_8657;
  assign _GEN_8752 = 6'h2 == _T_4025 ? _T_3372_2_dst_rtype : _GEN_8662;
  assign _GEN_8756 = 6'h2 == _T_4025 ? _T_3372_2_fp_val : _GEN_8666;
  assign _GEN_8816 = 6'h3 == _T_4025 ? _T_3372_3_pdst : _GEN_8726;
  assign _GEN_8823 = 6'h3 == _T_4025 ? _T_3372_3_stale_pdst : _GEN_8733;
  assign _GEN_8830 = 6'h3 == _T_4025 ? _T_3372_3_is_fencei : _GEN_8740;
  assign _GEN_8831 = 6'h3 == _T_4025 ? _T_3372_3_is_store : _GEN_8741;
  assign _GEN_8833 = 6'h3 == _T_4025 ? _T_3372_3_is_load : _GEN_8743;
  assign _GEN_8834 = 6'h3 == _T_4025 ? _T_3372_3_is_sys_pc2epc : _GEN_8744;
  assign _GEN_8836 = 6'h3 == _T_4025 ? _T_3372_3_flush_on_commit : _GEN_8746;
  assign _GEN_8837 = 6'h3 == _T_4025 ? _T_3372_3_ldst : _GEN_8747;
  assign _GEN_8842 = 6'h3 == _T_4025 ? _T_3372_3_dst_rtype : _GEN_8752;
  assign _GEN_8846 = 6'h3 == _T_4025 ? _T_3372_3_fp_val : _GEN_8756;
  assign _GEN_8906 = 6'h4 == _T_4025 ? _T_3372_4_pdst : _GEN_8816;
  assign _GEN_8913 = 6'h4 == _T_4025 ? _T_3372_4_stale_pdst : _GEN_8823;
  assign _GEN_8920 = 6'h4 == _T_4025 ? _T_3372_4_is_fencei : _GEN_8830;
  assign _GEN_8921 = 6'h4 == _T_4025 ? _T_3372_4_is_store : _GEN_8831;
  assign _GEN_8923 = 6'h4 == _T_4025 ? _T_3372_4_is_load : _GEN_8833;
  assign _GEN_8924 = 6'h4 == _T_4025 ? _T_3372_4_is_sys_pc2epc : _GEN_8834;
  assign _GEN_8926 = 6'h4 == _T_4025 ? _T_3372_4_flush_on_commit : _GEN_8836;
  assign _GEN_8927 = 6'h4 == _T_4025 ? _T_3372_4_ldst : _GEN_8837;
  assign _GEN_8932 = 6'h4 == _T_4025 ? _T_3372_4_dst_rtype : _GEN_8842;
  assign _GEN_8936 = 6'h4 == _T_4025 ? _T_3372_4_fp_val : _GEN_8846;
  assign _GEN_8996 = 6'h5 == _T_4025 ? _T_3372_5_pdst : _GEN_8906;
  assign _GEN_9003 = 6'h5 == _T_4025 ? _T_3372_5_stale_pdst : _GEN_8913;
  assign _GEN_9010 = 6'h5 == _T_4025 ? _T_3372_5_is_fencei : _GEN_8920;
  assign _GEN_9011 = 6'h5 == _T_4025 ? _T_3372_5_is_store : _GEN_8921;
  assign _GEN_9013 = 6'h5 == _T_4025 ? _T_3372_5_is_load : _GEN_8923;
  assign _GEN_9014 = 6'h5 == _T_4025 ? _T_3372_5_is_sys_pc2epc : _GEN_8924;
  assign _GEN_9016 = 6'h5 == _T_4025 ? _T_3372_5_flush_on_commit : _GEN_8926;
  assign _GEN_9017 = 6'h5 == _T_4025 ? _T_3372_5_ldst : _GEN_8927;
  assign _GEN_9022 = 6'h5 == _T_4025 ? _T_3372_5_dst_rtype : _GEN_8932;
  assign _GEN_9026 = 6'h5 == _T_4025 ? _T_3372_5_fp_val : _GEN_8936;
  assign _GEN_9086 = 6'h6 == _T_4025 ? _T_3372_6_pdst : _GEN_8996;
  assign _GEN_9093 = 6'h6 == _T_4025 ? _T_3372_6_stale_pdst : _GEN_9003;
  assign _GEN_9100 = 6'h6 == _T_4025 ? _T_3372_6_is_fencei : _GEN_9010;
  assign _GEN_9101 = 6'h6 == _T_4025 ? _T_3372_6_is_store : _GEN_9011;
  assign _GEN_9103 = 6'h6 == _T_4025 ? _T_3372_6_is_load : _GEN_9013;
  assign _GEN_9104 = 6'h6 == _T_4025 ? _T_3372_6_is_sys_pc2epc : _GEN_9014;
  assign _GEN_9106 = 6'h6 == _T_4025 ? _T_3372_6_flush_on_commit : _GEN_9016;
  assign _GEN_9107 = 6'h6 == _T_4025 ? _T_3372_6_ldst : _GEN_9017;
  assign _GEN_9112 = 6'h6 == _T_4025 ? _T_3372_6_dst_rtype : _GEN_9022;
  assign _GEN_9116 = 6'h6 == _T_4025 ? _T_3372_6_fp_val : _GEN_9026;
  assign _GEN_9176 = 6'h7 == _T_4025 ? _T_3372_7_pdst : _GEN_9086;
  assign _GEN_9183 = 6'h7 == _T_4025 ? _T_3372_7_stale_pdst : _GEN_9093;
  assign _GEN_9190 = 6'h7 == _T_4025 ? _T_3372_7_is_fencei : _GEN_9100;
  assign _GEN_9191 = 6'h7 == _T_4025 ? _T_3372_7_is_store : _GEN_9101;
  assign _GEN_9193 = 6'h7 == _T_4025 ? _T_3372_7_is_load : _GEN_9103;
  assign _GEN_9194 = 6'h7 == _T_4025 ? _T_3372_7_is_sys_pc2epc : _GEN_9104;
  assign _GEN_9196 = 6'h7 == _T_4025 ? _T_3372_7_flush_on_commit : _GEN_9106;
  assign _GEN_9197 = 6'h7 == _T_4025 ? _T_3372_7_ldst : _GEN_9107;
  assign _GEN_9202 = 6'h7 == _T_4025 ? _T_3372_7_dst_rtype : _GEN_9112;
  assign _GEN_9206 = 6'h7 == _T_4025 ? _T_3372_7_fp_val : _GEN_9116;
  assign _GEN_9266 = 6'h8 == _T_4025 ? _T_3372_8_pdst : _GEN_9176;
  assign _GEN_9273 = 6'h8 == _T_4025 ? _T_3372_8_stale_pdst : _GEN_9183;
  assign _GEN_9280 = 6'h8 == _T_4025 ? _T_3372_8_is_fencei : _GEN_9190;
  assign _GEN_9281 = 6'h8 == _T_4025 ? _T_3372_8_is_store : _GEN_9191;
  assign _GEN_9283 = 6'h8 == _T_4025 ? _T_3372_8_is_load : _GEN_9193;
  assign _GEN_9284 = 6'h8 == _T_4025 ? _T_3372_8_is_sys_pc2epc : _GEN_9194;
  assign _GEN_9286 = 6'h8 == _T_4025 ? _T_3372_8_flush_on_commit : _GEN_9196;
  assign _GEN_9287 = 6'h8 == _T_4025 ? _T_3372_8_ldst : _GEN_9197;
  assign _GEN_9292 = 6'h8 == _T_4025 ? _T_3372_8_dst_rtype : _GEN_9202;
  assign _GEN_9296 = 6'h8 == _T_4025 ? _T_3372_8_fp_val : _GEN_9206;
  assign _GEN_9356 = 6'h9 == _T_4025 ? _T_3372_9_pdst : _GEN_9266;
  assign _GEN_9363 = 6'h9 == _T_4025 ? _T_3372_9_stale_pdst : _GEN_9273;
  assign _GEN_9370 = 6'h9 == _T_4025 ? _T_3372_9_is_fencei : _GEN_9280;
  assign _GEN_9371 = 6'h9 == _T_4025 ? _T_3372_9_is_store : _GEN_9281;
  assign _GEN_9373 = 6'h9 == _T_4025 ? _T_3372_9_is_load : _GEN_9283;
  assign _GEN_9374 = 6'h9 == _T_4025 ? _T_3372_9_is_sys_pc2epc : _GEN_9284;
  assign _GEN_9376 = 6'h9 == _T_4025 ? _T_3372_9_flush_on_commit : _GEN_9286;
  assign _GEN_9377 = 6'h9 == _T_4025 ? _T_3372_9_ldst : _GEN_9287;
  assign _GEN_9382 = 6'h9 == _T_4025 ? _T_3372_9_dst_rtype : _GEN_9292;
  assign _GEN_9386 = 6'h9 == _T_4025 ? _T_3372_9_fp_val : _GEN_9296;
  assign _GEN_9446 = 6'ha == _T_4025 ? _T_3372_10_pdst : _GEN_9356;
  assign _GEN_9453 = 6'ha == _T_4025 ? _T_3372_10_stale_pdst : _GEN_9363;
  assign _GEN_9460 = 6'ha == _T_4025 ? _T_3372_10_is_fencei : _GEN_9370;
  assign _GEN_9461 = 6'ha == _T_4025 ? _T_3372_10_is_store : _GEN_9371;
  assign _GEN_9463 = 6'ha == _T_4025 ? _T_3372_10_is_load : _GEN_9373;
  assign _GEN_9464 = 6'ha == _T_4025 ? _T_3372_10_is_sys_pc2epc : _GEN_9374;
  assign _GEN_9466 = 6'ha == _T_4025 ? _T_3372_10_flush_on_commit : _GEN_9376;
  assign _GEN_9467 = 6'ha == _T_4025 ? _T_3372_10_ldst : _GEN_9377;
  assign _GEN_9472 = 6'ha == _T_4025 ? _T_3372_10_dst_rtype : _GEN_9382;
  assign _GEN_9476 = 6'ha == _T_4025 ? _T_3372_10_fp_val : _GEN_9386;
  assign _GEN_9536 = 6'hb == _T_4025 ? _T_3372_11_pdst : _GEN_9446;
  assign _GEN_9543 = 6'hb == _T_4025 ? _T_3372_11_stale_pdst : _GEN_9453;
  assign _GEN_9550 = 6'hb == _T_4025 ? _T_3372_11_is_fencei : _GEN_9460;
  assign _GEN_9551 = 6'hb == _T_4025 ? _T_3372_11_is_store : _GEN_9461;
  assign _GEN_9553 = 6'hb == _T_4025 ? _T_3372_11_is_load : _GEN_9463;
  assign _GEN_9554 = 6'hb == _T_4025 ? _T_3372_11_is_sys_pc2epc : _GEN_9464;
  assign _GEN_9556 = 6'hb == _T_4025 ? _T_3372_11_flush_on_commit : _GEN_9466;
  assign _GEN_9557 = 6'hb == _T_4025 ? _T_3372_11_ldst : _GEN_9467;
  assign _GEN_9562 = 6'hb == _T_4025 ? _T_3372_11_dst_rtype : _GEN_9472;
  assign _GEN_9566 = 6'hb == _T_4025 ? _T_3372_11_fp_val : _GEN_9476;
  assign _GEN_9626 = 6'hc == _T_4025 ? _T_3372_12_pdst : _GEN_9536;
  assign _GEN_9633 = 6'hc == _T_4025 ? _T_3372_12_stale_pdst : _GEN_9543;
  assign _GEN_9640 = 6'hc == _T_4025 ? _T_3372_12_is_fencei : _GEN_9550;
  assign _GEN_9641 = 6'hc == _T_4025 ? _T_3372_12_is_store : _GEN_9551;
  assign _GEN_9643 = 6'hc == _T_4025 ? _T_3372_12_is_load : _GEN_9553;
  assign _GEN_9644 = 6'hc == _T_4025 ? _T_3372_12_is_sys_pc2epc : _GEN_9554;
  assign _GEN_9646 = 6'hc == _T_4025 ? _T_3372_12_flush_on_commit : _GEN_9556;
  assign _GEN_9647 = 6'hc == _T_4025 ? _T_3372_12_ldst : _GEN_9557;
  assign _GEN_9652 = 6'hc == _T_4025 ? _T_3372_12_dst_rtype : _GEN_9562;
  assign _GEN_9656 = 6'hc == _T_4025 ? _T_3372_12_fp_val : _GEN_9566;
  assign _GEN_9716 = 6'hd == _T_4025 ? _T_3372_13_pdst : _GEN_9626;
  assign _GEN_9723 = 6'hd == _T_4025 ? _T_3372_13_stale_pdst : _GEN_9633;
  assign _GEN_9730 = 6'hd == _T_4025 ? _T_3372_13_is_fencei : _GEN_9640;
  assign _GEN_9731 = 6'hd == _T_4025 ? _T_3372_13_is_store : _GEN_9641;
  assign _GEN_9733 = 6'hd == _T_4025 ? _T_3372_13_is_load : _GEN_9643;
  assign _GEN_9734 = 6'hd == _T_4025 ? _T_3372_13_is_sys_pc2epc : _GEN_9644;
  assign _GEN_9736 = 6'hd == _T_4025 ? _T_3372_13_flush_on_commit : _GEN_9646;
  assign _GEN_9737 = 6'hd == _T_4025 ? _T_3372_13_ldst : _GEN_9647;
  assign _GEN_9742 = 6'hd == _T_4025 ? _T_3372_13_dst_rtype : _GEN_9652;
  assign _GEN_9746 = 6'hd == _T_4025 ? _T_3372_13_fp_val : _GEN_9656;
  assign _GEN_9806 = 6'he == _T_4025 ? _T_3372_14_pdst : _GEN_9716;
  assign _GEN_9813 = 6'he == _T_4025 ? _T_3372_14_stale_pdst : _GEN_9723;
  assign _GEN_9820 = 6'he == _T_4025 ? _T_3372_14_is_fencei : _GEN_9730;
  assign _GEN_9821 = 6'he == _T_4025 ? _T_3372_14_is_store : _GEN_9731;
  assign _GEN_9823 = 6'he == _T_4025 ? _T_3372_14_is_load : _GEN_9733;
  assign _GEN_9824 = 6'he == _T_4025 ? _T_3372_14_is_sys_pc2epc : _GEN_9734;
  assign _GEN_9826 = 6'he == _T_4025 ? _T_3372_14_flush_on_commit : _GEN_9736;
  assign _GEN_9827 = 6'he == _T_4025 ? _T_3372_14_ldst : _GEN_9737;
  assign _GEN_9832 = 6'he == _T_4025 ? _T_3372_14_dst_rtype : _GEN_9742;
  assign _GEN_9836 = 6'he == _T_4025 ? _T_3372_14_fp_val : _GEN_9746;
  assign _GEN_9896 = 6'hf == _T_4025 ? _T_3372_15_pdst : _GEN_9806;
  assign _GEN_9903 = 6'hf == _T_4025 ? _T_3372_15_stale_pdst : _GEN_9813;
  assign _GEN_9910 = 6'hf == _T_4025 ? _T_3372_15_is_fencei : _GEN_9820;
  assign _GEN_9911 = 6'hf == _T_4025 ? _T_3372_15_is_store : _GEN_9821;
  assign _GEN_9913 = 6'hf == _T_4025 ? _T_3372_15_is_load : _GEN_9823;
  assign _GEN_9914 = 6'hf == _T_4025 ? _T_3372_15_is_sys_pc2epc : _GEN_9824;
  assign _GEN_9916 = 6'hf == _T_4025 ? _T_3372_15_flush_on_commit : _GEN_9826;
  assign _GEN_9917 = 6'hf == _T_4025 ? _T_3372_15_ldst : _GEN_9827;
  assign _GEN_9922 = 6'hf == _T_4025 ? _T_3372_15_dst_rtype : _GEN_9832;
  assign _GEN_9926 = 6'hf == _T_4025 ? _T_3372_15_fp_val : _GEN_9836;
  assign _GEN_9986 = 6'h10 == _T_4025 ? _T_3372_16_pdst : _GEN_9896;
  assign _GEN_9993 = 6'h10 == _T_4025 ? _T_3372_16_stale_pdst : _GEN_9903;
  assign _GEN_10000 = 6'h10 == _T_4025 ? _T_3372_16_is_fencei : _GEN_9910;
  assign _GEN_10001 = 6'h10 == _T_4025 ? _T_3372_16_is_store : _GEN_9911;
  assign _GEN_10003 = 6'h10 == _T_4025 ? _T_3372_16_is_load : _GEN_9913;
  assign _GEN_10004 = 6'h10 == _T_4025 ? _T_3372_16_is_sys_pc2epc : _GEN_9914;
  assign _GEN_10006 = 6'h10 == _T_4025 ? _T_3372_16_flush_on_commit : _GEN_9916;
  assign _GEN_10007 = 6'h10 == _T_4025 ? _T_3372_16_ldst : _GEN_9917;
  assign _GEN_10012 = 6'h10 == _T_4025 ? _T_3372_16_dst_rtype : _GEN_9922;
  assign _GEN_10016 = 6'h10 == _T_4025 ? _T_3372_16_fp_val : _GEN_9926;
  assign _GEN_10076 = 6'h11 == _T_4025 ? _T_3372_17_pdst : _GEN_9986;
  assign _GEN_10083 = 6'h11 == _T_4025 ? _T_3372_17_stale_pdst : _GEN_9993;
  assign _GEN_10090 = 6'h11 == _T_4025 ? _T_3372_17_is_fencei : _GEN_10000;
  assign _GEN_10091 = 6'h11 == _T_4025 ? _T_3372_17_is_store : _GEN_10001;
  assign _GEN_10093 = 6'h11 == _T_4025 ? _T_3372_17_is_load : _GEN_10003;
  assign _GEN_10094 = 6'h11 == _T_4025 ? _T_3372_17_is_sys_pc2epc : _GEN_10004;
  assign _GEN_10096 = 6'h11 == _T_4025 ? _T_3372_17_flush_on_commit : _GEN_10006;
  assign _GEN_10097 = 6'h11 == _T_4025 ? _T_3372_17_ldst : _GEN_10007;
  assign _GEN_10102 = 6'h11 == _T_4025 ? _T_3372_17_dst_rtype : _GEN_10012;
  assign _GEN_10106 = 6'h11 == _T_4025 ? _T_3372_17_fp_val : _GEN_10016;
  assign _GEN_10166 = 6'h12 == _T_4025 ? _T_3372_18_pdst : _GEN_10076;
  assign _GEN_10173 = 6'h12 == _T_4025 ? _T_3372_18_stale_pdst : _GEN_10083;
  assign _GEN_10180 = 6'h12 == _T_4025 ? _T_3372_18_is_fencei : _GEN_10090;
  assign _GEN_10181 = 6'h12 == _T_4025 ? _T_3372_18_is_store : _GEN_10091;
  assign _GEN_10183 = 6'h12 == _T_4025 ? _T_3372_18_is_load : _GEN_10093;
  assign _GEN_10184 = 6'h12 == _T_4025 ? _T_3372_18_is_sys_pc2epc : _GEN_10094;
  assign _GEN_10186 = 6'h12 == _T_4025 ? _T_3372_18_flush_on_commit : _GEN_10096;
  assign _GEN_10187 = 6'h12 == _T_4025 ? _T_3372_18_ldst : _GEN_10097;
  assign _GEN_10192 = 6'h12 == _T_4025 ? _T_3372_18_dst_rtype : _GEN_10102;
  assign _GEN_10196 = 6'h12 == _T_4025 ? _T_3372_18_fp_val : _GEN_10106;
  assign _GEN_10256 = 6'h13 == _T_4025 ? _T_3372_19_pdst : _GEN_10166;
  assign _GEN_10263 = 6'h13 == _T_4025 ? _T_3372_19_stale_pdst : _GEN_10173;
  assign _GEN_10270 = 6'h13 == _T_4025 ? _T_3372_19_is_fencei : _GEN_10180;
  assign _GEN_10271 = 6'h13 == _T_4025 ? _T_3372_19_is_store : _GEN_10181;
  assign _GEN_10273 = 6'h13 == _T_4025 ? _T_3372_19_is_load : _GEN_10183;
  assign _GEN_10274 = 6'h13 == _T_4025 ? _T_3372_19_is_sys_pc2epc : _GEN_10184;
  assign _GEN_10276 = 6'h13 == _T_4025 ? _T_3372_19_flush_on_commit : _GEN_10186;
  assign _GEN_10277 = 6'h13 == _T_4025 ? _T_3372_19_ldst : _GEN_10187;
  assign _GEN_10282 = 6'h13 == _T_4025 ? _T_3372_19_dst_rtype : _GEN_10192;
  assign _GEN_10286 = 6'h13 == _T_4025 ? _T_3372_19_fp_val : _GEN_10196;
  assign _GEN_10346 = 6'h14 == _T_4025 ? _T_3372_20_pdst : _GEN_10256;
  assign _GEN_10353 = 6'h14 == _T_4025 ? _T_3372_20_stale_pdst : _GEN_10263;
  assign _GEN_10360 = 6'h14 == _T_4025 ? _T_3372_20_is_fencei : _GEN_10270;
  assign _GEN_10361 = 6'h14 == _T_4025 ? _T_3372_20_is_store : _GEN_10271;
  assign _GEN_10363 = 6'h14 == _T_4025 ? _T_3372_20_is_load : _GEN_10273;
  assign _GEN_10364 = 6'h14 == _T_4025 ? _T_3372_20_is_sys_pc2epc : _GEN_10274;
  assign _GEN_10366 = 6'h14 == _T_4025 ? _T_3372_20_flush_on_commit : _GEN_10276;
  assign _GEN_10367 = 6'h14 == _T_4025 ? _T_3372_20_ldst : _GEN_10277;
  assign _GEN_10372 = 6'h14 == _T_4025 ? _T_3372_20_dst_rtype : _GEN_10282;
  assign _GEN_10376 = 6'h14 == _T_4025 ? _T_3372_20_fp_val : _GEN_10286;
  assign _GEN_10436 = 6'h15 == _T_4025 ? _T_3372_21_pdst : _GEN_10346;
  assign _GEN_10443 = 6'h15 == _T_4025 ? _T_3372_21_stale_pdst : _GEN_10353;
  assign _GEN_10450 = 6'h15 == _T_4025 ? _T_3372_21_is_fencei : _GEN_10360;
  assign _GEN_10451 = 6'h15 == _T_4025 ? _T_3372_21_is_store : _GEN_10361;
  assign _GEN_10453 = 6'h15 == _T_4025 ? _T_3372_21_is_load : _GEN_10363;
  assign _GEN_10454 = 6'h15 == _T_4025 ? _T_3372_21_is_sys_pc2epc : _GEN_10364;
  assign _GEN_10456 = 6'h15 == _T_4025 ? _T_3372_21_flush_on_commit : _GEN_10366;
  assign _GEN_10457 = 6'h15 == _T_4025 ? _T_3372_21_ldst : _GEN_10367;
  assign _GEN_10462 = 6'h15 == _T_4025 ? _T_3372_21_dst_rtype : _GEN_10372;
  assign _GEN_10466 = 6'h15 == _T_4025 ? _T_3372_21_fp_val : _GEN_10376;
  assign _GEN_10526 = 6'h16 == _T_4025 ? _T_3372_22_pdst : _GEN_10436;
  assign _GEN_10533 = 6'h16 == _T_4025 ? _T_3372_22_stale_pdst : _GEN_10443;
  assign _GEN_10540 = 6'h16 == _T_4025 ? _T_3372_22_is_fencei : _GEN_10450;
  assign _GEN_10541 = 6'h16 == _T_4025 ? _T_3372_22_is_store : _GEN_10451;
  assign _GEN_10543 = 6'h16 == _T_4025 ? _T_3372_22_is_load : _GEN_10453;
  assign _GEN_10544 = 6'h16 == _T_4025 ? _T_3372_22_is_sys_pc2epc : _GEN_10454;
  assign _GEN_10546 = 6'h16 == _T_4025 ? _T_3372_22_flush_on_commit : _GEN_10456;
  assign _GEN_10547 = 6'h16 == _T_4025 ? _T_3372_22_ldst : _GEN_10457;
  assign _GEN_10552 = 6'h16 == _T_4025 ? _T_3372_22_dst_rtype : _GEN_10462;
  assign _GEN_10556 = 6'h16 == _T_4025 ? _T_3372_22_fp_val : _GEN_10466;
  assign _GEN_10616 = 6'h17 == _T_4025 ? _T_3372_23_pdst : _GEN_10526;
  assign _GEN_10623 = 6'h17 == _T_4025 ? _T_3372_23_stale_pdst : _GEN_10533;
  assign _GEN_10630 = 6'h17 == _T_4025 ? _T_3372_23_is_fencei : _GEN_10540;
  assign _GEN_10631 = 6'h17 == _T_4025 ? _T_3372_23_is_store : _GEN_10541;
  assign _GEN_10633 = 6'h17 == _T_4025 ? _T_3372_23_is_load : _GEN_10543;
  assign _GEN_10634 = 6'h17 == _T_4025 ? _T_3372_23_is_sys_pc2epc : _GEN_10544;
  assign _GEN_10636 = 6'h17 == _T_4025 ? _T_3372_23_flush_on_commit : _GEN_10546;
  assign _GEN_10637 = 6'h17 == _T_4025 ? _T_3372_23_ldst : _GEN_10547;
  assign _GEN_10642 = 6'h17 == _T_4025 ? _T_3372_23_dst_rtype : _GEN_10552;
  assign _GEN_10646 = 6'h17 == _T_4025 ? _T_3372_23_fp_val : _GEN_10556;
  assign _GEN_10706 = 6'h18 == _T_4025 ? _T_3372_24_pdst : _GEN_10616;
  assign _GEN_10713 = 6'h18 == _T_4025 ? _T_3372_24_stale_pdst : _GEN_10623;
  assign _GEN_10720 = 6'h18 == _T_4025 ? _T_3372_24_is_fencei : _GEN_10630;
  assign _GEN_10721 = 6'h18 == _T_4025 ? _T_3372_24_is_store : _GEN_10631;
  assign _GEN_10723 = 6'h18 == _T_4025 ? _T_3372_24_is_load : _GEN_10633;
  assign _GEN_10724 = 6'h18 == _T_4025 ? _T_3372_24_is_sys_pc2epc : _GEN_10634;
  assign _GEN_10726 = 6'h18 == _T_4025 ? _T_3372_24_flush_on_commit : _GEN_10636;
  assign _GEN_10727 = 6'h18 == _T_4025 ? _T_3372_24_ldst : _GEN_10637;
  assign _GEN_10732 = 6'h18 == _T_4025 ? _T_3372_24_dst_rtype : _GEN_10642;
  assign _GEN_10736 = 6'h18 == _T_4025 ? _T_3372_24_fp_val : _GEN_10646;
  assign _GEN_10796 = 6'h19 == _T_4025 ? _T_3372_25_pdst : _GEN_10706;
  assign _GEN_10803 = 6'h19 == _T_4025 ? _T_3372_25_stale_pdst : _GEN_10713;
  assign _GEN_10810 = 6'h19 == _T_4025 ? _T_3372_25_is_fencei : _GEN_10720;
  assign _GEN_10811 = 6'h19 == _T_4025 ? _T_3372_25_is_store : _GEN_10721;
  assign _GEN_10813 = 6'h19 == _T_4025 ? _T_3372_25_is_load : _GEN_10723;
  assign _GEN_10814 = 6'h19 == _T_4025 ? _T_3372_25_is_sys_pc2epc : _GEN_10724;
  assign _GEN_10816 = 6'h19 == _T_4025 ? _T_3372_25_flush_on_commit : _GEN_10726;
  assign _GEN_10817 = 6'h19 == _T_4025 ? _T_3372_25_ldst : _GEN_10727;
  assign _GEN_10822 = 6'h19 == _T_4025 ? _T_3372_25_dst_rtype : _GEN_10732;
  assign _GEN_10826 = 6'h19 == _T_4025 ? _T_3372_25_fp_val : _GEN_10736;
  assign _GEN_10886 = 6'h1a == _T_4025 ? _T_3372_26_pdst : _GEN_10796;
  assign _GEN_10893 = 6'h1a == _T_4025 ? _T_3372_26_stale_pdst : _GEN_10803;
  assign _GEN_10900 = 6'h1a == _T_4025 ? _T_3372_26_is_fencei : _GEN_10810;
  assign _GEN_10901 = 6'h1a == _T_4025 ? _T_3372_26_is_store : _GEN_10811;
  assign _GEN_10903 = 6'h1a == _T_4025 ? _T_3372_26_is_load : _GEN_10813;
  assign _GEN_10904 = 6'h1a == _T_4025 ? _T_3372_26_is_sys_pc2epc : _GEN_10814;
  assign _GEN_10906 = 6'h1a == _T_4025 ? _T_3372_26_flush_on_commit : _GEN_10816;
  assign _GEN_10907 = 6'h1a == _T_4025 ? _T_3372_26_ldst : _GEN_10817;
  assign _GEN_10912 = 6'h1a == _T_4025 ? _T_3372_26_dst_rtype : _GEN_10822;
  assign _GEN_10916 = 6'h1a == _T_4025 ? _T_3372_26_fp_val : _GEN_10826;
  assign _GEN_10976 = 6'h1b == _T_4025 ? _T_3372_27_pdst : _GEN_10886;
  assign _GEN_10983 = 6'h1b == _T_4025 ? _T_3372_27_stale_pdst : _GEN_10893;
  assign _GEN_10990 = 6'h1b == _T_4025 ? _T_3372_27_is_fencei : _GEN_10900;
  assign _GEN_10991 = 6'h1b == _T_4025 ? _T_3372_27_is_store : _GEN_10901;
  assign _GEN_10993 = 6'h1b == _T_4025 ? _T_3372_27_is_load : _GEN_10903;
  assign _GEN_10994 = 6'h1b == _T_4025 ? _T_3372_27_is_sys_pc2epc : _GEN_10904;
  assign _GEN_10996 = 6'h1b == _T_4025 ? _T_3372_27_flush_on_commit : _GEN_10906;
  assign _GEN_10997 = 6'h1b == _T_4025 ? _T_3372_27_ldst : _GEN_10907;
  assign _GEN_11002 = 6'h1b == _T_4025 ? _T_3372_27_dst_rtype : _GEN_10912;
  assign _GEN_11006 = 6'h1b == _T_4025 ? _T_3372_27_fp_val : _GEN_10916;
  assign _GEN_11066 = 6'h1c == _T_4025 ? _T_3372_28_pdst : _GEN_10976;
  assign _GEN_11073 = 6'h1c == _T_4025 ? _T_3372_28_stale_pdst : _GEN_10983;
  assign _GEN_11080 = 6'h1c == _T_4025 ? _T_3372_28_is_fencei : _GEN_10990;
  assign _GEN_11081 = 6'h1c == _T_4025 ? _T_3372_28_is_store : _GEN_10991;
  assign _GEN_11083 = 6'h1c == _T_4025 ? _T_3372_28_is_load : _GEN_10993;
  assign _GEN_11084 = 6'h1c == _T_4025 ? _T_3372_28_is_sys_pc2epc : _GEN_10994;
  assign _GEN_11086 = 6'h1c == _T_4025 ? _T_3372_28_flush_on_commit : _GEN_10996;
  assign _GEN_11087 = 6'h1c == _T_4025 ? _T_3372_28_ldst : _GEN_10997;
  assign _GEN_11092 = 6'h1c == _T_4025 ? _T_3372_28_dst_rtype : _GEN_11002;
  assign _GEN_11096 = 6'h1c == _T_4025 ? _T_3372_28_fp_val : _GEN_11006;
  assign _GEN_11156 = 6'h1d == _T_4025 ? _T_3372_29_pdst : _GEN_11066;
  assign _GEN_11163 = 6'h1d == _T_4025 ? _T_3372_29_stale_pdst : _GEN_11073;
  assign _GEN_11170 = 6'h1d == _T_4025 ? _T_3372_29_is_fencei : _GEN_11080;
  assign _GEN_11171 = 6'h1d == _T_4025 ? _T_3372_29_is_store : _GEN_11081;
  assign _GEN_11173 = 6'h1d == _T_4025 ? _T_3372_29_is_load : _GEN_11083;
  assign _GEN_11174 = 6'h1d == _T_4025 ? _T_3372_29_is_sys_pc2epc : _GEN_11084;
  assign _GEN_11176 = 6'h1d == _T_4025 ? _T_3372_29_flush_on_commit : _GEN_11086;
  assign _GEN_11177 = 6'h1d == _T_4025 ? _T_3372_29_ldst : _GEN_11087;
  assign _GEN_11182 = 6'h1d == _T_4025 ? _T_3372_29_dst_rtype : _GEN_11092;
  assign _GEN_11186 = 6'h1d == _T_4025 ? _T_3372_29_fp_val : _GEN_11096;
  assign _GEN_11246 = 6'h1e == _T_4025 ? _T_3372_30_pdst : _GEN_11156;
  assign _GEN_11253 = 6'h1e == _T_4025 ? _T_3372_30_stale_pdst : _GEN_11163;
  assign _GEN_11260 = 6'h1e == _T_4025 ? _T_3372_30_is_fencei : _GEN_11170;
  assign _GEN_11261 = 6'h1e == _T_4025 ? _T_3372_30_is_store : _GEN_11171;
  assign _GEN_11263 = 6'h1e == _T_4025 ? _T_3372_30_is_load : _GEN_11173;
  assign _GEN_11264 = 6'h1e == _T_4025 ? _T_3372_30_is_sys_pc2epc : _GEN_11174;
  assign _GEN_11266 = 6'h1e == _T_4025 ? _T_3372_30_flush_on_commit : _GEN_11176;
  assign _GEN_11267 = 6'h1e == _T_4025 ? _T_3372_30_ldst : _GEN_11177;
  assign _GEN_11272 = 6'h1e == _T_4025 ? _T_3372_30_dst_rtype : _GEN_11182;
  assign _GEN_11276 = 6'h1e == _T_4025 ? _T_3372_30_fp_val : _GEN_11186;
  assign _GEN_11336 = 6'h1f == _T_4025 ? _T_3372_31_pdst : _GEN_11246;
  assign _GEN_11343 = 6'h1f == _T_4025 ? _T_3372_31_stale_pdst : _GEN_11253;
  assign _GEN_11350 = 6'h1f == _T_4025 ? _T_3372_31_is_fencei : _GEN_11260;
  assign _GEN_11351 = 6'h1f == _T_4025 ? _T_3372_31_is_store : _GEN_11261;
  assign _GEN_11353 = 6'h1f == _T_4025 ? _T_3372_31_is_load : _GEN_11263;
  assign _GEN_11354 = 6'h1f == _T_4025 ? _T_3372_31_is_sys_pc2epc : _GEN_11264;
  assign _GEN_11356 = 6'h1f == _T_4025 ? _T_3372_31_flush_on_commit : _GEN_11266;
  assign _GEN_11357 = 6'h1f == _T_4025 ? _T_3372_31_ldst : _GEN_11267;
  assign _GEN_11362 = 6'h1f == _T_4025 ? _T_3372_31_dst_rtype : _GEN_11272;
  assign _GEN_11366 = 6'h1f == _T_4025 ? _T_3372_31_fp_val : _GEN_11276;
  assign _GEN_11426 = 6'h20 == _T_4025 ? _T_3372_32_pdst : _GEN_11336;
  assign _GEN_11433 = 6'h20 == _T_4025 ? _T_3372_32_stale_pdst : _GEN_11343;
  assign _GEN_11440 = 6'h20 == _T_4025 ? _T_3372_32_is_fencei : _GEN_11350;
  assign _GEN_11441 = 6'h20 == _T_4025 ? _T_3372_32_is_store : _GEN_11351;
  assign _GEN_11443 = 6'h20 == _T_4025 ? _T_3372_32_is_load : _GEN_11353;
  assign _GEN_11444 = 6'h20 == _T_4025 ? _T_3372_32_is_sys_pc2epc : _GEN_11354;
  assign _GEN_11446 = 6'h20 == _T_4025 ? _T_3372_32_flush_on_commit : _GEN_11356;
  assign _GEN_11447 = 6'h20 == _T_4025 ? _T_3372_32_ldst : _GEN_11357;
  assign _GEN_11452 = 6'h20 == _T_4025 ? _T_3372_32_dst_rtype : _GEN_11362;
  assign _GEN_11456 = 6'h20 == _T_4025 ? _T_3372_32_fp_val : _GEN_11366;
  assign _GEN_11516 = 6'h21 == _T_4025 ? _T_3372_33_pdst : _GEN_11426;
  assign _GEN_11523 = 6'h21 == _T_4025 ? _T_3372_33_stale_pdst : _GEN_11433;
  assign _GEN_11530 = 6'h21 == _T_4025 ? _T_3372_33_is_fencei : _GEN_11440;
  assign _GEN_11531 = 6'h21 == _T_4025 ? _T_3372_33_is_store : _GEN_11441;
  assign _GEN_11533 = 6'h21 == _T_4025 ? _T_3372_33_is_load : _GEN_11443;
  assign _GEN_11534 = 6'h21 == _T_4025 ? _T_3372_33_is_sys_pc2epc : _GEN_11444;
  assign _GEN_11536 = 6'h21 == _T_4025 ? _T_3372_33_flush_on_commit : _GEN_11446;
  assign _GEN_11537 = 6'h21 == _T_4025 ? _T_3372_33_ldst : _GEN_11447;
  assign _GEN_11542 = 6'h21 == _T_4025 ? _T_3372_33_dst_rtype : _GEN_11452;
  assign _GEN_11546 = 6'h21 == _T_4025 ? _T_3372_33_fp_val : _GEN_11456;
  assign _GEN_11606 = 6'h22 == _T_4025 ? _T_3372_34_pdst : _GEN_11516;
  assign _GEN_11613 = 6'h22 == _T_4025 ? _T_3372_34_stale_pdst : _GEN_11523;
  assign _GEN_11620 = 6'h22 == _T_4025 ? _T_3372_34_is_fencei : _GEN_11530;
  assign _GEN_11621 = 6'h22 == _T_4025 ? _T_3372_34_is_store : _GEN_11531;
  assign _GEN_11623 = 6'h22 == _T_4025 ? _T_3372_34_is_load : _GEN_11533;
  assign _GEN_11624 = 6'h22 == _T_4025 ? _T_3372_34_is_sys_pc2epc : _GEN_11534;
  assign _GEN_11626 = 6'h22 == _T_4025 ? _T_3372_34_flush_on_commit : _GEN_11536;
  assign _GEN_11627 = 6'h22 == _T_4025 ? _T_3372_34_ldst : _GEN_11537;
  assign _GEN_11632 = 6'h22 == _T_4025 ? _T_3372_34_dst_rtype : _GEN_11542;
  assign _GEN_11636 = 6'h22 == _T_4025 ? _T_3372_34_fp_val : _GEN_11546;
  assign _GEN_11696 = 6'h23 == _T_4025 ? _T_3372_35_pdst : _GEN_11606;
  assign _GEN_11703 = 6'h23 == _T_4025 ? _T_3372_35_stale_pdst : _GEN_11613;
  assign _GEN_11710 = 6'h23 == _T_4025 ? _T_3372_35_is_fencei : _GEN_11620;
  assign _GEN_11711 = 6'h23 == _T_4025 ? _T_3372_35_is_store : _GEN_11621;
  assign _GEN_11713 = 6'h23 == _T_4025 ? _T_3372_35_is_load : _GEN_11623;
  assign _GEN_11714 = 6'h23 == _T_4025 ? _T_3372_35_is_sys_pc2epc : _GEN_11624;
  assign _GEN_11716 = 6'h23 == _T_4025 ? _T_3372_35_flush_on_commit : _GEN_11626;
  assign _GEN_11717 = 6'h23 == _T_4025 ? _T_3372_35_ldst : _GEN_11627;
  assign _GEN_11722 = 6'h23 == _T_4025 ? _T_3372_35_dst_rtype : _GEN_11632;
  assign _GEN_11726 = 6'h23 == _T_4025 ? _T_3372_35_fp_val : _GEN_11636;
  assign _GEN_11786 = 6'h24 == _T_4025 ? _T_3372_36_pdst : _GEN_11696;
  assign _GEN_11793 = 6'h24 == _T_4025 ? _T_3372_36_stale_pdst : _GEN_11703;
  assign _GEN_11800 = 6'h24 == _T_4025 ? _T_3372_36_is_fencei : _GEN_11710;
  assign _GEN_11801 = 6'h24 == _T_4025 ? _T_3372_36_is_store : _GEN_11711;
  assign _GEN_11803 = 6'h24 == _T_4025 ? _T_3372_36_is_load : _GEN_11713;
  assign _GEN_11804 = 6'h24 == _T_4025 ? _T_3372_36_is_sys_pc2epc : _GEN_11714;
  assign _GEN_11806 = 6'h24 == _T_4025 ? _T_3372_36_flush_on_commit : _GEN_11716;
  assign _GEN_11807 = 6'h24 == _T_4025 ? _T_3372_36_ldst : _GEN_11717;
  assign _GEN_11812 = 6'h24 == _T_4025 ? _T_3372_36_dst_rtype : _GEN_11722;
  assign _GEN_11816 = 6'h24 == _T_4025 ? _T_3372_36_fp_val : _GEN_11726;
  assign _GEN_11876 = 6'h25 == _T_4025 ? _T_3372_37_pdst : _GEN_11786;
  assign _GEN_11883 = 6'h25 == _T_4025 ? _T_3372_37_stale_pdst : _GEN_11793;
  assign _GEN_11890 = 6'h25 == _T_4025 ? _T_3372_37_is_fencei : _GEN_11800;
  assign _GEN_11891 = 6'h25 == _T_4025 ? _T_3372_37_is_store : _GEN_11801;
  assign _GEN_11893 = 6'h25 == _T_4025 ? _T_3372_37_is_load : _GEN_11803;
  assign _GEN_11894 = 6'h25 == _T_4025 ? _T_3372_37_is_sys_pc2epc : _GEN_11804;
  assign _GEN_11896 = 6'h25 == _T_4025 ? _T_3372_37_flush_on_commit : _GEN_11806;
  assign _GEN_11897 = 6'h25 == _T_4025 ? _T_3372_37_ldst : _GEN_11807;
  assign _GEN_11902 = 6'h25 == _T_4025 ? _T_3372_37_dst_rtype : _GEN_11812;
  assign _GEN_11906 = 6'h25 == _T_4025 ? _T_3372_37_fp_val : _GEN_11816;
  assign _GEN_11966 = 6'h26 == _T_4025 ? _T_3372_38_pdst : _GEN_11876;
  assign _GEN_11973 = 6'h26 == _T_4025 ? _T_3372_38_stale_pdst : _GEN_11883;
  assign _GEN_11980 = 6'h26 == _T_4025 ? _T_3372_38_is_fencei : _GEN_11890;
  assign _GEN_11981 = 6'h26 == _T_4025 ? _T_3372_38_is_store : _GEN_11891;
  assign _GEN_11983 = 6'h26 == _T_4025 ? _T_3372_38_is_load : _GEN_11893;
  assign _GEN_11984 = 6'h26 == _T_4025 ? _T_3372_38_is_sys_pc2epc : _GEN_11894;
  assign _GEN_11986 = 6'h26 == _T_4025 ? _T_3372_38_flush_on_commit : _GEN_11896;
  assign _GEN_11987 = 6'h26 == _T_4025 ? _T_3372_38_ldst : _GEN_11897;
  assign _GEN_11992 = 6'h26 == _T_4025 ? _T_3372_38_dst_rtype : _GEN_11902;
  assign _GEN_11996 = 6'h26 == _T_4025 ? _T_3372_38_fp_val : _GEN_11906;
  assign _GEN_12056 = 6'h27 == _T_4025 ? _T_3372_39_pdst : _GEN_11966;
  assign _GEN_12063 = 6'h27 == _T_4025 ? _T_3372_39_stale_pdst : _GEN_11973;
  assign _GEN_12070 = 6'h27 == _T_4025 ? _T_3372_39_is_fencei : _GEN_11980;
  assign _GEN_12071 = 6'h27 == _T_4025 ? _T_3372_39_is_store : _GEN_11981;
  assign _GEN_12073 = 6'h27 == _T_4025 ? _T_3372_39_is_load : _GEN_11983;
  assign _GEN_12074 = 6'h27 == _T_4025 ? _T_3372_39_is_sys_pc2epc : _GEN_11984;
  assign _GEN_12076 = 6'h27 == _T_4025 ? _T_3372_39_flush_on_commit : _GEN_11986;
  assign _GEN_12077 = 6'h27 == _T_4025 ? _T_3372_39_ldst : _GEN_11987;
  assign _GEN_12082 = 6'h27 == _T_4025 ? _T_3372_39_dst_rtype : _GEN_11992;
  assign _GEN_12086 = 6'h27 == _T_4025 ? _T_3372_39_fp_val : _GEN_11996;
  assign _GEN_12094 = 6'h1 == _T_4025 ? _T_3073_1 : _T_3073_0;
  assign _GEN_12095 = 6'h2 == _T_4025 ? _T_3073_2 : _GEN_12094;
  assign _GEN_12096 = 6'h3 == _T_4025 ? _T_3073_3 : _GEN_12095;
  assign _GEN_12097 = 6'h4 == _T_4025 ? _T_3073_4 : _GEN_12096;
  assign _GEN_12098 = 6'h5 == _T_4025 ? _T_3073_5 : _GEN_12097;
  assign _GEN_12099 = 6'h6 == _T_4025 ? _T_3073_6 : _GEN_12098;
  assign _GEN_12100 = 6'h7 == _T_4025 ? _T_3073_7 : _GEN_12099;
  assign _GEN_12101 = 6'h8 == _T_4025 ? _T_3073_8 : _GEN_12100;
  assign _GEN_12102 = 6'h9 == _T_4025 ? _T_3073_9 : _GEN_12101;
  assign _GEN_12103 = 6'ha == _T_4025 ? _T_3073_10 : _GEN_12102;
  assign _GEN_12104 = 6'hb == _T_4025 ? _T_3073_11 : _GEN_12103;
  assign _GEN_12105 = 6'hc == _T_4025 ? _T_3073_12 : _GEN_12104;
  assign _GEN_12106 = 6'hd == _T_4025 ? _T_3073_13 : _GEN_12105;
  assign _GEN_12107 = 6'he == _T_4025 ? _T_3073_14 : _GEN_12106;
  assign _GEN_12108 = 6'hf == _T_4025 ? _T_3073_15 : _GEN_12107;
  assign _GEN_12109 = 6'h10 == _T_4025 ? _T_3073_16 : _GEN_12108;
  assign _GEN_12110 = 6'h11 == _T_4025 ? _T_3073_17 : _GEN_12109;
  assign _GEN_12111 = 6'h12 == _T_4025 ? _T_3073_18 : _GEN_12110;
  assign _GEN_12112 = 6'h13 == _T_4025 ? _T_3073_19 : _GEN_12111;
  assign _GEN_12113 = 6'h14 == _T_4025 ? _T_3073_20 : _GEN_12112;
  assign _GEN_12114 = 6'h15 == _T_4025 ? _T_3073_21 : _GEN_12113;
  assign _GEN_12115 = 6'h16 == _T_4025 ? _T_3073_22 : _GEN_12114;
  assign _GEN_12116 = 6'h17 == _T_4025 ? _T_3073_23 : _GEN_12115;
  assign _GEN_12117 = 6'h18 == _T_4025 ? _T_3073_24 : _GEN_12116;
  assign _GEN_12118 = 6'h19 == _T_4025 ? _T_3073_25 : _GEN_12117;
  assign _GEN_12119 = 6'h1a == _T_4025 ? _T_3073_26 : _GEN_12118;
  assign _GEN_12120 = 6'h1b == _T_4025 ? _T_3073_27 : _GEN_12119;
  assign _GEN_12121 = 6'h1c == _T_4025 ? _T_3073_28 : _GEN_12120;
  assign _GEN_12122 = 6'h1d == _T_4025 ? _T_3073_29 : _GEN_12121;
  assign _GEN_12123 = 6'h1e == _T_4025 ? _T_3073_30 : _GEN_12122;
  assign _GEN_12124 = 6'h1f == _T_4025 ? _T_3073_31 : _GEN_12123;
  assign _GEN_12125 = 6'h20 == _T_4025 ? _T_3073_32 : _GEN_12124;
  assign _GEN_12126 = 6'h21 == _T_4025 ? _T_3073_33 : _GEN_12125;
  assign _GEN_12127 = 6'h22 == _T_4025 ? _T_3073_34 : _GEN_12126;
  assign _GEN_12128 = 6'h23 == _T_4025 ? _T_3073_35 : _GEN_12127;
  assign _GEN_12129 = 6'h24 == _T_4025 ? _T_3073_36 : _GEN_12128;
  assign _GEN_12130 = 6'h25 == _T_4025 ? _T_3073_37 : _GEN_12129;
  assign _GEN_12131 = 6'h26 == _T_4025 ? _T_3073_38 : _GEN_12130;
  assign _GEN_12132 = 6'h27 == _T_4025 ? _T_3073_39 : _GEN_12131;
  assign _T_4046 = _T_4026 & _GEN_195;
  assign _T_4059 = _GEN_196_dst_rtype == 2'h0;
  assign _T_4072 = _GEN_197_dst_rtype == 2'h1;
  assign _T_4073 = _T_4059 | _T_4072;
  assign _T_4074 = _T_4046 & _T_4073;
  assign _T_4077 = rob_state == 2'h2;
  assign _GEN_19153 = 6'h0 == _T_4025 ? 1'h0 : _GEN_4374;
  assign _GEN_19154 = 6'h1 == _T_4025 ? 1'h0 : _GEN_4375;
  assign _GEN_19155 = 6'h2 == _T_4025 ? 1'h0 : _GEN_4376;
  assign _GEN_19156 = 6'h3 == _T_4025 ? 1'h0 : _GEN_4377;
  assign _GEN_19157 = 6'h4 == _T_4025 ? 1'h0 : _GEN_4378;
  assign _GEN_19158 = 6'h5 == _T_4025 ? 1'h0 : _GEN_4379;
  assign _GEN_19159 = 6'h6 == _T_4025 ? 1'h0 : _GEN_4380;
  assign _GEN_19160 = 6'h7 == _T_4025 ? 1'h0 : _GEN_4381;
  assign _GEN_19161 = 6'h8 == _T_4025 ? 1'h0 : _GEN_4382;
  assign _GEN_19162 = 6'h9 == _T_4025 ? 1'h0 : _GEN_4383;
  assign _GEN_19163 = 6'ha == _T_4025 ? 1'h0 : _GEN_4384;
  assign _GEN_19164 = 6'hb == _T_4025 ? 1'h0 : _GEN_4385;
  assign _GEN_19165 = 6'hc == _T_4025 ? 1'h0 : _GEN_4386;
  assign _GEN_19166 = 6'hd == _T_4025 ? 1'h0 : _GEN_4387;
  assign _GEN_19167 = 6'he == _T_4025 ? 1'h0 : _GEN_4388;
  assign _GEN_19168 = 6'hf == _T_4025 ? 1'h0 : _GEN_4389;
  assign _GEN_19169 = 6'h10 == _T_4025 ? 1'h0 : _GEN_4390;
  assign _GEN_19170 = 6'h11 == _T_4025 ? 1'h0 : _GEN_4391;
  assign _GEN_19171 = 6'h12 == _T_4025 ? 1'h0 : _GEN_4392;
  assign _GEN_19172 = 6'h13 == _T_4025 ? 1'h0 : _GEN_4393;
  assign _GEN_19173 = 6'h14 == _T_4025 ? 1'h0 : _GEN_4394;
  assign _GEN_19174 = 6'h15 == _T_4025 ? 1'h0 : _GEN_4395;
  assign _GEN_19175 = 6'h16 == _T_4025 ? 1'h0 : _GEN_4396;
  assign _GEN_19176 = 6'h17 == _T_4025 ? 1'h0 : _GEN_4397;
  assign _GEN_19177 = 6'h18 == _T_4025 ? 1'h0 : _GEN_4398;
  assign _GEN_19178 = 6'h19 == _T_4025 ? 1'h0 : _GEN_4399;
  assign _GEN_19179 = 6'h1a == _T_4025 ? 1'h0 : _GEN_4400;
  assign _GEN_19180 = 6'h1b == _T_4025 ? 1'h0 : _GEN_4401;
  assign _GEN_19181 = 6'h1c == _T_4025 ? 1'h0 : _GEN_4402;
  assign _GEN_19182 = 6'h1d == _T_4025 ? 1'h0 : _GEN_4403;
  assign _GEN_19183 = 6'h1e == _T_4025 ? 1'h0 : _GEN_4404;
  assign _GEN_19184 = 6'h1f == _T_4025 ? 1'h0 : _GEN_4405;
  assign _GEN_19185 = 6'h20 == _T_4025 ? 1'h0 : _GEN_4406;
  assign _GEN_19186 = 6'h21 == _T_4025 ? 1'h0 : _GEN_4407;
  assign _GEN_19187 = 6'h22 == _T_4025 ? 1'h0 : _GEN_4408;
  assign _GEN_19188 = 6'h23 == _T_4025 ? 1'h0 : _GEN_4409;
  assign _GEN_19189 = 6'h24 == _T_4025 ? 1'h0 : _GEN_4410;
  assign _GEN_19190 = 6'h25 == _T_4025 ? 1'h0 : _GEN_4411;
  assign _GEN_19191 = 6'h26 == _T_4025 ? 1'h0 : _GEN_4412;
  assign _GEN_19192 = 6'h27 == _T_4025 ? 1'h0 : _GEN_4413;
  assign _GEN_19193 = _T_4026 ? _GEN_19153 : _GEN_4374;
  assign _GEN_19194 = _T_4026 ? _GEN_19154 : _GEN_4375;
  assign _GEN_19195 = _T_4026 ? _GEN_19155 : _GEN_4376;
  assign _GEN_19196 = _T_4026 ? _GEN_19156 : _GEN_4377;
  assign _GEN_19197 = _T_4026 ? _GEN_19157 : _GEN_4378;
  assign _GEN_19198 = _T_4026 ? _GEN_19158 : _GEN_4379;
  assign _GEN_19199 = _T_4026 ? _GEN_19159 : _GEN_4380;
  assign _GEN_19200 = _T_4026 ? _GEN_19160 : _GEN_4381;
  assign _GEN_19201 = _T_4026 ? _GEN_19161 : _GEN_4382;
  assign _GEN_19202 = _T_4026 ? _GEN_19162 : _GEN_4383;
  assign _GEN_19203 = _T_4026 ? _GEN_19163 : _GEN_4384;
  assign _GEN_19204 = _T_4026 ? _GEN_19164 : _GEN_4385;
  assign _GEN_19205 = _T_4026 ? _GEN_19165 : _GEN_4386;
  assign _GEN_19206 = _T_4026 ? _GEN_19166 : _GEN_4387;
  assign _GEN_19207 = _T_4026 ? _GEN_19167 : _GEN_4388;
  assign _GEN_19208 = _T_4026 ? _GEN_19168 : _GEN_4389;
  assign _GEN_19209 = _T_4026 ? _GEN_19169 : _GEN_4390;
  assign _GEN_19210 = _T_4026 ? _GEN_19170 : _GEN_4391;
  assign _GEN_19211 = _T_4026 ? _GEN_19171 : _GEN_4392;
  assign _GEN_19212 = _T_4026 ? _GEN_19172 : _GEN_4393;
  assign _GEN_19213 = _T_4026 ? _GEN_19173 : _GEN_4394;
  assign _GEN_19214 = _T_4026 ? _GEN_19174 : _GEN_4395;
  assign _GEN_19215 = _T_4026 ? _GEN_19175 : _GEN_4396;
  assign _GEN_19216 = _T_4026 ? _GEN_19176 : _GEN_4397;
  assign _GEN_19217 = _T_4026 ? _GEN_19177 : _GEN_4398;
  assign _GEN_19218 = _T_4026 ? _GEN_19178 : _GEN_4399;
  assign _GEN_19219 = _T_4026 ? _GEN_19179 : _GEN_4400;
  assign _GEN_19220 = _T_4026 ? _GEN_19180 : _GEN_4401;
  assign _GEN_19221 = _T_4026 ? _GEN_19181 : _GEN_4402;
  assign _GEN_19222 = _T_4026 ? _GEN_19182 : _GEN_4403;
  assign _GEN_19223 = _T_4026 ? _GEN_19183 : _GEN_4404;
  assign _GEN_19224 = _T_4026 ? _GEN_19184 : _GEN_4405;
  assign _GEN_19225 = _T_4026 ? _GEN_19185 : _GEN_4406;
  assign _GEN_19226 = _T_4026 ? _GEN_19186 : _GEN_4407;
  assign _GEN_19227 = _T_4026 ? _GEN_19187 : _GEN_4408;
  assign _GEN_19228 = _T_4026 ? _GEN_19188 : _GEN_4409;
  assign _GEN_19229 = _T_4026 ? _GEN_19189 : _GEN_4410;
  assign _GEN_19230 = _T_4026 ? _GEN_19190 : _GEN_4411;
  assign _GEN_19231 = _T_4026 ? _GEN_19191 : _GEN_4412;
  assign _GEN_19232 = _T_4026 ? _GEN_19192 : _GEN_4413;
  assign _T_4090 = io_brinfo_mask & _T_3372_0_br_mask;
  assign _T_4092 = _T_4090 != 8'h0;
  assign _T_4093 = _T_3073_0 & _T_4092;
  assign _T_4094 = io_brinfo_valid & io_brinfo_mispredict;
  assign _T_4095 = _T_4094 & _T_4093;
  assign _T_4108 = io_brinfo_mispredict == 1'h0;
  assign _T_4109 = io_brinfo_valid & _T_4108;
  assign _T_4110 = _T_4109 & _T_4093;
  assign _T_4111 = ~ io_brinfo_mask;
  assign _T_4112 = _T_3372_0_br_mask & _T_4111;
  assign _GEN_19237 = _T_4110 ? _T_4112 : _GEN_5378;
  assign _GEN_19238 = _T_4095 ? 1'h0 : _GEN_19193;
  assign _GEN_19240 = _T_4095 ? _GEN_5378 : _GEN_19237;
  assign _T_4113 = io_brinfo_mask & _T_3372_1_br_mask;
  assign _T_4115 = _T_4113 != 8'h0;
  assign _T_4116 = _T_3073_1 & _T_4115;
  assign _T_4118 = _T_4094 & _T_4116;
  assign _T_4133 = _T_4109 & _T_4116;
  assign _T_4135 = _T_3372_1_br_mask & _T_4111;
  assign _GEN_19241 = _T_4133 ? _T_4135 : _GEN_5379;
  assign _GEN_19242 = _T_4118 ? 1'h0 : _GEN_19194;
  assign _GEN_19244 = _T_4118 ? _GEN_5379 : _GEN_19241;
  assign _T_4136 = io_brinfo_mask & _T_3372_2_br_mask;
  assign _T_4138 = _T_4136 != 8'h0;
  assign _T_4139 = _T_3073_2 & _T_4138;
  assign _T_4141 = _T_4094 & _T_4139;
  assign _T_4156 = _T_4109 & _T_4139;
  assign _T_4158 = _T_3372_2_br_mask & _T_4111;
  assign _GEN_19245 = _T_4156 ? _T_4158 : _GEN_5380;
  assign _GEN_19246 = _T_4141 ? 1'h0 : _GEN_19195;
  assign _GEN_19248 = _T_4141 ? _GEN_5380 : _GEN_19245;
  assign _T_4159 = io_brinfo_mask & _T_3372_3_br_mask;
  assign _T_4161 = _T_4159 != 8'h0;
  assign _T_4162 = _T_3073_3 & _T_4161;
  assign _T_4164 = _T_4094 & _T_4162;
  assign _T_4179 = _T_4109 & _T_4162;
  assign _T_4181 = _T_3372_3_br_mask & _T_4111;
  assign _GEN_19249 = _T_4179 ? _T_4181 : _GEN_5381;
  assign _GEN_19250 = _T_4164 ? 1'h0 : _GEN_19196;
  assign _GEN_19252 = _T_4164 ? _GEN_5381 : _GEN_19249;
  assign _T_4182 = io_brinfo_mask & _T_3372_4_br_mask;
  assign _T_4184 = _T_4182 != 8'h0;
  assign _T_4185 = _T_3073_4 & _T_4184;
  assign _T_4187 = _T_4094 & _T_4185;
  assign _T_4202 = _T_4109 & _T_4185;
  assign _T_4204 = _T_3372_4_br_mask & _T_4111;
  assign _GEN_19253 = _T_4202 ? _T_4204 : _GEN_5382;
  assign _GEN_19254 = _T_4187 ? 1'h0 : _GEN_19197;
  assign _GEN_19256 = _T_4187 ? _GEN_5382 : _GEN_19253;
  assign _T_4205 = io_brinfo_mask & _T_3372_5_br_mask;
  assign _T_4207 = _T_4205 != 8'h0;
  assign _T_4208 = _T_3073_5 & _T_4207;
  assign _T_4210 = _T_4094 & _T_4208;
  assign _T_4225 = _T_4109 & _T_4208;
  assign _T_4227 = _T_3372_5_br_mask & _T_4111;
  assign _GEN_19257 = _T_4225 ? _T_4227 : _GEN_5383;
  assign _GEN_19258 = _T_4210 ? 1'h0 : _GEN_19198;
  assign _GEN_19260 = _T_4210 ? _GEN_5383 : _GEN_19257;
  assign _T_4228 = io_brinfo_mask & _T_3372_6_br_mask;
  assign _T_4230 = _T_4228 != 8'h0;
  assign _T_4231 = _T_3073_6 & _T_4230;
  assign _T_4233 = _T_4094 & _T_4231;
  assign _T_4248 = _T_4109 & _T_4231;
  assign _T_4250 = _T_3372_6_br_mask & _T_4111;
  assign _GEN_19261 = _T_4248 ? _T_4250 : _GEN_5384;
  assign _GEN_19262 = _T_4233 ? 1'h0 : _GEN_19199;
  assign _GEN_19264 = _T_4233 ? _GEN_5384 : _GEN_19261;
  assign _T_4251 = io_brinfo_mask & _T_3372_7_br_mask;
  assign _T_4253 = _T_4251 != 8'h0;
  assign _T_4254 = _T_3073_7 & _T_4253;
  assign _T_4256 = _T_4094 & _T_4254;
  assign _T_4271 = _T_4109 & _T_4254;
  assign _T_4273 = _T_3372_7_br_mask & _T_4111;
  assign _GEN_19265 = _T_4271 ? _T_4273 : _GEN_5385;
  assign _GEN_19266 = _T_4256 ? 1'h0 : _GEN_19200;
  assign _GEN_19268 = _T_4256 ? _GEN_5385 : _GEN_19265;
  assign _T_4274 = io_brinfo_mask & _T_3372_8_br_mask;
  assign _T_4276 = _T_4274 != 8'h0;
  assign _T_4277 = _T_3073_8 & _T_4276;
  assign _T_4279 = _T_4094 & _T_4277;
  assign _T_4294 = _T_4109 & _T_4277;
  assign _T_4296 = _T_3372_8_br_mask & _T_4111;
  assign _GEN_19269 = _T_4294 ? _T_4296 : _GEN_5386;
  assign _GEN_19270 = _T_4279 ? 1'h0 : _GEN_19201;
  assign _GEN_19272 = _T_4279 ? _GEN_5386 : _GEN_19269;
  assign _T_4297 = io_brinfo_mask & _T_3372_9_br_mask;
  assign _T_4299 = _T_4297 != 8'h0;
  assign _T_4300 = _T_3073_9 & _T_4299;
  assign _T_4302 = _T_4094 & _T_4300;
  assign _T_4317 = _T_4109 & _T_4300;
  assign _T_4319 = _T_3372_9_br_mask & _T_4111;
  assign _GEN_19273 = _T_4317 ? _T_4319 : _GEN_5387;
  assign _GEN_19274 = _T_4302 ? 1'h0 : _GEN_19202;
  assign _GEN_19276 = _T_4302 ? _GEN_5387 : _GEN_19273;
  assign _T_4320 = io_brinfo_mask & _T_3372_10_br_mask;
  assign _T_4322 = _T_4320 != 8'h0;
  assign _T_4323 = _T_3073_10 & _T_4322;
  assign _T_4325 = _T_4094 & _T_4323;
  assign _T_4340 = _T_4109 & _T_4323;
  assign _T_4342 = _T_3372_10_br_mask & _T_4111;
  assign _GEN_19277 = _T_4340 ? _T_4342 : _GEN_5388;
  assign _GEN_19278 = _T_4325 ? 1'h0 : _GEN_19203;
  assign _GEN_19280 = _T_4325 ? _GEN_5388 : _GEN_19277;
  assign _T_4343 = io_brinfo_mask & _T_3372_11_br_mask;
  assign _T_4345 = _T_4343 != 8'h0;
  assign _T_4346 = _T_3073_11 & _T_4345;
  assign _T_4348 = _T_4094 & _T_4346;
  assign _T_4363 = _T_4109 & _T_4346;
  assign _T_4365 = _T_3372_11_br_mask & _T_4111;
  assign _GEN_19281 = _T_4363 ? _T_4365 : _GEN_5389;
  assign _GEN_19282 = _T_4348 ? 1'h0 : _GEN_19204;
  assign _GEN_19284 = _T_4348 ? _GEN_5389 : _GEN_19281;
  assign _T_4366 = io_brinfo_mask & _T_3372_12_br_mask;
  assign _T_4368 = _T_4366 != 8'h0;
  assign _T_4369 = _T_3073_12 & _T_4368;
  assign _T_4371 = _T_4094 & _T_4369;
  assign _T_4386 = _T_4109 & _T_4369;
  assign _T_4388 = _T_3372_12_br_mask & _T_4111;
  assign _GEN_19285 = _T_4386 ? _T_4388 : _GEN_5390;
  assign _GEN_19286 = _T_4371 ? 1'h0 : _GEN_19205;
  assign _GEN_19288 = _T_4371 ? _GEN_5390 : _GEN_19285;
  assign _T_4389 = io_brinfo_mask & _T_3372_13_br_mask;
  assign _T_4391 = _T_4389 != 8'h0;
  assign _T_4392 = _T_3073_13 & _T_4391;
  assign _T_4394 = _T_4094 & _T_4392;
  assign _T_4409 = _T_4109 & _T_4392;
  assign _T_4411 = _T_3372_13_br_mask & _T_4111;
  assign _GEN_19289 = _T_4409 ? _T_4411 : _GEN_5391;
  assign _GEN_19290 = _T_4394 ? 1'h0 : _GEN_19206;
  assign _GEN_19292 = _T_4394 ? _GEN_5391 : _GEN_19289;
  assign _T_4412 = io_brinfo_mask & _T_3372_14_br_mask;
  assign _T_4414 = _T_4412 != 8'h0;
  assign _T_4415 = _T_3073_14 & _T_4414;
  assign _T_4417 = _T_4094 & _T_4415;
  assign _T_4432 = _T_4109 & _T_4415;
  assign _T_4434 = _T_3372_14_br_mask & _T_4111;
  assign _GEN_19293 = _T_4432 ? _T_4434 : _GEN_5392;
  assign _GEN_19294 = _T_4417 ? 1'h0 : _GEN_19207;
  assign _GEN_19296 = _T_4417 ? _GEN_5392 : _GEN_19293;
  assign _T_4435 = io_brinfo_mask & _T_3372_15_br_mask;
  assign _T_4437 = _T_4435 != 8'h0;
  assign _T_4438 = _T_3073_15 & _T_4437;
  assign _T_4440 = _T_4094 & _T_4438;
  assign _T_4455 = _T_4109 & _T_4438;
  assign _T_4457 = _T_3372_15_br_mask & _T_4111;
  assign _GEN_19297 = _T_4455 ? _T_4457 : _GEN_5393;
  assign _GEN_19298 = _T_4440 ? 1'h0 : _GEN_19208;
  assign _GEN_19300 = _T_4440 ? _GEN_5393 : _GEN_19297;
  assign _T_4458 = io_brinfo_mask & _T_3372_16_br_mask;
  assign _T_4460 = _T_4458 != 8'h0;
  assign _T_4461 = _T_3073_16 & _T_4460;
  assign _T_4463 = _T_4094 & _T_4461;
  assign _T_4478 = _T_4109 & _T_4461;
  assign _T_4480 = _T_3372_16_br_mask & _T_4111;
  assign _GEN_19301 = _T_4478 ? _T_4480 : _GEN_5394;
  assign _GEN_19302 = _T_4463 ? 1'h0 : _GEN_19209;
  assign _GEN_19304 = _T_4463 ? _GEN_5394 : _GEN_19301;
  assign _T_4481 = io_brinfo_mask & _T_3372_17_br_mask;
  assign _T_4483 = _T_4481 != 8'h0;
  assign _T_4484 = _T_3073_17 & _T_4483;
  assign _T_4486 = _T_4094 & _T_4484;
  assign _T_4501 = _T_4109 & _T_4484;
  assign _T_4503 = _T_3372_17_br_mask & _T_4111;
  assign _GEN_19305 = _T_4501 ? _T_4503 : _GEN_5395;
  assign _GEN_19306 = _T_4486 ? 1'h0 : _GEN_19210;
  assign _GEN_19308 = _T_4486 ? _GEN_5395 : _GEN_19305;
  assign _T_4504 = io_brinfo_mask & _T_3372_18_br_mask;
  assign _T_4506 = _T_4504 != 8'h0;
  assign _T_4507 = _T_3073_18 & _T_4506;
  assign _T_4509 = _T_4094 & _T_4507;
  assign _T_4524 = _T_4109 & _T_4507;
  assign _T_4526 = _T_3372_18_br_mask & _T_4111;
  assign _GEN_19309 = _T_4524 ? _T_4526 : _GEN_5396;
  assign _GEN_19310 = _T_4509 ? 1'h0 : _GEN_19211;
  assign _GEN_19312 = _T_4509 ? _GEN_5396 : _GEN_19309;
  assign _T_4527 = io_brinfo_mask & _T_3372_19_br_mask;
  assign _T_4529 = _T_4527 != 8'h0;
  assign _T_4530 = _T_3073_19 & _T_4529;
  assign _T_4532 = _T_4094 & _T_4530;
  assign _T_4547 = _T_4109 & _T_4530;
  assign _T_4549 = _T_3372_19_br_mask & _T_4111;
  assign _GEN_19313 = _T_4547 ? _T_4549 : _GEN_5397;
  assign _GEN_19314 = _T_4532 ? 1'h0 : _GEN_19212;
  assign _GEN_19316 = _T_4532 ? _GEN_5397 : _GEN_19313;
  assign _T_4550 = io_brinfo_mask & _T_3372_20_br_mask;
  assign _T_4552 = _T_4550 != 8'h0;
  assign _T_4553 = _T_3073_20 & _T_4552;
  assign _T_4555 = _T_4094 & _T_4553;
  assign _T_4570 = _T_4109 & _T_4553;
  assign _T_4572 = _T_3372_20_br_mask & _T_4111;
  assign _GEN_19317 = _T_4570 ? _T_4572 : _GEN_5398;
  assign _GEN_19318 = _T_4555 ? 1'h0 : _GEN_19213;
  assign _GEN_19320 = _T_4555 ? _GEN_5398 : _GEN_19317;
  assign _T_4573 = io_brinfo_mask & _T_3372_21_br_mask;
  assign _T_4575 = _T_4573 != 8'h0;
  assign _T_4576 = _T_3073_21 & _T_4575;
  assign _T_4578 = _T_4094 & _T_4576;
  assign _T_4593 = _T_4109 & _T_4576;
  assign _T_4595 = _T_3372_21_br_mask & _T_4111;
  assign _GEN_19321 = _T_4593 ? _T_4595 : _GEN_5399;
  assign _GEN_19322 = _T_4578 ? 1'h0 : _GEN_19214;
  assign _GEN_19324 = _T_4578 ? _GEN_5399 : _GEN_19321;
  assign _T_4596 = io_brinfo_mask & _T_3372_22_br_mask;
  assign _T_4598 = _T_4596 != 8'h0;
  assign _T_4599 = _T_3073_22 & _T_4598;
  assign _T_4601 = _T_4094 & _T_4599;
  assign _T_4616 = _T_4109 & _T_4599;
  assign _T_4618 = _T_3372_22_br_mask & _T_4111;
  assign _GEN_19325 = _T_4616 ? _T_4618 : _GEN_5400;
  assign _GEN_19326 = _T_4601 ? 1'h0 : _GEN_19215;
  assign _GEN_19328 = _T_4601 ? _GEN_5400 : _GEN_19325;
  assign _T_4619 = io_brinfo_mask & _T_3372_23_br_mask;
  assign _T_4621 = _T_4619 != 8'h0;
  assign _T_4622 = _T_3073_23 & _T_4621;
  assign _T_4624 = _T_4094 & _T_4622;
  assign _T_4639 = _T_4109 & _T_4622;
  assign _T_4641 = _T_3372_23_br_mask & _T_4111;
  assign _GEN_19329 = _T_4639 ? _T_4641 : _GEN_5401;
  assign _GEN_19330 = _T_4624 ? 1'h0 : _GEN_19216;
  assign _GEN_19332 = _T_4624 ? _GEN_5401 : _GEN_19329;
  assign _T_4642 = io_brinfo_mask & _T_3372_24_br_mask;
  assign _T_4644 = _T_4642 != 8'h0;
  assign _T_4645 = _T_3073_24 & _T_4644;
  assign _T_4647 = _T_4094 & _T_4645;
  assign _T_4662 = _T_4109 & _T_4645;
  assign _T_4664 = _T_3372_24_br_mask & _T_4111;
  assign _GEN_19333 = _T_4662 ? _T_4664 : _GEN_5402;
  assign _GEN_19334 = _T_4647 ? 1'h0 : _GEN_19217;
  assign _GEN_19336 = _T_4647 ? _GEN_5402 : _GEN_19333;
  assign _T_4665 = io_brinfo_mask & _T_3372_25_br_mask;
  assign _T_4667 = _T_4665 != 8'h0;
  assign _T_4668 = _T_3073_25 & _T_4667;
  assign _T_4670 = _T_4094 & _T_4668;
  assign _T_4685 = _T_4109 & _T_4668;
  assign _T_4687 = _T_3372_25_br_mask & _T_4111;
  assign _GEN_19337 = _T_4685 ? _T_4687 : _GEN_5403;
  assign _GEN_19338 = _T_4670 ? 1'h0 : _GEN_19218;
  assign _GEN_19340 = _T_4670 ? _GEN_5403 : _GEN_19337;
  assign _T_4688 = io_brinfo_mask & _T_3372_26_br_mask;
  assign _T_4690 = _T_4688 != 8'h0;
  assign _T_4691 = _T_3073_26 & _T_4690;
  assign _T_4693 = _T_4094 & _T_4691;
  assign _T_4708 = _T_4109 & _T_4691;
  assign _T_4710 = _T_3372_26_br_mask & _T_4111;
  assign _GEN_19341 = _T_4708 ? _T_4710 : _GEN_5404;
  assign _GEN_19342 = _T_4693 ? 1'h0 : _GEN_19219;
  assign _GEN_19344 = _T_4693 ? _GEN_5404 : _GEN_19341;
  assign _T_4711 = io_brinfo_mask & _T_3372_27_br_mask;
  assign _T_4713 = _T_4711 != 8'h0;
  assign _T_4714 = _T_3073_27 & _T_4713;
  assign _T_4716 = _T_4094 & _T_4714;
  assign _T_4731 = _T_4109 & _T_4714;
  assign _T_4733 = _T_3372_27_br_mask & _T_4111;
  assign _GEN_19345 = _T_4731 ? _T_4733 : _GEN_5405;
  assign _GEN_19346 = _T_4716 ? 1'h0 : _GEN_19220;
  assign _GEN_19348 = _T_4716 ? _GEN_5405 : _GEN_19345;
  assign _T_4734 = io_brinfo_mask & _T_3372_28_br_mask;
  assign _T_4736 = _T_4734 != 8'h0;
  assign _T_4737 = _T_3073_28 & _T_4736;
  assign _T_4739 = _T_4094 & _T_4737;
  assign _T_4754 = _T_4109 & _T_4737;
  assign _T_4756 = _T_3372_28_br_mask & _T_4111;
  assign _GEN_19349 = _T_4754 ? _T_4756 : _GEN_5406;
  assign _GEN_19350 = _T_4739 ? 1'h0 : _GEN_19221;
  assign _GEN_19352 = _T_4739 ? _GEN_5406 : _GEN_19349;
  assign _T_4757 = io_brinfo_mask & _T_3372_29_br_mask;
  assign _T_4759 = _T_4757 != 8'h0;
  assign _T_4760 = _T_3073_29 & _T_4759;
  assign _T_4762 = _T_4094 & _T_4760;
  assign _T_4777 = _T_4109 & _T_4760;
  assign _T_4779 = _T_3372_29_br_mask & _T_4111;
  assign _GEN_19353 = _T_4777 ? _T_4779 : _GEN_5407;
  assign _GEN_19354 = _T_4762 ? 1'h0 : _GEN_19222;
  assign _GEN_19356 = _T_4762 ? _GEN_5407 : _GEN_19353;
  assign _T_4780 = io_brinfo_mask & _T_3372_30_br_mask;
  assign _T_4782 = _T_4780 != 8'h0;
  assign _T_4783 = _T_3073_30 & _T_4782;
  assign _T_4785 = _T_4094 & _T_4783;
  assign _T_4800 = _T_4109 & _T_4783;
  assign _T_4802 = _T_3372_30_br_mask & _T_4111;
  assign _GEN_19357 = _T_4800 ? _T_4802 : _GEN_5408;
  assign _GEN_19358 = _T_4785 ? 1'h0 : _GEN_19223;
  assign _GEN_19360 = _T_4785 ? _GEN_5408 : _GEN_19357;
  assign _T_4803 = io_brinfo_mask & _T_3372_31_br_mask;
  assign _T_4805 = _T_4803 != 8'h0;
  assign _T_4806 = _T_3073_31 & _T_4805;
  assign _T_4808 = _T_4094 & _T_4806;
  assign _T_4823 = _T_4109 & _T_4806;
  assign _T_4825 = _T_3372_31_br_mask & _T_4111;
  assign _GEN_19361 = _T_4823 ? _T_4825 : _GEN_5409;
  assign _GEN_19362 = _T_4808 ? 1'h0 : _GEN_19224;
  assign _GEN_19364 = _T_4808 ? _GEN_5409 : _GEN_19361;
  assign _T_4826 = io_brinfo_mask & _T_3372_32_br_mask;
  assign _T_4828 = _T_4826 != 8'h0;
  assign _T_4829 = _T_3073_32 & _T_4828;
  assign _T_4831 = _T_4094 & _T_4829;
  assign _T_4846 = _T_4109 & _T_4829;
  assign _T_4848 = _T_3372_32_br_mask & _T_4111;
  assign _GEN_19365 = _T_4846 ? _T_4848 : _GEN_5410;
  assign _GEN_19366 = _T_4831 ? 1'h0 : _GEN_19225;
  assign _GEN_19368 = _T_4831 ? _GEN_5410 : _GEN_19365;
  assign _T_4849 = io_brinfo_mask & _T_3372_33_br_mask;
  assign _T_4851 = _T_4849 != 8'h0;
  assign _T_4852 = _T_3073_33 & _T_4851;
  assign _T_4854 = _T_4094 & _T_4852;
  assign _T_4869 = _T_4109 & _T_4852;
  assign _T_4871 = _T_3372_33_br_mask & _T_4111;
  assign _GEN_19369 = _T_4869 ? _T_4871 : _GEN_5411;
  assign _GEN_19370 = _T_4854 ? 1'h0 : _GEN_19226;
  assign _GEN_19372 = _T_4854 ? _GEN_5411 : _GEN_19369;
  assign _T_4872 = io_brinfo_mask & _T_3372_34_br_mask;
  assign _T_4874 = _T_4872 != 8'h0;
  assign _T_4875 = _T_3073_34 & _T_4874;
  assign _T_4877 = _T_4094 & _T_4875;
  assign _T_4892 = _T_4109 & _T_4875;
  assign _T_4894 = _T_3372_34_br_mask & _T_4111;
  assign _GEN_19373 = _T_4892 ? _T_4894 : _GEN_5412;
  assign _GEN_19374 = _T_4877 ? 1'h0 : _GEN_19227;
  assign _GEN_19376 = _T_4877 ? _GEN_5412 : _GEN_19373;
  assign _T_4895 = io_brinfo_mask & _T_3372_35_br_mask;
  assign _T_4897 = _T_4895 != 8'h0;
  assign _T_4898 = _T_3073_35 & _T_4897;
  assign _T_4900 = _T_4094 & _T_4898;
  assign _T_4915 = _T_4109 & _T_4898;
  assign _T_4917 = _T_3372_35_br_mask & _T_4111;
  assign _GEN_19377 = _T_4915 ? _T_4917 : _GEN_5413;
  assign _GEN_19378 = _T_4900 ? 1'h0 : _GEN_19228;
  assign _GEN_19380 = _T_4900 ? _GEN_5413 : _GEN_19377;
  assign _T_4918 = io_brinfo_mask & _T_3372_36_br_mask;
  assign _T_4920 = _T_4918 != 8'h0;
  assign _T_4921 = _T_3073_36 & _T_4920;
  assign _T_4923 = _T_4094 & _T_4921;
  assign _T_4938 = _T_4109 & _T_4921;
  assign _T_4940 = _T_3372_36_br_mask & _T_4111;
  assign _GEN_19381 = _T_4938 ? _T_4940 : _GEN_5414;
  assign _GEN_19382 = _T_4923 ? 1'h0 : _GEN_19229;
  assign _GEN_19384 = _T_4923 ? _GEN_5414 : _GEN_19381;
  assign _T_4941 = io_brinfo_mask & _T_3372_37_br_mask;
  assign _T_4943 = _T_4941 != 8'h0;
  assign _T_4944 = _T_3073_37 & _T_4943;
  assign _T_4946 = _T_4094 & _T_4944;
  assign _T_4961 = _T_4109 & _T_4944;
  assign _T_4963 = _T_3372_37_br_mask & _T_4111;
  assign _GEN_19385 = _T_4961 ? _T_4963 : _GEN_5415;
  assign _GEN_19386 = _T_4946 ? 1'h0 : _GEN_19230;
  assign _GEN_19388 = _T_4946 ? _GEN_5415 : _GEN_19385;
  assign _T_4964 = io_brinfo_mask & _T_3372_38_br_mask;
  assign _T_4966 = _T_4964 != 8'h0;
  assign _T_4967 = _T_3073_38 & _T_4966;
  assign _T_4969 = _T_4094 & _T_4967;
  assign _T_4984 = _T_4109 & _T_4967;
  assign _T_4986 = _T_3372_38_br_mask & _T_4111;
  assign _GEN_19389 = _T_4984 ? _T_4986 : _GEN_5416;
  assign _GEN_19390 = _T_4969 ? 1'h0 : _GEN_19231;
  assign _GEN_19392 = _T_4969 ? _GEN_5416 : _GEN_19389;
  assign _T_4987 = io_brinfo_mask & _T_3372_39_br_mask;
  assign _T_4989 = _T_4987 != 8'h0;
  assign _T_4990 = _T_3073_39 & _T_4989;
  assign _T_4992 = _T_4094 & _T_4990;
  assign _T_5007 = _T_4109 & _T_4990;
  assign _T_5009 = _T_3372_39_br_mask & _T_4111;
  assign _GEN_19393 = _T_5007 ? _T_5009 : _GEN_5417;
  assign _GEN_19394 = _T_4992 ? 1'h0 : _GEN_19232;
  assign _GEN_19396 = _T_4992 ? _GEN_5417 : _GEN_19393;
  assign _GEN_19397 = 6'h0 == rob_head ? 1'h0 : _GEN_19238;
  assign _GEN_19398 = 6'h1 == rob_head ? 1'h0 : _GEN_19242;
  assign _GEN_19399 = 6'h2 == rob_head ? 1'h0 : _GEN_19246;
  assign _GEN_19400 = 6'h3 == rob_head ? 1'h0 : _GEN_19250;
  assign _GEN_19401 = 6'h4 == rob_head ? 1'h0 : _GEN_19254;
  assign _GEN_19402 = 6'h5 == rob_head ? 1'h0 : _GEN_19258;
  assign _GEN_19403 = 6'h6 == rob_head ? 1'h0 : _GEN_19262;
  assign _GEN_19404 = 6'h7 == rob_head ? 1'h0 : _GEN_19266;
  assign _GEN_19405 = 6'h8 == rob_head ? 1'h0 : _GEN_19270;
  assign _GEN_19406 = 6'h9 == rob_head ? 1'h0 : _GEN_19274;
  assign _GEN_19407 = 6'ha == rob_head ? 1'h0 : _GEN_19278;
  assign _GEN_19408 = 6'hb == rob_head ? 1'h0 : _GEN_19282;
  assign _GEN_19409 = 6'hc == rob_head ? 1'h0 : _GEN_19286;
  assign _GEN_19410 = 6'hd == rob_head ? 1'h0 : _GEN_19290;
  assign _GEN_19411 = 6'he == rob_head ? 1'h0 : _GEN_19294;
  assign _GEN_19412 = 6'hf == rob_head ? 1'h0 : _GEN_19298;
  assign _GEN_19413 = 6'h10 == rob_head ? 1'h0 : _GEN_19302;
  assign _GEN_19414 = 6'h11 == rob_head ? 1'h0 : _GEN_19306;
  assign _GEN_19415 = 6'h12 == rob_head ? 1'h0 : _GEN_19310;
  assign _GEN_19416 = 6'h13 == rob_head ? 1'h0 : _GEN_19314;
  assign _GEN_19417 = 6'h14 == rob_head ? 1'h0 : _GEN_19318;
  assign _GEN_19418 = 6'h15 == rob_head ? 1'h0 : _GEN_19322;
  assign _GEN_19419 = 6'h16 == rob_head ? 1'h0 : _GEN_19326;
  assign _GEN_19420 = 6'h17 == rob_head ? 1'h0 : _GEN_19330;
  assign _GEN_19421 = 6'h18 == rob_head ? 1'h0 : _GEN_19334;
  assign _GEN_19422 = 6'h19 == rob_head ? 1'h0 : _GEN_19338;
  assign _GEN_19423 = 6'h1a == rob_head ? 1'h0 : _GEN_19342;
  assign _GEN_19424 = 6'h1b == rob_head ? 1'h0 : _GEN_19346;
  assign _GEN_19425 = 6'h1c == rob_head ? 1'h0 : _GEN_19350;
  assign _GEN_19426 = 6'h1d == rob_head ? 1'h0 : _GEN_19354;
  assign _GEN_19427 = 6'h1e == rob_head ? 1'h0 : _GEN_19358;
  assign _GEN_19428 = 6'h1f == rob_head ? 1'h0 : _GEN_19362;
  assign _GEN_19429 = 6'h20 == rob_head ? 1'h0 : _GEN_19366;
  assign _GEN_19430 = 6'h21 == rob_head ? 1'h0 : _GEN_19370;
  assign _GEN_19431 = 6'h22 == rob_head ? 1'h0 : _GEN_19374;
  assign _GEN_19432 = 6'h23 == rob_head ? 1'h0 : _GEN_19378;
  assign _GEN_19433 = 6'h24 == rob_head ? 1'h0 : _GEN_19382;
  assign _GEN_19434 = 6'h25 == rob_head ? 1'h0 : _GEN_19386;
  assign _GEN_19435 = 6'h26 == rob_head ? 1'h0 : _GEN_19390;
  assign _GEN_19436 = 6'h27 == rob_head ? 1'h0 : _GEN_19394;
  assign _GEN_19437 = will_commit_0 ? _GEN_19397 : _GEN_19238;
  assign _GEN_19438 = will_commit_0 ? _GEN_19398 : _GEN_19242;
  assign _GEN_19439 = will_commit_0 ? _GEN_19399 : _GEN_19246;
  assign _GEN_19440 = will_commit_0 ? _GEN_19400 : _GEN_19250;
  assign _GEN_19441 = will_commit_0 ? _GEN_19401 : _GEN_19254;
  assign _GEN_19442 = will_commit_0 ? _GEN_19402 : _GEN_19258;
  assign _GEN_19443 = will_commit_0 ? _GEN_19403 : _GEN_19262;
  assign _GEN_19444 = will_commit_0 ? _GEN_19404 : _GEN_19266;
  assign _GEN_19445 = will_commit_0 ? _GEN_19405 : _GEN_19270;
  assign _GEN_19446 = will_commit_0 ? _GEN_19406 : _GEN_19274;
  assign _GEN_19447 = will_commit_0 ? _GEN_19407 : _GEN_19278;
  assign _GEN_19448 = will_commit_0 ? _GEN_19408 : _GEN_19282;
  assign _GEN_19449 = will_commit_0 ? _GEN_19409 : _GEN_19286;
  assign _GEN_19450 = will_commit_0 ? _GEN_19410 : _GEN_19290;
  assign _GEN_19451 = will_commit_0 ? _GEN_19411 : _GEN_19294;
  assign _GEN_19452 = will_commit_0 ? _GEN_19412 : _GEN_19298;
  assign _GEN_19453 = will_commit_0 ? _GEN_19413 : _GEN_19302;
  assign _GEN_19454 = will_commit_0 ? _GEN_19414 : _GEN_19306;
  assign _GEN_19455 = will_commit_0 ? _GEN_19415 : _GEN_19310;
  assign _GEN_19456 = will_commit_0 ? _GEN_19416 : _GEN_19314;
  assign _GEN_19457 = will_commit_0 ? _GEN_19417 : _GEN_19318;
  assign _GEN_19458 = will_commit_0 ? _GEN_19418 : _GEN_19322;
  assign _GEN_19459 = will_commit_0 ? _GEN_19419 : _GEN_19326;
  assign _GEN_19460 = will_commit_0 ? _GEN_19420 : _GEN_19330;
  assign _GEN_19461 = will_commit_0 ? _GEN_19421 : _GEN_19334;
  assign _GEN_19462 = will_commit_0 ? _GEN_19422 : _GEN_19338;
  assign _GEN_19463 = will_commit_0 ? _GEN_19423 : _GEN_19342;
  assign _GEN_19464 = will_commit_0 ? _GEN_19424 : _GEN_19346;
  assign _GEN_19465 = will_commit_0 ? _GEN_19425 : _GEN_19350;
  assign _GEN_19466 = will_commit_0 ? _GEN_19426 : _GEN_19354;
  assign _GEN_19467 = will_commit_0 ? _GEN_19427 : _GEN_19358;
  assign _GEN_19468 = will_commit_0 ? _GEN_19428 : _GEN_19362;
  assign _GEN_19469 = will_commit_0 ? _GEN_19429 : _GEN_19366;
  assign _GEN_19470 = will_commit_0 ? _GEN_19430 : _GEN_19370;
  assign _GEN_19471 = will_commit_0 ? _GEN_19431 : _GEN_19374;
  assign _GEN_19472 = will_commit_0 ? _GEN_19432 : _GEN_19378;
  assign _GEN_19473 = will_commit_0 ? _GEN_19433 : _GEN_19382;
  assign _GEN_19474 = will_commit_0 ? _GEN_19434 : _GEN_19386;
  assign _GEN_19475 = will_commit_0 ? _GEN_19435 : _GEN_19390;
  assign _GEN_19476 = will_commit_0 ? _GEN_19436 : _GEN_19394;
  assign _GEN_19544 = 6'h1 == rob_head ? _T_3372_1_is_store : _T_3372_0_is_store;
  assign _GEN_19546 = 6'h1 == rob_head ? _T_3372_1_is_load : _T_3372_0_is_load;
  assign _GEN_19634 = 6'h2 == rob_head ? _T_3372_2_is_store : _GEN_19544;
  assign _GEN_19636 = 6'h2 == rob_head ? _T_3372_2_is_load : _GEN_19546;
  assign _GEN_19724 = 6'h3 == rob_head ? _T_3372_3_is_store : _GEN_19634;
  assign _GEN_19726 = 6'h3 == rob_head ? _T_3372_3_is_load : _GEN_19636;
  assign _GEN_19814 = 6'h4 == rob_head ? _T_3372_4_is_store : _GEN_19724;
  assign _GEN_19816 = 6'h4 == rob_head ? _T_3372_4_is_load : _GEN_19726;
  assign _GEN_19904 = 6'h5 == rob_head ? _T_3372_5_is_store : _GEN_19814;
  assign _GEN_19906 = 6'h5 == rob_head ? _T_3372_5_is_load : _GEN_19816;
  assign _GEN_19994 = 6'h6 == rob_head ? _T_3372_6_is_store : _GEN_19904;
  assign _GEN_19996 = 6'h6 == rob_head ? _T_3372_6_is_load : _GEN_19906;
  assign _GEN_20084 = 6'h7 == rob_head ? _T_3372_7_is_store : _GEN_19994;
  assign _GEN_20086 = 6'h7 == rob_head ? _T_3372_7_is_load : _GEN_19996;
  assign _GEN_20174 = 6'h8 == rob_head ? _T_3372_8_is_store : _GEN_20084;
  assign _GEN_20176 = 6'h8 == rob_head ? _T_3372_8_is_load : _GEN_20086;
  assign _GEN_20264 = 6'h9 == rob_head ? _T_3372_9_is_store : _GEN_20174;
  assign _GEN_20266 = 6'h9 == rob_head ? _T_3372_9_is_load : _GEN_20176;
  assign _GEN_20354 = 6'ha == rob_head ? _T_3372_10_is_store : _GEN_20264;
  assign _GEN_20356 = 6'ha == rob_head ? _T_3372_10_is_load : _GEN_20266;
  assign _GEN_20444 = 6'hb == rob_head ? _T_3372_11_is_store : _GEN_20354;
  assign _GEN_20446 = 6'hb == rob_head ? _T_3372_11_is_load : _GEN_20356;
  assign _GEN_20534 = 6'hc == rob_head ? _T_3372_12_is_store : _GEN_20444;
  assign _GEN_20536 = 6'hc == rob_head ? _T_3372_12_is_load : _GEN_20446;
  assign _GEN_20624 = 6'hd == rob_head ? _T_3372_13_is_store : _GEN_20534;
  assign _GEN_20626 = 6'hd == rob_head ? _T_3372_13_is_load : _GEN_20536;
  assign _GEN_20714 = 6'he == rob_head ? _T_3372_14_is_store : _GEN_20624;
  assign _GEN_20716 = 6'he == rob_head ? _T_3372_14_is_load : _GEN_20626;
  assign _GEN_20804 = 6'hf == rob_head ? _T_3372_15_is_store : _GEN_20714;
  assign _GEN_20806 = 6'hf == rob_head ? _T_3372_15_is_load : _GEN_20716;
  assign _GEN_20894 = 6'h10 == rob_head ? _T_3372_16_is_store : _GEN_20804;
  assign _GEN_20896 = 6'h10 == rob_head ? _T_3372_16_is_load : _GEN_20806;
  assign _GEN_20984 = 6'h11 == rob_head ? _T_3372_17_is_store : _GEN_20894;
  assign _GEN_20986 = 6'h11 == rob_head ? _T_3372_17_is_load : _GEN_20896;
  assign _GEN_21074 = 6'h12 == rob_head ? _T_3372_18_is_store : _GEN_20984;
  assign _GEN_21076 = 6'h12 == rob_head ? _T_3372_18_is_load : _GEN_20986;
  assign _GEN_21164 = 6'h13 == rob_head ? _T_3372_19_is_store : _GEN_21074;
  assign _GEN_21166 = 6'h13 == rob_head ? _T_3372_19_is_load : _GEN_21076;
  assign _GEN_21254 = 6'h14 == rob_head ? _T_3372_20_is_store : _GEN_21164;
  assign _GEN_21256 = 6'h14 == rob_head ? _T_3372_20_is_load : _GEN_21166;
  assign _GEN_21344 = 6'h15 == rob_head ? _T_3372_21_is_store : _GEN_21254;
  assign _GEN_21346 = 6'h15 == rob_head ? _T_3372_21_is_load : _GEN_21256;
  assign _GEN_21434 = 6'h16 == rob_head ? _T_3372_22_is_store : _GEN_21344;
  assign _GEN_21436 = 6'h16 == rob_head ? _T_3372_22_is_load : _GEN_21346;
  assign _GEN_21524 = 6'h17 == rob_head ? _T_3372_23_is_store : _GEN_21434;
  assign _GEN_21526 = 6'h17 == rob_head ? _T_3372_23_is_load : _GEN_21436;
  assign _GEN_21614 = 6'h18 == rob_head ? _T_3372_24_is_store : _GEN_21524;
  assign _GEN_21616 = 6'h18 == rob_head ? _T_3372_24_is_load : _GEN_21526;
  assign _GEN_21704 = 6'h19 == rob_head ? _T_3372_25_is_store : _GEN_21614;
  assign _GEN_21706 = 6'h19 == rob_head ? _T_3372_25_is_load : _GEN_21616;
  assign _GEN_21794 = 6'h1a == rob_head ? _T_3372_26_is_store : _GEN_21704;
  assign _GEN_21796 = 6'h1a == rob_head ? _T_3372_26_is_load : _GEN_21706;
  assign _GEN_21884 = 6'h1b == rob_head ? _T_3372_27_is_store : _GEN_21794;
  assign _GEN_21886 = 6'h1b == rob_head ? _T_3372_27_is_load : _GEN_21796;
  assign _GEN_21974 = 6'h1c == rob_head ? _T_3372_28_is_store : _GEN_21884;
  assign _GEN_21976 = 6'h1c == rob_head ? _T_3372_28_is_load : _GEN_21886;
  assign _GEN_22064 = 6'h1d == rob_head ? _T_3372_29_is_store : _GEN_21974;
  assign _GEN_22066 = 6'h1d == rob_head ? _T_3372_29_is_load : _GEN_21976;
  assign _GEN_22154 = 6'h1e == rob_head ? _T_3372_30_is_store : _GEN_22064;
  assign _GEN_22156 = 6'h1e == rob_head ? _T_3372_30_is_load : _GEN_22066;
  assign _GEN_22244 = 6'h1f == rob_head ? _T_3372_31_is_store : _GEN_22154;
  assign _GEN_22246 = 6'h1f == rob_head ? _T_3372_31_is_load : _GEN_22156;
  assign _GEN_22334 = 6'h20 == rob_head ? _T_3372_32_is_store : _GEN_22244;
  assign _GEN_22336 = 6'h20 == rob_head ? _T_3372_32_is_load : _GEN_22246;
  assign _GEN_22424 = 6'h21 == rob_head ? _T_3372_33_is_store : _GEN_22334;
  assign _GEN_22426 = 6'h21 == rob_head ? _T_3372_33_is_load : _GEN_22336;
  assign _GEN_22514 = 6'h22 == rob_head ? _T_3372_34_is_store : _GEN_22424;
  assign _GEN_22516 = 6'h22 == rob_head ? _T_3372_34_is_load : _GEN_22426;
  assign _GEN_22604 = 6'h23 == rob_head ? _T_3372_35_is_store : _GEN_22514;
  assign _GEN_22606 = 6'h23 == rob_head ? _T_3372_35_is_load : _GEN_22516;
  assign _GEN_22694 = 6'h24 == rob_head ? _T_3372_36_is_store : _GEN_22604;
  assign _GEN_22696 = 6'h24 == rob_head ? _T_3372_36_is_load : _GEN_22606;
  assign _GEN_22784 = 6'h25 == rob_head ? _T_3372_37_is_store : _GEN_22694;
  assign _GEN_22786 = 6'h25 == rob_head ? _T_3372_37_is_load : _GEN_22696;
  assign _GEN_22874 = 6'h26 == rob_head ? _T_3372_38_is_store : _GEN_22784;
  assign _GEN_22876 = 6'h26 == rob_head ? _T_3372_38_is_load : _GEN_22786;
  assign _GEN_22964 = 6'h27 == rob_head ? _T_3372_39_is_store : _GEN_22874;
  assign _GEN_22966 = 6'h27 == rob_head ? _T_3372_39_is_load : _GEN_22876;
  assign _GEN_22987 = 6'h1 == _T_2899 ? _T_3073_1 : _T_3073_0;
  assign _GEN_22988 = 6'h2 == _T_2899 ? _T_3073_2 : _GEN_22987;
  assign _GEN_22989 = 6'h3 == _T_2899 ? _T_3073_3 : _GEN_22988;
  assign _GEN_22990 = 6'h4 == _T_2899 ? _T_3073_4 : _GEN_22989;
  assign _GEN_22991 = 6'h5 == _T_2899 ? _T_3073_5 : _GEN_22990;
  assign _GEN_22992 = 6'h6 == _T_2899 ? _T_3073_6 : _GEN_22991;
  assign _GEN_22993 = 6'h7 == _T_2899 ? _T_3073_7 : _GEN_22992;
  assign _GEN_22994 = 6'h8 == _T_2899 ? _T_3073_8 : _GEN_22993;
  assign _GEN_22995 = 6'h9 == _T_2899 ? _T_3073_9 : _GEN_22994;
  assign _GEN_22996 = 6'ha == _T_2899 ? _T_3073_10 : _GEN_22995;
  assign _GEN_22997 = 6'hb == _T_2899 ? _T_3073_11 : _GEN_22996;
  assign _GEN_22998 = 6'hc == _T_2899 ? _T_3073_12 : _GEN_22997;
  assign _GEN_22999 = 6'hd == _T_2899 ? _T_3073_13 : _GEN_22998;
  assign _GEN_23000 = 6'he == _T_2899 ? _T_3073_14 : _GEN_22999;
  assign _GEN_23001 = 6'hf == _T_2899 ? _T_3073_15 : _GEN_23000;
  assign _GEN_23002 = 6'h10 == _T_2899 ? _T_3073_16 : _GEN_23001;
  assign _GEN_23003 = 6'h11 == _T_2899 ? _T_3073_17 : _GEN_23002;
  assign _GEN_23004 = 6'h12 == _T_2899 ? _T_3073_18 : _GEN_23003;
  assign _GEN_23005 = 6'h13 == _T_2899 ? _T_3073_19 : _GEN_23004;
  assign _GEN_23006 = 6'h14 == _T_2899 ? _T_3073_20 : _GEN_23005;
  assign _GEN_23007 = 6'h15 == _T_2899 ? _T_3073_21 : _GEN_23006;
  assign _GEN_23008 = 6'h16 == _T_2899 ? _T_3073_22 : _GEN_23007;
  assign _GEN_23009 = 6'h17 == _T_2899 ? _T_3073_23 : _GEN_23008;
  assign _GEN_23010 = 6'h18 == _T_2899 ? _T_3073_24 : _GEN_23009;
  assign _GEN_23011 = 6'h19 == _T_2899 ? _T_3073_25 : _GEN_23010;
  assign _GEN_23012 = 6'h1a == _T_2899 ? _T_3073_26 : _GEN_23011;
  assign _GEN_23013 = 6'h1b == _T_2899 ? _T_3073_27 : _GEN_23012;
  assign _GEN_23014 = 6'h1c == _T_2899 ? _T_3073_28 : _GEN_23013;
  assign _GEN_23015 = 6'h1d == _T_2899 ? _T_3073_29 : _GEN_23014;
  assign _GEN_23016 = 6'h1e == _T_2899 ? _T_3073_30 : _GEN_23015;
  assign _GEN_23017 = 6'h1f == _T_2899 ? _T_3073_31 : _GEN_23016;
  assign _GEN_23018 = 6'h20 == _T_2899 ? _T_3073_32 : _GEN_23017;
  assign _GEN_23019 = 6'h21 == _T_2899 ? _T_3073_33 : _GEN_23018;
  assign _GEN_23020 = 6'h22 == _T_2899 ? _T_3073_34 : _GEN_23019;
  assign _GEN_23021 = 6'h23 == _T_2899 ? _T_3073_35 : _GEN_23020;
  assign _GEN_23022 = 6'h24 == _T_2899 ? _T_3073_36 : _GEN_23021;
  assign _GEN_23023 = 6'h25 == _T_2899 ? _T_3073_37 : _GEN_23022;
  assign _GEN_23024 = 6'h26 == _T_2899 ? _T_3073_38 : _GEN_23023;
  assign _GEN_23025 = 6'h27 == _T_2899 ? _T_3073_39 : _GEN_23024;
  assign _T_5045 = _T_2790 == 7'h27;
  assign _T_5048 = _T_2790 + 7'h1;
  assign _T_5049 = _T_5048[6:0];
  assign _T_5050 = _T_5045 ? 7'h0 : _T_5049;
  assign _T_5054 = _T_5050[5:0];
  assign _GEN_23026 = 6'h1 == _T_5054 ? _T_3073_1 : _T_3073_0;
  assign _GEN_23027 = 6'h2 == _T_5054 ? _T_3073_2 : _GEN_23026;
  assign _GEN_23028 = 6'h3 == _T_5054 ? _T_3073_3 : _GEN_23027;
  assign _GEN_23029 = 6'h4 == _T_5054 ? _T_3073_4 : _GEN_23028;
  assign _GEN_23030 = 6'h5 == _T_5054 ? _T_3073_5 : _GEN_23029;
  assign _GEN_23031 = 6'h6 == _T_5054 ? _T_3073_6 : _GEN_23030;
  assign _GEN_23032 = 6'h7 == _T_5054 ? _T_3073_7 : _GEN_23031;
  assign _GEN_23033 = 6'h8 == _T_5054 ? _T_3073_8 : _GEN_23032;
  assign _GEN_23034 = 6'h9 == _T_5054 ? _T_3073_9 : _GEN_23033;
  assign _GEN_23035 = 6'ha == _T_5054 ? _T_3073_10 : _GEN_23034;
  assign _GEN_23036 = 6'hb == _T_5054 ? _T_3073_11 : _GEN_23035;
  assign _GEN_23037 = 6'hc == _T_5054 ? _T_3073_12 : _GEN_23036;
  assign _GEN_23038 = 6'hd == _T_5054 ? _T_3073_13 : _GEN_23037;
  assign _GEN_23039 = 6'he == _T_5054 ? _T_3073_14 : _GEN_23038;
  assign _GEN_23040 = 6'hf == _T_5054 ? _T_3073_15 : _GEN_23039;
  assign _GEN_23041 = 6'h10 == _T_5054 ? _T_3073_16 : _GEN_23040;
  assign _GEN_23042 = 6'h11 == _T_5054 ? _T_3073_17 : _GEN_23041;
  assign _GEN_23043 = 6'h12 == _T_5054 ? _T_3073_18 : _GEN_23042;
  assign _GEN_23044 = 6'h13 == _T_5054 ? _T_3073_19 : _GEN_23043;
  assign _GEN_23045 = 6'h14 == _T_5054 ? _T_3073_20 : _GEN_23044;
  assign _GEN_23046 = 6'h15 == _T_5054 ? _T_3073_21 : _GEN_23045;
  assign _GEN_23047 = 6'h16 == _T_5054 ? _T_3073_22 : _GEN_23046;
  assign _GEN_23048 = 6'h17 == _T_5054 ? _T_3073_23 : _GEN_23047;
  assign _GEN_23049 = 6'h18 == _T_5054 ? _T_3073_24 : _GEN_23048;
  assign _GEN_23050 = 6'h19 == _T_5054 ? _T_3073_25 : _GEN_23049;
  assign _GEN_23051 = 6'h1a == _T_5054 ? _T_3073_26 : _GEN_23050;
  assign _GEN_23052 = 6'h1b == _T_5054 ? _T_3073_27 : _GEN_23051;
  assign _GEN_23053 = 6'h1c == _T_5054 ? _T_3073_28 : _GEN_23052;
  assign _GEN_23054 = 6'h1d == _T_5054 ? _T_3073_29 : _GEN_23053;
  assign _GEN_23055 = 6'h1e == _T_5054 ? _T_3073_30 : _GEN_23054;
  assign _GEN_23056 = 6'h1f == _T_5054 ? _T_3073_31 : _GEN_23055;
  assign _GEN_23057 = 6'h20 == _T_5054 ? _T_3073_32 : _GEN_23056;
  assign _GEN_23058 = 6'h21 == _T_5054 ? _T_3073_33 : _GEN_23057;
  assign _GEN_23059 = 6'h22 == _T_5054 ? _T_3073_34 : _GEN_23058;
  assign _GEN_23060 = 6'h23 == _T_5054 ? _T_3073_35 : _GEN_23059;
  assign _GEN_23061 = 6'h24 == _T_5054 ? _T_3073_36 : _GEN_23060;
  assign _GEN_23062 = 6'h25 == _T_5054 ? _T_3073_37 : _GEN_23061;
  assign _GEN_23063 = 6'h26 == _T_5054 ? _T_3073_38 : _GEN_23062;
  assign _GEN_23064 = 6'h27 == _T_5054 ? _T_3073_39 : _GEN_23063;
  assign _GEN_23305 = 6'h1 == _T_3818 ? _T_3073_1 : _T_3073_0;
  assign _GEN_23306 = 6'h2 == _T_3818 ? _T_3073_2 : _GEN_23305;
  assign _GEN_23307 = 6'h3 == _T_3818 ? _T_3073_3 : _GEN_23306;
  assign _GEN_23308 = 6'h4 == _T_3818 ? _T_3073_4 : _GEN_23307;
  assign _GEN_23309 = 6'h5 == _T_3818 ? _T_3073_5 : _GEN_23308;
  assign _GEN_23310 = 6'h6 == _T_3818 ? _T_3073_6 : _GEN_23309;
  assign _GEN_23311 = 6'h7 == _T_3818 ? _T_3073_7 : _GEN_23310;
  assign _GEN_23312 = 6'h8 == _T_3818 ? _T_3073_8 : _GEN_23311;
  assign _GEN_23313 = 6'h9 == _T_3818 ? _T_3073_9 : _GEN_23312;
  assign _GEN_23314 = 6'ha == _T_3818 ? _T_3073_10 : _GEN_23313;
  assign _GEN_23315 = 6'hb == _T_3818 ? _T_3073_11 : _GEN_23314;
  assign _GEN_23316 = 6'hc == _T_3818 ? _T_3073_12 : _GEN_23315;
  assign _GEN_23317 = 6'hd == _T_3818 ? _T_3073_13 : _GEN_23316;
  assign _GEN_23318 = 6'he == _T_3818 ? _T_3073_14 : _GEN_23317;
  assign _GEN_23319 = 6'hf == _T_3818 ? _T_3073_15 : _GEN_23318;
  assign _GEN_23320 = 6'h10 == _T_3818 ? _T_3073_16 : _GEN_23319;
  assign _GEN_23321 = 6'h11 == _T_3818 ? _T_3073_17 : _GEN_23320;
  assign _GEN_23322 = 6'h12 == _T_3818 ? _T_3073_18 : _GEN_23321;
  assign _GEN_23323 = 6'h13 == _T_3818 ? _T_3073_19 : _GEN_23322;
  assign _GEN_23324 = 6'h14 == _T_3818 ? _T_3073_20 : _GEN_23323;
  assign _GEN_23325 = 6'h15 == _T_3818 ? _T_3073_21 : _GEN_23324;
  assign _GEN_23326 = 6'h16 == _T_3818 ? _T_3073_22 : _GEN_23325;
  assign _GEN_23327 = 6'h17 == _T_3818 ? _T_3073_23 : _GEN_23326;
  assign _GEN_23328 = 6'h18 == _T_3818 ? _T_3073_24 : _GEN_23327;
  assign _GEN_23329 = 6'h19 == _T_3818 ? _T_3073_25 : _GEN_23328;
  assign _GEN_23330 = 6'h1a == _T_3818 ? _T_3073_26 : _GEN_23329;
  assign _GEN_23331 = 6'h1b == _T_3818 ? _T_3073_27 : _GEN_23330;
  assign _GEN_23332 = 6'h1c == _T_3818 ? _T_3073_28 : _GEN_23331;
  assign _GEN_23333 = 6'h1d == _T_3818 ? _T_3073_29 : _GEN_23332;
  assign _GEN_23334 = 6'h1e == _T_3818 ? _T_3073_30 : _GEN_23333;
  assign _GEN_23335 = 6'h1f == _T_3818 ? _T_3073_31 : _GEN_23334;
  assign _GEN_23336 = 6'h20 == _T_3818 ? _T_3073_32 : _GEN_23335;
  assign _GEN_23337 = 6'h21 == _T_3818 ? _T_3073_33 : _GEN_23336;
  assign _GEN_23338 = 6'h22 == _T_3818 ? _T_3073_34 : _GEN_23337;
  assign _GEN_23339 = 6'h23 == _T_3818 ? _T_3073_35 : _GEN_23338;
  assign _GEN_23340 = 6'h24 == _T_3818 ? _T_3073_36 : _GEN_23339;
  assign _GEN_23341 = 6'h25 == _T_3818 ? _T_3073_37 : _GEN_23340;
  assign _GEN_23342 = 6'h26 == _T_3818 ? _T_3073_38 : _GEN_23341;
  assign _GEN_23343 = 6'h27 == _T_3818 ? _T_3073_39 : _GEN_23342;
  assign _T_5113 = _GEN_208 == 1'h0;
  assign _T_5114 = _T_3817 & _T_5113;
  assign _T_5116 = _T_5114 == 1'h0;
  assign _T_5118 = _T_5116 | reset;
  assign _T_5120 = _T_5118 == 1'h0;
  assign _T_5127 = _T_3813[5:0];
  assign _T_5130 = _T_3200__T_5128_data == 1'h0;
  assign _T_5131 = _T_3817 & _T_5130;
  assign _T_5133 = _T_5131 == 1'h0;
  assign _T_5135 = _T_5133 | reset;
  assign _T_5137 = _T_5135 == 1'h0;
  assign _GEN_23396 = 6'h1 == _T_3818 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_23421 = 6'h1 == _T_3818 ? _T_3372_1_ldst_val : _T_3372_0_ldst_val;
  assign _GEN_23486 = 6'h2 == _T_3818 ? _T_3372_2_pdst : _GEN_23396;
  assign _GEN_23511 = 6'h2 == _T_3818 ? _T_3372_2_ldst_val : _GEN_23421;
  assign _GEN_23576 = 6'h3 == _T_3818 ? _T_3372_3_pdst : _GEN_23486;
  assign _GEN_23601 = 6'h3 == _T_3818 ? _T_3372_3_ldst_val : _GEN_23511;
  assign _GEN_23666 = 6'h4 == _T_3818 ? _T_3372_4_pdst : _GEN_23576;
  assign _GEN_23691 = 6'h4 == _T_3818 ? _T_3372_4_ldst_val : _GEN_23601;
  assign _GEN_23756 = 6'h5 == _T_3818 ? _T_3372_5_pdst : _GEN_23666;
  assign _GEN_23781 = 6'h5 == _T_3818 ? _T_3372_5_ldst_val : _GEN_23691;
  assign _GEN_23846 = 6'h6 == _T_3818 ? _T_3372_6_pdst : _GEN_23756;
  assign _GEN_23871 = 6'h6 == _T_3818 ? _T_3372_6_ldst_val : _GEN_23781;
  assign _GEN_23936 = 6'h7 == _T_3818 ? _T_3372_7_pdst : _GEN_23846;
  assign _GEN_23961 = 6'h7 == _T_3818 ? _T_3372_7_ldst_val : _GEN_23871;
  assign _GEN_24026 = 6'h8 == _T_3818 ? _T_3372_8_pdst : _GEN_23936;
  assign _GEN_24051 = 6'h8 == _T_3818 ? _T_3372_8_ldst_val : _GEN_23961;
  assign _GEN_24116 = 6'h9 == _T_3818 ? _T_3372_9_pdst : _GEN_24026;
  assign _GEN_24141 = 6'h9 == _T_3818 ? _T_3372_9_ldst_val : _GEN_24051;
  assign _GEN_24206 = 6'ha == _T_3818 ? _T_3372_10_pdst : _GEN_24116;
  assign _GEN_24231 = 6'ha == _T_3818 ? _T_3372_10_ldst_val : _GEN_24141;
  assign _GEN_24296 = 6'hb == _T_3818 ? _T_3372_11_pdst : _GEN_24206;
  assign _GEN_24321 = 6'hb == _T_3818 ? _T_3372_11_ldst_val : _GEN_24231;
  assign _GEN_24386 = 6'hc == _T_3818 ? _T_3372_12_pdst : _GEN_24296;
  assign _GEN_24411 = 6'hc == _T_3818 ? _T_3372_12_ldst_val : _GEN_24321;
  assign _GEN_24476 = 6'hd == _T_3818 ? _T_3372_13_pdst : _GEN_24386;
  assign _GEN_24501 = 6'hd == _T_3818 ? _T_3372_13_ldst_val : _GEN_24411;
  assign _GEN_24566 = 6'he == _T_3818 ? _T_3372_14_pdst : _GEN_24476;
  assign _GEN_24591 = 6'he == _T_3818 ? _T_3372_14_ldst_val : _GEN_24501;
  assign _GEN_24656 = 6'hf == _T_3818 ? _T_3372_15_pdst : _GEN_24566;
  assign _GEN_24681 = 6'hf == _T_3818 ? _T_3372_15_ldst_val : _GEN_24591;
  assign _GEN_24746 = 6'h10 == _T_3818 ? _T_3372_16_pdst : _GEN_24656;
  assign _GEN_24771 = 6'h10 == _T_3818 ? _T_3372_16_ldst_val : _GEN_24681;
  assign _GEN_24836 = 6'h11 == _T_3818 ? _T_3372_17_pdst : _GEN_24746;
  assign _GEN_24861 = 6'h11 == _T_3818 ? _T_3372_17_ldst_val : _GEN_24771;
  assign _GEN_24926 = 6'h12 == _T_3818 ? _T_3372_18_pdst : _GEN_24836;
  assign _GEN_24951 = 6'h12 == _T_3818 ? _T_3372_18_ldst_val : _GEN_24861;
  assign _GEN_25016 = 6'h13 == _T_3818 ? _T_3372_19_pdst : _GEN_24926;
  assign _GEN_25041 = 6'h13 == _T_3818 ? _T_3372_19_ldst_val : _GEN_24951;
  assign _GEN_25106 = 6'h14 == _T_3818 ? _T_3372_20_pdst : _GEN_25016;
  assign _GEN_25131 = 6'h14 == _T_3818 ? _T_3372_20_ldst_val : _GEN_25041;
  assign _GEN_25196 = 6'h15 == _T_3818 ? _T_3372_21_pdst : _GEN_25106;
  assign _GEN_25221 = 6'h15 == _T_3818 ? _T_3372_21_ldst_val : _GEN_25131;
  assign _GEN_25286 = 6'h16 == _T_3818 ? _T_3372_22_pdst : _GEN_25196;
  assign _GEN_25311 = 6'h16 == _T_3818 ? _T_3372_22_ldst_val : _GEN_25221;
  assign _GEN_25376 = 6'h17 == _T_3818 ? _T_3372_23_pdst : _GEN_25286;
  assign _GEN_25401 = 6'h17 == _T_3818 ? _T_3372_23_ldst_val : _GEN_25311;
  assign _GEN_25466 = 6'h18 == _T_3818 ? _T_3372_24_pdst : _GEN_25376;
  assign _GEN_25491 = 6'h18 == _T_3818 ? _T_3372_24_ldst_val : _GEN_25401;
  assign _GEN_25556 = 6'h19 == _T_3818 ? _T_3372_25_pdst : _GEN_25466;
  assign _GEN_25581 = 6'h19 == _T_3818 ? _T_3372_25_ldst_val : _GEN_25491;
  assign _GEN_25646 = 6'h1a == _T_3818 ? _T_3372_26_pdst : _GEN_25556;
  assign _GEN_25671 = 6'h1a == _T_3818 ? _T_3372_26_ldst_val : _GEN_25581;
  assign _GEN_25736 = 6'h1b == _T_3818 ? _T_3372_27_pdst : _GEN_25646;
  assign _GEN_25761 = 6'h1b == _T_3818 ? _T_3372_27_ldst_val : _GEN_25671;
  assign _GEN_25826 = 6'h1c == _T_3818 ? _T_3372_28_pdst : _GEN_25736;
  assign _GEN_25851 = 6'h1c == _T_3818 ? _T_3372_28_ldst_val : _GEN_25761;
  assign _GEN_25916 = 6'h1d == _T_3818 ? _T_3372_29_pdst : _GEN_25826;
  assign _GEN_25941 = 6'h1d == _T_3818 ? _T_3372_29_ldst_val : _GEN_25851;
  assign _GEN_26006 = 6'h1e == _T_3818 ? _T_3372_30_pdst : _GEN_25916;
  assign _GEN_26031 = 6'h1e == _T_3818 ? _T_3372_30_ldst_val : _GEN_25941;
  assign _GEN_26096 = 6'h1f == _T_3818 ? _T_3372_31_pdst : _GEN_26006;
  assign _GEN_26121 = 6'h1f == _T_3818 ? _T_3372_31_ldst_val : _GEN_26031;
  assign _GEN_26186 = 6'h20 == _T_3818 ? _T_3372_32_pdst : _GEN_26096;
  assign _GEN_26211 = 6'h20 == _T_3818 ? _T_3372_32_ldst_val : _GEN_26121;
  assign _GEN_26276 = 6'h21 == _T_3818 ? _T_3372_33_pdst : _GEN_26186;
  assign _GEN_26301 = 6'h21 == _T_3818 ? _T_3372_33_ldst_val : _GEN_26211;
  assign _GEN_26366 = 6'h22 == _T_3818 ? _T_3372_34_pdst : _GEN_26276;
  assign _GEN_26391 = 6'h22 == _T_3818 ? _T_3372_34_ldst_val : _GEN_26301;
  assign _GEN_26456 = 6'h23 == _T_3818 ? _T_3372_35_pdst : _GEN_26366;
  assign _GEN_26481 = 6'h23 == _T_3818 ? _T_3372_35_ldst_val : _GEN_26391;
  assign _GEN_26546 = 6'h24 == _T_3818 ? _T_3372_36_pdst : _GEN_26456;
  assign _GEN_26571 = 6'h24 == _T_3818 ? _T_3372_36_ldst_val : _GEN_26481;
  assign _GEN_26636 = 6'h25 == _T_3818 ? _T_3372_37_pdst : _GEN_26546;
  assign _GEN_26661 = 6'h25 == _T_3818 ? _T_3372_37_ldst_val : _GEN_26571;
  assign _GEN_26726 = 6'h26 == _T_3818 ? _T_3372_38_pdst : _GEN_26636;
  assign _GEN_26751 = 6'h26 == _T_3818 ? _T_3372_38_ldst_val : _GEN_26661;
  assign _GEN_26816 = 6'h27 == _T_3818 ? _T_3372_39_pdst : _GEN_26726;
  assign _GEN_26841 = 6'h27 == _T_3818 ? _T_3372_39_ldst_val : _GEN_26751;
  assign _T_5142 = _T_3817 & _GEN_209_ldst_val;
  assign _T_5143 = _GEN_210_pdst != io_wb_resps_0_bits_uop_pdst;
  assign _T_5144 = _T_5142 & _T_5143;
  assign _T_5146 = _T_5144 == 1'h0;
  assign _T_5148 = _T_5146 | reset;
  assign _T_5150 = _T_5148 == 1'h0;
  assign _GEN_26934 = 6'h1 == _T_3827 ? _T_3073_1 : _T_3073_0;
  assign _GEN_26935 = 6'h2 == _T_3827 ? _T_3073_2 : _GEN_26934;
  assign _GEN_26936 = 6'h3 == _T_3827 ? _T_3073_3 : _GEN_26935;
  assign _GEN_26937 = 6'h4 == _T_3827 ? _T_3073_4 : _GEN_26936;
  assign _GEN_26938 = 6'h5 == _T_3827 ? _T_3073_5 : _GEN_26937;
  assign _GEN_26939 = 6'h6 == _T_3827 ? _T_3073_6 : _GEN_26938;
  assign _GEN_26940 = 6'h7 == _T_3827 ? _T_3073_7 : _GEN_26939;
  assign _GEN_26941 = 6'h8 == _T_3827 ? _T_3073_8 : _GEN_26940;
  assign _GEN_26942 = 6'h9 == _T_3827 ? _T_3073_9 : _GEN_26941;
  assign _GEN_26943 = 6'ha == _T_3827 ? _T_3073_10 : _GEN_26942;
  assign _GEN_26944 = 6'hb == _T_3827 ? _T_3073_11 : _GEN_26943;
  assign _GEN_26945 = 6'hc == _T_3827 ? _T_3073_12 : _GEN_26944;
  assign _GEN_26946 = 6'hd == _T_3827 ? _T_3073_13 : _GEN_26945;
  assign _GEN_26947 = 6'he == _T_3827 ? _T_3073_14 : _GEN_26946;
  assign _GEN_26948 = 6'hf == _T_3827 ? _T_3073_15 : _GEN_26947;
  assign _GEN_26949 = 6'h10 == _T_3827 ? _T_3073_16 : _GEN_26948;
  assign _GEN_26950 = 6'h11 == _T_3827 ? _T_3073_17 : _GEN_26949;
  assign _GEN_26951 = 6'h12 == _T_3827 ? _T_3073_18 : _GEN_26950;
  assign _GEN_26952 = 6'h13 == _T_3827 ? _T_3073_19 : _GEN_26951;
  assign _GEN_26953 = 6'h14 == _T_3827 ? _T_3073_20 : _GEN_26952;
  assign _GEN_26954 = 6'h15 == _T_3827 ? _T_3073_21 : _GEN_26953;
  assign _GEN_26955 = 6'h16 == _T_3827 ? _T_3073_22 : _GEN_26954;
  assign _GEN_26956 = 6'h17 == _T_3827 ? _T_3073_23 : _GEN_26955;
  assign _GEN_26957 = 6'h18 == _T_3827 ? _T_3073_24 : _GEN_26956;
  assign _GEN_26958 = 6'h19 == _T_3827 ? _T_3073_25 : _GEN_26957;
  assign _GEN_26959 = 6'h1a == _T_3827 ? _T_3073_26 : _GEN_26958;
  assign _GEN_26960 = 6'h1b == _T_3827 ? _T_3073_27 : _GEN_26959;
  assign _GEN_26961 = 6'h1c == _T_3827 ? _T_3073_28 : _GEN_26960;
  assign _GEN_26962 = 6'h1d == _T_3827 ? _T_3073_29 : _GEN_26961;
  assign _GEN_26963 = 6'h1e == _T_3827 ? _T_3073_30 : _GEN_26962;
  assign _GEN_26964 = 6'h1f == _T_3827 ? _T_3073_31 : _GEN_26963;
  assign _GEN_26965 = 6'h20 == _T_3827 ? _T_3073_32 : _GEN_26964;
  assign _GEN_26966 = 6'h21 == _T_3827 ? _T_3073_33 : _GEN_26965;
  assign _GEN_26967 = 6'h22 == _T_3827 ? _T_3073_34 : _GEN_26966;
  assign _GEN_26968 = 6'h23 == _T_3827 ? _T_3073_35 : _GEN_26967;
  assign _GEN_26969 = 6'h24 == _T_3827 ? _T_3073_36 : _GEN_26968;
  assign _GEN_26970 = 6'h25 == _T_3827 ? _T_3073_37 : _GEN_26969;
  assign _GEN_26971 = 6'h26 == _T_3827 ? _T_3073_38 : _GEN_26970;
  assign _GEN_26972 = 6'h27 == _T_3827 ? _T_3073_39 : _GEN_26971;
  assign _T_5190 = _GEN_212 == 1'h0;
  assign _T_5191 = _T_3826 & _T_5190;
  assign _T_5193 = _T_5191 == 1'h0;
  assign _T_5195 = _T_5193 | reset;
  assign _T_5197 = _T_5195 == 1'h0;
  assign _T_5204 = _T_3822[5:0];
  assign _T_5207 = _T_3200__T_5205_data == 1'h0;
  assign _T_5208 = _T_3826 & _T_5207;
  assign _T_5210 = _T_5208 == 1'h0;
  assign _T_5212 = _T_5210 | reset;
  assign _T_5214 = _T_5212 == 1'h0;
  assign _GEN_27025 = 6'h1 == _T_3827 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_27050 = 6'h1 == _T_3827 ? _T_3372_1_ldst_val : _T_3372_0_ldst_val;
  assign _GEN_27115 = 6'h2 == _T_3827 ? _T_3372_2_pdst : _GEN_27025;
  assign _GEN_27140 = 6'h2 == _T_3827 ? _T_3372_2_ldst_val : _GEN_27050;
  assign _GEN_27205 = 6'h3 == _T_3827 ? _T_3372_3_pdst : _GEN_27115;
  assign _GEN_27230 = 6'h3 == _T_3827 ? _T_3372_3_ldst_val : _GEN_27140;
  assign _GEN_27295 = 6'h4 == _T_3827 ? _T_3372_4_pdst : _GEN_27205;
  assign _GEN_27320 = 6'h4 == _T_3827 ? _T_3372_4_ldst_val : _GEN_27230;
  assign _GEN_27385 = 6'h5 == _T_3827 ? _T_3372_5_pdst : _GEN_27295;
  assign _GEN_27410 = 6'h5 == _T_3827 ? _T_3372_5_ldst_val : _GEN_27320;
  assign _GEN_27475 = 6'h6 == _T_3827 ? _T_3372_6_pdst : _GEN_27385;
  assign _GEN_27500 = 6'h6 == _T_3827 ? _T_3372_6_ldst_val : _GEN_27410;
  assign _GEN_27565 = 6'h7 == _T_3827 ? _T_3372_7_pdst : _GEN_27475;
  assign _GEN_27590 = 6'h7 == _T_3827 ? _T_3372_7_ldst_val : _GEN_27500;
  assign _GEN_27655 = 6'h8 == _T_3827 ? _T_3372_8_pdst : _GEN_27565;
  assign _GEN_27680 = 6'h8 == _T_3827 ? _T_3372_8_ldst_val : _GEN_27590;
  assign _GEN_27745 = 6'h9 == _T_3827 ? _T_3372_9_pdst : _GEN_27655;
  assign _GEN_27770 = 6'h9 == _T_3827 ? _T_3372_9_ldst_val : _GEN_27680;
  assign _GEN_27835 = 6'ha == _T_3827 ? _T_3372_10_pdst : _GEN_27745;
  assign _GEN_27860 = 6'ha == _T_3827 ? _T_3372_10_ldst_val : _GEN_27770;
  assign _GEN_27925 = 6'hb == _T_3827 ? _T_3372_11_pdst : _GEN_27835;
  assign _GEN_27950 = 6'hb == _T_3827 ? _T_3372_11_ldst_val : _GEN_27860;
  assign _GEN_28015 = 6'hc == _T_3827 ? _T_3372_12_pdst : _GEN_27925;
  assign _GEN_28040 = 6'hc == _T_3827 ? _T_3372_12_ldst_val : _GEN_27950;
  assign _GEN_28105 = 6'hd == _T_3827 ? _T_3372_13_pdst : _GEN_28015;
  assign _GEN_28130 = 6'hd == _T_3827 ? _T_3372_13_ldst_val : _GEN_28040;
  assign _GEN_28195 = 6'he == _T_3827 ? _T_3372_14_pdst : _GEN_28105;
  assign _GEN_28220 = 6'he == _T_3827 ? _T_3372_14_ldst_val : _GEN_28130;
  assign _GEN_28285 = 6'hf == _T_3827 ? _T_3372_15_pdst : _GEN_28195;
  assign _GEN_28310 = 6'hf == _T_3827 ? _T_3372_15_ldst_val : _GEN_28220;
  assign _GEN_28375 = 6'h10 == _T_3827 ? _T_3372_16_pdst : _GEN_28285;
  assign _GEN_28400 = 6'h10 == _T_3827 ? _T_3372_16_ldst_val : _GEN_28310;
  assign _GEN_28465 = 6'h11 == _T_3827 ? _T_3372_17_pdst : _GEN_28375;
  assign _GEN_28490 = 6'h11 == _T_3827 ? _T_3372_17_ldst_val : _GEN_28400;
  assign _GEN_28555 = 6'h12 == _T_3827 ? _T_3372_18_pdst : _GEN_28465;
  assign _GEN_28580 = 6'h12 == _T_3827 ? _T_3372_18_ldst_val : _GEN_28490;
  assign _GEN_28645 = 6'h13 == _T_3827 ? _T_3372_19_pdst : _GEN_28555;
  assign _GEN_28670 = 6'h13 == _T_3827 ? _T_3372_19_ldst_val : _GEN_28580;
  assign _GEN_28735 = 6'h14 == _T_3827 ? _T_3372_20_pdst : _GEN_28645;
  assign _GEN_28760 = 6'h14 == _T_3827 ? _T_3372_20_ldst_val : _GEN_28670;
  assign _GEN_28825 = 6'h15 == _T_3827 ? _T_3372_21_pdst : _GEN_28735;
  assign _GEN_28850 = 6'h15 == _T_3827 ? _T_3372_21_ldst_val : _GEN_28760;
  assign _GEN_28915 = 6'h16 == _T_3827 ? _T_3372_22_pdst : _GEN_28825;
  assign _GEN_28940 = 6'h16 == _T_3827 ? _T_3372_22_ldst_val : _GEN_28850;
  assign _GEN_29005 = 6'h17 == _T_3827 ? _T_3372_23_pdst : _GEN_28915;
  assign _GEN_29030 = 6'h17 == _T_3827 ? _T_3372_23_ldst_val : _GEN_28940;
  assign _GEN_29095 = 6'h18 == _T_3827 ? _T_3372_24_pdst : _GEN_29005;
  assign _GEN_29120 = 6'h18 == _T_3827 ? _T_3372_24_ldst_val : _GEN_29030;
  assign _GEN_29185 = 6'h19 == _T_3827 ? _T_3372_25_pdst : _GEN_29095;
  assign _GEN_29210 = 6'h19 == _T_3827 ? _T_3372_25_ldst_val : _GEN_29120;
  assign _GEN_29275 = 6'h1a == _T_3827 ? _T_3372_26_pdst : _GEN_29185;
  assign _GEN_29300 = 6'h1a == _T_3827 ? _T_3372_26_ldst_val : _GEN_29210;
  assign _GEN_29365 = 6'h1b == _T_3827 ? _T_3372_27_pdst : _GEN_29275;
  assign _GEN_29390 = 6'h1b == _T_3827 ? _T_3372_27_ldst_val : _GEN_29300;
  assign _GEN_29455 = 6'h1c == _T_3827 ? _T_3372_28_pdst : _GEN_29365;
  assign _GEN_29480 = 6'h1c == _T_3827 ? _T_3372_28_ldst_val : _GEN_29390;
  assign _GEN_29545 = 6'h1d == _T_3827 ? _T_3372_29_pdst : _GEN_29455;
  assign _GEN_29570 = 6'h1d == _T_3827 ? _T_3372_29_ldst_val : _GEN_29480;
  assign _GEN_29635 = 6'h1e == _T_3827 ? _T_3372_30_pdst : _GEN_29545;
  assign _GEN_29660 = 6'h1e == _T_3827 ? _T_3372_30_ldst_val : _GEN_29570;
  assign _GEN_29725 = 6'h1f == _T_3827 ? _T_3372_31_pdst : _GEN_29635;
  assign _GEN_29750 = 6'h1f == _T_3827 ? _T_3372_31_ldst_val : _GEN_29660;
  assign _GEN_29815 = 6'h20 == _T_3827 ? _T_3372_32_pdst : _GEN_29725;
  assign _GEN_29840 = 6'h20 == _T_3827 ? _T_3372_32_ldst_val : _GEN_29750;
  assign _GEN_29905 = 6'h21 == _T_3827 ? _T_3372_33_pdst : _GEN_29815;
  assign _GEN_29930 = 6'h21 == _T_3827 ? _T_3372_33_ldst_val : _GEN_29840;
  assign _GEN_29995 = 6'h22 == _T_3827 ? _T_3372_34_pdst : _GEN_29905;
  assign _GEN_30020 = 6'h22 == _T_3827 ? _T_3372_34_ldst_val : _GEN_29930;
  assign _GEN_30085 = 6'h23 == _T_3827 ? _T_3372_35_pdst : _GEN_29995;
  assign _GEN_30110 = 6'h23 == _T_3827 ? _T_3372_35_ldst_val : _GEN_30020;
  assign _GEN_30175 = 6'h24 == _T_3827 ? _T_3372_36_pdst : _GEN_30085;
  assign _GEN_30200 = 6'h24 == _T_3827 ? _T_3372_36_ldst_val : _GEN_30110;
  assign _GEN_30265 = 6'h25 == _T_3827 ? _T_3372_37_pdst : _GEN_30175;
  assign _GEN_30290 = 6'h25 == _T_3827 ? _T_3372_37_ldst_val : _GEN_30200;
  assign _GEN_30355 = 6'h26 == _T_3827 ? _T_3372_38_pdst : _GEN_30265;
  assign _GEN_30380 = 6'h26 == _T_3827 ? _T_3372_38_ldst_val : _GEN_30290;
  assign _GEN_30445 = 6'h27 == _T_3827 ? _T_3372_39_pdst : _GEN_30355;
  assign _GEN_30470 = 6'h27 == _T_3827 ? _T_3372_39_ldst_val : _GEN_30380;
  assign _T_5219 = _T_3826 & _GEN_213_ldst_val;
  assign _T_5220 = _GEN_214_pdst != io_wb_resps_1_bits_uop_pdst;
  assign _T_5221 = _T_5219 & _T_5220;
  assign _T_5223 = _T_5221 == 1'h0;
  assign _T_5225 = _T_5223 | reset;
  assign _T_5227 = _T_5225 == 1'h0;
  assign _GEN_30563 = 6'h1 == _T_3836 ? _T_3073_1 : _T_3073_0;
  assign _GEN_30564 = 6'h2 == _T_3836 ? _T_3073_2 : _GEN_30563;
  assign _GEN_30565 = 6'h3 == _T_3836 ? _T_3073_3 : _GEN_30564;
  assign _GEN_30566 = 6'h4 == _T_3836 ? _T_3073_4 : _GEN_30565;
  assign _GEN_30567 = 6'h5 == _T_3836 ? _T_3073_5 : _GEN_30566;
  assign _GEN_30568 = 6'h6 == _T_3836 ? _T_3073_6 : _GEN_30567;
  assign _GEN_30569 = 6'h7 == _T_3836 ? _T_3073_7 : _GEN_30568;
  assign _GEN_30570 = 6'h8 == _T_3836 ? _T_3073_8 : _GEN_30569;
  assign _GEN_30571 = 6'h9 == _T_3836 ? _T_3073_9 : _GEN_30570;
  assign _GEN_30572 = 6'ha == _T_3836 ? _T_3073_10 : _GEN_30571;
  assign _GEN_30573 = 6'hb == _T_3836 ? _T_3073_11 : _GEN_30572;
  assign _GEN_30574 = 6'hc == _T_3836 ? _T_3073_12 : _GEN_30573;
  assign _GEN_30575 = 6'hd == _T_3836 ? _T_3073_13 : _GEN_30574;
  assign _GEN_30576 = 6'he == _T_3836 ? _T_3073_14 : _GEN_30575;
  assign _GEN_30577 = 6'hf == _T_3836 ? _T_3073_15 : _GEN_30576;
  assign _GEN_30578 = 6'h10 == _T_3836 ? _T_3073_16 : _GEN_30577;
  assign _GEN_30579 = 6'h11 == _T_3836 ? _T_3073_17 : _GEN_30578;
  assign _GEN_30580 = 6'h12 == _T_3836 ? _T_3073_18 : _GEN_30579;
  assign _GEN_30581 = 6'h13 == _T_3836 ? _T_3073_19 : _GEN_30580;
  assign _GEN_30582 = 6'h14 == _T_3836 ? _T_3073_20 : _GEN_30581;
  assign _GEN_30583 = 6'h15 == _T_3836 ? _T_3073_21 : _GEN_30582;
  assign _GEN_30584 = 6'h16 == _T_3836 ? _T_3073_22 : _GEN_30583;
  assign _GEN_30585 = 6'h17 == _T_3836 ? _T_3073_23 : _GEN_30584;
  assign _GEN_30586 = 6'h18 == _T_3836 ? _T_3073_24 : _GEN_30585;
  assign _GEN_30587 = 6'h19 == _T_3836 ? _T_3073_25 : _GEN_30586;
  assign _GEN_30588 = 6'h1a == _T_3836 ? _T_3073_26 : _GEN_30587;
  assign _GEN_30589 = 6'h1b == _T_3836 ? _T_3073_27 : _GEN_30588;
  assign _GEN_30590 = 6'h1c == _T_3836 ? _T_3073_28 : _GEN_30589;
  assign _GEN_30591 = 6'h1d == _T_3836 ? _T_3073_29 : _GEN_30590;
  assign _GEN_30592 = 6'h1e == _T_3836 ? _T_3073_30 : _GEN_30591;
  assign _GEN_30593 = 6'h1f == _T_3836 ? _T_3073_31 : _GEN_30592;
  assign _GEN_30594 = 6'h20 == _T_3836 ? _T_3073_32 : _GEN_30593;
  assign _GEN_30595 = 6'h21 == _T_3836 ? _T_3073_33 : _GEN_30594;
  assign _GEN_30596 = 6'h22 == _T_3836 ? _T_3073_34 : _GEN_30595;
  assign _GEN_30597 = 6'h23 == _T_3836 ? _T_3073_35 : _GEN_30596;
  assign _GEN_30598 = 6'h24 == _T_3836 ? _T_3073_36 : _GEN_30597;
  assign _GEN_30599 = 6'h25 == _T_3836 ? _T_3073_37 : _GEN_30598;
  assign _GEN_30600 = 6'h26 == _T_3836 ? _T_3073_38 : _GEN_30599;
  assign _GEN_30601 = 6'h27 == _T_3836 ? _T_3073_39 : _GEN_30600;
  assign _T_5267 = _GEN_216 == 1'h0;
  assign _T_5268 = _T_3835 & _T_5267;
  assign _T_5270 = _T_5268 == 1'h0;
  assign _T_5272 = _T_5270 | reset;
  assign _T_5274 = _T_5272 == 1'h0;
  assign _T_5281 = _T_3831[5:0];
  assign _T_5284 = _T_3200__T_5282_data == 1'h0;
  assign _T_5285 = _T_3835 & _T_5284;
  assign _T_5287 = _T_5285 == 1'h0;
  assign _T_5289 = _T_5287 | reset;
  assign _T_5291 = _T_5289 == 1'h0;
  assign _GEN_30654 = 6'h1 == _T_3836 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_30679 = 6'h1 == _T_3836 ? _T_3372_1_ldst_val : _T_3372_0_ldst_val;
  assign _GEN_30744 = 6'h2 == _T_3836 ? _T_3372_2_pdst : _GEN_30654;
  assign _GEN_30769 = 6'h2 == _T_3836 ? _T_3372_2_ldst_val : _GEN_30679;
  assign _GEN_30834 = 6'h3 == _T_3836 ? _T_3372_3_pdst : _GEN_30744;
  assign _GEN_30859 = 6'h3 == _T_3836 ? _T_3372_3_ldst_val : _GEN_30769;
  assign _GEN_30924 = 6'h4 == _T_3836 ? _T_3372_4_pdst : _GEN_30834;
  assign _GEN_30949 = 6'h4 == _T_3836 ? _T_3372_4_ldst_val : _GEN_30859;
  assign _GEN_31014 = 6'h5 == _T_3836 ? _T_3372_5_pdst : _GEN_30924;
  assign _GEN_31039 = 6'h5 == _T_3836 ? _T_3372_5_ldst_val : _GEN_30949;
  assign _GEN_31104 = 6'h6 == _T_3836 ? _T_3372_6_pdst : _GEN_31014;
  assign _GEN_31129 = 6'h6 == _T_3836 ? _T_3372_6_ldst_val : _GEN_31039;
  assign _GEN_31194 = 6'h7 == _T_3836 ? _T_3372_7_pdst : _GEN_31104;
  assign _GEN_31219 = 6'h7 == _T_3836 ? _T_3372_7_ldst_val : _GEN_31129;
  assign _GEN_31284 = 6'h8 == _T_3836 ? _T_3372_8_pdst : _GEN_31194;
  assign _GEN_31309 = 6'h8 == _T_3836 ? _T_3372_8_ldst_val : _GEN_31219;
  assign _GEN_31374 = 6'h9 == _T_3836 ? _T_3372_9_pdst : _GEN_31284;
  assign _GEN_31399 = 6'h9 == _T_3836 ? _T_3372_9_ldst_val : _GEN_31309;
  assign _GEN_31464 = 6'ha == _T_3836 ? _T_3372_10_pdst : _GEN_31374;
  assign _GEN_31489 = 6'ha == _T_3836 ? _T_3372_10_ldst_val : _GEN_31399;
  assign _GEN_31554 = 6'hb == _T_3836 ? _T_3372_11_pdst : _GEN_31464;
  assign _GEN_31579 = 6'hb == _T_3836 ? _T_3372_11_ldst_val : _GEN_31489;
  assign _GEN_31644 = 6'hc == _T_3836 ? _T_3372_12_pdst : _GEN_31554;
  assign _GEN_31669 = 6'hc == _T_3836 ? _T_3372_12_ldst_val : _GEN_31579;
  assign _GEN_31734 = 6'hd == _T_3836 ? _T_3372_13_pdst : _GEN_31644;
  assign _GEN_31759 = 6'hd == _T_3836 ? _T_3372_13_ldst_val : _GEN_31669;
  assign _GEN_31824 = 6'he == _T_3836 ? _T_3372_14_pdst : _GEN_31734;
  assign _GEN_31849 = 6'he == _T_3836 ? _T_3372_14_ldst_val : _GEN_31759;
  assign _GEN_31914 = 6'hf == _T_3836 ? _T_3372_15_pdst : _GEN_31824;
  assign _GEN_31939 = 6'hf == _T_3836 ? _T_3372_15_ldst_val : _GEN_31849;
  assign _GEN_32004 = 6'h10 == _T_3836 ? _T_3372_16_pdst : _GEN_31914;
  assign _GEN_32029 = 6'h10 == _T_3836 ? _T_3372_16_ldst_val : _GEN_31939;
  assign _GEN_32094 = 6'h11 == _T_3836 ? _T_3372_17_pdst : _GEN_32004;
  assign _GEN_32119 = 6'h11 == _T_3836 ? _T_3372_17_ldst_val : _GEN_32029;
  assign _GEN_32184 = 6'h12 == _T_3836 ? _T_3372_18_pdst : _GEN_32094;
  assign _GEN_32209 = 6'h12 == _T_3836 ? _T_3372_18_ldst_val : _GEN_32119;
  assign _GEN_32274 = 6'h13 == _T_3836 ? _T_3372_19_pdst : _GEN_32184;
  assign _GEN_32299 = 6'h13 == _T_3836 ? _T_3372_19_ldst_val : _GEN_32209;
  assign _GEN_32364 = 6'h14 == _T_3836 ? _T_3372_20_pdst : _GEN_32274;
  assign _GEN_32389 = 6'h14 == _T_3836 ? _T_3372_20_ldst_val : _GEN_32299;
  assign _GEN_32454 = 6'h15 == _T_3836 ? _T_3372_21_pdst : _GEN_32364;
  assign _GEN_32479 = 6'h15 == _T_3836 ? _T_3372_21_ldst_val : _GEN_32389;
  assign _GEN_32544 = 6'h16 == _T_3836 ? _T_3372_22_pdst : _GEN_32454;
  assign _GEN_32569 = 6'h16 == _T_3836 ? _T_3372_22_ldst_val : _GEN_32479;
  assign _GEN_32634 = 6'h17 == _T_3836 ? _T_3372_23_pdst : _GEN_32544;
  assign _GEN_32659 = 6'h17 == _T_3836 ? _T_3372_23_ldst_val : _GEN_32569;
  assign _GEN_32724 = 6'h18 == _T_3836 ? _T_3372_24_pdst : _GEN_32634;
  assign _GEN_32749 = 6'h18 == _T_3836 ? _T_3372_24_ldst_val : _GEN_32659;
  assign _GEN_32814 = 6'h19 == _T_3836 ? _T_3372_25_pdst : _GEN_32724;
  assign _GEN_32839 = 6'h19 == _T_3836 ? _T_3372_25_ldst_val : _GEN_32749;
  assign _GEN_32904 = 6'h1a == _T_3836 ? _T_3372_26_pdst : _GEN_32814;
  assign _GEN_32929 = 6'h1a == _T_3836 ? _T_3372_26_ldst_val : _GEN_32839;
  assign _GEN_32994 = 6'h1b == _T_3836 ? _T_3372_27_pdst : _GEN_32904;
  assign _GEN_33019 = 6'h1b == _T_3836 ? _T_3372_27_ldst_val : _GEN_32929;
  assign _GEN_33084 = 6'h1c == _T_3836 ? _T_3372_28_pdst : _GEN_32994;
  assign _GEN_33109 = 6'h1c == _T_3836 ? _T_3372_28_ldst_val : _GEN_33019;
  assign _GEN_33174 = 6'h1d == _T_3836 ? _T_3372_29_pdst : _GEN_33084;
  assign _GEN_33199 = 6'h1d == _T_3836 ? _T_3372_29_ldst_val : _GEN_33109;
  assign _GEN_33264 = 6'h1e == _T_3836 ? _T_3372_30_pdst : _GEN_33174;
  assign _GEN_33289 = 6'h1e == _T_3836 ? _T_3372_30_ldst_val : _GEN_33199;
  assign _GEN_33354 = 6'h1f == _T_3836 ? _T_3372_31_pdst : _GEN_33264;
  assign _GEN_33379 = 6'h1f == _T_3836 ? _T_3372_31_ldst_val : _GEN_33289;
  assign _GEN_33444 = 6'h20 == _T_3836 ? _T_3372_32_pdst : _GEN_33354;
  assign _GEN_33469 = 6'h20 == _T_3836 ? _T_3372_32_ldst_val : _GEN_33379;
  assign _GEN_33534 = 6'h21 == _T_3836 ? _T_3372_33_pdst : _GEN_33444;
  assign _GEN_33559 = 6'h21 == _T_3836 ? _T_3372_33_ldst_val : _GEN_33469;
  assign _GEN_33624 = 6'h22 == _T_3836 ? _T_3372_34_pdst : _GEN_33534;
  assign _GEN_33649 = 6'h22 == _T_3836 ? _T_3372_34_ldst_val : _GEN_33559;
  assign _GEN_33714 = 6'h23 == _T_3836 ? _T_3372_35_pdst : _GEN_33624;
  assign _GEN_33739 = 6'h23 == _T_3836 ? _T_3372_35_ldst_val : _GEN_33649;
  assign _GEN_33804 = 6'h24 == _T_3836 ? _T_3372_36_pdst : _GEN_33714;
  assign _GEN_33829 = 6'h24 == _T_3836 ? _T_3372_36_ldst_val : _GEN_33739;
  assign _GEN_33894 = 6'h25 == _T_3836 ? _T_3372_37_pdst : _GEN_33804;
  assign _GEN_33919 = 6'h25 == _T_3836 ? _T_3372_37_ldst_val : _GEN_33829;
  assign _GEN_33984 = 6'h26 == _T_3836 ? _T_3372_38_pdst : _GEN_33894;
  assign _GEN_34009 = 6'h26 == _T_3836 ? _T_3372_38_ldst_val : _GEN_33919;
  assign _GEN_34074 = 6'h27 == _T_3836 ? _T_3372_39_pdst : _GEN_33984;
  assign _GEN_34099 = 6'h27 == _T_3836 ? _T_3372_39_ldst_val : _GEN_34009;
  assign _T_5296 = _T_3835 & _GEN_217_ldst_val;
  assign _T_5297 = _GEN_218_pdst != io_wb_resps_2_bits_uop_pdst;
  assign _T_5298 = _T_5296 & _T_5297;
  assign _T_5300 = _T_5298 == 1'h0;
  assign _T_5302 = _T_5300 | reset;
  assign _T_5304 = _T_5302 == 1'h0;
  assign _GEN_34192 = 6'h1 == _T_3845 ? _T_3073_1 : _T_3073_0;
  assign _GEN_34193 = 6'h2 == _T_3845 ? _T_3073_2 : _GEN_34192;
  assign _GEN_34194 = 6'h3 == _T_3845 ? _T_3073_3 : _GEN_34193;
  assign _GEN_34195 = 6'h4 == _T_3845 ? _T_3073_4 : _GEN_34194;
  assign _GEN_34196 = 6'h5 == _T_3845 ? _T_3073_5 : _GEN_34195;
  assign _GEN_34197 = 6'h6 == _T_3845 ? _T_3073_6 : _GEN_34196;
  assign _GEN_34198 = 6'h7 == _T_3845 ? _T_3073_7 : _GEN_34197;
  assign _GEN_34199 = 6'h8 == _T_3845 ? _T_3073_8 : _GEN_34198;
  assign _GEN_34200 = 6'h9 == _T_3845 ? _T_3073_9 : _GEN_34199;
  assign _GEN_34201 = 6'ha == _T_3845 ? _T_3073_10 : _GEN_34200;
  assign _GEN_34202 = 6'hb == _T_3845 ? _T_3073_11 : _GEN_34201;
  assign _GEN_34203 = 6'hc == _T_3845 ? _T_3073_12 : _GEN_34202;
  assign _GEN_34204 = 6'hd == _T_3845 ? _T_3073_13 : _GEN_34203;
  assign _GEN_34205 = 6'he == _T_3845 ? _T_3073_14 : _GEN_34204;
  assign _GEN_34206 = 6'hf == _T_3845 ? _T_3073_15 : _GEN_34205;
  assign _GEN_34207 = 6'h10 == _T_3845 ? _T_3073_16 : _GEN_34206;
  assign _GEN_34208 = 6'h11 == _T_3845 ? _T_3073_17 : _GEN_34207;
  assign _GEN_34209 = 6'h12 == _T_3845 ? _T_3073_18 : _GEN_34208;
  assign _GEN_34210 = 6'h13 == _T_3845 ? _T_3073_19 : _GEN_34209;
  assign _GEN_34211 = 6'h14 == _T_3845 ? _T_3073_20 : _GEN_34210;
  assign _GEN_34212 = 6'h15 == _T_3845 ? _T_3073_21 : _GEN_34211;
  assign _GEN_34213 = 6'h16 == _T_3845 ? _T_3073_22 : _GEN_34212;
  assign _GEN_34214 = 6'h17 == _T_3845 ? _T_3073_23 : _GEN_34213;
  assign _GEN_34215 = 6'h18 == _T_3845 ? _T_3073_24 : _GEN_34214;
  assign _GEN_34216 = 6'h19 == _T_3845 ? _T_3073_25 : _GEN_34215;
  assign _GEN_34217 = 6'h1a == _T_3845 ? _T_3073_26 : _GEN_34216;
  assign _GEN_34218 = 6'h1b == _T_3845 ? _T_3073_27 : _GEN_34217;
  assign _GEN_34219 = 6'h1c == _T_3845 ? _T_3073_28 : _GEN_34218;
  assign _GEN_34220 = 6'h1d == _T_3845 ? _T_3073_29 : _GEN_34219;
  assign _GEN_34221 = 6'h1e == _T_3845 ? _T_3073_30 : _GEN_34220;
  assign _GEN_34222 = 6'h1f == _T_3845 ? _T_3073_31 : _GEN_34221;
  assign _GEN_34223 = 6'h20 == _T_3845 ? _T_3073_32 : _GEN_34222;
  assign _GEN_34224 = 6'h21 == _T_3845 ? _T_3073_33 : _GEN_34223;
  assign _GEN_34225 = 6'h22 == _T_3845 ? _T_3073_34 : _GEN_34224;
  assign _GEN_34226 = 6'h23 == _T_3845 ? _T_3073_35 : _GEN_34225;
  assign _GEN_34227 = 6'h24 == _T_3845 ? _T_3073_36 : _GEN_34226;
  assign _GEN_34228 = 6'h25 == _T_3845 ? _T_3073_37 : _GEN_34227;
  assign _GEN_34229 = 6'h26 == _T_3845 ? _T_3073_38 : _GEN_34228;
  assign _GEN_34230 = 6'h27 == _T_3845 ? _T_3073_39 : _GEN_34229;
  assign _T_5344 = _GEN_220 == 1'h0;
  assign _T_5345 = _T_3844 & _T_5344;
  assign _T_5347 = _T_5345 == 1'h0;
  assign _T_5349 = _T_5347 | reset;
  assign _T_5351 = _T_5349 == 1'h0;
  assign _T_5358 = _T_3840[5:0];
  assign _T_5361 = _T_3200__T_5359_data == 1'h0;
  assign _T_5362 = _T_3844 & _T_5361;
  assign _T_5364 = _T_5362 == 1'h0;
  assign _T_5366 = _T_5364 | reset;
  assign _T_5368 = _T_5366 == 1'h0;
  assign _GEN_34283 = 6'h1 == _T_3845 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_34308 = 6'h1 == _T_3845 ? _T_3372_1_ldst_val : _T_3372_0_ldst_val;
  assign _GEN_34373 = 6'h2 == _T_3845 ? _T_3372_2_pdst : _GEN_34283;
  assign _GEN_34398 = 6'h2 == _T_3845 ? _T_3372_2_ldst_val : _GEN_34308;
  assign _GEN_34463 = 6'h3 == _T_3845 ? _T_3372_3_pdst : _GEN_34373;
  assign _GEN_34488 = 6'h3 == _T_3845 ? _T_3372_3_ldst_val : _GEN_34398;
  assign _GEN_34553 = 6'h4 == _T_3845 ? _T_3372_4_pdst : _GEN_34463;
  assign _GEN_34578 = 6'h4 == _T_3845 ? _T_3372_4_ldst_val : _GEN_34488;
  assign _GEN_34643 = 6'h5 == _T_3845 ? _T_3372_5_pdst : _GEN_34553;
  assign _GEN_34668 = 6'h5 == _T_3845 ? _T_3372_5_ldst_val : _GEN_34578;
  assign _GEN_34733 = 6'h6 == _T_3845 ? _T_3372_6_pdst : _GEN_34643;
  assign _GEN_34758 = 6'h6 == _T_3845 ? _T_3372_6_ldst_val : _GEN_34668;
  assign _GEN_34823 = 6'h7 == _T_3845 ? _T_3372_7_pdst : _GEN_34733;
  assign _GEN_34848 = 6'h7 == _T_3845 ? _T_3372_7_ldst_val : _GEN_34758;
  assign _GEN_34913 = 6'h8 == _T_3845 ? _T_3372_8_pdst : _GEN_34823;
  assign _GEN_34938 = 6'h8 == _T_3845 ? _T_3372_8_ldst_val : _GEN_34848;
  assign _GEN_35003 = 6'h9 == _T_3845 ? _T_3372_9_pdst : _GEN_34913;
  assign _GEN_35028 = 6'h9 == _T_3845 ? _T_3372_9_ldst_val : _GEN_34938;
  assign _GEN_35093 = 6'ha == _T_3845 ? _T_3372_10_pdst : _GEN_35003;
  assign _GEN_35118 = 6'ha == _T_3845 ? _T_3372_10_ldst_val : _GEN_35028;
  assign _GEN_35183 = 6'hb == _T_3845 ? _T_3372_11_pdst : _GEN_35093;
  assign _GEN_35208 = 6'hb == _T_3845 ? _T_3372_11_ldst_val : _GEN_35118;
  assign _GEN_35273 = 6'hc == _T_3845 ? _T_3372_12_pdst : _GEN_35183;
  assign _GEN_35298 = 6'hc == _T_3845 ? _T_3372_12_ldst_val : _GEN_35208;
  assign _GEN_35363 = 6'hd == _T_3845 ? _T_3372_13_pdst : _GEN_35273;
  assign _GEN_35388 = 6'hd == _T_3845 ? _T_3372_13_ldst_val : _GEN_35298;
  assign _GEN_35453 = 6'he == _T_3845 ? _T_3372_14_pdst : _GEN_35363;
  assign _GEN_35478 = 6'he == _T_3845 ? _T_3372_14_ldst_val : _GEN_35388;
  assign _GEN_35543 = 6'hf == _T_3845 ? _T_3372_15_pdst : _GEN_35453;
  assign _GEN_35568 = 6'hf == _T_3845 ? _T_3372_15_ldst_val : _GEN_35478;
  assign _GEN_35633 = 6'h10 == _T_3845 ? _T_3372_16_pdst : _GEN_35543;
  assign _GEN_35658 = 6'h10 == _T_3845 ? _T_3372_16_ldst_val : _GEN_35568;
  assign _GEN_35723 = 6'h11 == _T_3845 ? _T_3372_17_pdst : _GEN_35633;
  assign _GEN_35748 = 6'h11 == _T_3845 ? _T_3372_17_ldst_val : _GEN_35658;
  assign _GEN_35813 = 6'h12 == _T_3845 ? _T_3372_18_pdst : _GEN_35723;
  assign _GEN_35838 = 6'h12 == _T_3845 ? _T_3372_18_ldst_val : _GEN_35748;
  assign _GEN_35903 = 6'h13 == _T_3845 ? _T_3372_19_pdst : _GEN_35813;
  assign _GEN_35928 = 6'h13 == _T_3845 ? _T_3372_19_ldst_val : _GEN_35838;
  assign _GEN_35993 = 6'h14 == _T_3845 ? _T_3372_20_pdst : _GEN_35903;
  assign _GEN_36018 = 6'h14 == _T_3845 ? _T_3372_20_ldst_val : _GEN_35928;
  assign _GEN_36083 = 6'h15 == _T_3845 ? _T_3372_21_pdst : _GEN_35993;
  assign _GEN_36108 = 6'h15 == _T_3845 ? _T_3372_21_ldst_val : _GEN_36018;
  assign _GEN_36173 = 6'h16 == _T_3845 ? _T_3372_22_pdst : _GEN_36083;
  assign _GEN_36198 = 6'h16 == _T_3845 ? _T_3372_22_ldst_val : _GEN_36108;
  assign _GEN_36263 = 6'h17 == _T_3845 ? _T_3372_23_pdst : _GEN_36173;
  assign _GEN_36288 = 6'h17 == _T_3845 ? _T_3372_23_ldst_val : _GEN_36198;
  assign _GEN_36353 = 6'h18 == _T_3845 ? _T_3372_24_pdst : _GEN_36263;
  assign _GEN_36378 = 6'h18 == _T_3845 ? _T_3372_24_ldst_val : _GEN_36288;
  assign _GEN_36443 = 6'h19 == _T_3845 ? _T_3372_25_pdst : _GEN_36353;
  assign _GEN_36468 = 6'h19 == _T_3845 ? _T_3372_25_ldst_val : _GEN_36378;
  assign _GEN_36533 = 6'h1a == _T_3845 ? _T_3372_26_pdst : _GEN_36443;
  assign _GEN_36558 = 6'h1a == _T_3845 ? _T_3372_26_ldst_val : _GEN_36468;
  assign _GEN_36623 = 6'h1b == _T_3845 ? _T_3372_27_pdst : _GEN_36533;
  assign _GEN_36648 = 6'h1b == _T_3845 ? _T_3372_27_ldst_val : _GEN_36558;
  assign _GEN_36713 = 6'h1c == _T_3845 ? _T_3372_28_pdst : _GEN_36623;
  assign _GEN_36738 = 6'h1c == _T_3845 ? _T_3372_28_ldst_val : _GEN_36648;
  assign _GEN_36803 = 6'h1d == _T_3845 ? _T_3372_29_pdst : _GEN_36713;
  assign _GEN_36828 = 6'h1d == _T_3845 ? _T_3372_29_ldst_val : _GEN_36738;
  assign _GEN_36893 = 6'h1e == _T_3845 ? _T_3372_30_pdst : _GEN_36803;
  assign _GEN_36918 = 6'h1e == _T_3845 ? _T_3372_30_ldst_val : _GEN_36828;
  assign _GEN_36983 = 6'h1f == _T_3845 ? _T_3372_31_pdst : _GEN_36893;
  assign _GEN_37008 = 6'h1f == _T_3845 ? _T_3372_31_ldst_val : _GEN_36918;
  assign _GEN_37073 = 6'h20 == _T_3845 ? _T_3372_32_pdst : _GEN_36983;
  assign _GEN_37098 = 6'h20 == _T_3845 ? _T_3372_32_ldst_val : _GEN_37008;
  assign _GEN_37163 = 6'h21 == _T_3845 ? _T_3372_33_pdst : _GEN_37073;
  assign _GEN_37188 = 6'h21 == _T_3845 ? _T_3372_33_ldst_val : _GEN_37098;
  assign _GEN_37253 = 6'h22 == _T_3845 ? _T_3372_34_pdst : _GEN_37163;
  assign _GEN_37278 = 6'h22 == _T_3845 ? _T_3372_34_ldst_val : _GEN_37188;
  assign _GEN_37343 = 6'h23 == _T_3845 ? _T_3372_35_pdst : _GEN_37253;
  assign _GEN_37368 = 6'h23 == _T_3845 ? _T_3372_35_ldst_val : _GEN_37278;
  assign _GEN_37433 = 6'h24 == _T_3845 ? _T_3372_36_pdst : _GEN_37343;
  assign _GEN_37458 = 6'h24 == _T_3845 ? _T_3372_36_ldst_val : _GEN_37368;
  assign _GEN_37523 = 6'h25 == _T_3845 ? _T_3372_37_pdst : _GEN_37433;
  assign _GEN_37548 = 6'h25 == _T_3845 ? _T_3372_37_ldst_val : _GEN_37458;
  assign _GEN_37613 = 6'h26 == _T_3845 ? _T_3372_38_pdst : _GEN_37523;
  assign _GEN_37638 = 6'h26 == _T_3845 ? _T_3372_38_ldst_val : _GEN_37548;
  assign _GEN_37703 = 6'h27 == _T_3845 ? _T_3372_39_pdst : _GEN_37613;
  assign _GEN_37728 = 6'h27 == _T_3845 ? _T_3372_39_ldst_val : _GEN_37638;
  assign _T_5373 = _T_3844 & _GEN_221_ldst_val;
  assign _T_5374 = _GEN_222_pdst != io_wb_resps_3_bits_uop_pdst;
  assign _T_5375 = _T_5373 & _T_5374;
  assign _T_5377 = _T_5375 == 1'h0;
  assign _T_5379 = _T_5377 | reset;
  assign _T_5381 = _T_5379 == 1'h0;
  assign _GEN_37821 = 6'h1 == _T_3854 ? _T_3073_1 : _T_3073_0;
  assign _GEN_37822 = 6'h2 == _T_3854 ? _T_3073_2 : _GEN_37821;
  assign _GEN_37823 = 6'h3 == _T_3854 ? _T_3073_3 : _GEN_37822;
  assign _GEN_37824 = 6'h4 == _T_3854 ? _T_3073_4 : _GEN_37823;
  assign _GEN_37825 = 6'h5 == _T_3854 ? _T_3073_5 : _GEN_37824;
  assign _GEN_37826 = 6'h6 == _T_3854 ? _T_3073_6 : _GEN_37825;
  assign _GEN_37827 = 6'h7 == _T_3854 ? _T_3073_7 : _GEN_37826;
  assign _GEN_37828 = 6'h8 == _T_3854 ? _T_3073_8 : _GEN_37827;
  assign _GEN_37829 = 6'h9 == _T_3854 ? _T_3073_9 : _GEN_37828;
  assign _GEN_37830 = 6'ha == _T_3854 ? _T_3073_10 : _GEN_37829;
  assign _GEN_37831 = 6'hb == _T_3854 ? _T_3073_11 : _GEN_37830;
  assign _GEN_37832 = 6'hc == _T_3854 ? _T_3073_12 : _GEN_37831;
  assign _GEN_37833 = 6'hd == _T_3854 ? _T_3073_13 : _GEN_37832;
  assign _GEN_37834 = 6'he == _T_3854 ? _T_3073_14 : _GEN_37833;
  assign _GEN_37835 = 6'hf == _T_3854 ? _T_3073_15 : _GEN_37834;
  assign _GEN_37836 = 6'h10 == _T_3854 ? _T_3073_16 : _GEN_37835;
  assign _GEN_37837 = 6'h11 == _T_3854 ? _T_3073_17 : _GEN_37836;
  assign _GEN_37838 = 6'h12 == _T_3854 ? _T_3073_18 : _GEN_37837;
  assign _GEN_37839 = 6'h13 == _T_3854 ? _T_3073_19 : _GEN_37838;
  assign _GEN_37840 = 6'h14 == _T_3854 ? _T_3073_20 : _GEN_37839;
  assign _GEN_37841 = 6'h15 == _T_3854 ? _T_3073_21 : _GEN_37840;
  assign _GEN_37842 = 6'h16 == _T_3854 ? _T_3073_22 : _GEN_37841;
  assign _GEN_37843 = 6'h17 == _T_3854 ? _T_3073_23 : _GEN_37842;
  assign _GEN_37844 = 6'h18 == _T_3854 ? _T_3073_24 : _GEN_37843;
  assign _GEN_37845 = 6'h19 == _T_3854 ? _T_3073_25 : _GEN_37844;
  assign _GEN_37846 = 6'h1a == _T_3854 ? _T_3073_26 : _GEN_37845;
  assign _GEN_37847 = 6'h1b == _T_3854 ? _T_3073_27 : _GEN_37846;
  assign _GEN_37848 = 6'h1c == _T_3854 ? _T_3073_28 : _GEN_37847;
  assign _GEN_37849 = 6'h1d == _T_3854 ? _T_3073_29 : _GEN_37848;
  assign _GEN_37850 = 6'h1e == _T_3854 ? _T_3073_30 : _GEN_37849;
  assign _GEN_37851 = 6'h1f == _T_3854 ? _T_3073_31 : _GEN_37850;
  assign _GEN_37852 = 6'h20 == _T_3854 ? _T_3073_32 : _GEN_37851;
  assign _GEN_37853 = 6'h21 == _T_3854 ? _T_3073_33 : _GEN_37852;
  assign _GEN_37854 = 6'h22 == _T_3854 ? _T_3073_34 : _GEN_37853;
  assign _GEN_37855 = 6'h23 == _T_3854 ? _T_3073_35 : _GEN_37854;
  assign _GEN_37856 = 6'h24 == _T_3854 ? _T_3073_36 : _GEN_37855;
  assign _GEN_37857 = 6'h25 == _T_3854 ? _T_3073_37 : _GEN_37856;
  assign _GEN_37858 = 6'h26 == _T_3854 ? _T_3073_38 : _GEN_37857;
  assign _GEN_37859 = 6'h27 == _T_3854 ? _T_3073_39 : _GEN_37858;
  assign _T_5421 = _GEN_224 == 1'h0;
  assign _T_5422 = _T_3853 & _T_5421;
  assign _T_5424 = _T_5422 == 1'h0;
  assign _T_5426 = _T_5424 | reset;
  assign _T_5428 = _T_5426 == 1'h0;
  assign _T_5435 = _T_3849[5:0];
  assign _T_5438 = _T_3200__T_5436_data == 1'h0;
  assign _T_5439 = _T_3853 & _T_5438;
  assign _T_5441 = _T_5439 == 1'h0;
  assign _T_5443 = _T_5441 | reset;
  assign _T_5445 = _T_5443 == 1'h0;
  assign _GEN_37912 = 6'h1 == _T_3854 ? _T_3372_1_pdst : _T_3372_0_pdst;
  assign _GEN_37937 = 6'h1 == _T_3854 ? _T_3372_1_ldst_val : _T_3372_0_ldst_val;
  assign _GEN_38002 = 6'h2 == _T_3854 ? _T_3372_2_pdst : _GEN_37912;
  assign _GEN_38027 = 6'h2 == _T_3854 ? _T_3372_2_ldst_val : _GEN_37937;
  assign _GEN_38092 = 6'h3 == _T_3854 ? _T_3372_3_pdst : _GEN_38002;
  assign _GEN_38117 = 6'h3 == _T_3854 ? _T_3372_3_ldst_val : _GEN_38027;
  assign _GEN_38182 = 6'h4 == _T_3854 ? _T_3372_4_pdst : _GEN_38092;
  assign _GEN_38207 = 6'h4 == _T_3854 ? _T_3372_4_ldst_val : _GEN_38117;
  assign _GEN_38272 = 6'h5 == _T_3854 ? _T_3372_5_pdst : _GEN_38182;
  assign _GEN_38297 = 6'h5 == _T_3854 ? _T_3372_5_ldst_val : _GEN_38207;
  assign _GEN_38362 = 6'h6 == _T_3854 ? _T_3372_6_pdst : _GEN_38272;
  assign _GEN_38387 = 6'h6 == _T_3854 ? _T_3372_6_ldst_val : _GEN_38297;
  assign _GEN_38452 = 6'h7 == _T_3854 ? _T_3372_7_pdst : _GEN_38362;
  assign _GEN_38477 = 6'h7 == _T_3854 ? _T_3372_7_ldst_val : _GEN_38387;
  assign _GEN_38542 = 6'h8 == _T_3854 ? _T_3372_8_pdst : _GEN_38452;
  assign _GEN_38567 = 6'h8 == _T_3854 ? _T_3372_8_ldst_val : _GEN_38477;
  assign _GEN_38632 = 6'h9 == _T_3854 ? _T_3372_9_pdst : _GEN_38542;
  assign _GEN_38657 = 6'h9 == _T_3854 ? _T_3372_9_ldst_val : _GEN_38567;
  assign _GEN_38722 = 6'ha == _T_3854 ? _T_3372_10_pdst : _GEN_38632;
  assign _GEN_38747 = 6'ha == _T_3854 ? _T_3372_10_ldst_val : _GEN_38657;
  assign _GEN_38812 = 6'hb == _T_3854 ? _T_3372_11_pdst : _GEN_38722;
  assign _GEN_38837 = 6'hb == _T_3854 ? _T_3372_11_ldst_val : _GEN_38747;
  assign _GEN_38902 = 6'hc == _T_3854 ? _T_3372_12_pdst : _GEN_38812;
  assign _GEN_38927 = 6'hc == _T_3854 ? _T_3372_12_ldst_val : _GEN_38837;
  assign _GEN_38992 = 6'hd == _T_3854 ? _T_3372_13_pdst : _GEN_38902;
  assign _GEN_39017 = 6'hd == _T_3854 ? _T_3372_13_ldst_val : _GEN_38927;
  assign _GEN_39082 = 6'he == _T_3854 ? _T_3372_14_pdst : _GEN_38992;
  assign _GEN_39107 = 6'he == _T_3854 ? _T_3372_14_ldst_val : _GEN_39017;
  assign _GEN_39172 = 6'hf == _T_3854 ? _T_3372_15_pdst : _GEN_39082;
  assign _GEN_39197 = 6'hf == _T_3854 ? _T_3372_15_ldst_val : _GEN_39107;
  assign _GEN_39262 = 6'h10 == _T_3854 ? _T_3372_16_pdst : _GEN_39172;
  assign _GEN_39287 = 6'h10 == _T_3854 ? _T_3372_16_ldst_val : _GEN_39197;
  assign _GEN_39352 = 6'h11 == _T_3854 ? _T_3372_17_pdst : _GEN_39262;
  assign _GEN_39377 = 6'h11 == _T_3854 ? _T_3372_17_ldst_val : _GEN_39287;
  assign _GEN_39442 = 6'h12 == _T_3854 ? _T_3372_18_pdst : _GEN_39352;
  assign _GEN_39467 = 6'h12 == _T_3854 ? _T_3372_18_ldst_val : _GEN_39377;
  assign _GEN_39532 = 6'h13 == _T_3854 ? _T_3372_19_pdst : _GEN_39442;
  assign _GEN_39557 = 6'h13 == _T_3854 ? _T_3372_19_ldst_val : _GEN_39467;
  assign _GEN_39622 = 6'h14 == _T_3854 ? _T_3372_20_pdst : _GEN_39532;
  assign _GEN_39647 = 6'h14 == _T_3854 ? _T_3372_20_ldst_val : _GEN_39557;
  assign _GEN_39712 = 6'h15 == _T_3854 ? _T_3372_21_pdst : _GEN_39622;
  assign _GEN_39737 = 6'h15 == _T_3854 ? _T_3372_21_ldst_val : _GEN_39647;
  assign _GEN_39802 = 6'h16 == _T_3854 ? _T_3372_22_pdst : _GEN_39712;
  assign _GEN_39827 = 6'h16 == _T_3854 ? _T_3372_22_ldst_val : _GEN_39737;
  assign _GEN_39892 = 6'h17 == _T_3854 ? _T_3372_23_pdst : _GEN_39802;
  assign _GEN_39917 = 6'h17 == _T_3854 ? _T_3372_23_ldst_val : _GEN_39827;
  assign _GEN_39982 = 6'h18 == _T_3854 ? _T_3372_24_pdst : _GEN_39892;
  assign _GEN_40007 = 6'h18 == _T_3854 ? _T_3372_24_ldst_val : _GEN_39917;
  assign _GEN_40072 = 6'h19 == _T_3854 ? _T_3372_25_pdst : _GEN_39982;
  assign _GEN_40097 = 6'h19 == _T_3854 ? _T_3372_25_ldst_val : _GEN_40007;
  assign _GEN_40162 = 6'h1a == _T_3854 ? _T_3372_26_pdst : _GEN_40072;
  assign _GEN_40187 = 6'h1a == _T_3854 ? _T_3372_26_ldst_val : _GEN_40097;
  assign _GEN_40252 = 6'h1b == _T_3854 ? _T_3372_27_pdst : _GEN_40162;
  assign _GEN_40277 = 6'h1b == _T_3854 ? _T_3372_27_ldst_val : _GEN_40187;
  assign _GEN_40342 = 6'h1c == _T_3854 ? _T_3372_28_pdst : _GEN_40252;
  assign _GEN_40367 = 6'h1c == _T_3854 ? _T_3372_28_ldst_val : _GEN_40277;
  assign _GEN_40432 = 6'h1d == _T_3854 ? _T_3372_29_pdst : _GEN_40342;
  assign _GEN_40457 = 6'h1d == _T_3854 ? _T_3372_29_ldst_val : _GEN_40367;
  assign _GEN_40522 = 6'h1e == _T_3854 ? _T_3372_30_pdst : _GEN_40432;
  assign _GEN_40547 = 6'h1e == _T_3854 ? _T_3372_30_ldst_val : _GEN_40457;
  assign _GEN_40612 = 6'h1f == _T_3854 ? _T_3372_31_pdst : _GEN_40522;
  assign _GEN_40637 = 6'h1f == _T_3854 ? _T_3372_31_ldst_val : _GEN_40547;
  assign _GEN_40702 = 6'h20 == _T_3854 ? _T_3372_32_pdst : _GEN_40612;
  assign _GEN_40727 = 6'h20 == _T_3854 ? _T_3372_32_ldst_val : _GEN_40637;
  assign _GEN_40792 = 6'h21 == _T_3854 ? _T_3372_33_pdst : _GEN_40702;
  assign _GEN_40817 = 6'h21 == _T_3854 ? _T_3372_33_ldst_val : _GEN_40727;
  assign _GEN_40882 = 6'h22 == _T_3854 ? _T_3372_34_pdst : _GEN_40792;
  assign _GEN_40907 = 6'h22 == _T_3854 ? _T_3372_34_ldst_val : _GEN_40817;
  assign _GEN_40972 = 6'h23 == _T_3854 ? _T_3372_35_pdst : _GEN_40882;
  assign _GEN_40997 = 6'h23 == _T_3854 ? _T_3372_35_ldst_val : _GEN_40907;
  assign _GEN_41062 = 6'h24 == _T_3854 ? _T_3372_36_pdst : _GEN_40972;
  assign _GEN_41087 = 6'h24 == _T_3854 ? _T_3372_36_ldst_val : _GEN_40997;
  assign _GEN_41152 = 6'h25 == _T_3854 ? _T_3372_37_pdst : _GEN_41062;
  assign _GEN_41177 = 6'h25 == _T_3854 ? _T_3372_37_ldst_val : _GEN_41087;
  assign _GEN_41242 = 6'h26 == _T_3854 ? _T_3372_38_pdst : _GEN_41152;
  assign _GEN_41267 = 6'h26 == _T_3854 ? _T_3372_38_ldst_val : _GEN_41177;
  assign _GEN_41332 = 6'h27 == _T_3854 ? _T_3372_39_pdst : _GEN_41242;
  assign _GEN_41357 = 6'h27 == _T_3854 ? _T_3372_39_ldst_val : _GEN_41267;
  assign _T_5450 = _T_3853 & _GEN_225_ldst_val;
  assign _T_5451 = _GEN_226_pdst != io_wb_resps_4_bits_uop_pdst;
  assign _T_5452 = _T_5450 & _T_5451;
  assign _T_5454 = _T_5452 == 1'h0;
  assign _T_5456 = _T_5454 | reset;
  assign _T_5458 = _T_5456 == 1'h0;
  assign _T_5764__T_6441_addr = _T_6440;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6441_data = _T_5764[_T_5764__T_6441_addr];
  `else
  assign _T_5764__T_6441_data = _T_5764__T_6441_addr >= 6'h28 ? _RAND_594[0:0] : _T_5764[_T_5764__T_6441_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6468_addr = _T_6467;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6468_data = _T_5764[_T_5764__T_6468_addr];
  `else
  assign _T_5764__T_6468_data = _T_5764__T_6468_addr >= 6'h28 ? _RAND_595[0:0] : _T_5764[_T_5764__T_6468_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6581_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6581_data = _T_5764[_T_5764__T_6581_addr];
  `else
  assign _T_5764__T_6581_data = _T_5764__T_6581_addr >= 6'h28 ? _RAND_596[0:0] : _T_5764[_T_5764__T_6581_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7692_addr = _T_7691;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7692_data = _T_5764[_T_5764__T_7692_addr];
  `else
  assign _T_5764__T_7692_data = _T_5764__T_7692_addr >= 6'h28 ? _RAND_597[0:0] : _T_5764[_T_5764__T_7692_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7769_addr = _T_7768;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7769_data = _T_5764[_T_5764__T_7769_addr];
  `else
  assign _T_5764__T_7769_data = _T_5764__T_7769_addr >= 6'h28 ? _RAND_598[0:0] : _T_5764[_T_5764__T_7769_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7846_addr = _T_7845;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7846_data = _T_5764[_T_5764__T_7846_addr];
  `else
  assign _T_5764__T_7846_data = _T_5764__T_7846_addr >= 6'h28 ? _RAND_599[0:0] : _T_5764[_T_5764__T_7846_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7923_addr = _T_7922;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_7923_data = _T_5764[_T_5764__T_7923_addr];
  `else
  assign _T_5764__T_7923_data = _T_5764__T_7923_addr >= 6'h28 ? _RAND_600[0:0] : _T_5764[_T_5764__T_7923_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_8000_addr = _T_7999;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_8000_data = _T_5764[_T_5764__T_8000_addr];
  `else
  assign _T_5764__T_8000_data = _T_5764__T_8000_addr >= 6'h28 ? _RAND_601[0:0] : _T_5764[_T_5764__T_8000_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5764__T_6317_data = _T_6322;
  assign _T_5764__T_6317_addr = rob_tail;
  assign _T_5764__T_6317_mask = io_enq_valids_1;
  assign _T_5764__T_6317_en = io_enq_valids_1;
  assign _T_5764__T_6383_data = 1'h0;
  assign _T_5764__T_6383_addr = _T_6382;
  assign _T_5764__T_6383_mask = _T_6381;
  assign _T_5764__T_6383_en = _T_6381;
  assign _T_5764__T_6392_data = 1'h0;
  assign _T_5764__T_6392_addr = _T_6391;
  assign _T_5764__T_6392_mask = _T_6390;
  assign _T_5764__T_6392_en = _T_6390;
  assign _T_5764__T_6401_data = 1'h0;
  assign _T_5764__T_6401_addr = _T_6400;
  assign _T_5764__T_6401_mask = _T_6399;
  assign _T_5764__T_6401_en = _T_6399;
  assign _T_5764__T_6410_data = 1'h0;
  assign _T_5764__T_6410_addr = _T_6409;
  assign _T_5764__T_6410_mask = _T_6408;
  assign _T_5764__T_6410_en = _T_6408;
  assign _T_5764__T_6419_data = 1'h0;
  assign _T_5764__T_6419_addr = _T_6418;
  assign _T_5764__T_6419_mask = _T_6417;
  assign _T_5764__T_6419_en = _T_6417;
  assign _T_5764__T_6428_data = 1'h0;
  assign _T_5764__T_6428_addr = _T_6427;
  assign _T_5764__T_6428_mask = _T_6424;
  assign _T_5764__T_6428_en = _T_6424;
  assign _T_5764__T_6455_data = 1'h0;
  assign _T_5764__T_6455_addr = _T_6454;
  assign _T_5764__T_6455_mask = _T_6451;
  assign _T_5764__T_6455_en = _T_6451;
  assign _T_6309__T_6576_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6309__T_6576_data = _T_6309[_T_6309__T_6576_addr];
  `else
  assign _T_6309__T_6576_data = _T_6309__T_6576_addr >= 6'h28 ? _RAND_1083[0:0] : _T_6309[_T_6309__T_6576_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6309__T_6332_data = io_enq_uops_1_exception;
  assign _T_6309__T_6332_addr = rob_tail;
  assign _T_6309__T_6332_mask = io_enq_valids_1;
  assign _T_6309__T_6332_en = io_enq_valids_1;
  assign _T_6309__T_6562_data = 1'h1;
  assign _T_6309__T_6562_addr = _T_6561;
  assign _T_6309__T_6562_mask = _T_6558;
  assign _T_6309__T_6562_en = _T_6558;
  assign _T_6309__T_6571_data = 1'h1;
  assign _T_6309__T_6571_addr = _T_6570;
  assign _T_6309__T_6571_mask = _T_6567;
  assign _T_6309__T_6571_en = _T_6567;
  assign _T_6309__T_6652_data = 1'h0;
  assign _T_6309__T_6652_addr = _T_6589;
  assign _T_6309__T_6652_mask = _T_6641;
  assign _T_6309__T_6652_en = _T_6641;
  assign _T_6312__T_7581_addr = rob_head;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6312__T_7581_data = _T_6312[_T_6312__T_7581_addr];
  `else
  assign _T_6312__T_7581_data = _T_6312__T_7581_addr >= 6'h28 ? _RAND_1085[4:0] : _T_6312[_T_6312__T_7581_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6312__T_6333_data = 5'h0;
  assign _T_6312__T_6333_addr = rob_tail;
  assign _T_6312__T_6333_mask = io_enq_valids_1;
  assign _T_6312__T_6333_en = io_enq_valids_1;
  assign _T_6312__T_6546_data = io_fflags_0_bits_flags;
  assign _T_6312__T_6546_addr = _T_6545;
  assign _T_6312__T_6546_mask = _T_6542;
  assign _T_6312__T_6546_en = _T_6542;
  assign _T_6312__T_6554_data = io_fflags_1_bits_flags;
  assign _T_6312__T_6554_addr = _T_6553;
  assign _T_6312__T_6554_mask = _T_6550;
  assign _T_6312__T_6554_en = _T_6550;
  assign _GEN_41370 = 6'h0 == rob_tail ? 1'h1 : _T_5637_0;
  assign _GEN_41371 = 6'h1 == rob_tail ? 1'h1 : _T_5637_1;
  assign _GEN_41372 = 6'h2 == rob_tail ? 1'h1 : _T_5637_2;
  assign _GEN_41373 = 6'h3 == rob_tail ? 1'h1 : _T_5637_3;
  assign _GEN_41374 = 6'h4 == rob_tail ? 1'h1 : _T_5637_4;
  assign _GEN_41375 = 6'h5 == rob_tail ? 1'h1 : _T_5637_5;
  assign _GEN_41376 = 6'h6 == rob_tail ? 1'h1 : _T_5637_6;
  assign _GEN_41377 = 6'h7 == rob_tail ? 1'h1 : _T_5637_7;
  assign _GEN_41378 = 6'h8 == rob_tail ? 1'h1 : _T_5637_8;
  assign _GEN_41379 = 6'h9 == rob_tail ? 1'h1 : _T_5637_9;
  assign _GEN_41380 = 6'ha == rob_tail ? 1'h1 : _T_5637_10;
  assign _GEN_41381 = 6'hb == rob_tail ? 1'h1 : _T_5637_11;
  assign _GEN_41382 = 6'hc == rob_tail ? 1'h1 : _T_5637_12;
  assign _GEN_41383 = 6'hd == rob_tail ? 1'h1 : _T_5637_13;
  assign _GEN_41384 = 6'he == rob_tail ? 1'h1 : _T_5637_14;
  assign _GEN_41385 = 6'hf == rob_tail ? 1'h1 : _T_5637_15;
  assign _GEN_41386 = 6'h10 == rob_tail ? 1'h1 : _T_5637_16;
  assign _GEN_41387 = 6'h11 == rob_tail ? 1'h1 : _T_5637_17;
  assign _GEN_41388 = 6'h12 == rob_tail ? 1'h1 : _T_5637_18;
  assign _GEN_41389 = 6'h13 == rob_tail ? 1'h1 : _T_5637_19;
  assign _GEN_41390 = 6'h14 == rob_tail ? 1'h1 : _T_5637_20;
  assign _GEN_41391 = 6'h15 == rob_tail ? 1'h1 : _T_5637_21;
  assign _GEN_41392 = 6'h16 == rob_tail ? 1'h1 : _T_5637_22;
  assign _GEN_41393 = 6'h17 == rob_tail ? 1'h1 : _T_5637_23;
  assign _GEN_41394 = 6'h18 == rob_tail ? 1'h1 : _T_5637_24;
  assign _GEN_41395 = 6'h19 == rob_tail ? 1'h1 : _T_5637_25;
  assign _GEN_41396 = 6'h1a == rob_tail ? 1'h1 : _T_5637_26;
  assign _GEN_41397 = 6'h1b == rob_tail ? 1'h1 : _T_5637_27;
  assign _GEN_41398 = 6'h1c == rob_tail ? 1'h1 : _T_5637_28;
  assign _GEN_41399 = 6'h1d == rob_tail ? 1'h1 : _T_5637_29;
  assign _GEN_41400 = 6'h1e == rob_tail ? 1'h1 : _T_5637_30;
  assign _GEN_41401 = 6'h1f == rob_tail ? 1'h1 : _T_5637_31;
  assign _GEN_41402 = 6'h20 == rob_tail ? 1'h1 : _T_5637_32;
  assign _GEN_41403 = 6'h21 == rob_tail ? 1'h1 : _T_5637_33;
  assign _GEN_41404 = 6'h22 == rob_tail ? 1'h1 : _T_5637_34;
  assign _GEN_41405 = 6'h23 == rob_tail ? 1'h1 : _T_5637_35;
  assign _GEN_41406 = 6'h24 == rob_tail ? 1'h1 : _T_5637_36;
  assign _GEN_41407 = 6'h25 == rob_tail ? 1'h1 : _T_5637_37;
  assign _GEN_41408 = 6'h26 == rob_tail ? 1'h1 : _T_5637_38;
  assign _GEN_41409 = 6'h27 == rob_tail ? 1'h1 : _T_5637_39;
  assign _T_6319 = io_enq_uops_1_is_fence == 1'h0;
  assign _T_6321 = io_enq_uops_1_is_fencei == 1'h0;
  assign _T_6322 = _T_6319 & _T_6321;
  assign _GEN_42370 = 6'h0 == rob_tail ? _GEN_253 : _T_5936_0_br_mask;
  assign _GEN_42371 = 6'h1 == rob_tail ? _GEN_253 : _T_5936_1_br_mask;
  assign _GEN_42372 = 6'h2 == rob_tail ? _GEN_253 : _T_5936_2_br_mask;
  assign _GEN_42373 = 6'h3 == rob_tail ? _GEN_253 : _T_5936_3_br_mask;
  assign _GEN_42374 = 6'h4 == rob_tail ? _GEN_253 : _T_5936_4_br_mask;
  assign _GEN_42375 = 6'h5 == rob_tail ? _GEN_253 : _T_5936_5_br_mask;
  assign _GEN_42376 = 6'h6 == rob_tail ? _GEN_253 : _T_5936_6_br_mask;
  assign _GEN_42377 = 6'h7 == rob_tail ? _GEN_253 : _T_5936_7_br_mask;
  assign _GEN_42378 = 6'h8 == rob_tail ? _GEN_253 : _T_5936_8_br_mask;
  assign _GEN_42379 = 6'h9 == rob_tail ? _GEN_253 : _T_5936_9_br_mask;
  assign _GEN_42380 = 6'ha == rob_tail ? _GEN_253 : _T_5936_10_br_mask;
  assign _GEN_42381 = 6'hb == rob_tail ? _GEN_253 : _T_5936_11_br_mask;
  assign _GEN_42382 = 6'hc == rob_tail ? _GEN_253 : _T_5936_12_br_mask;
  assign _GEN_42383 = 6'hd == rob_tail ? _GEN_253 : _T_5936_13_br_mask;
  assign _GEN_42384 = 6'he == rob_tail ? _GEN_253 : _T_5936_14_br_mask;
  assign _GEN_42385 = 6'hf == rob_tail ? _GEN_253 : _T_5936_15_br_mask;
  assign _GEN_42386 = 6'h10 == rob_tail ? _GEN_253 : _T_5936_16_br_mask;
  assign _GEN_42387 = 6'h11 == rob_tail ? _GEN_253 : _T_5936_17_br_mask;
  assign _GEN_42388 = 6'h12 == rob_tail ? _GEN_253 : _T_5936_18_br_mask;
  assign _GEN_42389 = 6'h13 == rob_tail ? _GEN_253 : _T_5936_19_br_mask;
  assign _GEN_42390 = 6'h14 == rob_tail ? _GEN_253 : _T_5936_20_br_mask;
  assign _GEN_42391 = 6'h15 == rob_tail ? _GEN_253 : _T_5936_21_br_mask;
  assign _GEN_42392 = 6'h16 == rob_tail ? _GEN_253 : _T_5936_22_br_mask;
  assign _GEN_42393 = 6'h17 == rob_tail ? _GEN_253 : _T_5936_23_br_mask;
  assign _GEN_42394 = 6'h18 == rob_tail ? _GEN_253 : _T_5936_24_br_mask;
  assign _GEN_42395 = 6'h19 == rob_tail ? _GEN_253 : _T_5936_25_br_mask;
  assign _GEN_42396 = 6'h1a == rob_tail ? _GEN_253 : _T_5936_26_br_mask;
  assign _GEN_42397 = 6'h1b == rob_tail ? _GEN_253 : _T_5936_27_br_mask;
  assign _GEN_42398 = 6'h1c == rob_tail ? _GEN_253 : _T_5936_28_br_mask;
  assign _GEN_42399 = 6'h1d == rob_tail ? _GEN_253 : _T_5936_29_br_mask;
  assign _GEN_42400 = 6'h1e == rob_tail ? _GEN_253 : _T_5936_30_br_mask;
  assign _GEN_42401 = 6'h1f == rob_tail ? _GEN_253 : _T_5936_31_br_mask;
  assign _GEN_42402 = 6'h20 == rob_tail ? _GEN_253 : _T_5936_32_br_mask;
  assign _GEN_42403 = 6'h21 == rob_tail ? _GEN_253 : _T_5936_33_br_mask;
  assign _GEN_42404 = 6'h22 == rob_tail ? _GEN_253 : _T_5936_34_br_mask;
  assign _GEN_42405 = 6'h23 == rob_tail ? _GEN_253 : _T_5936_35_br_mask;
  assign _GEN_42406 = 6'h24 == rob_tail ? _GEN_253 : _T_5936_36_br_mask;
  assign _GEN_42407 = 6'h25 == rob_tail ? _GEN_253 : _T_5936_37_br_mask;
  assign _GEN_42408 = 6'h26 == rob_tail ? _GEN_253 : _T_5936_38_br_mask;
  assign _GEN_42409 = 6'h27 == rob_tail ? _GEN_253 : _T_5936_39_br_mask;
  assign _GEN_43490 = 6'h0 == rob_tail ? _GEN_281 : _T_5936_0_pdst;
  assign _GEN_43491 = 6'h1 == rob_tail ? _GEN_281 : _T_5936_1_pdst;
  assign _GEN_43492 = 6'h2 == rob_tail ? _GEN_281 : _T_5936_2_pdst;
  assign _GEN_43493 = 6'h3 == rob_tail ? _GEN_281 : _T_5936_3_pdst;
  assign _GEN_43494 = 6'h4 == rob_tail ? _GEN_281 : _T_5936_4_pdst;
  assign _GEN_43495 = 6'h5 == rob_tail ? _GEN_281 : _T_5936_5_pdst;
  assign _GEN_43496 = 6'h6 == rob_tail ? _GEN_281 : _T_5936_6_pdst;
  assign _GEN_43497 = 6'h7 == rob_tail ? _GEN_281 : _T_5936_7_pdst;
  assign _GEN_43498 = 6'h8 == rob_tail ? _GEN_281 : _T_5936_8_pdst;
  assign _GEN_43499 = 6'h9 == rob_tail ? _GEN_281 : _T_5936_9_pdst;
  assign _GEN_43500 = 6'ha == rob_tail ? _GEN_281 : _T_5936_10_pdst;
  assign _GEN_43501 = 6'hb == rob_tail ? _GEN_281 : _T_5936_11_pdst;
  assign _GEN_43502 = 6'hc == rob_tail ? _GEN_281 : _T_5936_12_pdst;
  assign _GEN_43503 = 6'hd == rob_tail ? _GEN_281 : _T_5936_13_pdst;
  assign _GEN_43504 = 6'he == rob_tail ? _GEN_281 : _T_5936_14_pdst;
  assign _GEN_43505 = 6'hf == rob_tail ? _GEN_281 : _T_5936_15_pdst;
  assign _GEN_43506 = 6'h10 == rob_tail ? _GEN_281 : _T_5936_16_pdst;
  assign _GEN_43507 = 6'h11 == rob_tail ? _GEN_281 : _T_5936_17_pdst;
  assign _GEN_43508 = 6'h12 == rob_tail ? _GEN_281 : _T_5936_18_pdst;
  assign _GEN_43509 = 6'h13 == rob_tail ? _GEN_281 : _T_5936_19_pdst;
  assign _GEN_43510 = 6'h14 == rob_tail ? _GEN_281 : _T_5936_20_pdst;
  assign _GEN_43511 = 6'h15 == rob_tail ? _GEN_281 : _T_5936_21_pdst;
  assign _GEN_43512 = 6'h16 == rob_tail ? _GEN_281 : _T_5936_22_pdst;
  assign _GEN_43513 = 6'h17 == rob_tail ? _GEN_281 : _T_5936_23_pdst;
  assign _GEN_43514 = 6'h18 == rob_tail ? _GEN_281 : _T_5936_24_pdst;
  assign _GEN_43515 = 6'h19 == rob_tail ? _GEN_281 : _T_5936_25_pdst;
  assign _GEN_43516 = 6'h1a == rob_tail ? _GEN_281 : _T_5936_26_pdst;
  assign _GEN_43517 = 6'h1b == rob_tail ? _GEN_281 : _T_5936_27_pdst;
  assign _GEN_43518 = 6'h1c == rob_tail ? _GEN_281 : _T_5936_28_pdst;
  assign _GEN_43519 = 6'h1d == rob_tail ? _GEN_281 : _T_5936_29_pdst;
  assign _GEN_43520 = 6'h1e == rob_tail ? _GEN_281 : _T_5936_30_pdst;
  assign _GEN_43521 = 6'h1f == rob_tail ? _GEN_281 : _T_5936_31_pdst;
  assign _GEN_43522 = 6'h20 == rob_tail ? _GEN_281 : _T_5936_32_pdst;
  assign _GEN_43523 = 6'h21 == rob_tail ? _GEN_281 : _T_5936_33_pdst;
  assign _GEN_43524 = 6'h22 == rob_tail ? _GEN_281 : _T_5936_34_pdst;
  assign _GEN_43525 = 6'h23 == rob_tail ? _GEN_281 : _T_5936_35_pdst;
  assign _GEN_43526 = 6'h24 == rob_tail ? _GEN_281 : _T_5936_36_pdst;
  assign _GEN_43527 = 6'h25 == rob_tail ? _GEN_281 : _T_5936_37_pdst;
  assign _GEN_43528 = 6'h26 == rob_tail ? _GEN_281 : _T_5936_38_pdst;
  assign _GEN_43529 = 6'h27 == rob_tail ? _GEN_281 : _T_5936_39_pdst;
  assign _GEN_43770 = 6'h0 == rob_tail ? _GEN_288 : _T_5936_0_stale_pdst;
  assign _GEN_43771 = 6'h1 == rob_tail ? _GEN_288 : _T_5936_1_stale_pdst;
  assign _GEN_43772 = 6'h2 == rob_tail ? _GEN_288 : _T_5936_2_stale_pdst;
  assign _GEN_43773 = 6'h3 == rob_tail ? _GEN_288 : _T_5936_3_stale_pdst;
  assign _GEN_43774 = 6'h4 == rob_tail ? _GEN_288 : _T_5936_4_stale_pdst;
  assign _GEN_43775 = 6'h5 == rob_tail ? _GEN_288 : _T_5936_5_stale_pdst;
  assign _GEN_43776 = 6'h6 == rob_tail ? _GEN_288 : _T_5936_6_stale_pdst;
  assign _GEN_43777 = 6'h7 == rob_tail ? _GEN_288 : _T_5936_7_stale_pdst;
  assign _GEN_43778 = 6'h8 == rob_tail ? _GEN_288 : _T_5936_8_stale_pdst;
  assign _GEN_43779 = 6'h9 == rob_tail ? _GEN_288 : _T_5936_9_stale_pdst;
  assign _GEN_43780 = 6'ha == rob_tail ? _GEN_288 : _T_5936_10_stale_pdst;
  assign _GEN_43781 = 6'hb == rob_tail ? _GEN_288 : _T_5936_11_stale_pdst;
  assign _GEN_43782 = 6'hc == rob_tail ? _GEN_288 : _T_5936_12_stale_pdst;
  assign _GEN_43783 = 6'hd == rob_tail ? _GEN_288 : _T_5936_13_stale_pdst;
  assign _GEN_43784 = 6'he == rob_tail ? _GEN_288 : _T_5936_14_stale_pdst;
  assign _GEN_43785 = 6'hf == rob_tail ? _GEN_288 : _T_5936_15_stale_pdst;
  assign _GEN_43786 = 6'h10 == rob_tail ? _GEN_288 : _T_5936_16_stale_pdst;
  assign _GEN_43787 = 6'h11 == rob_tail ? _GEN_288 : _T_5936_17_stale_pdst;
  assign _GEN_43788 = 6'h12 == rob_tail ? _GEN_288 : _T_5936_18_stale_pdst;
  assign _GEN_43789 = 6'h13 == rob_tail ? _GEN_288 : _T_5936_19_stale_pdst;
  assign _GEN_43790 = 6'h14 == rob_tail ? _GEN_288 : _T_5936_20_stale_pdst;
  assign _GEN_43791 = 6'h15 == rob_tail ? _GEN_288 : _T_5936_21_stale_pdst;
  assign _GEN_43792 = 6'h16 == rob_tail ? _GEN_288 : _T_5936_22_stale_pdst;
  assign _GEN_43793 = 6'h17 == rob_tail ? _GEN_288 : _T_5936_23_stale_pdst;
  assign _GEN_43794 = 6'h18 == rob_tail ? _GEN_288 : _T_5936_24_stale_pdst;
  assign _GEN_43795 = 6'h19 == rob_tail ? _GEN_288 : _T_5936_25_stale_pdst;
  assign _GEN_43796 = 6'h1a == rob_tail ? _GEN_288 : _T_5936_26_stale_pdst;
  assign _GEN_43797 = 6'h1b == rob_tail ? _GEN_288 : _T_5936_27_stale_pdst;
  assign _GEN_43798 = 6'h1c == rob_tail ? _GEN_288 : _T_5936_28_stale_pdst;
  assign _GEN_43799 = 6'h1d == rob_tail ? _GEN_288 : _T_5936_29_stale_pdst;
  assign _GEN_43800 = 6'h1e == rob_tail ? _GEN_288 : _T_5936_30_stale_pdst;
  assign _GEN_43801 = 6'h1f == rob_tail ? _GEN_288 : _T_5936_31_stale_pdst;
  assign _GEN_43802 = 6'h20 == rob_tail ? _GEN_288 : _T_5936_32_stale_pdst;
  assign _GEN_43803 = 6'h21 == rob_tail ? _GEN_288 : _T_5936_33_stale_pdst;
  assign _GEN_43804 = 6'h22 == rob_tail ? _GEN_288 : _T_5936_34_stale_pdst;
  assign _GEN_43805 = 6'h23 == rob_tail ? _GEN_288 : _T_5936_35_stale_pdst;
  assign _GEN_43806 = 6'h24 == rob_tail ? _GEN_288 : _T_5936_36_stale_pdst;
  assign _GEN_43807 = 6'h25 == rob_tail ? _GEN_288 : _T_5936_37_stale_pdst;
  assign _GEN_43808 = 6'h26 == rob_tail ? _GEN_288 : _T_5936_38_stale_pdst;
  assign _GEN_43809 = 6'h27 == rob_tail ? _GEN_288 : _T_5936_39_stale_pdst;
  assign _GEN_44050 = 6'h0 == rob_tail ? _GEN_295 : _T_5936_0_is_fencei;
  assign _GEN_44051 = 6'h1 == rob_tail ? _GEN_295 : _T_5936_1_is_fencei;
  assign _GEN_44052 = 6'h2 == rob_tail ? _GEN_295 : _T_5936_2_is_fencei;
  assign _GEN_44053 = 6'h3 == rob_tail ? _GEN_295 : _T_5936_3_is_fencei;
  assign _GEN_44054 = 6'h4 == rob_tail ? _GEN_295 : _T_5936_4_is_fencei;
  assign _GEN_44055 = 6'h5 == rob_tail ? _GEN_295 : _T_5936_5_is_fencei;
  assign _GEN_44056 = 6'h6 == rob_tail ? _GEN_295 : _T_5936_6_is_fencei;
  assign _GEN_44057 = 6'h7 == rob_tail ? _GEN_295 : _T_5936_7_is_fencei;
  assign _GEN_44058 = 6'h8 == rob_tail ? _GEN_295 : _T_5936_8_is_fencei;
  assign _GEN_44059 = 6'h9 == rob_tail ? _GEN_295 : _T_5936_9_is_fencei;
  assign _GEN_44060 = 6'ha == rob_tail ? _GEN_295 : _T_5936_10_is_fencei;
  assign _GEN_44061 = 6'hb == rob_tail ? _GEN_295 : _T_5936_11_is_fencei;
  assign _GEN_44062 = 6'hc == rob_tail ? _GEN_295 : _T_5936_12_is_fencei;
  assign _GEN_44063 = 6'hd == rob_tail ? _GEN_295 : _T_5936_13_is_fencei;
  assign _GEN_44064 = 6'he == rob_tail ? _GEN_295 : _T_5936_14_is_fencei;
  assign _GEN_44065 = 6'hf == rob_tail ? _GEN_295 : _T_5936_15_is_fencei;
  assign _GEN_44066 = 6'h10 == rob_tail ? _GEN_295 : _T_5936_16_is_fencei;
  assign _GEN_44067 = 6'h11 == rob_tail ? _GEN_295 : _T_5936_17_is_fencei;
  assign _GEN_44068 = 6'h12 == rob_tail ? _GEN_295 : _T_5936_18_is_fencei;
  assign _GEN_44069 = 6'h13 == rob_tail ? _GEN_295 : _T_5936_19_is_fencei;
  assign _GEN_44070 = 6'h14 == rob_tail ? _GEN_295 : _T_5936_20_is_fencei;
  assign _GEN_44071 = 6'h15 == rob_tail ? _GEN_295 : _T_5936_21_is_fencei;
  assign _GEN_44072 = 6'h16 == rob_tail ? _GEN_295 : _T_5936_22_is_fencei;
  assign _GEN_44073 = 6'h17 == rob_tail ? _GEN_295 : _T_5936_23_is_fencei;
  assign _GEN_44074 = 6'h18 == rob_tail ? _GEN_295 : _T_5936_24_is_fencei;
  assign _GEN_44075 = 6'h19 == rob_tail ? _GEN_295 : _T_5936_25_is_fencei;
  assign _GEN_44076 = 6'h1a == rob_tail ? _GEN_295 : _T_5936_26_is_fencei;
  assign _GEN_44077 = 6'h1b == rob_tail ? _GEN_295 : _T_5936_27_is_fencei;
  assign _GEN_44078 = 6'h1c == rob_tail ? _GEN_295 : _T_5936_28_is_fencei;
  assign _GEN_44079 = 6'h1d == rob_tail ? _GEN_295 : _T_5936_29_is_fencei;
  assign _GEN_44080 = 6'h1e == rob_tail ? _GEN_295 : _T_5936_30_is_fencei;
  assign _GEN_44081 = 6'h1f == rob_tail ? _GEN_295 : _T_5936_31_is_fencei;
  assign _GEN_44082 = 6'h20 == rob_tail ? _GEN_295 : _T_5936_32_is_fencei;
  assign _GEN_44083 = 6'h21 == rob_tail ? _GEN_295 : _T_5936_33_is_fencei;
  assign _GEN_44084 = 6'h22 == rob_tail ? _GEN_295 : _T_5936_34_is_fencei;
  assign _GEN_44085 = 6'h23 == rob_tail ? _GEN_295 : _T_5936_35_is_fencei;
  assign _GEN_44086 = 6'h24 == rob_tail ? _GEN_295 : _T_5936_36_is_fencei;
  assign _GEN_44087 = 6'h25 == rob_tail ? _GEN_295 : _T_5936_37_is_fencei;
  assign _GEN_44088 = 6'h26 == rob_tail ? _GEN_295 : _T_5936_38_is_fencei;
  assign _GEN_44089 = 6'h27 == rob_tail ? _GEN_295 : _T_5936_39_is_fencei;
  assign _GEN_44090 = 6'h0 == rob_tail ? _GEN_296 : _T_5936_0_is_store;
  assign _GEN_44091 = 6'h1 == rob_tail ? _GEN_296 : _T_5936_1_is_store;
  assign _GEN_44092 = 6'h2 == rob_tail ? _GEN_296 : _T_5936_2_is_store;
  assign _GEN_44093 = 6'h3 == rob_tail ? _GEN_296 : _T_5936_3_is_store;
  assign _GEN_44094 = 6'h4 == rob_tail ? _GEN_296 : _T_5936_4_is_store;
  assign _GEN_44095 = 6'h5 == rob_tail ? _GEN_296 : _T_5936_5_is_store;
  assign _GEN_44096 = 6'h6 == rob_tail ? _GEN_296 : _T_5936_6_is_store;
  assign _GEN_44097 = 6'h7 == rob_tail ? _GEN_296 : _T_5936_7_is_store;
  assign _GEN_44098 = 6'h8 == rob_tail ? _GEN_296 : _T_5936_8_is_store;
  assign _GEN_44099 = 6'h9 == rob_tail ? _GEN_296 : _T_5936_9_is_store;
  assign _GEN_44100 = 6'ha == rob_tail ? _GEN_296 : _T_5936_10_is_store;
  assign _GEN_44101 = 6'hb == rob_tail ? _GEN_296 : _T_5936_11_is_store;
  assign _GEN_44102 = 6'hc == rob_tail ? _GEN_296 : _T_5936_12_is_store;
  assign _GEN_44103 = 6'hd == rob_tail ? _GEN_296 : _T_5936_13_is_store;
  assign _GEN_44104 = 6'he == rob_tail ? _GEN_296 : _T_5936_14_is_store;
  assign _GEN_44105 = 6'hf == rob_tail ? _GEN_296 : _T_5936_15_is_store;
  assign _GEN_44106 = 6'h10 == rob_tail ? _GEN_296 : _T_5936_16_is_store;
  assign _GEN_44107 = 6'h11 == rob_tail ? _GEN_296 : _T_5936_17_is_store;
  assign _GEN_44108 = 6'h12 == rob_tail ? _GEN_296 : _T_5936_18_is_store;
  assign _GEN_44109 = 6'h13 == rob_tail ? _GEN_296 : _T_5936_19_is_store;
  assign _GEN_44110 = 6'h14 == rob_tail ? _GEN_296 : _T_5936_20_is_store;
  assign _GEN_44111 = 6'h15 == rob_tail ? _GEN_296 : _T_5936_21_is_store;
  assign _GEN_44112 = 6'h16 == rob_tail ? _GEN_296 : _T_5936_22_is_store;
  assign _GEN_44113 = 6'h17 == rob_tail ? _GEN_296 : _T_5936_23_is_store;
  assign _GEN_44114 = 6'h18 == rob_tail ? _GEN_296 : _T_5936_24_is_store;
  assign _GEN_44115 = 6'h19 == rob_tail ? _GEN_296 : _T_5936_25_is_store;
  assign _GEN_44116 = 6'h1a == rob_tail ? _GEN_296 : _T_5936_26_is_store;
  assign _GEN_44117 = 6'h1b == rob_tail ? _GEN_296 : _T_5936_27_is_store;
  assign _GEN_44118 = 6'h1c == rob_tail ? _GEN_296 : _T_5936_28_is_store;
  assign _GEN_44119 = 6'h1d == rob_tail ? _GEN_296 : _T_5936_29_is_store;
  assign _GEN_44120 = 6'h1e == rob_tail ? _GEN_296 : _T_5936_30_is_store;
  assign _GEN_44121 = 6'h1f == rob_tail ? _GEN_296 : _T_5936_31_is_store;
  assign _GEN_44122 = 6'h20 == rob_tail ? _GEN_296 : _T_5936_32_is_store;
  assign _GEN_44123 = 6'h21 == rob_tail ? _GEN_296 : _T_5936_33_is_store;
  assign _GEN_44124 = 6'h22 == rob_tail ? _GEN_296 : _T_5936_34_is_store;
  assign _GEN_44125 = 6'h23 == rob_tail ? _GEN_296 : _T_5936_35_is_store;
  assign _GEN_44126 = 6'h24 == rob_tail ? _GEN_296 : _T_5936_36_is_store;
  assign _GEN_44127 = 6'h25 == rob_tail ? _GEN_296 : _T_5936_37_is_store;
  assign _GEN_44128 = 6'h26 == rob_tail ? _GEN_296 : _T_5936_38_is_store;
  assign _GEN_44129 = 6'h27 == rob_tail ? _GEN_296 : _T_5936_39_is_store;
  assign _GEN_44170 = 6'h0 == rob_tail ? _GEN_298 : _T_5936_0_is_load;
  assign _GEN_44171 = 6'h1 == rob_tail ? _GEN_298 : _T_5936_1_is_load;
  assign _GEN_44172 = 6'h2 == rob_tail ? _GEN_298 : _T_5936_2_is_load;
  assign _GEN_44173 = 6'h3 == rob_tail ? _GEN_298 : _T_5936_3_is_load;
  assign _GEN_44174 = 6'h4 == rob_tail ? _GEN_298 : _T_5936_4_is_load;
  assign _GEN_44175 = 6'h5 == rob_tail ? _GEN_298 : _T_5936_5_is_load;
  assign _GEN_44176 = 6'h6 == rob_tail ? _GEN_298 : _T_5936_6_is_load;
  assign _GEN_44177 = 6'h7 == rob_tail ? _GEN_298 : _T_5936_7_is_load;
  assign _GEN_44178 = 6'h8 == rob_tail ? _GEN_298 : _T_5936_8_is_load;
  assign _GEN_44179 = 6'h9 == rob_tail ? _GEN_298 : _T_5936_9_is_load;
  assign _GEN_44180 = 6'ha == rob_tail ? _GEN_298 : _T_5936_10_is_load;
  assign _GEN_44181 = 6'hb == rob_tail ? _GEN_298 : _T_5936_11_is_load;
  assign _GEN_44182 = 6'hc == rob_tail ? _GEN_298 : _T_5936_12_is_load;
  assign _GEN_44183 = 6'hd == rob_tail ? _GEN_298 : _T_5936_13_is_load;
  assign _GEN_44184 = 6'he == rob_tail ? _GEN_298 : _T_5936_14_is_load;
  assign _GEN_44185 = 6'hf == rob_tail ? _GEN_298 : _T_5936_15_is_load;
  assign _GEN_44186 = 6'h10 == rob_tail ? _GEN_298 : _T_5936_16_is_load;
  assign _GEN_44187 = 6'h11 == rob_tail ? _GEN_298 : _T_5936_17_is_load;
  assign _GEN_44188 = 6'h12 == rob_tail ? _GEN_298 : _T_5936_18_is_load;
  assign _GEN_44189 = 6'h13 == rob_tail ? _GEN_298 : _T_5936_19_is_load;
  assign _GEN_44190 = 6'h14 == rob_tail ? _GEN_298 : _T_5936_20_is_load;
  assign _GEN_44191 = 6'h15 == rob_tail ? _GEN_298 : _T_5936_21_is_load;
  assign _GEN_44192 = 6'h16 == rob_tail ? _GEN_298 : _T_5936_22_is_load;
  assign _GEN_44193 = 6'h17 == rob_tail ? _GEN_298 : _T_5936_23_is_load;
  assign _GEN_44194 = 6'h18 == rob_tail ? _GEN_298 : _T_5936_24_is_load;
  assign _GEN_44195 = 6'h19 == rob_tail ? _GEN_298 : _T_5936_25_is_load;
  assign _GEN_44196 = 6'h1a == rob_tail ? _GEN_298 : _T_5936_26_is_load;
  assign _GEN_44197 = 6'h1b == rob_tail ? _GEN_298 : _T_5936_27_is_load;
  assign _GEN_44198 = 6'h1c == rob_tail ? _GEN_298 : _T_5936_28_is_load;
  assign _GEN_44199 = 6'h1d == rob_tail ? _GEN_298 : _T_5936_29_is_load;
  assign _GEN_44200 = 6'h1e == rob_tail ? _GEN_298 : _T_5936_30_is_load;
  assign _GEN_44201 = 6'h1f == rob_tail ? _GEN_298 : _T_5936_31_is_load;
  assign _GEN_44202 = 6'h20 == rob_tail ? _GEN_298 : _T_5936_32_is_load;
  assign _GEN_44203 = 6'h21 == rob_tail ? _GEN_298 : _T_5936_33_is_load;
  assign _GEN_44204 = 6'h22 == rob_tail ? _GEN_298 : _T_5936_34_is_load;
  assign _GEN_44205 = 6'h23 == rob_tail ? _GEN_298 : _T_5936_35_is_load;
  assign _GEN_44206 = 6'h24 == rob_tail ? _GEN_298 : _T_5936_36_is_load;
  assign _GEN_44207 = 6'h25 == rob_tail ? _GEN_298 : _T_5936_37_is_load;
  assign _GEN_44208 = 6'h26 == rob_tail ? _GEN_298 : _T_5936_38_is_load;
  assign _GEN_44209 = 6'h27 == rob_tail ? _GEN_298 : _T_5936_39_is_load;
  assign _GEN_44210 = 6'h0 == rob_tail ? _GEN_299 : _T_5936_0_is_sys_pc2epc;
  assign _GEN_44211 = 6'h1 == rob_tail ? _GEN_299 : _T_5936_1_is_sys_pc2epc;
  assign _GEN_44212 = 6'h2 == rob_tail ? _GEN_299 : _T_5936_2_is_sys_pc2epc;
  assign _GEN_44213 = 6'h3 == rob_tail ? _GEN_299 : _T_5936_3_is_sys_pc2epc;
  assign _GEN_44214 = 6'h4 == rob_tail ? _GEN_299 : _T_5936_4_is_sys_pc2epc;
  assign _GEN_44215 = 6'h5 == rob_tail ? _GEN_299 : _T_5936_5_is_sys_pc2epc;
  assign _GEN_44216 = 6'h6 == rob_tail ? _GEN_299 : _T_5936_6_is_sys_pc2epc;
  assign _GEN_44217 = 6'h7 == rob_tail ? _GEN_299 : _T_5936_7_is_sys_pc2epc;
  assign _GEN_44218 = 6'h8 == rob_tail ? _GEN_299 : _T_5936_8_is_sys_pc2epc;
  assign _GEN_44219 = 6'h9 == rob_tail ? _GEN_299 : _T_5936_9_is_sys_pc2epc;
  assign _GEN_44220 = 6'ha == rob_tail ? _GEN_299 : _T_5936_10_is_sys_pc2epc;
  assign _GEN_44221 = 6'hb == rob_tail ? _GEN_299 : _T_5936_11_is_sys_pc2epc;
  assign _GEN_44222 = 6'hc == rob_tail ? _GEN_299 : _T_5936_12_is_sys_pc2epc;
  assign _GEN_44223 = 6'hd == rob_tail ? _GEN_299 : _T_5936_13_is_sys_pc2epc;
  assign _GEN_44224 = 6'he == rob_tail ? _GEN_299 : _T_5936_14_is_sys_pc2epc;
  assign _GEN_44225 = 6'hf == rob_tail ? _GEN_299 : _T_5936_15_is_sys_pc2epc;
  assign _GEN_44226 = 6'h10 == rob_tail ? _GEN_299 : _T_5936_16_is_sys_pc2epc;
  assign _GEN_44227 = 6'h11 == rob_tail ? _GEN_299 : _T_5936_17_is_sys_pc2epc;
  assign _GEN_44228 = 6'h12 == rob_tail ? _GEN_299 : _T_5936_18_is_sys_pc2epc;
  assign _GEN_44229 = 6'h13 == rob_tail ? _GEN_299 : _T_5936_19_is_sys_pc2epc;
  assign _GEN_44230 = 6'h14 == rob_tail ? _GEN_299 : _T_5936_20_is_sys_pc2epc;
  assign _GEN_44231 = 6'h15 == rob_tail ? _GEN_299 : _T_5936_21_is_sys_pc2epc;
  assign _GEN_44232 = 6'h16 == rob_tail ? _GEN_299 : _T_5936_22_is_sys_pc2epc;
  assign _GEN_44233 = 6'h17 == rob_tail ? _GEN_299 : _T_5936_23_is_sys_pc2epc;
  assign _GEN_44234 = 6'h18 == rob_tail ? _GEN_299 : _T_5936_24_is_sys_pc2epc;
  assign _GEN_44235 = 6'h19 == rob_tail ? _GEN_299 : _T_5936_25_is_sys_pc2epc;
  assign _GEN_44236 = 6'h1a == rob_tail ? _GEN_299 : _T_5936_26_is_sys_pc2epc;
  assign _GEN_44237 = 6'h1b == rob_tail ? _GEN_299 : _T_5936_27_is_sys_pc2epc;
  assign _GEN_44238 = 6'h1c == rob_tail ? _GEN_299 : _T_5936_28_is_sys_pc2epc;
  assign _GEN_44239 = 6'h1d == rob_tail ? _GEN_299 : _T_5936_29_is_sys_pc2epc;
  assign _GEN_44240 = 6'h1e == rob_tail ? _GEN_299 : _T_5936_30_is_sys_pc2epc;
  assign _GEN_44241 = 6'h1f == rob_tail ? _GEN_299 : _T_5936_31_is_sys_pc2epc;
  assign _GEN_44242 = 6'h20 == rob_tail ? _GEN_299 : _T_5936_32_is_sys_pc2epc;
  assign _GEN_44243 = 6'h21 == rob_tail ? _GEN_299 : _T_5936_33_is_sys_pc2epc;
  assign _GEN_44244 = 6'h22 == rob_tail ? _GEN_299 : _T_5936_34_is_sys_pc2epc;
  assign _GEN_44245 = 6'h23 == rob_tail ? _GEN_299 : _T_5936_35_is_sys_pc2epc;
  assign _GEN_44246 = 6'h24 == rob_tail ? _GEN_299 : _T_5936_36_is_sys_pc2epc;
  assign _GEN_44247 = 6'h25 == rob_tail ? _GEN_299 : _T_5936_37_is_sys_pc2epc;
  assign _GEN_44248 = 6'h26 == rob_tail ? _GEN_299 : _T_5936_38_is_sys_pc2epc;
  assign _GEN_44249 = 6'h27 == rob_tail ? _GEN_299 : _T_5936_39_is_sys_pc2epc;
  assign _GEN_44290 = 6'h0 == rob_tail ? _GEN_301 : _T_5936_0_flush_on_commit;
  assign _GEN_44291 = 6'h1 == rob_tail ? _GEN_301 : _T_5936_1_flush_on_commit;
  assign _GEN_44292 = 6'h2 == rob_tail ? _GEN_301 : _T_5936_2_flush_on_commit;
  assign _GEN_44293 = 6'h3 == rob_tail ? _GEN_301 : _T_5936_3_flush_on_commit;
  assign _GEN_44294 = 6'h4 == rob_tail ? _GEN_301 : _T_5936_4_flush_on_commit;
  assign _GEN_44295 = 6'h5 == rob_tail ? _GEN_301 : _T_5936_5_flush_on_commit;
  assign _GEN_44296 = 6'h6 == rob_tail ? _GEN_301 : _T_5936_6_flush_on_commit;
  assign _GEN_44297 = 6'h7 == rob_tail ? _GEN_301 : _T_5936_7_flush_on_commit;
  assign _GEN_44298 = 6'h8 == rob_tail ? _GEN_301 : _T_5936_8_flush_on_commit;
  assign _GEN_44299 = 6'h9 == rob_tail ? _GEN_301 : _T_5936_9_flush_on_commit;
  assign _GEN_44300 = 6'ha == rob_tail ? _GEN_301 : _T_5936_10_flush_on_commit;
  assign _GEN_44301 = 6'hb == rob_tail ? _GEN_301 : _T_5936_11_flush_on_commit;
  assign _GEN_44302 = 6'hc == rob_tail ? _GEN_301 : _T_5936_12_flush_on_commit;
  assign _GEN_44303 = 6'hd == rob_tail ? _GEN_301 : _T_5936_13_flush_on_commit;
  assign _GEN_44304 = 6'he == rob_tail ? _GEN_301 : _T_5936_14_flush_on_commit;
  assign _GEN_44305 = 6'hf == rob_tail ? _GEN_301 : _T_5936_15_flush_on_commit;
  assign _GEN_44306 = 6'h10 == rob_tail ? _GEN_301 : _T_5936_16_flush_on_commit;
  assign _GEN_44307 = 6'h11 == rob_tail ? _GEN_301 : _T_5936_17_flush_on_commit;
  assign _GEN_44308 = 6'h12 == rob_tail ? _GEN_301 : _T_5936_18_flush_on_commit;
  assign _GEN_44309 = 6'h13 == rob_tail ? _GEN_301 : _T_5936_19_flush_on_commit;
  assign _GEN_44310 = 6'h14 == rob_tail ? _GEN_301 : _T_5936_20_flush_on_commit;
  assign _GEN_44311 = 6'h15 == rob_tail ? _GEN_301 : _T_5936_21_flush_on_commit;
  assign _GEN_44312 = 6'h16 == rob_tail ? _GEN_301 : _T_5936_22_flush_on_commit;
  assign _GEN_44313 = 6'h17 == rob_tail ? _GEN_301 : _T_5936_23_flush_on_commit;
  assign _GEN_44314 = 6'h18 == rob_tail ? _GEN_301 : _T_5936_24_flush_on_commit;
  assign _GEN_44315 = 6'h19 == rob_tail ? _GEN_301 : _T_5936_25_flush_on_commit;
  assign _GEN_44316 = 6'h1a == rob_tail ? _GEN_301 : _T_5936_26_flush_on_commit;
  assign _GEN_44317 = 6'h1b == rob_tail ? _GEN_301 : _T_5936_27_flush_on_commit;
  assign _GEN_44318 = 6'h1c == rob_tail ? _GEN_301 : _T_5936_28_flush_on_commit;
  assign _GEN_44319 = 6'h1d == rob_tail ? _GEN_301 : _T_5936_29_flush_on_commit;
  assign _GEN_44320 = 6'h1e == rob_tail ? _GEN_301 : _T_5936_30_flush_on_commit;
  assign _GEN_44321 = 6'h1f == rob_tail ? _GEN_301 : _T_5936_31_flush_on_commit;
  assign _GEN_44322 = 6'h20 == rob_tail ? _GEN_301 : _T_5936_32_flush_on_commit;
  assign _GEN_44323 = 6'h21 == rob_tail ? _GEN_301 : _T_5936_33_flush_on_commit;
  assign _GEN_44324 = 6'h22 == rob_tail ? _GEN_301 : _T_5936_34_flush_on_commit;
  assign _GEN_44325 = 6'h23 == rob_tail ? _GEN_301 : _T_5936_35_flush_on_commit;
  assign _GEN_44326 = 6'h24 == rob_tail ? _GEN_301 : _T_5936_36_flush_on_commit;
  assign _GEN_44327 = 6'h25 == rob_tail ? _GEN_301 : _T_5936_37_flush_on_commit;
  assign _GEN_44328 = 6'h26 == rob_tail ? _GEN_301 : _T_5936_38_flush_on_commit;
  assign _GEN_44329 = 6'h27 == rob_tail ? _GEN_301 : _T_5936_39_flush_on_commit;
  assign _GEN_44330 = 6'h0 == rob_tail ? _GEN_302 : _T_5936_0_ldst;
  assign _GEN_44331 = 6'h1 == rob_tail ? _GEN_302 : _T_5936_1_ldst;
  assign _GEN_44332 = 6'h2 == rob_tail ? _GEN_302 : _T_5936_2_ldst;
  assign _GEN_44333 = 6'h3 == rob_tail ? _GEN_302 : _T_5936_3_ldst;
  assign _GEN_44334 = 6'h4 == rob_tail ? _GEN_302 : _T_5936_4_ldst;
  assign _GEN_44335 = 6'h5 == rob_tail ? _GEN_302 : _T_5936_5_ldst;
  assign _GEN_44336 = 6'h6 == rob_tail ? _GEN_302 : _T_5936_6_ldst;
  assign _GEN_44337 = 6'h7 == rob_tail ? _GEN_302 : _T_5936_7_ldst;
  assign _GEN_44338 = 6'h8 == rob_tail ? _GEN_302 : _T_5936_8_ldst;
  assign _GEN_44339 = 6'h9 == rob_tail ? _GEN_302 : _T_5936_9_ldst;
  assign _GEN_44340 = 6'ha == rob_tail ? _GEN_302 : _T_5936_10_ldst;
  assign _GEN_44341 = 6'hb == rob_tail ? _GEN_302 : _T_5936_11_ldst;
  assign _GEN_44342 = 6'hc == rob_tail ? _GEN_302 : _T_5936_12_ldst;
  assign _GEN_44343 = 6'hd == rob_tail ? _GEN_302 : _T_5936_13_ldst;
  assign _GEN_44344 = 6'he == rob_tail ? _GEN_302 : _T_5936_14_ldst;
  assign _GEN_44345 = 6'hf == rob_tail ? _GEN_302 : _T_5936_15_ldst;
  assign _GEN_44346 = 6'h10 == rob_tail ? _GEN_302 : _T_5936_16_ldst;
  assign _GEN_44347 = 6'h11 == rob_tail ? _GEN_302 : _T_5936_17_ldst;
  assign _GEN_44348 = 6'h12 == rob_tail ? _GEN_302 : _T_5936_18_ldst;
  assign _GEN_44349 = 6'h13 == rob_tail ? _GEN_302 : _T_5936_19_ldst;
  assign _GEN_44350 = 6'h14 == rob_tail ? _GEN_302 : _T_5936_20_ldst;
  assign _GEN_44351 = 6'h15 == rob_tail ? _GEN_302 : _T_5936_21_ldst;
  assign _GEN_44352 = 6'h16 == rob_tail ? _GEN_302 : _T_5936_22_ldst;
  assign _GEN_44353 = 6'h17 == rob_tail ? _GEN_302 : _T_5936_23_ldst;
  assign _GEN_44354 = 6'h18 == rob_tail ? _GEN_302 : _T_5936_24_ldst;
  assign _GEN_44355 = 6'h19 == rob_tail ? _GEN_302 : _T_5936_25_ldst;
  assign _GEN_44356 = 6'h1a == rob_tail ? _GEN_302 : _T_5936_26_ldst;
  assign _GEN_44357 = 6'h1b == rob_tail ? _GEN_302 : _T_5936_27_ldst;
  assign _GEN_44358 = 6'h1c == rob_tail ? _GEN_302 : _T_5936_28_ldst;
  assign _GEN_44359 = 6'h1d == rob_tail ? _GEN_302 : _T_5936_29_ldst;
  assign _GEN_44360 = 6'h1e == rob_tail ? _GEN_302 : _T_5936_30_ldst;
  assign _GEN_44361 = 6'h1f == rob_tail ? _GEN_302 : _T_5936_31_ldst;
  assign _GEN_44362 = 6'h20 == rob_tail ? _GEN_302 : _T_5936_32_ldst;
  assign _GEN_44363 = 6'h21 == rob_tail ? _GEN_302 : _T_5936_33_ldst;
  assign _GEN_44364 = 6'h22 == rob_tail ? _GEN_302 : _T_5936_34_ldst;
  assign _GEN_44365 = 6'h23 == rob_tail ? _GEN_302 : _T_5936_35_ldst;
  assign _GEN_44366 = 6'h24 == rob_tail ? _GEN_302 : _T_5936_36_ldst;
  assign _GEN_44367 = 6'h25 == rob_tail ? _GEN_302 : _T_5936_37_ldst;
  assign _GEN_44368 = 6'h26 == rob_tail ? _GEN_302 : _T_5936_38_ldst;
  assign _GEN_44369 = 6'h27 == rob_tail ? _GEN_302 : _T_5936_39_ldst;
  assign _GEN_44490 = 6'h0 == rob_tail ? _GEN_306 : _T_5936_0_ldst_val;
  assign _GEN_44491 = 6'h1 == rob_tail ? _GEN_306 : _T_5936_1_ldst_val;
  assign _GEN_44492 = 6'h2 == rob_tail ? _GEN_306 : _T_5936_2_ldst_val;
  assign _GEN_44493 = 6'h3 == rob_tail ? _GEN_306 : _T_5936_3_ldst_val;
  assign _GEN_44494 = 6'h4 == rob_tail ? _GEN_306 : _T_5936_4_ldst_val;
  assign _GEN_44495 = 6'h5 == rob_tail ? _GEN_306 : _T_5936_5_ldst_val;
  assign _GEN_44496 = 6'h6 == rob_tail ? _GEN_306 : _T_5936_6_ldst_val;
  assign _GEN_44497 = 6'h7 == rob_tail ? _GEN_306 : _T_5936_7_ldst_val;
  assign _GEN_44498 = 6'h8 == rob_tail ? _GEN_306 : _T_5936_8_ldst_val;
  assign _GEN_44499 = 6'h9 == rob_tail ? _GEN_306 : _T_5936_9_ldst_val;
  assign _GEN_44500 = 6'ha == rob_tail ? _GEN_306 : _T_5936_10_ldst_val;
  assign _GEN_44501 = 6'hb == rob_tail ? _GEN_306 : _T_5936_11_ldst_val;
  assign _GEN_44502 = 6'hc == rob_tail ? _GEN_306 : _T_5936_12_ldst_val;
  assign _GEN_44503 = 6'hd == rob_tail ? _GEN_306 : _T_5936_13_ldst_val;
  assign _GEN_44504 = 6'he == rob_tail ? _GEN_306 : _T_5936_14_ldst_val;
  assign _GEN_44505 = 6'hf == rob_tail ? _GEN_306 : _T_5936_15_ldst_val;
  assign _GEN_44506 = 6'h10 == rob_tail ? _GEN_306 : _T_5936_16_ldst_val;
  assign _GEN_44507 = 6'h11 == rob_tail ? _GEN_306 : _T_5936_17_ldst_val;
  assign _GEN_44508 = 6'h12 == rob_tail ? _GEN_306 : _T_5936_18_ldst_val;
  assign _GEN_44509 = 6'h13 == rob_tail ? _GEN_306 : _T_5936_19_ldst_val;
  assign _GEN_44510 = 6'h14 == rob_tail ? _GEN_306 : _T_5936_20_ldst_val;
  assign _GEN_44511 = 6'h15 == rob_tail ? _GEN_306 : _T_5936_21_ldst_val;
  assign _GEN_44512 = 6'h16 == rob_tail ? _GEN_306 : _T_5936_22_ldst_val;
  assign _GEN_44513 = 6'h17 == rob_tail ? _GEN_306 : _T_5936_23_ldst_val;
  assign _GEN_44514 = 6'h18 == rob_tail ? _GEN_306 : _T_5936_24_ldst_val;
  assign _GEN_44515 = 6'h19 == rob_tail ? _GEN_306 : _T_5936_25_ldst_val;
  assign _GEN_44516 = 6'h1a == rob_tail ? _GEN_306 : _T_5936_26_ldst_val;
  assign _GEN_44517 = 6'h1b == rob_tail ? _GEN_306 : _T_5936_27_ldst_val;
  assign _GEN_44518 = 6'h1c == rob_tail ? _GEN_306 : _T_5936_28_ldst_val;
  assign _GEN_44519 = 6'h1d == rob_tail ? _GEN_306 : _T_5936_29_ldst_val;
  assign _GEN_44520 = 6'h1e == rob_tail ? _GEN_306 : _T_5936_30_ldst_val;
  assign _GEN_44521 = 6'h1f == rob_tail ? _GEN_306 : _T_5936_31_ldst_val;
  assign _GEN_44522 = 6'h20 == rob_tail ? _GEN_306 : _T_5936_32_ldst_val;
  assign _GEN_44523 = 6'h21 == rob_tail ? _GEN_306 : _T_5936_33_ldst_val;
  assign _GEN_44524 = 6'h22 == rob_tail ? _GEN_306 : _T_5936_34_ldst_val;
  assign _GEN_44525 = 6'h23 == rob_tail ? _GEN_306 : _T_5936_35_ldst_val;
  assign _GEN_44526 = 6'h24 == rob_tail ? _GEN_306 : _T_5936_36_ldst_val;
  assign _GEN_44527 = 6'h25 == rob_tail ? _GEN_306 : _T_5936_37_ldst_val;
  assign _GEN_44528 = 6'h26 == rob_tail ? _GEN_306 : _T_5936_38_ldst_val;
  assign _GEN_44529 = 6'h27 == rob_tail ? _GEN_306 : _T_5936_39_ldst_val;
  assign _GEN_44530 = 6'h0 == rob_tail ? _GEN_307 : _T_5936_0_dst_rtype;
  assign _GEN_44531 = 6'h1 == rob_tail ? _GEN_307 : _T_5936_1_dst_rtype;
  assign _GEN_44532 = 6'h2 == rob_tail ? _GEN_307 : _T_5936_2_dst_rtype;
  assign _GEN_44533 = 6'h3 == rob_tail ? _GEN_307 : _T_5936_3_dst_rtype;
  assign _GEN_44534 = 6'h4 == rob_tail ? _GEN_307 : _T_5936_4_dst_rtype;
  assign _GEN_44535 = 6'h5 == rob_tail ? _GEN_307 : _T_5936_5_dst_rtype;
  assign _GEN_44536 = 6'h6 == rob_tail ? _GEN_307 : _T_5936_6_dst_rtype;
  assign _GEN_44537 = 6'h7 == rob_tail ? _GEN_307 : _T_5936_7_dst_rtype;
  assign _GEN_44538 = 6'h8 == rob_tail ? _GEN_307 : _T_5936_8_dst_rtype;
  assign _GEN_44539 = 6'h9 == rob_tail ? _GEN_307 : _T_5936_9_dst_rtype;
  assign _GEN_44540 = 6'ha == rob_tail ? _GEN_307 : _T_5936_10_dst_rtype;
  assign _GEN_44541 = 6'hb == rob_tail ? _GEN_307 : _T_5936_11_dst_rtype;
  assign _GEN_44542 = 6'hc == rob_tail ? _GEN_307 : _T_5936_12_dst_rtype;
  assign _GEN_44543 = 6'hd == rob_tail ? _GEN_307 : _T_5936_13_dst_rtype;
  assign _GEN_44544 = 6'he == rob_tail ? _GEN_307 : _T_5936_14_dst_rtype;
  assign _GEN_44545 = 6'hf == rob_tail ? _GEN_307 : _T_5936_15_dst_rtype;
  assign _GEN_44546 = 6'h10 == rob_tail ? _GEN_307 : _T_5936_16_dst_rtype;
  assign _GEN_44547 = 6'h11 == rob_tail ? _GEN_307 : _T_5936_17_dst_rtype;
  assign _GEN_44548 = 6'h12 == rob_tail ? _GEN_307 : _T_5936_18_dst_rtype;
  assign _GEN_44549 = 6'h13 == rob_tail ? _GEN_307 : _T_5936_19_dst_rtype;
  assign _GEN_44550 = 6'h14 == rob_tail ? _GEN_307 : _T_5936_20_dst_rtype;
  assign _GEN_44551 = 6'h15 == rob_tail ? _GEN_307 : _T_5936_21_dst_rtype;
  assign _GEN_44552 = 6'h16 == rob_tail ? _GEN_307 : _T_5936_22_dst_rtype;
  assign _GEN_44553 = 6'h17 == rob_tail ? _GEN_307 : _T_5936_23_dst_rtype;
  assign _GEN_44554 = 6'h18 == rob_tail ? _GEN_307 : _T_5936_24_dst_rtype;
  assign _GEN_44555 = 6'h19 == rob_tail ? _GEN_307 : _T_5936_25_dst_rtype;
  assign _GEN_44556 = 6'h1a == rob_tail ? _GEN_307 : _T_5936_26_dst_rtype;
  assign _GEN_44557 = 6'h1b == rob_tail ? _GEN_307 : _T_5936_27_dst_rtype;
  assign _GEN_44558 = 6'h1c == rob_tail ? _GEN_307 : _T_5936_28_dst_rtype;
  assign _GEN_44559 = 6'h1d == rob_tail ? _GEN_307 : _T_5936_29_dst_rtype;
  assign _GEN_44560 = 6'h1e == rob_tail ? _GEN_307 : _T_5936_30_dst_rtype;
  assign _GEN_44561 = 6'h1f == rob_tail ? _GEN_307 : _T_5936_31_dst_rtype;
  assign _GEN_44562 = 6'h20 == rob_tail ? _GEN_307 : _T_5936_32_dst_rtype;
  assign _GEN_44563 = 6'h21 == rob_tail ? _GEN_307 : _T_5936_33_dst_rtype;
  assign _GEN_44564 = 6'h22 == rob_tail ? _GEN_307 : _T_5936_34_dst_rtype;
  assign _GEN_44565 = 6'h23 == rob_tail ? _GEN_307 : _T_5936_35_dst_rtype;
  assign _GEN_44566 = 6'h24 == rob_tail ? _GEN_307 : _T_5936_36_dst_rtype;
  assign _GEN_44567 = 6'h25 == rob_tail ? _GEN_307 : _T_5936_37_dst_rtype;
  assign _GEN_44568 = 6'h26 == rob_tail ? _GEN_307 : _T_5936_38_dst_rtype;
  assign _GEN_44569 = 6'h27 == rob_tail ? _GEN_307 : _T_5936_39_dst_rtype;
  assign _GEN_44690 = 6'h0 == rob_tail ? _GEN_311 : _T_5936_0_fp_val;
  assign _GEN_44691 = 6'h1 == rob_tail ? _GEN_311 : _T_5936_1_fp_val;
  assign _GEN_44692 = 6'h2 == rob_tail ? _GEN_311 : _T_5936_2_fp_val;
  assign _GEN_44693 = 6'h3 == rob_tail ? _GEN_311 : _T_5936_3_fp_val;
  assign _GEN_44694 = 6'h4 == rob_tail ? _GEN_311 : _T_5936_4_fp_val;
  assign _GEN_44695 = 6'h5 == rob_tail ? _GEN_311 : _T_5936_5_fp_val;
  assign _GEN_44696 = 6'h6 == rob_tail ? _GEN_311 : _T_5936_6_fp_val;
  assign _GEN_44697 = 6'h7 == rob_tail ? _GEN_311 : _T_5936_7_fp_val;
  assign _GEN_44698 = 6'h8 == rob_tail ? _GEN_311 : _T_5936_8_fp_val;
  assign _GEN_44699 = 6'h9 == rob_tail ? _GEN_311 : _T_5936_9_fp_val;
  assign _GEN_44700 = 6'ha == rob_tail ? _GEN_311 : _T_5936_10_fp_val;
  assign _GEN_44701 = 6'hb == rob_tail ? _GEN_311 : _T_5936_11_fp_val;
  assign _GEN_44702 = 6'hc == rob_tail ? _GEN_311 : _T_5936_12_fp_val;
  assign _GEN_44703 = 6'hd == rob_tail ? _GEN_311 : _T_5936_13_fp_val;
  assign _GEN_44704 = 6'he == rob_tail ? _GEN_311 : _T_5936_14_fp_val;
  assign _GEN_44705 = 6'hf == rob_tail ? _GEN_311 : _T_5936_15_fp_val;
  assign _GEN_44706 = 6'h10 == rob_tail ? _GEN_311 : _T_5936_16_fp_val;
  assign _GEN_44707 = 6'h11 == rob_tail ? _GEN_311 : _T_5936_17_fp_val;
  assign _GEN_44708 = 6'h12 == rob_tail ? _GEN_311 : _T_5936_18_fp_val;
  assign _GEN_44709 = 6'h13 == rob_tail ? _GEN_311 : _T_5936_19_fp_val;
  assign _GEN_44710 = 6'h14 == rob_tail ? _GEN_311 : _T_5936_20_fp_val;
  assign _GEN_44711 = 6'h15 == rob_tail ? _GEN_311 : _T_5936_21_fp_val;
  assign _GEN_44712 = 6'h16 == rob_tail ? _GEN_311 : _T_5936_22_fp_val;
  assign _GEN_44713 = 6'h17 == rob_tail ? _GEN_311 : _T_5936_23_fp_val;
  assign _GEN_44714 = 6'h18 == rob_tail ? _GEN_311 : _T_5936_24_fp_val;
  assign _GEN_44715 = 6'h19 == rob_tail ? _GEN_311 : _T_5936_25_fp_val;
  assign _GEN_44716 = 6'h1a == rob_tail ? _GEN_311 : _T_5936_26_fp_val;
  assign _GEN_44717 = 6'h1b == rob_tail ? _GEN_311 : _T_5936_27_fp_val;
  assign _GEN_44718 = 6'h1c == rob_tail ? _GEN_311 : _T_5936_28_fp_val;
  assign _GEN_44719 = 6'h1d == rob_tail ? _GEN_311 : _T_5936_29_fp_val;
  assign _GEN_44720 = 6'h1e == rob_tail ? _GEN_311 : _T_5936_30_fp_val;
  assign _GEN_44721 = 6'h1f == rob_tail ? _GEN_311 : _T_5936_31_fp_val;
  assign _GEN_44722 = 6'h20 == rob_tail ? _GEN_311 : _T_5936_32_fp_val;
  assign _GEN_44723 = 6'h21 == rob_tail ? _GEN_311 : _T_5936_33_fp_val;
  assign _GEN_44724 = 6'h22 == rob_tail ? _GEN_311 : _T_5936_34_fp_val;
  assign _GEN_44725 = 6'h23 == rob_tail ? _GEN_311 : _T_5936_35_fp_val;
  assign _GEN_44726 = 6'h24 == rob_tail ? _GEN_311 : _T_5936_36_fp_val;
  assign _GEN_44727 = 6'h25 == rob_tail ? _GEN_311 : _T_5936_37_fp_val;
  assign _GEN_44728 = 6'h26 == rob_tail ? _GEN_311 : _T_5936_38_fp_val;
  assign _GEN_44729 = 6'h27 == rob_tail ? _GEN_311 : _T_5936_39_fp_val;
  assign _GEN_45050 = 6'h1 == rob_tail ? _T_5637_1 : _T_5637_0;
  assign _GEN_45051 = 6'h2 == rob_tail ? _T_5637_2 : _GEN_45050;
  assign _GEN_45052 = 6'h3 == rob_tail ? _T_5637_3 : _GEN_45051;
  assign _GEN_45053 = 6'h4 == rob_tail ? _T_5637_4 : _GEN_45052;
  assign _GEN_45054 = 6'h5 == rob_tail ? _T_5637_5 : _GEN_45053;
  assign _GEN_45055 = 6'h6 == rob_tail ? _T_5637_6 : _GEN_45054;
  assign _GEN_45056 = 6'h7 == rob_tail ? _T_5637_7 : _GEN_45055;
  assign _GEN_45057 = 6'h8 == rob_tail ? _T_5637_8 : _GEN_45056;
  assign _GEN_45058 = 6'h9 == rob_tail ? _T_5637_9 : _GEN_45057;
  assign _GEN_45059 = 6'ha == rob_tail ? _T_5637_10 : _GEN_45058;
  assign _GEN_45060 = 6'hb == rob_tail ? _T_5637_11 : _GEN_45059;
  assign _GEN_45061 = 6'hc == rob_tail ? _T_5637_12 : _GEN_45060;
  assign _GEN_45062 = 6'hd == rob_tail ? _T_5637_13 : _GEN_45061;
  assign _GEN_45063 = 6'he == rob_tail ? _T_5637_14 : _GEN_45062;
  assign _GEN_45064 = 6'hf == rob_tail ? _T_5637_15 : _GEN_45063;
  assign _GEN_45065 = 6'h10 == rob_tail ? _T_5637_16 : _GEN_45064;
  assign _GEN_45066 = 6'h11 == rob_tail ? _T_5637_17 : _GEN_45065;
  assign _GEN_45067 = 6'h12 == rob_tail ? _T_5637_18 : _GEN_45066;
  assign _GEN_45068 = 6'h13 == rob_tail ? _T_5637_19 : _GEN_45067;
  assign _GEN_45069 = 6'h14 == rob_tail ? _T_5637_20 : _GEN_45068;
  assign _GEN_45070 = 6'h15 == rob_tail ? _T_5637_21 : _GEN_45069;
  assign _GEN_45071 = 6'h16 == rob_tail ? _T_5637_22 : _GEN_45070;
  assign _GEN_45072 = 6'h17 == rob_tail ? _T_5637_23 : _GEN_45071;
  assign _GEN_45073 = 6'h18 == rob_tail ? _T_5637_24 : _GEN_45072;
  assign _GEN_45074 = 6'h19 == rob_tail ? _T_5637_25 : _GEN_45073;
  assign _GEN_45075 = 6'h1a == rob_tail ? _T_5637_26 : _GEN_45074;
  assign _GEN_45076 = 6'h1b == rob_tail ? _T_5637_27 : _GEN_45075;
  assign _GEN_45077 = 6'h1c == rob_tail ? _T_5637_28 : _GEN_45076;
  assign _GEN_45078 = 6'h1d == rob_tail ? _T_5637_29 : _GEN_45077;
  assign _GEN_45079 = 6'h1e == rob_tail ? _T_5637_30 : _GEN_45078;
  assign _GEN_45080 = 6'h1f == rob_tail ? _T_5637_31 : _GEN_45079;
  assign _GEN_45081 = 6'h20 == rob_tail ? _T_5637_32 : _GEN_45080;
  assign _GEN_45082 = 6'h21 == rob_tail ? _T_5637_33 : _GEN_45081;
  assign _GEN_45083 = 6'h22 == rob_tail ? _T_5637_34 : _GEN_45082;
  assign _GEN_45084 = 6'h23 == rob_tail ? _T_5637_35 : _GEN_45083;
  assign _GEN_45085 = 6'h24 == rob_tail ? _T_5637_36 : _GEN_45084;
  assign _GEN_45086 = 6'h25 == rob_tail ? _T_5637_37 : _GEN_45085;
  assign _GEN_45087 = 6'h26 == rob_tail ? _T_5637_38 : _GEN_45086;
  assign _GEN_45088 = 6'h27 == rob_tail ? _T_5637_39 : _GEN_45087;
  assign _T_6349 = _GEN_320 == 1'h0;
  assign _T_6351 = _T_6349 | reset;
  assign _T_6353 = _T_6351 == 1'h0;
  assign _T_6354 = io_enq_uops_1_rob_idx[6:1];
  assign _T_6355 = _T_6354 == rob_tail;
  assign _T_6357 = _T_6355 | reset;
  assign _T_6359 = _T_6357 == 1'h0;
  assign _GEN_45169 = io_enq_valids_1 ? _GEN_41370 : _T_5637_0;
  assign _GEN_45170 = io_enq_valids_1 ? _GEN_41371 : _T_5637_1;
  assign _GEN_45171 = io_enq_valids_1 ? _GEN_41372 : _T_5637_2;
  assign _GEN_45172 = io_enq_valids_1 ? _GEN_41373 : _T_5637_3;
  assign _GEN_45173 = io_enq_valids_1 ? _GEN_41374 : _T_5637_4;
  assign _GEN_45174 = io_enq_valids_1 ? _GEN_41375 : _T_5637_5;
  assign _GEN_45175 = io_enq_valids_1 ? _GEN_41376 : _T_5637_6;
  assign _GEN_45176 = io_enq_valids_1 ? _GEN_41377 : _T_5637_7;
  assign _GEN_45177 = io_enq_valids_1 ? _GEN_41378 : _T_5637_8;
  assign _GEN_45178 = io_enq_valids_1 ? _GEN_41379 : _T_5637_9;
  assign _GEN_45179 = io_enq_valids_1 ? _GEN_41380 : _T_5637_10;
  assign _GEN_45180 = io_enq_valids_1 ? _GEN_41381 : _T_5637_11;
  assign _GEN_45181 = io_enq_valids_1 ? _GEN_41382 : _T_5637_12;
  assign _GEN_45182 = io_enq_valids_1 ? _GEN_41383 : _T_5637_13;
  assign _GEN_45183 = io_enq_valids_1 ? _GEN_41384 : _T_5637_14;
  assign _GEN_45184 = io_enq_valids_1 ? _GEN_41385 : _T_5637_15;
  assign _GEN_45185 = io_enq_valids_1 ? _GEN_41386 : _T_5637_16;
  assign _GEN_45186 = io_enq_valids_1 ? _GEN_41387 : _T_5637_17;
  assign _GEN_45187 = io_enq_valids_1 ? _GEN_41388 : _T_5637_18;
  assign _GEN_45188 = io_enq_valids_1 ? _GEN_41389 : _T_5637_19;
  assign _GEN_45189 = io_enq_valids_1 ? _GEN_41390 : _T_5637_20;
  assign _GEN_45190 = io_enq_valids_1 ? _GEN_41391 : _T_5637_21;
  assign _GEN_45191 = io_enq_valids_1 ? _GEN_41392 : _T_5637_22;
  assign _GEN_45192 = io_enq_valids_1 ? _GEN_41393 : _T_5637_23;
  assign _GEN_45193 = io_enq_valids_1 ? _GEN_41394 : _T_5637_24;
  assign _GEN_45194 = io_enq_valids_1 ? _GEN_41395 : _T_5637_25;
  assign _GEN_45195 = io_enq_valids_1 ? _GEN_41396 : _T_5637_26;
  assign _GEN_45196 = io_enq_valids_1 ? _GEN_41397 : _T_5637_27;
  assign _GEN_45197 = io_enq_valids_1 ? _GEN_41398 : _T_5637_28;
  assign _GEN_45198 = io_enq_valids_1 ? _GEN_41399 : _T_5637_29;
  assign _GEN_45199 = io_enq_valids_1 ? _GEN_41400 : _T_5637_30;
  assign _GEN_45200 = io_enq_valids_1 ? _GEN_41401 : _T_5637_31;
  assign _GEN_45201 = io_enq_valids_1 ? _GEN_41402 : _T_5637_32;
  assign _GEN_45202 = io_enq_valids_1 ? _GEN_41403 : _T_5637_33;
  assign _GEN_45203 = io_enq_valids_1 ? _GEN_41404 : _T_5637_34;
  assign _GEN_45204 = io_enq_valids_1 ? _GEN_41405 : _T_5637_35;
  assign _GEN_45205 = io_enq_valids_1 ? _GEN_41406 : _T_5637_36;
  assign _GEN_45206 = io_enq_valids_1 ? _GEN_41407 : _T_5637_37;
  assign _GEN_45207 = io_enq_valids_1 ? _GEN_41408 : _T_5637_38;
  assign _GEN_45208 = io_enq_valids_1 ? _GEN_41409 : _T_5637_39;
  assign _GEN_46173 = io_enq_valids_1 ? _GEN_42370 : _T_5936_0_br_mask;
  assign _GEN_46174 = io_enq_valids_1 ? _GEN_42371 : _T_5936_1_br_mask;
  assign _GEN_46175 = io_enq_valids_1 ? _GEN_42372 : _T_5936_2_br_mask;
  assign _GEN_46176 = io_enq_valids_1 ? _GEN_42373 : _T_5936_3_br_mask;
  assign _GEN_46177 = io_enq_valids_1 ? _GEN_42374 : _T_5936_4_br_mask;
  assign _GEN_46178 = io_enq_valids_1 ? _GEN_42375 : _T_5936_5_br_mask;
  assign _GEN_46179 = io_enq_valids_1 ? _GEN_42376 : _T_5936_6_br_mask;
  assign _GEN_46180 = io_enq_valids_1 ? _GEN_42377 : _T_5936_7_br_mask;
  assign _GEN_46181 = io_enq_valids_1 ? _GEN_42378 : _T_5936_8_br_mask;
  assign _GEN_46182 = io_enq_valids_1 ? _GEN_42379 : _T_5936_9_br_mask;
  assign _GEN_46183 = io_enq_valids_1 ? _GEN_42380 : _T_5936_10_br_mask;
  assign _GEN_46184 = io_enq_valids_1 ? _GEN_42381 : _T_5936_11_br_mask;
  assign _GEN_46185 = io_enq_valids_1 ? _GEN_42382 : _T_5936_12_br_mask;
  assign _GEN_46186 = io_enq_valids_1 ? _GEN_42383 : _T_5936_13_br_mask;
  assign _GEN_46187 = io_enq_valids_1 ? _GEN_42384 : _T_5936_14_br_mask;
  assign _GEN_46188 = io_enq_valids_1 ? _GEN_42385 : _T_5936_15_br_mask;
  assign _GEN_46189 = io_enq_valids_1 ? _GEN_42386 : _T_5936_16_br_mask;
  assign _GEN_46190 = io_enq_valids_1 ? _GEN_42387 : _T_5936_17_br_mask;
  assign _GEN_46191 = io_enq_valids_1 ? _GEN_42388 : _T_5936_18_br_mask;
  assign _GEN_46192 = io_enq_valids_1 ? _GEN_42389 : _T_5936_19_br_mask;
  assign _GEN_46193 = io_enq_valids_1 ? _GEN_42390 : _T_5936_20_br_mask;
  assign _GEN_46194 = io_enq_valids_1 ? _GEN_42391 : _T_5936_21_br_mask;
  assign _GEN_46195 = io_enq_valids_1 ? _GEN_42392 : _T_5936_22_br_mask;
  assign _GEN_46196 = io_enq_valids_1 ? _GEN_42393 : _T_5936_23_br_mask;
  assign _GEN_46197 = io_enq_valids_1 ? _GEN_42394 : _T_5936_24_br_mask;
  assign _GEN_46198 = io_enq_valids_1 ? _GEN_42395 : _T_5936_25_br_mask;
  assign _GEN_46199 = io_enq_valids_1 ? _GEN_42396 : _T_5936_26_br_mask;
  assign _GEN_46200 = io_enq_valids_1 ? _GEN_42397 : _T_5936_27_br_mask;
  assign _GEN_46201 = io_enq_valids_1 ? _GEN_42398 : _T_5936_28_br_mask;
  assign _GEN_46202 = io_enq_valids_1 ? _GEN_42399 : _T_5936_29_br_mask;
  assign _GEN_46203 = io_enq_valids_1 ? _GEN_42400 : _T_5936_30_br_mask;
  assign _GEN_46204 = io_enq_valids_1 ? _GEN_42401 : _T_5936_31_br_mask;
  assign _GEN_46205 = io_enq_valids_1 ? _GEN_42402 : _T_5936_32_br_mask;
  assign _GEN_46206 = io_enq_valids_1 ? _GEN_42403 : _T_5936_33_br_mask;
  assign _GEN_46207 = io_enq_valids_1 ? _GEN_42404 : _T_5936_34_br_mask;
  assign _GEN_46208 = io_enq_valids_1 ? _GEN_42405 : _T_5936_35_br_mask;
  assign _GEN_46209 = io_enq_valids_1 ? _GEN_42406 : _T_5936_36_br_mask;
  assign _GEN_46210 = io_enq_valids_1 ? _GEN_42407 : _T_5936_37_br_mask;
  assign _GEN_46211 = io_enq_valids_1 ? _GEN_42408 : _T_5936_38_br_mask;
  assign _GEN_46212 = io_enq_valids_1 ? _GEN_42409 : _T_5936_39_br_mask;
  assign _GEN_47293 = io_enq_valids_1 ? _GEN_43490 : _T_5936_0_pdst;
  assign _GEN_47294 = io_enq_valids_1 ? _GEN_43491 : _T_5936_1_pdst;
  assign _GEN_47295 = io_enq_valids_1 ? _GEN_43492 : _T_5936_2_pdst;
  assign _GEN_47296 = io_enq_valids_1 ? _GEN_43493 : _T_5936_3_pdst;
  assign _GEN_47297 = io_enq_valids_1 ? _GEN_43494 : _T_5936_4_pdst;
  assign _GEN_47298 = io_enq_valids_1 ? _GEN_43495 : _T_5936_5_pdst;
  assign _GEN_47299 = io_enq_valids_1 ? _GEN_43496 : _T_5936_6_pdst;
  assign _GEN_47300 = io_enq_valids_1 ? _GEN_43497 : _T_5936_7_pdst;
  assign _GEN_47301 = io_enq_valids_1 ? _GEN_43498 : _T_5936_8_pdst;
  assign _GEN_47302 = io_enq_valids_1 ? _GEN_43499 : _T_5936_9_pdst;
  assign _GEN_47303 = io_enq_valids_1 ? _GEN_43500 : _T_5936_10_pdst;
  assign _GEN_47304 = io_enq_valids_1 ? _GEN_43501 : _T_5936_11_pdst;
  assign _GEN_47305 = io_enq_valids_1 ? _GEN_43502 : _T_5936_12_pdst;
  assign _GEN_47306 = io_enq_valids_1 ? _GEN_43503 : _T_5936_13_pdst;
  assign _GEN_47307 = io_enq_valids_1 ? _GEN_43504 : _T_5936_14_pdst;
  assign _GEN_47308 = io_enq_valids_1 ? _GEN_43505 : _T_5936_15_pdst;
  assign _GEN_47309 = io_enq_valids_1 ? _GEN_43506 : _T_5936_16_pdst;
  assign _GEN_47310 = io_enq_valids_1 ? _GEN_43507 : _T_5936_17_pdst;
  assign _GEN_47311 = io_enq_valids_1 ? _GEN_43508 : _T_5936_18_pdst;
  assign _GEN_47312 = io_enq_valids_1 ? _GEN_43509 : _T_5936_19_pdst;
  assign _GEN_47313 = io_enq_valids_1 ? _GEN_43510 : _T_5936_20_pdst;
  assign _GEN_47314 = io_enq_valids_1 ? _GEN_43511 : _T_5936_21_pdst;
  assign _GEN_47315 = io_enq_valids_1 ? _GEN_43512 : _T_5936_22_pdst;
  assign _GEN_47316 = io_enq_valids_1 ? _GEN_43513 : _T_5936_23_pdst;
  assign _GEN_47317 = io_enq_valids_1 ? _GEN_43514 : _T_5936_24_pdst;
  assign _GEN_47318 = io_enq_valids_1 ? _GEN_43515 : _T_5936_25_pdst;
  assign _GEN_47319 = io_enq_valids_1 ? _GEN_43516 : _T_5936_26_pdst;
  assign _GEN_47320 = io_enq_valids_1 ? _GEN_43517 : _T_5936_27_pdst;
  assign _GEN_47321 = io_enq_valids_1 ? _GEN_43518 : _T_5936_28_pdst;
  assign _GEN_47322 = io_enq_valids_1 ? _GEN_43519 : _T_5936_29_pdst;
  assign _GEN_47323 = io_enq_valids_1 ? _GEN_43520 : _T_5936_30_pdst;
  assign _GEN_47324 = io_enq_valids_1 ? _GEN_43521 : _T_5936_31_pdst;
  assign _GEN_47325 = io_enq_valids_1 ? _GEN_43522 : _T_5936_32_pdst;
  assign _GEN_47326 = io_enq_valids_1 ? _GEN_43523 : _T_5936_33_pdst;
  assign _GEN_47327 = io_enq_valids_1 ? _GEN_43524 : _T_5936_34_pdst;
  assign _GEN_47328 = io_enq_valids_1 ? _GEN_43525 : _T_5936_35_pdst;
  assign _GEN_47329 = io_enq_valids_1 ? _GEN_43526 : _T_5936_36_pdst;
  assign _GEN_47330 = io_enq_valids_1 ? _GEN_43527 : _T_5936_37_pdst;
  assign _GEN_47331 = io_enq_valids_1 ? _GEN_43528 : _T_5936_38_pdst;
  assign _GEN_47332 = io_enq_valids_1 ? _GEN_43529 : _T_5936_39_pdst;
  assign _GEN_47573 = io_enq_valids_1 ? _GEN_43770 : _T_5936_0_stale_pdst;
  assign _GEN_47574 = io_enq_valids_1 ? _GEN_43771 : _T_5936_1_stale_pdst;
  assign _GEN_47575 = io_enq_valids_1 ? _GEN_43772 : _T_5936_2_stale_pdst;
  assign _GEN_47576 = io_enq_valids_1 ? _GEN_43773 : _T_5936_3_stale_pdst;
  assign _GEN_47577 = io_enq_valids_1 ? _GEN_43774 : _T_5936_4_stale_pdst;
  assign _GEN_47578 = io_enq_valids_1 ? _GEN_43775 : _T_5936_5_stale_pdst;
  assign _GEN_47579 = io_enq_valids_1 ? _GEN_43776 : _T_5936_6_stale_pdst;
  assign _GEN_47580 = io_enq_valids_1 ? _GEN_43777 : _T_5936_7_stale_pdst;
  assign _GEN_47581 = io_enq_valids_1 ? _GEN_43778 : _T_5936_8_stale_pdst;
  assign _GEN_47582 = io_enq_valids_1 ? _GEN_43779 : _T_5936_9_stale_pdst;
  assign _GEN_47583 = io_enq_valids_1 ? _GEN_43780 : _T_5936_10_stale_pdst;
  assign _GEN_47584 = io_enq_valids_1 ? _GEN_43781 : _T_5936_11_stale_pdst;
  assign _GEN_47585 = io_enq_valids_1 ? _GEN_43782 : _T_5936_12_stale_pdst;
  assign _GEN_47586 = io_enq_valids_1 ? _GEN_43783 : _T_5936_13_stale_pdst;
  assign _GEN_47587 = io_enq_valids_1 ? _GEN_43784 : _T_5936_14_stale_pdst;
  assign _GEN_47588 = io_enq_valids_1 ? _GEN_43785 : _T_5936_15_stale_pdst;
  assign _GEN_47589 = io_enq_valids_1 ? _GEN_43786 : _T_5936_16_stale_pdst;
  assign _GEN_47590 = io_enq_valids_1 ? _GEN_43787 : _T_5936_17_stale_pdst;
  assign _GEN_47591 = io_enq_valids_1 ? _GEN_43788 : _T_5936_18_stale_pdst;
  assign _GEN_47592 = io_enq_valids_1 ? _GEN_43789 : _T_5936_19_stale_pdst;
  assign _GEN_47593 = io_enq_valids_1 ? _GEN_43790 : _T_5936_20_stale_pdst;
  assign _GEN_47594 = io_enq_valids_1 ? _GEN_43791 : _T_5936_21_stale_pdst;
  assign _GEN_47595 = io_enq_valids_1 ? _GEN_43792 : _T_5936_22_stale_pdst;
  assign _GEN_47596 = io_enq_valids_1 ? _GEN_43793 : _T_5936_23_stale_pdst;
  assign _GEN_47597 = io_enq_valids_1 ? _GEN_43794 : _T_5936_24_stale_pdst;
  assign _GEN_47598 = io_enq_valids_1 ? _GEN_43795 : _T_5936_25_stale_pdst;
  assign _GEN_47599 = io_enq_valids_1 ? _GEN_43796 : _T_5936_26_stale_pdst;
  assign _GEN_47600 = io_enq_valids_1 ? _GEN_43797 : _T_5936_27_stale_pdst;
  assign _GEN_47601 = io_enq_valids_1 ? _GEN_43798 : _T_5936_28_stale_pdst;
  assign _GEN_47602 = io_enq_valids_1 ? _GEN_43799 : _T_5936_29_stale_pdst;
  assign _GEN_47603 = io_enq_valids_1 ? _GEN_43800 : _T_5936_30_stale_pdst;
  assign _GEN_47604 = io_enq_valids_1 ? _GEN_43801 : _T_5936_31_stale_pdst;
  assign _GEN_47605 = io_enq_valids_1 ? _GEN_43802 : _T_5936_32_stale_pdst;
  assign _GEN_47606 = io_enq_valids_1 ? _GEN_43803 : _T_5936_33_stale_pdst;
  assign _GEN_47607 = io_enq_valids_1 ? _GEN_43804 : _T_5936_34_stale_pdst;
  assign _GEN_47608 = io_enq_valids_1 ? _GEN_43805 : _T_5936_35_stale_pdst;
  assign _GEN_47609 = io_enq_valids_1 ? _GEN_43806 : _T_5936_36_stale_pdst;
  assign _GEN_47610 = io_enq_valids_1 ? _GEN_43807 : _T_5936_37_stale_pdst;
  assign _GEN_47611 = io_enq_valids_1 ? _GEN_43808 : _T_5936_38_stale_pdst;
  assign _GEN_47612 = io_enq_valids_1 ? _GEN_43809 : _T_5936_39_stale_pdst;
  assign _GEN_47853 = io_enq_valids_1 ? _GEN_44050 : _T_5936_0_is_fencei;
  assign _GEN_47854 = io_enq_valids_1 ? _GEN_44051 : _T_5936_1_is_fencei;
  assign _GEN_47855 = io_enq_valids_1 ? _GEN_44052 : _T_5936_2_is_fencei;
  assign _GEN_47856 = io_enq_valids_1 ? _GEN_44053 : _T_5936_3_is_fencei;
  assign _GEN_47857 = io_enq_valids_1 ? _GEN_44054 : _T_5936_4_is_fencei;
  assign _GEN_47858 = io_enq_valids_1 ? _GEN_44055 : _T_5936_5_is_fencei;
  assign _GEN_47859 = io_enq_valids_1 ? _GEN_44056 : _T_5936_6_is_fencei;
  assign _GEN_47860 = io_enq_valids_1 ? _GEN_44057 : _T_5936_7_is_fencei;
  assign _GEN_47861 = io_enq_valids_1 ? _GEN_44058 : _T_5936_8_is_fencei;
  assign _GEN_47862 = io_enq_valids_1 ? _GEN_44059 : _T_5936_9_is_fencei;
  assign _GEN_47863 = io_enq_valids_1 ? _GEN_44060 : _T_5936_10_is_fencei;
  assign _GEN_47864 = io_enq_valids_1 ? _GEN_44061 : _T_5936_11_is_fencei;
  assign _GEN_47865 = io_enq_valids_1 ? _GEN_44062 : _T_5936_12_is_fencei;
  assign _GEN_47866 = io_enq_valids_1 ? _GEN_44063 : _T_5936_13_is_fencei;
  assign _GEN_47867 = io_enq_valids_1 ? _GEN_44064 : _T_5936_14_is_fencei;
  assign _GEN_47868 = io_enq_valids_1 ? _GEN_44065 : _T_5936_15_is_fencei;
  assign _GEN_47869 = io_enq_valids_1 ? _GEN_44066 : _T_5936_16_is_fencei;
  assign _GEN_47870 = io_enq_valids_1 ? _GEN_44067 : _T_5936_17_is_fencei;
  assign _GEN_47871 = io_enq_valids_1 ? _GEN_44068 : _T_5936_18_is_fencei;
  assign _GEN_47872 = io_enq_valids_1 ? _GEN_44069 : _T_5936_19_is_fencei;
  assign _GEN_47873 = io_enq_valids_1 ? _GEN_44070 : _T_5936_20_is_fencei;
  assign _GEN_47874 = io_enq_valids_1 ? _GEN_44071 : _T_5936_21_is_fencei;
  assign _GEN_47875 = io_enq_valids_1 ? _GEN_44072 : _T_5936_22_is_fencei;
  assign _GEN_47876 = io_enq_valids_1 ? _GEN_44073 : _T_5936_23_is_fencei;
  assign _GEN_47877 = io_enq_valids_1 ? _GEN_44074 : _T_5936_24_is_fencei;
  assign _GEN_47878 = io_enq_valids_1 ? _GEN_44075 : _T_5936_25_is_fencei;
  assign _GEN_47879 = io_enq_valids_1 ? _GEN_44076 : _T_5936_26_is_fencei;
  assign _GEN_47880 = io_enq_valids_1 ? _GEN_44077 : _T_5936_27_is_fencei;
  assign _GEN_47881 = io_enq_valids_1 ? _GEN_44078 : _T_5936_28_is_fencei;
  assign _GEN_47882 = io_enq_valids_1 ? _GEN_44079 : _T_5936_29_is_fencei;
  assign _GEN_47883 = io_enq_valids_1 ? _GEN_44080 : _T_5936_30_is_fencei;
  assign _GEN_47884 = io_enq_valids_1 ? _GEN_44081 : _T_5936_31_is_fencei;
  assign _GEN_47885 = io_enq_valids_1 ? _GEN_44082 : _T_5936_32_is_fencei;
  assign _GEN_47886 = io_enq_valids_1 ? _GEN_44083 : _T_5936_33_is_fencei;
  assign _GEN_47887 = io_enq_valids_1 ? _GEN_44084 : _T_5936_34_is_fencei;
  assign _GEN_47888 = io_enq_valids_1 ? _GEN_44085 : _T_5936_35_is_fencei;
  assign _GEN_47889 = io_enq_valids_1 ? _GEN_44086 : _T_5936_36_is_fencei;
  assign _GEN_47890 = io_enq_valids_1 ? _GEN_44087 : _T_5936_37_is_fencei;
  assign _GEN_47891 = io_enq_valids_1 ? _GEN_44088 : _T_5936_38_is_fencei;
  assign _GEN_47892 = io_enq_valids_1 ? _GEN_44089 : _T_5936_39_is_fencei;
  assign _GEN_47893 = io_enq_valids_1 ? _GEN_44090 : _T_5936_0_is_store;
  assign _GEN_47894 = io_enq_valids_1 ? _GEN_44091 : _T_5936_1_is_store;
  assign _GEN_47895 = io_enq_valids_1 ? _GEN_44092 : _T_5936_2_is_store;
  assign _GEN_47896 = io_enq_valids_1 ? _GEN_44093 : _T_5936_3_is_store;
  assign _GEN_47897 = io_enq_valids_1 ? _GEN_44094 : _T_5936_4_is_store;
  assign _GEN_47898 = io_enq_valids_1 ? _GEN_44095 : _T_5936_5_is_store;
  assign _GEN_47899 = io_enq_valids_1 ? _GEN_44096 : _T_5936_6_is_store;
  assign _GEN_47900 = io_enq_valids_1 ? _GEN_44097 : _T_5936_7_is_store;
  assign _GEN_47901 = io_enq_valids_1 ? _GEN_44098 : _T_5936_8_is_store;
  assign _GEN_47902 = io_enq_valids_1 ? _GEN_44099 : _T_5936_9_is_store;
  assign _GEN_47903 = io_enq_valids_1 ? _GEN_44100 : _T_5936_10_is_store;
  assign _GEN_47904 = io_enq_valids_1 ? _GEN_44101 : _T_5936_11_is_store;
  assign _GEN_47905 = io_enq_valids_1 ? _GEN_44102 : _T_5936_12_is_store;
  assign _GEN_47906 = io_enq_valids_1 ? _GEN_44103 : _T_5936_13_is_store;
  assign _GEN_47907 = io_enq_valids_1 ? _GEN_44104 : _T_5936_14_is_store;
  assign _GEN_47908 = io_enq_valids_1 ? _GEN_44105 : _T_5936_15_is_store;
  assign _GEN_47909 = io_enq_valids_1 ? _GEN_44106 : _T_5936_16_is_store;
  assign _GEN_47910 = io_enq_valids_1 ? _GEN_44107 : _T_5936_17_is_store;
  assign _GEN_47911 = io_enq_valids_1 ? _GEN_44108 : _T_5936_18_is_store;
  assign _GEN_47912 = io_enq_valids_1 ? _GEN_44109 : _T_5936_19_is_store;
  assign _GEN_47913 = io_enq_valids_1 ? _GEN_44110 : _T_5936_20_is_store;
  assign _GEN_47914 = io_enq_valids_1 ? _GEN_44111 : _T_5936_21_is_store;
  assign _GEN_47915 = io_enq_valids_1 ? _GEN_44112 : _T_5936_22_is_store;
  assign _GEN_47916 = io_enq_valids_1 ? _GEN_44113 : _T_5936_23_is_store;
  assign _GEN_47917 = io_enq_valids_1 ? _GEN_44114 : _T_5936_24_is_store;
  assign _GEN_47918 = io_enq_valids_1 ? _GEN_44115 : _T_5936_25_is_store;
  assign _GEN_47919 = io_enq_valids_1 ? _GEN_44116 : _T_5936_26_is_store;
  assign _GEN_47920 = io_enq_valids_1 ? _GEN_44117 : _T_5936_27_is_store;
  assign _GEN_47921 = io_enq_valids_1 ? _GEN_44118 : _T_5936_28_is_store;
  assign _GEN_47922 = io_enq_valids_1 ? _GEN_44119 : _T_5936_29_is_store;
  assign _GEN_47923 = io_enq_valids_1 ? _GEN_44120 : _T_5936_30_is_store;
  assign _GEN_47924 = io_enq_valids_1 ? _GEN_44121 : _T_5936_31_is_store;
  assign _GEN_47925 = io_enq_valids_1 ? _GEN_44122 : _T_5936_32_is_store;
  assign _GEN_47926 = io_enq_valids_1 ? _GEN_44123 : _T_5936_33_is_store;
  assign _GEN_47927 = io_enq_valids_1 ? _GEN_44124 : _T_5936_34_is_store;
  assign _GEN_47928 = io_enq_valids_1 ? _GEN_44125 : _T_5936_35_is_store;
  assign _GEN_47929 = io_enq_valids_1 ? _GEN_44126 : _T_5936_36_is_store;
  assign _GEN_47930 = io_enq_valids_1 ? _GEN_44127 : _T_5936_37_is_store;
  assign _GEN_47931 = io_enq_valids_1 ? _GEN_44128 : _T_5936_38_is_store;
  assign _GEN_47932 = io_enq_valids_1 ? _GEN_44129 : _T_5936_39_is_store;
  assign _GEN_47973 = io_enq_valids_1 ? _GEN_44170 : _T_5936_0_is_load;
  assign _GEN_47974 = io_enq_valids_1 ? _GEN_44171 : _T_5936_1_is_load;
  assign _GEN_47975 = io_enq_valids_1 ? _GEN_44172 : _T_5936_2_is_load;
  assign _GEN_47976 = io_enq_valids_1 ? _GEN_44173 : _T_5936_3_is_load;
  assign _GEN_47977 = io_enq_valids_1 ? _GEN_44174 : _T_5936_4_is_load;
  assign _GEN_47978 = io_enq_valids_1 ? _GEN_44175 : _T_5936_5_is_load;
  assign _GEN_47979 = io_enq_valids_1 ? _GEN_44176 : _T_5936_6_is_load;
  assign _GEN_47980 = io_enq_valids_1 ? _GEN_44177 : _T_5936_7_is_load;
  assign _GEN_47981 = io_enq_valids_1 ? _GEN_44178 : _T_5936_8_is_load;
  assign _GEN_47982 = io_enq_valids_1 ? _GEN_44179 : _T_5936_9_is_load;
  assign _GEN_47983 = io_enq_valids_1 ? _GEN_44180 : _T_5936_10_is_load;
  assign _GEN_47984 = io_enq_valids_1 ? _GEN_44181 : _T_5936_11_is_load;
  assign _GEN_47985 = io_enq_valids_1 ? _GEN_44182 : _T_5936_12_is_load;
  assign _GEN_47986 = io_enq_valids_1 ? _GEN_44183 : _T_5936_13_is_load;
  assign _GEN_47987 = io_enq_valids_1 ? _GEN_44184 : _T_5936_14_is_load;
  assign _GEN_47988 = io_enq_valids_1 ? _GEN_44185 : _T_5936_15_is_load;
  assign _GEN_47989 = io_enq_valids_1 ? _GEN_44186 : _T_5936_16_is_load;
  assign _GEN_47990 = io_enq_valids_1 ? _GEN_44187 : _T_5936_17_is_load;
  assign _GEN_47991 = io_enq_valids_1 ? _GEN_44188 : _T_5936_18_is_load;
  assign _GEN_47992 = io_enq_valids_1 ? _GEN_44189 : _T_5936_19_is_load;
  assign _GEN_47993 = io_enq_valids_1 ? _GEN_44190 : _T_5936_20_is_load;
  assign _GEN_47994 = io_enq_valids_1 ? _GEN_44191 : _T_5936_21_is_load;
  assign _GEN_47995 = io_enq_valids_1 ? _GEN_44192 : _T_5936_22_is_load;
  assign _GEN_47996 = io_enq_valids_1 ? _GEN_44193 : _T_5936_23_is_load;
  assign _GEN_47997 = io_enq_valids_1 ? _GEN_44194 : _T_5936_24_is_load;
  assign _GEN_47998 = io_enq_valids_1 ? _GEN_44195 : _T_5936_25_is_load;
  assign _GEN_47999 = io_enq_valids_1 ? _GEN_44196 : _T_5936_26_is_load;
  assign _GEN_48000 = io_enq_valids_1 ? _GEN_44197 : _T_5936_27_is_load;
  assign _GEN_48001 = io_enq_valids_1 ? _GEN_44198 : _T_5936_28_is_load;
  assign _GEN_48002 = io_enq_valids_1 ? _GEN_44199 : _T_5936_29_is_load;
  assign _GEN_48003 = io_enq_valids_1 ? _GEN_44200 : _T_5936_30_is_load;
  assign _GEN_48004 = io_enq_valids_1 ? _GEN_44201 : _T_5936_31_is_load;
  assign _GEN_48005 = io_enq_valids_1 ? _GEN_44202 : _T_5936_32_is_load;
  assign _GEN_48006 = io_enq_valids_1 ? _GEN_44203 : _T_5936_33_is_load;
  assign _GEN_48007 = io_enq_valids_1 ? _GEN_44204 : _T_5936_34_is_load;
  assign _GEN_48008 = io_enq_valids_1 ? _GEN_44205 : _T_5936_35_is_load;
  assign _GEN_48009 = io_enq_valids_1 ? _GEN_44206 : _T_5936_36_is_load;
  assign _GEN_48010 = io_enq_valids_1 ? _GEN_44207 : _T_5936_37_is_load;
  assign _GEN_48011 = io_enq_valids_1 ? _GEN_44208 : _T_5936_38_is_load;
  assign _GEN_48012 = io_enq_valids_1 ? _GEN_44209 : _T_5936_39_is_load;
  assign _GEN_48013 = io_enq_valids_1 ? _GEN_44210 : _T_5936_0_is_sys_pc2epc;
  assign _GEN_48014 = io_enq_valids_1 ? _GEN_44211 : _T_5936_1_is_sys_pc2epc;
  assign _GEN_48015 = io_enq_valids_1 ? _GEN_44212 : _T_5936_2_is_sys_pc2epc;
  assign _GEN_48016 = io_enq_valids_1 ? _GEN_44213 : _T_5936_3_is_sys_pc2epc;
  assign _GEN_48017 = io_enq_valids_1 ? _GEN_44214 : _T_5936_4_is_sys_pc2epc;
  assign _GEN_48018 = io_enq_valids_1 ? _GEN_44215 : _T_5936_5_is_sys_pc2epc;
  assign _GEN_48019 = io_enq_valids_1 ? _GEN_44216 : _T_5936_6_is_sys_pc2epc;
  assign _GEN_48020 = io_enq_valids_1 ? _GEN_44217 : _T_5936_7_is_sys_pc2epc;
  assign _GEN_48021 = io_enq_valids_1 ? _GEN_44218 : _T_5936_8_is_sys_pc2epc;
  assign _GEN_48022 = io_enq_valids_1 ? _GEN_44219 : _T_5936_9_is_sys_pc2epc;
  assign _GEN_48023 = io_enq_valids_1 ? _GEN_44220 : _T_5936_10_is_sys_pc2epc;
  assign _GEN_48024 = io_enq_valids_1 ? _GEN_44221 : _T_5936_11_is_sys_pc2epc;
  assign _GEN_48025 = io_enq_valids_1 ? _GEN_44222 : _T_5936_12_is_sys_pc2epc;
  assign _GEN_48026 = io_enq_valids_1 ? _GEN_44223 : _T_5936_13_is_sys_pc2epc;
  assign _GEN_48027 = io_enq_valids_1 ? _GEN_44224 : _T_5936_14_is_sys_pc2epc;
  assign _GEN_48028 = io_enq_valids_1 ? _GEN_44225 : _T_5936_15_is_sys_pc2epc;
  assign _GEN_48029 = io_enq_valids_1 ? _GEN_44226 : _T_5936_16_is_sys_pc2epc;
  assign _GEN_48030 = io_enq_valids_1 ? _GEN_44227 : _T_5936_17_is_sys_pc2epc;
  assign _GEN_48031 = io_enq_valids_1 ? _GEN_44228 : _T_5936_18_is_sys_pc2epc;
  assign _GEN_48032 = io_enq_valids_1 ? _GEN_44229 : _T_5936_19_is_sys_pc2epc;
  assign _GEN_48033 = io_enq_valids_1 ? _GEN_44230 : _T_5936_20_is_sys_pc2epc;
  assign _GEN_48034 = io_enq_valids_1 ? _GEN_44231 : _T_5936_21_is_sys_pc2epc;
  assign _GEN_48035 = io_enq_valids_1 ? _GEN_44232 : _T_5936_22_is_sys_pc2epc;
  assign _GEN_48036 = io_enq_valids_1 ? _GEN_44233 : _T_5936_23_is_sys_pc2epc;
  assign _GEN_48037 = io_enq_valids_1 ? _GEN_44234 : _T_5936_24_is_sys_pc2epc;
  assign _GEN_48038 = io_enq_valids_1 ? _GEN_44235 : _T_5936_25_is_sys_pc2epc;
  assign _GEN_48039 = io_enq_valids_1 ? _GEN_44236 : _T_5936_26_is_sys_pc2epc;
  assign _GEN_48040 = io_enq_valids_1 ? _GEN_44237 : _T_5936_27_is_sys_pc2epc;
  assign _GEN_48041 = io_enq_valids_1 ? _GEN_44238 : _T_5936_28_is_sys_pc2epc;
  assign _GEN_48042 = io_enq_valids_1 ? _GEN_44239 : _T_5936_29_is_sys_pc2epc;
  assign _GEN_48043 = io_enq_valids_1 ? _GEN_44240 : _T_5936_30_is_sys_pc2epc;
  assign _GEN_48044 = io_enq_valids_1 ? _GEN_44241 : _T_5936_31_is_sys_pc2epc;
  assign _GEN_48045 = io_enq_valids_1 ? _GEN_44242 : _T_5936_32_is_sys_pc2epc;
  assign _GEN_48046 = io_enq_valids_1 ? _GEN_44243 : _T_5936_33_is_sys_pc2epc;
  assign _GEN_48047 = io_enq_valids_1 ? _GEN_44244 : _T_5936_34_is_sys_pc2epc;
  assign _GEN_48048 = io_enq_valids_1 ? _GEN_44245 : _T_5936_35_is_sys_pc2epc;
  assign _GEN_48049 = io_enq_valids_1 ? _GEN_44246 : _T_5936_36_is_sys_pc2epc;
  assign _GEN_48050 = io_enq_valids_1 ? _GEN_44247 : _T_5936_37_is_sys_pc2epc;
  assign _GEN_48051 = io_enq_valids_1 ? _GEN_44248 : _T_5936_38_is_sys_pc2epc;
  assign _GEN_48052 = io_enq_valids_1 ? _GEN_44249 : _T_5936_39_is_sys_pc2epc;
  assign _GEN_48093 = io_enq_valids_1 ? _GEN_44290 : _T_5936_0_flush_on_commit;
  assign _GEN_48094 = io_enq_valids_1 ? _GEN_44291 : _T_5936_1_flush_on_commit;
  assign _GEN_48095 = io_enq_valids_1 ? _GEN_44292 : _T_5936_2_flush_on_commit;
  assign _GEN_48096 = io_enq_valids_1 ? _GEN_44293 : _T_5936_3_flush_on_commit;
  assign _GEN_48097 = io_enq_valids_1 ? _GEN_44294 : _T_5936_4_flush_on_commit;
  assign _GEN_48098 = io_enq_valids_1 ? _GEN_44295 : _T_5936_5_flush_on_commit;
  assign _GEN_48099 = io_enq_valids_1 ? _GEN_44296 : _T_5936_6_flush_on_commit;
  assign _GEN_48100 = io_enq_valids_1 ? _GEN_44297 : _T_5936_7_flush_on_commit;
  assign _GEN_48101 = io_enq_valids_1 ? _GEN_44298 : _T_5936_8_flush_on_commit;
  assign _GEN_48102 = io_enq_valids_1 ? _GEN_44299 : _T_5936_9_flush_on_commit;
  assign _GEN_48103 = io_enq_valids_1 ? _GEN_44300 : _T_5936_10_flush_on_commit;
  assign _GEN_48104 = io_enq_valids_1 ? _GEN_44301 : _T_5936_11_flush_on_commit;
  assign _GEN_48105 = io_enq_valids_1 ? _GEN_44302 : _T_5936_12_flush_on_commit;
  assign _GEN_48106 = io_enq_valids_1 ? _GEN_44303 : _T_5936_13_flush_on_commit;
  assign _GEN_48107 = io_enq_valids_1 ? _GEN_44304 : _T_5936_14_flush_on_commit;
  assign _GEN_48108 = io_enq_valids_1 ? _GEN_44305 : _T_5936_15_flush_on_commit;
  assign _GEN_48109 = io_enq_valids_1 ? _GEN_44306 : _T_5936_16_flush_on_commit;
  assign _GEN_48110 = io_enq_valids_1 ? _GEN_44307 : _T_5936_17_flush_on_commit;
  assign _GEN_48111 = io_enq_valids_1 ? _GEN_44308 : _T_5936_18_flush_on_commit;
  assign _GEN_48112 = io_enq_valids_1 ? _GEN_44309 : _T_5936_19_flush_on_commit;
  assign _GEN_48113 = io_enq_valids_1 ? _GEN_44310 : _T_5936_20_flush_on_commit;
  assign _GEN_48114 = io_enq_valids_1 ? _GEN_44311 : _T_5936_21_flush_on_commit;
  assign _GEN_48115 = io_enq_valids_1 ? _GEN_44312 : _T_5936_22_flush_on_commit;
  assign _GEN_48116 = io_enq_valids_1 ? _GEN_44313 : _T_5936_23_flush_on_commit;
  assign _GEN_48117 = io_enq_valids_1 ? _GEN_44314 : _T_5936_24_flush_on_commit;
  assign _GEN_48118 = io_enq_valids_1 ? _GEN_44315 : _T_5936_25_flush_on_commit;
  assign _GEN_48119 = io_enq_valids_1 ? _GEN_44316 : _T_5936_26_flush_on_commit;
  assign _GEN_48120 = io_enq_valids_1 ? _GEN_44317 : _T_5936_27_flush_on_commit;
  assign _GEN_48121 = io_enq_valids_1 ? _GEN_44318 : _T_5936_28_flush_on_commit;
  assign _GEN_48122 = io_enq_valids_1 ? _GEN_44319 : _T_5936_29_flush_on_commit;
  assign _GEN_48123 = io_enq_valids_1 ? _GEN_44320 : _T_5936_30_flush_on_commit;
  assign _GEN_48124 = io_enq_valids_1 ? _GEN_44321 : _T_5936_31_flush_on_commit;
  assign _GEN_48125 = io_enq_valids_1 ? _GEN_44322 : _T_5936_32_flush_on_commit;
  assign _GEN_48126 = io_enq_valids_1 ? _GEN_44323 : _T_5936_33_flush_on_commit;
  assign _GEN_48127 = io_enq_valids_1 ? _GEN_44324 : _T_5936_34_flush_on_commit;
  assign _GEN_48128 = io_enq_valids_1 ? _GEN_44325 : _T_5936_35_flush_on_commit;
  assign _GEN_48129 = io_enq_valids_1 ? _GEN_44326 : _T_5936_36_flush_on_commit;
  assign _GEN_48130 = io_enq_valids_1 ? _GEN_44327 : _T_5936_37_flush_on_commit;
  assign _GEN_48131 = io_enq_valids_1 ? _GEN_44328 : _T_5936_38_flush_on_commit;
  assign _GEN_48132 = io_enq_valids_1 ? _GEN_44329 : _T_5936_39_flush_on_commit;
  assign _GEN_48133 = io_enq_valids_1 ? _GEN_44330 : _T_5936_0_ldst;
  assign _GEN_48134 = io_enq_valids_1 ? _GEN_44331 : _T_5936_1_ldst;
  assign _GEN_48135 = io_enq_valids_1 ? _GEN_44332 : _T_5936_2_ldst;
  assign _GEN_48136 = io_enq_valids_1 ? _GEN_44333 : _T_5936_3_ldst;
  assign _GEN_48137 = io_enq_valids_1 ? _GEN_44334 : _T_5936_4_ldst;
  assign _GEN_48138 = io_enq_valids_1 ? _GEN_44335 : _T_5936_5_ldst;
  assign _GEN_48139 = io_enq_valids_1 ? _GEN_44336 : _T_5936_6_ldst;
  assign _GEN_48140 = io_enq_valids_1 ? _GEN_44337 : _T_5936_7_ldst;
  assign _GEN_48141 = io_enq_valids_1 ? _GEN_44338 : _T_5936_8_ldst;
  assign _GEN_48142 = io_enq_valids_1 ? _GEN_44339 : _T_5936_9_ldst;
  assign _GEN_48143 = io_enq_valids_1 ? _GEN_44340 : _T_5936_10_ldst;
  assign _GEN_48144 = io_enq_valids_1 ? _GEN_44341 : _T_5936_11_ldst;
  assign _GEN_48145 = io_enq_valids_1 ? _GEN_44342 : _T_5936_12_ldst;
  assign _GEN_48146 = io_enq_valids_1 ? _GEN_44343 : _T_5936_13_ldst;
  assign _GEN_48147 = io_enq_valids_1 ? _GEN_44344 : _T_5936_14_ldst;
  assign _GEN_48148 = io_enq_valids_1 ? _GEN_44345 : _T_5936_15_ldst;
  assign _GEN_48149 = io_enq_valids_1 ? _GEN_44346 : _T_5936_16_ldst;
  assign _GEN_48150 = io_enq_valids_1 ? _GEN_44347 : _T_5936_17_ldst;
  assign _GEN_48151 = io_enq_valids_1 ? _GEN_44348 : _T_5936_18_ldst;
  assign _GEN_48152 = io_enq_valids_1 ? _GEN_44349 : _T_5936_19_ldst;
  assign _GEN_48153 = io_enq_valids_1 ? _GEN_44350 : _T_5936_20_ldst;
  assign _GEN_48154 = io_enq_valids_1 ? _GEN_44351 : _T_5936_21_ldst;
  assign _GEN_48155 = io_enq_valids_1 ? _GEN_44352 : _T_5936_22_ldst;
  assign _GEN_48156 = io_enq_valids_1 ? _GEN_44353 : _T_5936_23_ldst;
  assign _GEN_48157 = io_enq_valids_1 ? _GEN_44354 : _T_5936_24_ldst;
  assign _GEN_48158 = io_enq_valids_1 ? _GEN_44355 : _T_5936_25_ldst;
  assign _GEN_48159 = io_enq_valids_1 ? _GEN_44356 : _T_5936_26_ldst;
  assign _GEN_48160 = io_enq_valids_1 ? _GEN_44357 : _T_5936_27_ldst;
  assign _GEN_48161 = io_enq_valids_1 ? _GEN_44358 : _T_5936_28_ldst;
  assign _GEN_48162 = io_enq_valids_1 ? _GEN_44359 : _T_5936_29_ldst;
  assign _GEN_48163 = io_enq_valids_1 ? _GEN_44360 : _T_5936_30_ldst;
  assign _GEN_48164 = io_enq_valids_1 ? _GEN_44361 : _T_5936_31_ldst;
  assign _GEN_48165 = io_enq_valids_1 ? _GEN_44362 : _T_5936_32_ldst;
  assign _GEN_48166 = io_enq_valids_1 ? _GEN_44363 : _T_5936_33_ldst;
  assign _GEN_48167 = io_enq_valids_1 ? _GEN_44364 : _T_5936_34_ldst;
  assign _GEN_48168 = io_enq_valids_1 ? _GEN_44365 : _T_5936_35_ldst;
  assign _GEN_48169 = io_enq_valids_1 ? _GEN_44366 : _T_5936_36_ldst;
  assign _GEN_48170 = io_enq_valids_1 ? _GEN_44367 : _T_5936_37_ldst;
  assign _GEN_48171 = io_enq_valids_1 ? _GEN_44368 : _T_5936_38_ldst;
  assign _GEN_48172 = io_enq_valids_1 ? _GEN_44369 : _T_5936_39_ldst;
  assign _GEN_48293 = io_enq_valids_1 ? _GEN_44490 : _T_5936_0_ldst_val;
  assign _GEN_48294 = io_enq_valids_1 ? _GEN_44491 : _T_5936_1_ldst_val;
  assign _GEN_48295 = io_enq_valids_1 ? _GEN_44492 : _T_5936_2_ldst_val;
  assign _GEN_48296 = io_enq_valids_1 ? _GEN_44493 : _T_5936_3_ldst_val;
  assign _GEN_48297 = io_enq_valids_1 ? _GEN_44494 : _T_5936_4_ldst_val;
  assign _GEN_48298 = io_enq_valids_1 ? _GEN_44495 : _T_5936_5_ldst_val;
  assign _GEN_48299 = io_enq_valids_1 ? _GEN_44496 : _T_5936_6_ldst_val;
  assign _GEN_48300 = io_enq_valids_1 ? _GEN_44497 : _T_5936_7_ldst_val;
  assign _GEN_48301 = io_enq_valids_1 ? _GEN_44498 : _T_5936_8_ldst_val;
  assign _GEN_48302 = io_enq_valids_1 ? _GEN_44499 : _T_5936_9_ldst_val;
  assign _GEN_48303 = io_enq_valids_1 ? _GEN_44500 : _T_5936_10_ldst_val;
  assign _GEN_48304 = io_enq_valids_1 ? _GEN_44501 : _T_5936_11_ldst_val;
  assign _GEN_48305 = io_enq_valids_1 ? _GEN_44502 : _T_5936_12_ldst_val;
  assign _GEN_48306 = io_enq_valids_1 ? _GEN_44503 : _T_5936_13_ldst_val;
  assign _GEN_48307 = io_enq_valids_1 ? _GEN_44504 : _T_5936_14_ldst_val;
  assign _GEN_48308 = io_enq_valids_1 ? _GEN_44505 : _T_5936_15_ldst_val;
  assign _GEN_48309 = io_enq_valids_1 ? _GEN_44506 : _T_5936_16_ldst_val;
  assign _GEN_48310 = io_enq_valids_1 ? _GEN_44507 : _T_5936_17_ldst_val;
  assign _GEN_48311 = io_enq_valids_1 ? _GEN_44508 : _T_5936_18_ldst_val;
  assign _GEN_48312 = io_enq_valids_1 ? _GEN_44509 : _T_5936_19_ldst_val;
  assign _GEN_48313 = io_enq_valids_1 ? _GEN_44510 : _T_5936_20_ldst_val;
  assign _GEN_48314 = io_enq_valids_1 ? _GEN_44511 : _T_5936_21_ldst_val;
  assign _GEN_48315 = io_enq_valids_1 ? _GEN_44512 : _T_5936_22_ldst_val;
  assign _GEN_48316 = io_enq_valids_1 ? _GEN_44513 : _T_5936_23_ldst_val;
  assign _GEN_48317 = io_enq_valids_1 ? _GEN_44514 : _T_5936_24_ldst_val;
  assign _GEN_48318 = io_enq_valids_1 ? _GEN_44515 : _T_5936_25_ldst_val;
  assign _GEN_48319 = io_enq_valids_1 ? _GEN_44516 : _T_5936_26_ldst_val;
  assign _GEN_48320 = io_enq_valids_1 ? _GEN_44517 : _T_5936_27_ldst_val;
  assign _GEN_48321 = io_enq_valids_1 ? _GEN_44518 : _T_5936_28_ldst_val;
  assign _GEN_48322 = io_enq_valids_1 ? _GEN_44519 : _T_5936_29_ldst_val;
  assign _GEN_48323 = io_enq_valids_1 ? _GEN_44520 : _T_5936_30_ldst_val;
  assign _GEN_48324 = io_enq_valids_1 ? _GEN_44521 : _T_5936_31_ldst_val;
  assign _GEN_48325 = io_enq_valids_1 ? _GEN_44522 : _T_5936_32_ldst_val;
  assign _GEN_48326 = io_enq_valids_1 ? _GEN_44523 : _T_5936_33_ldst_val;
  assign _GEN_48327 = io_enq_valids_1 ? _GEN_44524 : _T_5936_34_ldst_val;
  assign _GEN_48328 = io_enq_valids_1 ? _GEN_44525 : _T_5936_35_ldst_val;
  assign _GEN_48329 = io_enq_valids_1 ? _GEN_44526 : _T_5936_36_ldst_val;
  assign _GEN_48330 = io_enq_valids_1 ? _GEN_44527 : _T_5936_37_ldst_val;
  assign _GEN_48331 = io_enq_valids_1 ? _GEN_44528 : _T_5936_38_ldst_val;
  assign _GEN_48332 = io_enq_valids_1 ? _GEN_44529 : _T_5936_39_ldst_val;
  assign _GEN_48333 = io_enq_valids_1 ? _GEN_44530 : _T_5936_0_dst_rtype;
  assign _GEN_48334 = io_enq_valids_1 ? _GEN_44531 : _T_5936_1_dst_rtype;
  assign _GEN_48335 = io_enq_valids_1 ? _GEN_44532 : _T_5936_2_dst_rtype;
  assign _GEN_48336 = io_enq_valids_1 ? _GEN_44533 : _T_5936_3_dst_rtype;
  assign _GEN_48337 = io_enq_valids_1 ? _GEN_44534 : _T_5936_4_dst_rtype;
  assign _GEN_48338 = io_enq_valids_1 ? _GEN_44535 : _T_5936_5_dst_rtype;
  assign _GEN_48339 = io_enq_valids_1 ? _GEN_44536 : _T_5936_6_dst_rtype;
  assign _GEN_48340 = io_enq_valids_1 ? _GEN_44537 : _T_5936_7_dst_rtype;
  assign _GEN_48341 = io_enq_valids_1 ? _GEN_44538 : _T_5936_8_dst_rtype;
  assign _GEN_48342 = io_enq_valids_1 ? _GEN_44539 : _T_5936_9_dst_rtype;
  assign _GEN_48343 = io_enq_valids_1 ? _GEN_44540 : _T_5936_10_dst_rtype;
  assign _GEN_48344 = io_enq_valids_1 ? _GEN_44541 : _T_5936_11_dst_rtype;
  assign _GEN_48345 = io_enq_valids_1 ? _GEN_44542 : _T_5936_12_dst_rtype;
  assign _GEN_48346 = io_enq_valids_1 ? _GEN_44543 : _T_5936_13_dst_rtype;
  assign _GEN_48347 = io_enq_valids_1 ? _GEN_44544 : _T_5936_14_dst_rtype;
  assign _GEN_48348 = io_enq_valids_1 ? _GEN_44545 : _T_5936_15_dst_rtype;
  assign _GEN_48349 = io_enq_valids_1 ? _GEN_44546 : _T_5936_16_dst_rtype;
  assign _GEN_48350 = io_enq_valids_1 ? _GEN_44547 : _T_5936_17_dst_rtype;
  assign _GEN_48351 = io_enq_valids_1 ? _GEN_44548 : _T_5936_18_dst_rtype;
  assign _GEN_48352 = io_enq_valids_1 ? _GEN_44549 : _T_5936_19_dst_rtype;
  assign _GEN_48353 = io_enq_valids_1 ? _GEN_44550 : _T_5936_20_dst_rtype;
  assign _GEN_48354 = io_enq_valids_1 ? _GEN_44551 : _T_5936_21_dst_rtype;
  assign _GEN_48355 = io_enq_valids_1 ? _GEN_44552 : _T_5936_22_dst_rtype;
  assign _GEN_48356 = io_enq_valids_1 ? _GEN_44553 : _T_5936_23_dst_rtype;
  assign _GEN_48357 = io_enq_valids_1 ? _GEN_44554 : _T_5936_24_dst_rtype;
  assign _GEN_48358 = io_enq_valids_1 ? _GEN_44555 : _T_5936_25_dst_rtype;
  assign _GEN_48359 = io_enq_valids_1 ? _GEN_44556 : _T_5936_26_dst_rtype;
  assign _GEN_48360 = io_enq_valids_1 ? _GEN_44557 : _T_5936_27_dst_rtype;
  assign _GEN_48361 = io_enq_valids_1 ? _GEN_44558 : _T_5936_28_dst_rtype;
  assign _GEN_48362 = io_enq_valids_1 ? _GEN_44559 : _T_5936_29_dst_rtype;
  assign _GEN_48363 = io_enq_valids_1 ? _GEN_44560 : _T_5936_30_dst_rtype;
  assign _GEN_48364 = io_enq_valids_1 ? _GEN_44561 : _T_5936_31_dst_rtype;
  assign _GEN_48365 = io_enq_valids_1 ? _GEN_44562 : _T_5936_32_dst_rtype;
  assign _GEN_48366 = io_enq_valids_1 ? _GEN_44563 : _T_5936_33_dst_rtype;
  assign _GEN_48367 = io_enq_valids_1 ? _GEN_44564 : _T_5936_34_dst_rtype;
  assign _GEN_48368 = io_enq_valids_1 ? _GEN_44565 : _T_5936_35_dst_rtype;
  assign _GEN_48369 = io_enq_valids_1 ? _GEN_44566 : _T_5936_36_dst_rtype;
  assign _GEN_48370 = io_enq_valids_1 ? _GEN_44567 : _T_5936_37_dst_rtype;
  assign _GEN_48371 = io_enq_valids_1 ? _GEN_44568 : _T_5936_38_dst_rtype;
  assign _GEN_48372 = io_enq_valids_1 ? _GEN_44569 : _T_5936_39_dst_rtype;
  assign _GEN_48493 = io_enq_valids_1 ? _GEN_44690 : _T_5936_0_fp_val;
  assign _GEN_48494 = io_enq_valids_1 ? _GEN_44691 : _T_5936_1_fp_val;
  assign _GEN_48495 = io_enq_valids_1 ? _GEN_44692 : _T_5936_2_fp_val;
  assign _GEN_48496 = io_enq_valids_1 ? _GEN_44693 : _T_5936_3_fp_val;
  assign _GEN_48497 = io_enq_valids_1 ? _GEN_44694 : _T_5936_4_fp_val;
  assign _GEN_48498 = io_enq_valids_1 ? _GEN_44695 : _T_5936_5_fp_val;
  assign _GEN_48499 = io_enq_valids_1 ? _GEN_44696 : _T_5936_6_fp_val;
  assign _GEN_48500 = io_enq_valids_1 ? _GEN_44697 : _T_5936_7_fp_val;
  assign _GEN_48501 = io_enq_valids_1 ? _GEN_44698 : _T_5936_8_fp_val;
  assign _GEN_48502 = io_enq_valids_1 ? _GEN_44699 : _T_5936_9_fp_val;
  assign _GEN_48503 = io_enq_valids_1 ? _GEN_44700 : _T_5936_10_fp_val;
  assign _GEN_48504 = io_enq_valids_1 ? _GEN_44701 : _T_5936_11_fp_val;
  assign _GEN_48505 = io_enq_valids_1 ? _GEN_44702 : _T_5936_12_fp_val;
  assign _GEN_48506 = io_enq_valids_1 ? _GEN_44703 : _T_5936_13_fp_val;
  assign _GEN_48507 = io_enq_valids_1 ? _GEN_44704 : _T_5936_14_fp_val;
  assign _GEN_48508 = io_enq_valids_1 ? _GEN_44705 : _T_5936_15_fp_val;
  assign _GEN_48509 = io_enq_valids_1 ? _GEN_44706 : _T_5936_16_fp_val;
  assign _GEN_48510 = io_enq_valids_1 ? _GEN_44707 : _T_5936_17_fp_val;
  assign _GEN_48511 = io_enq_valids_1 ? _GEN_44708 : _T_5936_18_fp_val;
  assign _GEN_48512 = io_enq_valids_1 ? _GEN_44709 : _T_5936_19_fp_val;
  assign _GEN_48513 = io_enq_valids_1 ? _GEN_44710 : _T_5936_20_fp_val;
  assign _GEN_48514 = io_enq_valids_1 ? _GEN_44711 : _T_5936_21_fp_val;
  assign _GEN_48515 = io_enq_valids_1 ? _GEN_44712 : _T_5936_22_fp_val;
  assign _GEN_48516 = io_enq_valids_1 ? _GEN_44713 : _T_5936_23_fp_val;
  assign _GEN_48517 = io_enq_valids_1 ? _GEN_44714 : _T_5936_24_fp_val;
  assign _GEN_48518 = io_enq_valids_1 ? _GEN_44715 : _T_5936_25_fp_val;
  assign _GEN_48519 = io_enq_valids_1 ? _GEN_44716 : _T_5936_26_fp_val;
  assign _GEN_48520 = io_enq_valids_1 ? _GEN_44717 : _T_5936_27_fp_val;
  assign _GEN_48521 = io_enq_valids_1 ? _GEN_44718 : _T_5936_28_fp_val;
  assign _GEN_48522 = io_enq_valids_1 ? _GEN_44719 : _T_5936_29_fp_val;
  assign _GEN_48523 = io_enq_valids_1 ? _GEN_44720 : _T_5936_30_fp_val;
  assign _GEN_48524 = io_enq_valids_1 ? _GEN_44721 : _T_5936_31_fp_val;
  assign _GEN_48525 = io_enq_valids_1 ? _GEN_44722 : _T_5936_32_fp_val;
  assign _GEN_48526 = io_enq_valids_1 ? _GEN_44723 : _T_5936_33_fp_val;
  assign _GEN_48527 = io_enq_valids_1 ? _GEN_44724 : _T_5936_34_fp_val;
  assign _GEN_48528 = io_enq_valids_1 ? _GEN_44725 : _T_5936_35_fp_val;
  assign _GEN_48529 = io_enq_valids_1 ? _GEN_44726 : _T_5936_36_fp_val;
  assign _GEN_48530 = io_enq_valids_1 ? _GEN_44727 : _T_5936_37_fp_val;
  assign _GEN_48531 = io_enq_valids_1 ? _GEN_44728 : _T_5936_38_fp_val;
  assign _GEN_48532 = io_enq_valids_1 ? _GEN_44729 : _T_5936_39_fp_val;
  assign _T_6381 = io_wb_resps_0_valid & _T_3814;
  assign _T_6382 = _T_3813[5:0];
  assign _T_6390 = io_wb_resps_1_valid & _T_3823;
  assign _T_6391 = _T_3822[5:0];
  assign _T_6399 = io_wb_resps_2_valid & _T_3832;
  assign _T_6400 = _T_3831[5:0];
  assign _T_6408 = io_wb_resps_3_valid & _T_3841;
  assign _T_6409 = _T_3840[5:0];
  assign _T_6417 = io_wb_resps_4_valid & _T_3850;
  assign _T_6418 = _T_3849[5:0];
  assign _T_6424 = io_lsu_clr_bsy_valid_0 & _T_3857;
  assign _T_6427 = _T_3862[5:0];
  assign _GEN_48835 = 6'h1 == _T_3863 ? _T_5637_1 : _T_5637_0;
  assign _GEN_48836 = 6'h2 == _T_3863 ? _T_5637_2 : _GEN_48835;
  assign _GEN_48837 = 6'h3 == _T_3863 ? _T_5637_3 : _GEN_48836;
  assign _GEN_48838 = 6'h4 == _T_3863 ? _T_5637_4 : _GEN_48837;
  assign _GEN_48839 = 6'h5 == _T_3863 ? _T_5637_5 : _GEN_48838;
  assign _GEN_48840 = 6'h6 == _T_3863 ? _T_5637_6 : _GEN_48839;
  assign _GEN_48841 = 6'h7 == _T_3863 ? _T_5637_7 : _GEN_48840;
  assign _GEN_48842 = 6'h8 == _T_3863 ? _T_5637_8 : _GEN_48841;
  assign _GEN_48843 = 6'h9 == _T_3863 ? _T_5637_9 : _GEN_48842;
  assign _GEN_48844 = 6'ha == _T_3863 ? _T_5637_10 : _GEN_48843;
  assign _GEN_48845 = 6'hb == _T_3863 ? _T_5637_11 : _GEN_48844;
  assign _GEN_48846 = 6'hc == _T_3863 ? _T_5637_12 : _GEN_48845;
  assign _GEN_48847 = 6'hd == _T_3863 ? _T_5637_13 : _GEN_48846;
  assign _GEN_48848 = 6'he == _T_3863 ? _T_5637_14 : _GEN_48847;
  assign _GEN_48849 = 6'hf == _T_3863 ? _T_5637_15 : _GEN_48848;
  assign _GEN_48850 = 6'h10 == _T_3863 ? _T_5637_16 : _GEN_48849;
  assign _GEN_48851 = 6'h11 == _T_3863 ? _T_5637_17 : _GEN_48850;
  assign _GEN_48852 = 6'h12 == _T_3863 ? _T_5637_18 : _GEN_48851;
  assign _GEN_48853 = 6'h13 == _T_3863 ? _T_5637_19 : _GEN_48852;
  assign _GEN_48854 = 6'h14 == _T_3863 ? _T_5637_20 : _GEN_48853;
  assign _GEN_48855 = 6'h15 == _T_3863 ? _T_5637_21 : _GEN_48854;
  assign _GEN_48856 = 6'h16 == _T_3863 ? _T_5637_22 : _GEN_48855;
  assign _GEN_48857 = 6'h17 == _T_3863 ? _T_5637_23 : _GEN_48856;
  assign _GEN_48858 = 6'h18 == _T_3863 ? _T_5637_24 : _GEN_48857;
  assign _GEN_48859 = 6'h19 == _T_3863 ? _T_5637_25 : _GEN_48858;
  assign _GEN_48860 = 6'h1a == _T_3863 ? _T_5637_26 : _GEN_48859;
  assign _GEN_48861 = 6'h1b == _T_3863 ? _T_5637_27 : _GEN_48860;
  assign _GEN_48862 = 6'h1c == _T_3863 ? _T_5637_28 : _GEN_48861;
  assign _GEN_48863 = 6'h1d == _T_3863 ? _T_5637_29 : _GEN_48862;
  assign _GEN_48864 = 6'h1e == _T_3863 ? _T_5637_30 : _GEN_48863;
  assign _GEN_48865 = 6'h1f == _T_3863 ? _T_5637_31 : _GEN_48864;
  assign _GEN_48866 = 6'h20 == _T_3863 ? _T_5637_32 : _GEN_48865;
  assign _GEN_48867 = 6'h21 == _T_3863 ? _T_5637_33 : _GEN_48866;
  assign _GEN_48868 = 6'h22 == _T_3863 ? _T_5637_34 : _GEN_48867;
  assign _GEN_48869 = 6'h23 == _T_3863 ? _T_5637_35 : _GEN_48868;
  assign _GEN_48870 = 6'h24 == _T_3863 ? _T_5637_36 : _GEN_48869;
  assign _GEN_48871 = 6'h25 == _T_3863 ? _T_5637_37 : _GEN_48870;
  assign _GEN_48872 = 6'h26 == _T_3863 ? _T_5637_38 : _GEN_48871;
  assign _GEN_48873 = 6'h27 == _T_3863 ? _T_5637_39 : _GEN_48872;
  assign _T_6437 = _GEN_323 | reset;
  assign _T_6439 = _T_6437 == 1'h0;
  assign _T_6440 = _T_3862[5:0];
  assign _T_6443 = _T_5764__T_6441_data;
  assign _T_6445 = _T_6443 | reset;
  assign _T_6447 = _T_6445 == 1'h0;
  assign _T_6451 = io_lsu_clr_bsy_valid_1 & _T_3884;
  assign _T_6454 = _T_3889[5:0];
  assign _GEN_48879 = 6'h1 == _T_3890 ? _T_5637_1 : _T_5637_0;
  assign _GEN_48880 = 6'h2 == _T_3890 ? _T_5637_2 : _GEN_48879;
  assign _GEN_48881 = 6'h3 == _T_3890 ? _T_5637_3 : _GEN_48880;
  assign _GEN_48882 = 6'h4 == _T_3890 ? _T_5637_4 : _GEN_48881;
  assign _GEN_48883 = 6'h5 == _T_3890 ? _T_5637_5 : _GEN_48882;
  assign _GEN_48884 = 6'h6 == _T_3890 ? _T_5637_6 : _GEN_48883;
  assign _GEN_48885 = 6'h7 == _T_3890 ? _T_5637_7 : _GEN_48884;
  assign _GEN_48886 = 6'h8 == _T_3890 ? _T_5637_8 : _GEN_48885;
  assign _GEN_48887 = 6'h9 == _T_3890 ? _T_5637_9 : _GEN_48886;
  assign _GEN_48888 = 6'ha == _T_3890 ? _T_5637_10 : _GEN_48887;
  assign _GEN_48889 = 6'hb == _T_3890 ? _T_5637_11 : _GEN_48888;
  assign _GEN_48890 = 6'hc == _T_3890 ? _T_5637_12 : _GEN_48889;
  assign _GEN_48891 = 6'hd == _T_3890 ? _T_5637_13 : _GEN_48890;
  assign _GEN_48892 = 6'he == _T_3890 ? _T_5637_14 : _GEN_48891;
  assign _GEN_48893 = 6'hf == _T_3890 ? _T_5637_15 : _GEN_48892;
  assign _GEN_48894 = 6'h10 == _T_3890 ? _T_5637_16 : _GEN_48893;
  assign _GEN_48895 = 6'h11 == _T_3890 ? _T_5637_17 : _GEN_48894;
  assign _GEN_48896 = 6'h12 == _T_3890 ? _T_5637_18 : _GEN_48895;
  assign _GEN_48897 = 6'h13 == _T_3890 ? _T_5637_19 : _GEN_48896;
  assign _GEN_48898 = 6'h14 == _T_3890 ? _T_5637_20 : _GEN_48897;
  assign _GEN_48899 = 6'h15 == _T_3890 ? _T_5637_21 : _GEN_48898;
  assign _GEN_48900 = 6'h16 == _T_3890 ? _T_5637_22 : _GEN_48899;
  assign _GEN_48901 = 6'h17 == _T_3890 ? _T_5637_23 : _GEN_48900;
  assign _GEN_48902 = 6'h18 == _T_3890 ? _T_5637_24 : _GEN_48901;
  assign _GEN_48903 = 6'h19 == _T_3890 ? _T_5637_25 : _GEN_48902;
  assign _GEN_48904 = 6'h1a == _T_3890 ? _T_5637_26 : _GEN_48903;
  assign _GEN_48905 = 6'h1b == _T_3890 ? _T_5637_27 : _GEN_48904;
  assign _GEN_48906 = 6'h1c == _T_3890 ? _T_5637_28 : _GEN_48905;
  assign _GEN_48907 = 6'h1d == _T_3890 ? _T_5637_29 : _GEN_48906;
  assign _GEN_48908 = 6'h1e == _T_3890 ? _T_5637_30 : _GEN_48907;
  assign _GEN_48909 = 6'h1f == _T_3890 ? _T_5637_31 : _GEN_48908;
  assign _GEN_48910 = 6'h20 == _T_3890 ? _T_5637_32 : _GEN_48909;
  assign _GEN_48911 = 6'h21 == _T_3890 ? _T_5637_33 : _GEN_48910;
  assign _GEN_48912 = 6'h22 == _T_3890 ? _T_5637_34 : _GEN_48911;
  assign _GEN_48913 = 6'h23 == _T_3890 ? _T_5637_35 : _GEN_48912;
  assign _GEN_48914 = 6'h24 == _T_3890 ? _T_5637_36 : _GEN_48913;
  assign _GEN_48915 = 6'h25 == _T_3890 ? _T_5637_37 : _GEN_48914;
  assign _GEN_48916 = 6'h26 == _T_3890 ? _T_5637_38 : _GEN_48915;
  assign _GEN_48917 = 6'h27 == _T_3890 ? _T_5637_39 : _GEN_48916;
  assign _T_6464 = _GEN_324 | reset;
  assign _T_6466 = _T_6464 == 1'h0;
  assign _T_6467 = _T_3889[5:0];
  assign _T_6470 = _T_5764__T_6468_data;
  assign _T_6472 = _T_6470 | reset;
  assign _T_6474 = _T_6472 == 1'h0;
  assign _T_6542 = io_fflags_0_valid & _T_3975;
  assign _T_6545 = _T_3980[5:0];
  assign _T_6550 = io_fflags_1_valid & _T_3983;
  assign _T_6553 = _T_3988[5:0];
  assign _T_6558 = io_lxcpt_valid & _T_3991;
  assign _T_6561 = _T_3996[5:0];
  assign _T_6567 = io_bxcpt_valid & _T_4000;
  assign _T_6570 = _T_4005[5:0];
  assign _GEN_49339 = 6'h1 == rob_head ? _T_5637_1 : _T_5637_0;
  assign _GEN_49340 = 6'h2 == rob_head ? _T_5637_2 : _GEN_49339;
  assign _GEN_49341 = 6'h3 == rob_head ? _T_5637_3 : _GEN_49340;
  assign _GEN_49342 = 6'h4 == rob_head ? _T_5637_4 : _GEN_49341;
  assign _GEN_49343 = 6'h5 == rob_head ? _T_5637_5 : _GEN_49342;
  assign _GEN_49344 = 6'h6 == rob_head ? _T_5637_6 : _GEN_49343;
  assign _GEN_49345 = 6'h7 == rob_head ? _T_5637_7 : _GEN_49344;
  assign _GEN_49346 = 6'h8 == rob_head ? _T_5637_8 : _GEN_49345;
  assign _GEN_49347 = 6'h9 == rob_head ? _T_5637_9 : _GEN_49346;
  assign _GEN_49348 = 6'ha == rob_head ? _T_5637_10 : _GEN_49347;
  assign _GEN_49349 = 6'hb == rob_head ? _T_5637_11 : _GEN_49348;
  assign _GEN_49350 = 6'hc == rob_head ? _T_5637_12 : _GEN_49349;
  assign _GEN_49351 = 6'hd == rob_head ? _T_5637_13 : _GEN_49350;
  assign _GEN_49352 = 6'he == rob_head ? _T_5637_14 : _GEN_49351;
  assign _GEN_49353 = 6'hf == rob_head ? _T_5637_15 : _GEN_49352;
  assign _GEN_49354 = 6'h10 == rob_head ? _T_5637_16 : _GEN_49353;
  assign _GEN_49355 = 6'h11 == rob_head ? _T_5637_17 : _GEN_49354;
  assign _GEN_49356 = 6'h12 == rob_head ? _T_5637_18 : _GEN_49355;
  assign _GEN_49357 = 6'h13 == rob_head ? _T_5637_19 : _GEN_49356;
  assign _GEN_49358 = 6'h14 == rob_head ? _T_5637_20 : _GEN_49357;
  assign _GEN_49359 = 6'h15 == rob_head ? _T_5637_21 : _GEN_49358;
  assign _GEN_49360 = 6'h16 == rob_head ? _T_5637_22 : _GEN_49359;
  assign _GEN_49361 = 6'h17 == rob_head ? _T_5637_23 : _GEN_49360;
  assign _GEN_49362 = 6'h18 == rob_head ? _T_5637_24 : _GEN_49361;
  assign _GEN_49363 = 6'h19 == rob_head ? _T_5637_25 : _GEN_49362;
  assign _GEN_49364 = 6'h1a == rob_head ? _T_5637_26 : _GEN_49363;
  assign _GEN_49365 = 6'h1b == rob_head ? _T_5637_27 : _GEN_49364;
  assign _GEN_49366 = 6'h1c == rob_head ? _T_5637_28 : _GEN_49365;
  assign _GEN_49367 = 6'h1d == rob_head ? _T_5637_29 : _GEN_49366;
  assign _GEN_49368 = 6'h1e == rob_head ? _T_5637_30 : _GEN_49367;
  assign _GEN_49369 = 6'h1f == rob_head ? _T_5637_31 : _GEN_49368;
  assign _GEN_49370 = 6'h20 == rob_head ? _T_5637_32 : _GEN_49369;
  assign _GEN_49371 = 6'h21 == rob_head ? _T_5637_33 : _GEN_49370;
  assign _GEN_49372 = 6'h22 == rob_head ? _T_5637_34 : _GEN_49371;
  assign _GEN_49373 = 6'h23 == rob_head ? _T_5637_35 : _GEN_49372;
  assign _GEN_49374 = 6'h24 == rob_head ? _T_5637_36 : _GEN_49373;
  assign _GEN_49375 = 6'h25 == rob_head ? _T_5637_37 : _GEN_49374;
  assign _GEN_49376 = 6'h26 == rob_head ? _T_5637_38 : _GEN_49375;
  assign _GEN_49377 = 6'h27 == rob_head ? _T_5637_39 : _GEN_49376;
  assign _T_6577 = _GEN_330 & _T_6309__T_6576_data;
  assign _T_6583 = _T_5764__T_6581_data == 1'h0;
  assign _T_6584 = _GEN_331 & _T_6583;
  assign _T_6587 = _T_6584 & _T_4022;
  assign _GEN_49431 = 6'h1 == _T_6589 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_49438 = 6'h1 == _T_6589 ? _T_5936_1_stale_pdst : _T_5936_0_stale_pdst;
  assign _GEN_49445 = 6'h1 == _T_6589 ? _T_5936_1_is_fencei : _T_5936_0_is_fencei;
  assign _GEN_49446 = 6'h1 == _T_6589 ? _T_5936_1_is_store : _T_5936_0_is_store;
  assign _GEN_49448 = 6'h1 == _T_6589 ? _T_5936_1_is_load : _T_5936_0_is_load;
  assign _GEN_49449 = 6'h1 == _T_6589 ? _T_5936_1_is_sys_pc2epc : _T_5936_0_is_sys_pc2epc;
  assign _GEN_49451 = 6'h1 == _T_6589 ? _T_5936_1_flush_on_commit : _T_5936_0_flush_on_commit;
  assign _GEN_49452 = 6'h1 == _T_6589 ? _T_5936_1_ldst : _T_5936_0_ldst;
  assign _GEN_49457 = 6'h1 == _T_6589 ? _T_5936_1_dst_rtype : _T_5936_0_dst_rtype;
  assign _GEN_49461 = 6'h1 == _T_6589 ? _T_5936_1_fp_val : _T_5936_0_fp_val;
  assign _GEN_49521 = 6'h2 == _T_6589 ? _T_5936_2_pdst : _GEN_49431;
  assign _GEN_49528 = 6'h2 == _T_6589 ? _T_5936_2_stale_pdst : _GEN_49438;
  assign _GEN_49535 = 6'h2 == _T_6589 ? _T_5936_2_is_fencei : _GEN_49445;
  assign _GEN_49536 = 6'h2 == _T_6589 ? _T_5936_2_is_store : _GEN_49446;
  assign _GEN_49538 = 6'h2 == _T_6589 ? _T_5936_2_is_load : _GEN_49448;
  assign _GEN_49539 = 6'h2 == _T_6589 ? _T_5936_2_is_sys_pc2epc : _GEN_49449;
  assign _GEN_49541 = 6'h2 == _T_6589 ? _T_5936_2_flush_on_commit : _GEN_49451;
  assign _GEN_49542 = 6'h2 == _T_6589 ? _T_5936_2_ldst : _GEN_49452;
  assign _GEN_49547 = 6'h2 == _T_6589 ? _T_5936_2_dst_rtype : _GEN_49457;
  assign _GEN_49551 = 6'h2 == _T_6589 ? _T_5936_2_fp_val : _GEN_49461;
  assign _GEN_49611 = 6'h3 == _T_6589 ? _T_5936_3_pdst : _GEN_49521;
  assign _GEN_49618 = 6'h3 == _T_6589 ? _T_5936_3_stale_pdst : _GEN_49528;
  assign _GEN_49625 = 6'h3 == _T_6589 ? _T_5936_3_is_fencei : _GEN_49535;
  assign _GEN_49626 = 6'h3 == _T_6589 ? _T_5936_3_is_store : _GEN_49536;
  assign _GEN_49628 = 6'h3 == _T_6589 ? _T_5936_3_is_load : _GEN_49538;
  assign _GEN_49629 = 6'h3 == _T_6589 ? _T_5936_3_is_sys_pc2epc : _GEN_49539;
  assign _GEN_49631 = 6'h3 == _T_6589 ? _T_5936_3_flush_on_commit : _GEN_49541;
  assign _GEN_49632 = 6'h3 == _T_6589 ? _T_5936_3_ldst : _GEN_49542;
  assign _GEN_49637 = 6'h3 == _T_6589 ? _T_5936_3_dst_rtype : _GEN_49547;
  assign _GEN_49641 = 6'h3 == _T_6589 ? _T_5936_3_fp_val : _GEN_49551;
  assign _GEN_49701 = 6'h4 == _T_6589 ? _T_5936_4_pdst : _GEN_49611;
  assign _GEN_49708 = 6'h4 == _T_6589 ? _T_5936_4_stale_pdst : _GEN_49618;
  assign _GEN_49715 = 6'h4 == _T_6589 ? _T_5936_4_is_fencei : _GEN_49625;
  assign _GEN_49716 = 6'h4 == _T_6589 ? _T_5936_4_is_store : _GEN_49626;
  assign _GEN_49718 = 6'h4 == _T_6589 ? _T_5936_4_is_load : _GEN_49628;
  assign _GEN_49719 = 6'h4 == _T_6589 ? _T_5936_4_is_sys_pc2epc : _GEN_49629;
  assign _GEN_49721 = 6'h4 == _T_6589 ? _T_5936_4_flush_on_commit : _GEN_49631;
  assign _GEN_49722 = 6'h4 == _T_6589 ? _T_5936_4_ldst : _GEN_49632;
  assign _GEN_49727 = 6'h4 == _T_6589 ? _T_5936_4_dst_rtype : _GEN_49637;
  assign _GEN_49731 = 6'h4 == _T_6589 ? _T_5936_4_fp_val : _GEN_49641;
  assign _GEN_49791 = 6'h5 == _T_6589 ? _T_5936_5_pdst : _GEN_49701;
  assign _GEN_49798 = 6'h5 == _T_6589 ? _T_5936_5_stale_pdst : _GEN_49708;
  assign _GEN_49805 = 6'h5 == _T_6589 ? _T_5936_5_is_fencei : _GEN_49715;
  assign _GEN_49806 = 6'h5 == _T_6589 ? _T_5936_5_is_store : _GEN_49716;
  assign _GEN_49808 = 6'h5 == _T_6589 ? _T_5936_5_is_load : _GEN_49718;
  assign _GEN_49809 = 6'h5 == _T_6589 ? _T_5936_5_is_sys_pc2epc : _GEN_49719;
  assign _GEN_49811 = 6'h5 == _T_6589 ? _T_5936_5_flush_on_commit : _GEN_49721;
  assign _GEN_49812 = 6'h5 == _T_6589 ? _T_5936_5_ldst : _GEN_49722;
  assign _GEN_49817 = 6'h5 == _T_6589 ? _T_5936_5_dst_rtype : _GEN_49727;
  assign _GEN_49821 = 6'h5 == _T_6589 ? _T_5936_5_fp_val : _GEN_49731;
  assign _GEN_49881 = 6'h6 == _T_6589 ? _T_5936_6_pdst : _GEN_49791;
  assign _GEN_49888 = 6'h6 == _T_6589 ? _T_5936_6_stale_pdst : _GEN_49798;
  assign _GEN_49895 = 6'h6 == _T_6589 ? _T_5936_6_is_fencei : _GEN_49805;
  assign _GEN_49896 = 6'h6 == _T_6589 ? _T_5936_6_is_store : _GEN_49806;
  assign _GEN_49898 = 6'h6 == _T_6589 ? _T_5936_6_is_load : _GEN_49808;
  assign _GEN_49899 = 6'h6 == _T_6589 ? _T_5936_6_is_sys_pc2epc : _GEN_49809;
  assign _GEN_49901 = 6'h6 == _T_6589 ? _T_5936_6_flush_on_commit : _GEN_49811;
  assign _GEN_49902 = 6'h6 == _T_6589 ? _T_5936_6_ldst : _GEN_49812;
  assign _GEN_49907 = 6'h6 == _T_6589 ? _T_5936_6_dst_rtype : _GEN_49817;
  assign _GEN_49911 = 6'h6 == _T_6589 ? _T_5936_6_fp_val : _GEN_49821;
  assign _GEN_49971 = 6'h7 == _T_6589 ? _T_5936_7_pdst : _GEN_49881;
  assign _GEN_49978 = 6'h7 == _T_6589 ? _T_5936_7_stale_pdst : _GEN_49888;
  assign _GEN_49985 = 6'h7 == _T_6589 ? _T_5936_7_is_fencei : _GEN_49895;
  assign _GEN_49986 = 6'h7 == _T_6589 ? _T_5936_7_is_store : _GEN_49896;
  assign _GEN_49988 = 6'h7 == _T_6589 ? _T_5936_7_is_load : _GEN_49898;
  assign _GEN_49989 = 6'h7 == _T_6589 ? _T_5936_7_is_sys_pc2epc : _GEN_49899;
  assign _GEN_49991 = 6'h7 == _T_6589 ? _T_5936_7_flush_on_commit : _GEN_49901;
  assign _GEN_49992 = 6'h7 == _T_6589 ? _T_5936_7_ldst : _GEN_49902;
  assign _GEN_49997 = 6'h7 == _T_6589 ? _T_5936_7_dst_rtype : _GEN_49907;
  assign _GEN_50001 = 6'h7 == _T_6589 ? _T_5936_7_fp_val : _GEN_49911;
  assign _GEN_50061 = 6'h8 == _T_6589 ? _T_5936_8_pdst : _GEN_49971;
  assign _GEN_50068 = 6'h8 == _T_6589 ? _T_5936_8_stale_pdst : _GEN_49978;
  assign _GEN_50075 = 6'h8 == _T_6589 ? _T_5936_8_is_fencei : _GEN_49985;
  assign _GEN_50076 = 6'h8 == _T_6589 ? _T_5936_8_is_store : _GEN_49986;
  assign _GEN_50078 = 6'h8 == _T_6589 ? _T_5936_8_is_load : _GEN_49988;
  assign _GEN_50079 = 6'h8 == _T_6589 ? _T_5936_8_is_sys_pc2epc : _GEN_49989;
  assign _GEN_50081 = 6'h8 == _T_6589 ? _T_5936_8_flush_on_commit : _GEN_49991;
  assign _GEN_50082 = 6'h8 == _T_6589 ? _T_5936_8_ldst : _GEN_49992;
  assign _GEN_50087 = 6'h8 == _T_6589 ? _T_5936_8_dst_rtype : _GEN_49997;
  assign _GEN_50091 = 6'h8 == _T_6589 ? _T_5936_8_fp_val : _GEN_50001;
  assign _GEN_50151 = 6'h9 == _T_6589 ? _T_5936_9_pdst : _GEN_50061;
  assign _GEN_50158 = 6'h9 == _T_6589 ? _T_5936_9_stale_pdst : _GEN_50068;
  assign _GEN_50165 = 6'h9 == _T_6589 ? _T_5936_9_is_fencei : _GEN_50075;
  assign _GEN_50166 = 6'h9 == _T_6589 ? _T_5936_9_is_store : _GEN_50076;
  assign _GEN_50168 = 6'h9 == _T_6589 ? _T_5936_9_is_load : _GEN_50078;
  assign _GEN_50169 = 6'h9 == _T_6589 ? _T_5936_9_is_sys_pc2epc : _GEN_50079;
  assign _GEN_50171 = 6'h9 == _T_6589 ? _T_5936_9_flush_on_commit : _GEN_50081;
  assign _GEN_50172 = 6'h9 == _T_6589 ? _T_5936_9_ldst : _GEN_50082;
  assign _GEN_50177 = 6'h9 == _T_6589 ? _T_5936_9_dst_rtype : _GEN_50087;
  assign _GEN_50181 = 6'h9 == _T_6589 ? _T_5936_9_fp_val : _GEN_50091;
  assign _GEN_50241 = 6'ha == _T_6589 ? _T_5936_10_pdst : _GEN_50151;
  assign _GEN_50248 = 6'ha == _T_6589 ? _T_5936_10_stale_pdst : _GEN_50158;
  assign _GEN_50255 = 6'ha == _T_6589 ? _T_5936_10_is_fencei : _GEN_50165;
  assign _GEN_50256 = 6'ha == _T_6589 ? _T_5936_10_is_store : _GEN_50166;
  assign _GEN_50258 = 6'ha == _T_6589 ? _T_5936_10_is_load : _GEN_50168;
  assign _GEN_50259 = 6'ha == _T_6589 ? _T_5936_10_is_sys_pc2epc : _GEN_50169;
  assign _GEN_50261 = 6'ha == _T_6589 ? _T_5936_10_flush_on_commit : _GEN_50171;
  assign _GEN_50262 = 6'ha == _T_6589 ? _T_5936_10_ldst : _GEN_50172;
  assign _GEN_50267 = 6'ha == _T_6589 ? _T_5936_10_dst_rtype : _GEN_50177;
  assign _GEN_50271 = 6'ha == _T_6589 ? _T_5936_10_fp_val : _GEN_50181;
  assign _GEN_50331 = 6'hb == _T_6589 ? _T_5936_11_pdst : _GEN_50241;
  assign _GEN_50338 = 6'hb == _T_6589 ? _T_5936_11_stale_pdst : _GEN_50248;
  assign _GEN_50345 = 6'hb == _T_6589 ? _T_5936_11_is_fencei : _GEN_50255;
  assign _GEN_50346 = 6'hb == _T_6589 ? _T_5936_11_is_store : _GEN_50256;
  assign _GEN_50348 = 6'hb == _T_6589 ? _T_5936_11_is_load : _GEN_50258;
  assign _GEN_50349 = 6'hb == _T_6589 ? _T_5936_11_is_sys_pc2epc : _GEN_50259;
  assign _GEN_50351 = 6'hb == _T_6589 ? _T_5936_11_flush_on_commit : _GEN_50261;
  assign _GEN_50352 = 6'hb == _T_6589 ? _T_5936_11_ldst : _GEN_50262;
  assign _GEN_50357 = 6'hb == _T_6589 ? _T_5936_11_dst_rtype : _GEN_50267;
  assign _GEN_50361 = 6'hb == _T_6589 ? _T_5936_11_fp_val : _GEN_50271;
  assign _GEN_50421 = 6'hc == _T_6589 ? _T_5936_12_pdst : _GEN_50331;
  assign _GEN_50428 = 6'hc == _T_6589 ? _T_5936_12_stale_pdst : _GEN_50338;
  assign _GEN_50435 = 6'hc == _T_6589 ? _T_5936_12_is_fencei : _GEN_50345;
  assign _GEN_50436 = 6'hc == _T_6589 ? _T_5936_12_is_store : _GEN_50346;
  assign _GEN_50438 = 6'hc == _T_6589 ? _T_5936_12_is_load : _GEN_50348;
  assign _GEN_50439 = 6'hc == _T_6589 ? _T_5936_12_is_sys_pc2epc : _GEN_50349;
  assign _GEN_50441 = 6'hc == _T_6589 ? _T_5936_12_flush_on_commit : _GEN_50351;
  assign _GEN_50442 = 6'hc == _T_6589 ? _T_5936_12_ldst : _GEN_50352;
  assign _GEN_50447 = 6'hc == _T_6589 ? _T_5936_12_dst_rtype : _GEN_50357;
  assign _GEN_50451 = 6'hc == _T_6589 ? _T_5936_12_fp_val : _GEN_50361;
  assign _GEN_50511 = 6'hd == _T_6589 ? _T_5936_13_pdst : _GEN_50421;
  assign _GEN_50518 = 6'hd == _T_6589 ? _T_5936_13_stale_pdst : _GEN_50428;
  assign _GEN_50525 = 6'hd == _T_6589 ? _T_5936_13_is_fencei : _GEN_50435;
  assign _GEN_50526 = 6'hd == _T_6589 ? _T_5936_13_is_store : _GEN_50436;
  assign _GEN_50528 = 6'hd == _T_6589 ? _T_5936_13_is_load : _GEN_50438;
  assign _GEN_50529 = 6'hd == _T_6589 ? _T_5936_13_is_sys_pc2epc : _GEN_50439;
  assign _GEN_50531 = 6'hd == _T_6589 ? _T_5936_13_flush_on_commit : _GEN_50441;
  assign _GEN_50532 = 6'hd == _T_6589 ? _T_5936_13_ldst : _GEN_50442;
  assign _GEN_50537 = 6'hd == _T_6589 ? _T_5936_13_dst_rtype : _GEN_50447;
  assign _GEN_50541 = 6'hd == _T_6589 ? _T_5936_13_fp_val : _GEN_50451;
  assign _GEN_50601 = 6'he == _T_6589 ? _T_5936_14_pdst : _GEN_50511;
  assign _GEN_50608 = 6'he == _T_6589 ? _T_5936_14_stale_pdst : _GEN_50518;
  assign _GEN_50615 = 6'he == _T_6589 ? _T_5936_14_is_fencei : _GEN_50525;
  assign _GEN_50616 = 6'he == _T_6589 ? _T_5936_14_is_store : _GEN_50526;
  assign _GEN_50618 = 6'he == _T_6589 ? _T_5936_14_is_load : _GEN_50528;
  assign _GEN_50619 = 6'he == _T_6589 ? _T_5936_14_is_sys_pc2epc : _GEN_50529;
  assign _GEN_50621 = 6'he == _T_6589 ? _T_5936_14_flush_on_commit : _GEN_50531;
  assign _GEN_50622 = 6'he == _T_6589 ? _T_5936_14_ldst : _GEN_50532;
  assign _GEN_50627 = 6'he == _T_6589 ? _T_5936_14_dst_rtype : _GEN_50537;
  assign _GEN_50631 = 6'he == _T_6589 ? _T_5936_14_fp_val : _GEN_50541;
  assign _GEN_50691 = 6'hf == _T_6589 ? _T_5936_15_pdst : _GEN_50601;
  assign _GEN_50698 = 6'hf == _T_6589 ? _T_5936_15_stale_pdst : _GEN_50608;
  assign _GEN_50705 = 6'hf == _T_6589 ? _T_5936_15_is_fencei : _GEN_50615;
  assign _GEN_50706 = 6'hf == _T_6589 ? _T_5936_15_is_store : _GEN_50616;
  assign _GEN_50708 = 6'hf == _T_6589 ? _T_5936_15_is_load : _GEN_50618;
  assign _GEN_50709 = 6'hf == _T_6589 ? _T_5936_15_is_sys_pc2epc : _GEN_50619;
  assign _GEN_50711 = 6'hf == _T_6589 ? _T_5936_15_flush_on_commit : _GEN_50621;
  assign _GEN_50712 = 6'hf == _T_6589 ? _T_5936_15_ldst : _GEN_50622;
  assign _GEN_50717 = 6'hf == _T_6589 ? _T_5936_15_dst_rtype : _GEN_50627;
  assign _GEN_50721 = 6'hf == _T_6589 ? _T_5936_15_fp_val : _GEN_50631;
  assign _GEN_50781 = 6'h10 == _T_6589 ? _T_5936_16_pdst : _GEN_50691;
  assign _GEN_50788 = 6'h10 == _T_6589 ? _T_5936_16_stale_pdst : _GEN_50698;
  assign _GEN_50795 = 6'h10 == _T_6589 ? _T_5936_16_is_fencei : _GEN_50705;
  assign _GEN_50796 = 6'h10 == _T_6589 ? _T_5936_16_is_store : _GEN_50706;
  assign _GEN_50798 = 6'h10 == _T_6589 ? _T_5936_16_is_load : _GEN_50708;
  assign _GEN_50799 = 6'h10 == _T_6589 ? _T_5936_16_is_sys_pc2epc : _GEN_50709;
  assign _GEN_50801 = 6'h10 == _T_6589 ? _T_5936_16_flush_on_commit : _GEN_50711;
  assign _GEN_50802 = 6'h10 == _T_6589 ? _T_5936_16_ldst : _GEN_50712;
  assign _GEN_50807 = 6'h10 == _T_6589 ? _T_5936_16_dst_rtype : _GEN_50717;
  assign _GEN_50811 = 6'h10 == _T_6589 ? _T_5936_16_fp_val : _GEN_50721;
  assign _GEN_50871 = 6'h11 == _T_6589 ? _T_5936_17_pdst : _GEN_50781;
  assign _GEN_50878 = 6'h11 == _T_6589 ? _T_5936_17_stale_pdst : _GEN_50788;
  assign _GEN_50885 = 6'h11 == _T_6589 ? _T_5936_17_is_fencei : _GEN_50795;
  assign _GEN_50886 = 6'h11 == _T_6589 ? _T_5936_17_is_store : _GEN_50796;
  assign _GEN_50888 = 6'h11 == _T_6589 ? _T_5936_17_is_load : _GEN_50798;
  assign _GEN_50889 = 6'h11 == _T_6589 ? _T_5936_17_is_sys_pc2epc : _GEN_50799;
  assign _GEN_50891 = 6'h11 == _T_6589 ? _T_5936_17_flush_on_commit : _GEN_50801;
  assign _GEN_50892 = 6'h11 == _T_6589 ? _T_5936_17_ldst : _GEN_50802;
  assign _GEN_50897 = 6'h11 == _T_6589 ? _T_5936_17_dst_rtype : _GEN_50807;
  assign _GEN_50901 = 6'h11 == _T_6589 ? _T_5936_17_fp_val : _GEN_50811;
  assign _GEN_50961 = 6'h12 == _T_6589 ? _T_5936_18_pdst : _GEN_50871;
  assign _GEN_50968 = 6'h12 == _T_6589 ? _T_5936_18_stale_pdst : _GEN_50878;
  assign _GEN_50975 = 6'h12 == _T_6589 ? _T_5936_18_is_fencei : _GEN_50885;
  assign _GEN_50976 = 6'h12 == _T_6589 ? _T_5936_18_is_store : _GEN_50886;
  assign _GEN_50978 = 6'h12 == _T_6589 ? _T_5936_18_is_load : _GEN_50888;
  assign _GEN_50979 = 6'h12 == _T_6589 ? _T_5936_18_is_sys_pc2epc : _GEN_50889;
  assign _GEN_50981 = 6'h12 == _T_6589 ? _T_5936_18_flush_on_commit : _GEN_50891;
  assign _GEN_50982 = 6'h12 == _T_6589 ? _T_5936_18_ldst : _GEN_50892;
  assign _GEN_50987 = 6'h12 == _T_6589 ? _T_5936_18_dst_rtype : _GEN_50897;
  assign _GEN_50991 = 6'h12 == _T_6589 ? _T_5936_18_fp_val : _GEN_50901;
  assign _GEN_51051 = 6'h13 == _T_6589 ? _T_5936_19_pdst : _GEN_50961;
  assign _GEN_51058 = 6'h13 == _T_6589 ? _T_5936_19_stale_pdst : _GEN_50968;
  assign _GEN_51065 = 6'h13 == _T_6589 ? _T_5936_19_is_fencei : _GEN_50975;
  assign _GEN_51066 = 6'h13 == _T_6589 ? _T_5936_19_is_store : _GEN_50976;
  assign _GEN_51068 = 6'h13 == _T_6589 ? _T_5936_19_is_load : _GEN_50978;
  assign _GEN_51069 = 6'h13 == _T_6589 ? _T_5936_19_is_sys_pc2epc : _GEN_50979;
  assign _GEN_51071 = 6'h13 == _T_6589 ? _T_5936_19_flush_on_commit : _GEN_50981;
  assign _GEN_51072 = 6'h13 == _T_6589 ? _T_5936_19_ldst : _GEN_50982;
  assign _GEN_51077 = 6'h13 == _T_6589 ? _T_5936_19_dst_rtype : _GEN_50987;
  assign _GEN_51081 = 6'h13 == _T_6589 ? _T_5936_19_fp_val : _GEN_50991;
  assign _GEN_51141 = 6'h14 == _T_6589 ? _T_5936_20_pdst : _GEN_51051;
  assign _GEN_51148 = 6'h14 == _T_6589 ? _T_5936_20_stale_pdst : _GEN_51058;
  assign _GEN_51155 = 6'h14 == _T_6589 ? _T_5936_20_is_fencei : _GEN_51065;
  assign _GEN_51156 = 6'h14 == _T_6589 ? _T_5936_20_is_store : _GEN_51066;
  assign _GEN_51158 = 6'h14 == _T_6589 ? _T_5936_20_is_load : _GEN_51068;
  assign _GEN_51159 = 6'h14 == _T_6589 ? _T_5936_20_is_sys_pc2epc : _GEN_51069;
  assign _GEN_51161 = 6'h14 == _T_6589 ? _T_5936_20_flush_on_commit : _GEN_51071;
  assign _GEN_51162 = 6'h14 == _T_6589 ? _T_5936_20_ldst : _GEN_51072;
  assign _GEN_51167 = 6'h14 == _T_6589 ? _T_5936_20_dst_rtype : _GEN_51077;
  assign _GEN_51171 = 6'h14 == _T_6589 ? _T_5936_20_fp_val : _GEN_51081;
  assign _GEN_51231 = 6'h15 == _T_6589 ? _T_5936_21_pdst : _GEN_51141;
  assign _GEN_51238 = 6'h15 == _T_6589 ? _T_5936_21_stale_pdst : _GEN_51148;
  assign _GEN_51245 = 6'h15 == _T_6589 ? _T_5936_21_is_fencei : _GEN_51155;
  assign _GEN_51246 = 6'h15 == _T_6589 ? _T_5936_21_is_store : _GEN_51156;
  assign _GEN_51248 = 6'h15 == _T_6589 ? _T_5936_21_is_load : _GEN_51158;
  assign _GEN_51249 = 6'h15 == _T_6589 ? _T_5936_21_is_sys_pc2epc : _GEN_51159;
  assign _GEN_51251 = 6'h15 == _T_6589 ? _T_5936_21_flush_on_commit : _GEN_51161;
  assign _GEN_51252 = 6'h15 == _T_6589 ? _T_5936_21_ldst : _GEN_51162;
  assign _GEN_51257 = 6'h15 == _T_6589 ? _T_5936_21_dst_rtype : _GEN_51167;
  assign _GEN_51261 = 6'h15 == _T_6589 ? _T_5936_21_fp_val : _GEN_51171;
  assign _GEN_51321 = 6'h16 == _T_6589 ? _T_5936_22_pdst : _GEN_51231;
  assign _GEN_51328 = 6'h16 == _T_6589 ? _T_5936_22_stale_pdst : _GEN_51238;
  assign _GEN_51335 = 6'h16 == _T_6589 ? _T_5936_22_is_fencei : _GEN_51245;
  assign _GEN_51336 = 6'h16 == _T_6589 ? _T_5936_22_is_store : _GEN_51246;
  assign _GEN_51338 = 6'h16 == _T_6589 ? _T_5936_22_is_load : _GEN_51248;
  assign _GEN_51339 = 6'h16 == _T_6589 ? _T_5936_22_is_sys_pc2epc : _GEN_51249;
  assign _GEN_51341 = 6'h16 == _T_6589 ? _T_5936_22_flush_on_commit : _GEN_51251;
  assign _GEN_51342 = 6'h16 == _T_6589 ? _T_5936_22_ldst : _GEN_51252;
  assign _GEN_51347 = 6'h16 == _T_6589 ? _T_5936_22_dst_rtype : _GEN_51257;
  assign _GEN_51351 = 6'h16 == _T_6589 ? _T_5936_22_fp_val : _GEN_51261;
  assign _GEN_51411 = 6'h17 == _T_6589 ? _T_5936_23_pdst : _GEN_51321;
  assign _GEN_51418 = 6'h17 == _T_6589 ? _T_5936_23_stale_pdst : _GEN_51328;
  assign _GEN_51425 = 6'h17 == _T_6589 ? _T_5936_23_is_fencei : _GEN_51335;
  assign _GEN_51426 = 6'h17 == _T_6589 ? _T_5936_23_is_store : _GEN_51336;
  assign _GEN_51428 = 6'h17 == _T_6589 ? _T_5936_23_is_load : _GEN_51338;
  assign _GEN_51429 = 6'h17 == _T_6589 ? _T_5936_23_is_sys_pc2epc : _GEN_51339;
  assign _GEN_51431 = 6'h17 == _T_6589 ? _T_5936_23_flush_on_commit : _GEN_51341;
  assign _GEN_51432 = 6'h17 == _T_6589 ? _T_5936_23_ldst : _GEN_51342;
  assign _GEN_51437 = 6'h17 == _T_6589 ? _T_5936_23_dst_rtype : _GEN_51347;
  assign _GEN_51441 = 6'h17 == _T_6589 ? _T_5936_23_fp_val : _GEN_51351;
  assign _GEN_51501 = 6'h18 == _T_6589 ? _T_5936_24_pdst : _GEN_51411;
  assign _GEN_51508 = 6'h18 == _T_6589 ? _T_5936_24_stale_pdst : _GEN_51418;
  assign _GEN_51515 = 6'h18 == _T_6589 ? _T_5936_24_is_fencei : _GEN_51425;
  assign _GEN_51516 = 6'h18 == _T_6589 ? _T_5936_24_is_store : _GEN_51426;
  assign _GEN_51518 = 6'h18 == _T_6589 ? _T_5936_24_is_load : _GEN_51428;
  assign _GEN_51519 = 6'h18 == _T_6589 ? _T_5936_24_is_sys_pc2epc : _GEN_51429;
  assign _GEN_51521 = 6'h18 == _T_6589 ? _T_5936_24_flush_on_commit : _GEN_51431;
  assign _GEN_51522 = 6'h18 == _T_6589 ? _T_5936_24_ldst : _GEN_51432;
  assign _GEN_51527 = 6'h18 == _T_6589 ? _T_5936_24_dst_rtype : _GEN_51437;
  assign _GEN_51531 = 6'h18 == _T_6589 ? _T_5936_24_fp_val : _GEN_51441;
  assign _GEN_51591 = 6'h19 == _T_6589 ? _T_5936_25_pdst : _GEN_51501;
  assign _GEN_51598 = 6'h19 == _T_6589 ? _T_5936_25_stale_pdst : _GEN_51508;
  assign _GEN_51605 = 6'h19 == _T_6589 ? _T_5936_25_is_fencei : _GEN_51515;
  assign _GEN_51606 = 6'h19 == _T_6589 ? _T_5936_25_is_store : _GEN_51516;
  assign _GEN_51608 = 6'h19 == _T_6589 ? _T_5936_25_is_load : _GEN_51518;
  assign _GEN_51609 = 6'h19 == _T_6589 ? _T_5936_25_is_sys_pc2epc : _GEN_51519;
  assign _GEN_51611 = 6'h19 == _T_6589 ? _T_5936_25_flush_on_commit : _GEN_51521;
  assign _GEN_51612 = 6'h19 == _T_6589 ? _T_5936_25_ldst : _GEN_51522;
  assign _GEN_51617 = 6'h19 == _T_6589 ? _T_5936_25_dst_rtype : _GEN_51527;
  assign _GEN_51621 = 6'h19 == _T_6589 ? _T_5936_25_fp_val : _GEN_51531;
  assign _GEN_51681 = 6'h1a == _T_6589 ? _T_5936_26_pdst : _GEN_51591;
  assign _GEN_51688 = 6'h1a == _T_6589 ? _T_5936_26_stale_pdst : _GEN_51598;
  assign _GEN_51695 = 6'h1a == _T_6589 ? _T_5936_26_is_fencei : _GEN_51605;
  assign _GEN_51696 = 6'h1a == _T_6589 ? _T_5936_26_is_store : _GEN_51606;
  assign _GEN_51698 = 6'h1a == _T_6589 ? _T_5936_26_is_load : _GEN_51608;
  assign _GEN_51699 = 6'h1a == _T_6589 ? _T_5936_26_is_sys_pc2epc : _GEN_51609;
  assign _GEN_51701 = 6'h1a == _T_6589 ? _T_5936_26_flush_on_commit : _GEN_51611;
  assign _GEN_51702 = 6'h1a == _T_6589 ? _T_5936_26_ldst : _GEN_51612;
  assign _GEN_51707 = 6'h1a == _T_6589 ? _T_5936_26_dst_rtype : _GEN_51617;
  assign _GEN_51711 = 6'h1a == _T_6589 ? _T_5936_26_fp_val : _GEN_51621;
  assign _GEN_51771 = 6'h1b == _T_6589 ? _T_5936_27_pdst : _GEN_51681;
  assign _GEN_51778 = 6'h1b == _T_6589 ? _T_5936_27_stale_pdst : _GEN_51688;
  assign _GEN_51785 = 6'h1b == _T_6589 ? _T_5936_27_is_fencei : _GEN_51695;
  assign _GEN_51786 = 6'h1b == _T_6589 ? _T_5936_27_is_store : _GEN_51696;
  assign _GEN_51788 = 6'h1b == _T_6589 ? _T_5936_27_is_load : _GEN_51698;
  assign _GEN_51789 = 6'h1b == _T_6589 ? _T_5936_27_is_sys_pc2epc : _GEN_51699;
  assign _GEN_51791 = 6'h1b == _T_6589 ? _T_5936_27_flush_on_commit : _GEN_51701;
  assign _GEN_51792 = 6'h1b == _T_6589 ? _T_5936_27_ldst : _GEN_51702;
  assign _GEN_51797 = 6'h1b == _T_6589 ? _T_5936_27_dst_rtype : _GEN_51707;
  assign _GEN_51801 = 6'h1b == _T_6589 ? _T_5936_27_fp_val : _GEN_51711;
  assign _GEN_51861 = 6'h1c == _T_6589 ? _T_5936_28_pdst : _GEN_51771;
  assign _GEN_51868 = 6'h1c == _T_6589 ? _T_5936_28_stale_pdst : _GEN_51778;
  assign _GEN_51875 = 6'h1c == _T_6589 ? _T_5936_28_is_fencei : _GEN_51785;
  assign _GEN_51876 = 6'h1c == _T_6589 ? _T_5936_28_is_store : _GEN_51786;
  assign _GEN_51878 = 6'h1c == _T_6589 ? _T_5936_28_is_load : _GEN_51788;
  assign _GEN_51879 = 6'h1c == _T_6589 ? _T_5936_28_is_sys_pc2epc : _GEN_51789;
  assign _GEN_51881 = 6'h1c == _T_6589 ? _T_5936_28_flush_on_commit : _GEN_51791;
  assign _GEN_51882 = 6'h1c == _T_6589 ? _T_5936_28_ldst : _GEN_51792;
  assign _GEN_51887 = 6'h1c == _T_6589 ? _T_5936_28_dst_rtype : _GEN_51797;
  assign _GEN_51891 = 6'h1c == _T_6589 ? _T_5936_28_fp_val : _GEN_51801;
  assign _GEN_51951 = 6'h1d == _T_6589 ? _T_5936_29_pdst : _GEN_51861;
  assign _GEN_51958 = 6'h1d == _T_6589 ? _T_5936_29_stale_pdst : _GEN_51868;
  assign _GEN_51965 = 6'h1d == _T_6589 ? _T_5936_29_is_fencei : _GEN_51875;
  assign _GEN_51966 = 6'h1d == _T_6589 ? _T_5936_29_is_store : _GEN_51876;
  assign _GEN_51968 = 6'h1d == _T_6589 ? _T_5936_29_is_load : _GEN_51878;
  assign _GEN_51969 = 6'h1d == _T_6589 ? _T_5936_29_is_sys_pc2epc : _GEN_51879;
  assign _GEN_51971 = 6'h1d == _T_6589 ? _T_5936_29_flush_on_commit : _GEN_51881;
  assign _GEN_51972 = 6'h1d == _T_6589 ? _T_5936_29_ldst : _GEN_51882;
  assign _GEN_51977 = 6'h1d == _T_6589 ? _T_5936_29_dst_rtype : _GEN_51887;
  assign _GEN_51981 = 6'h1d == _T_6589 ? _T_5936_29_fp_val : _GEN_51891;
  assign _GEN_52041 = 6'h1e == _T_6589 ? _T_5936_30_pdst : _GEN_51951;
  assign _GEN_52048 = 6'h1e == _T_6589 ? _T_5936_30_stale_pdst : _GEN_51958;
  assign _GEN_52055 = 6'h1e == _T_6589 ? _T_5936_30_is_fencei : _GEN_51965;
  assign _GEN_52056 = 6'h1e == _T_6589 ? _T_5936_30_is_store : _GEN_51966;
  assign _GEN_52058 = 6'h1e == _T_6589 ? _T_5936_30_is_load : _GEN_51968;
  assign _GEN_52059 = 6'h1e == _T_6589 ? _T_5936_30_is_sys_pc2epc : _GEN_51969;
  assign _GEN_52061 = 6'h1e == _T_6589 ? _T_5936_30_flush_on_commit : _GEN_51971;
  assign _GEN_52062 = 6'h1e == _T_6589 ? _T_5936_30_ldst : _GEN_51972;
  assign _GEN_52067 = 6'h1e == _T_6589 ? _T_5936_30_dst_rtype : _GEN_51977;
  assign _GEN_52071 = 6'h1e == _T_6589 ? _T_5936_30_fp_val : _GEN_51981;
  assign _GEN_52131 = 6'h1f == _T_6589 ? _T_5936_31_pdst : _GEN_52041;
  assign _GEN_52138 = 6'h1f == _T_6589 ? _T_5936_31_stale_pdst : _GEN_52048;
  assign _GEN_52145 = 6'h1f == _T_6589 ? _T_5936_31_is_fencei : _GEN_52055;
  assign _GEN_52146 = 6'h1f == _T_6589 ? _T_5936_31_is_store : _GEN_52056;
  assign _GEN_52148 = 6'h1f == _T_6589 ? _T_5936_31_is_load : _GEN_52058;
  assign _GEN_52149 = 6'h1f == _T_6589 ? _T_5936_31_is_sys_pc2epc : _GEN_52059;
  assign _GEN_52151 = 6'h1f == _T_6589 ? _T_5936_31_flush_on_commit : _GEN_52061;
  assign _GEN_52152 = 6'h1f == _T_6589 ? _T_5936_31_ldst : _GEN_52062;
  assign _GEN_52157 = 6'h1f == _T_6589 ? _T_5936_31_dst_rtype : _GEN_52067;
  assign _GEN_52161 = 6'h1f == _T_6589 ? _T_5936_31_fp_val : _GEN_52071;
  assign _GEN_52221 = 6'h20 == _T_6589 ? _T_5936_32_pdst : _GEN_52131;
  assign _GEN_52228 = 6'h20 == _T_6589 ? _T_5936_32_stale_pdst : _GEN_52138;
  assign _GEN_52235 = 6'h20 == _T_6589 ? _T_5936_32_is_fencei : _GEN_52145;
  assign _GEN_52236 = 6'h20 == _T_6589 ? _T_5936_32_is_store : _GEN_52146;
  assign _GEN_52238 = 6'h20 == _T_6589 ? _T_5936_32_is_load : _GEN_52148;
  assign _GEN_52239 = 6'h20 == _T_6589 ? _T_5936_32_is_sys_pc2epc : _GEN_52149;
  assign _GEN_52241 = 6'h20 == _T_6589 ? _T_5936_32_flush_on_commit : _GEN_52151;
  assign _GEN_52242 = 6'h20 == _T_6589 ? _T_5936_32_ldst : _GEN_52152;
  assign _GEN_52247 = 6'h20 == _T_6589 ? _T_5936_32_dst_rtype : _GEN_52157;
  assign _GEN_52251 = 6'h20 == _T_6589 ? _T_5936_32_fp_val : _GEN_52161;
  assign _GEN_52311 = 6'h21 == _T_6589 ? _T_5936_33_pdst : _GEN_52221;
  assign _GEN_52318 = 6'h21 == _T_6589 ? _T_5936_33_stale_pdst : _GEN_52228;
  assign _GEN_52325 = 6'h21 == _T_6589 ? _T_5936_33_is_fencei : _GEN_52235;
  assign _GEN_52326 = 6'h21 == _T_6589 ? _T_5936_33_is_store : _GEN_52236;
  assign _GEN_52328 = 6'h21 == _T_6589 ? _T_5936_33_is_load : _GEN_52238;
  assign _GEN_52329 = 6'h21 == _T_6589 ? _T_5936_33_is_sys_pc2epc : _GEN_52239;
  assign _GEN_52331 = 6'h21 == _T_6589 ? _T_5936_33_flush_on_commit : _GEN_52241;
  assign _GEN_52332 = 6'h21 == _T_6589 ? _T_5936_33_ldst : _GEN_52242;
  assign _GEN_52337 = 6'h21 == _T_6589 ? _T_5936_33_dst_rtype : _GEN_52247;
  assign _GEN_52341 = 6'h21 == _T_6589 ? _T_5936_33_fp_val : _GEN_52251;
  assign _GEN_52401 = 6'h22 == _T_6589 ? _T_5936_34_pdst : _GEN_52311;
  assign _GEN_52408 = 6'h22 == _T_6589 ? _T_5936_34_stale_pdst : _GEN_52318;
  assign _GEN_52415 = 6'h22 == _T_6589 ? _T_5936_34_is_fencei : _GEN_52325;
  assign _GEN_52416 = 6'h22 == _T_6589 ? _T_5936_34_is_store : _GEN_52326;
  assign _GEN_52418 = 6'h22 == _T_6589 ? _T_5936_34_is_load : _GEN_52328;
  assign _GEN_52419 = 6'h22 == _T_6589 ? _T_5936_34_is_sys_pc2epc : _GEN_52329;
  assign _GEN_52421 = 6'h22 == _T_6589 ? _T_5936_34_flush_on_commit : _GEN_52331;
  assign _GEN_52422 = 6'h22 == _T_6589 ? _T_5936_34_ldst : _GEN_52332;
  assign _GEN_52427 = 6'h22 == _T_6589 ? _T_5936_34_dst_rtype : _GEN_52337;
  assign _GEN_52431 = 6'h22 == _T_6589 ? _T_5936_34_fp_val : _GEN_52341;
  assign _GEN_52491 = 6'h23 == _T_6589 ? _T_5936_35_pdst : _GEN_52401;
  assign _GEN_52498 = 6'h23 == _T_6589 ? _T_5936_35_stale_pdst : _GEN_52408;
  assign _GEN_52505 = 6'h23 == _T_6589 ? _T_5936_35_is_fencei : _GEN_52415;
  assign _GEN_52506 = 6'h23 == _T_6589 ? _T_5936_35_is_store : _GEN_52416;
  assign _GEN_52508 = 6'h23 == _T_6589 ? _T_5936_35_is_load : _GEN_52418;
  assign _GEN_52509 = 6'h23 == _T_6589 ? _T_5936_35_is_sys_pc2epc : _GEN_52419;
  assign _GEN_52511 = 6'h23 == _T_6589 ? _T_5936_35_flush_on_commit : _GEN_52421;
  assign _GEN_52512 = 6'h23 == _T_6589 ? _T_5936_35_ldst : _GEN_52422;
  assign _GEN_52517 = 6'h23 == _T_6589 ? _T_5936_35_dst_rtype : _GEN_52427;
  assign _GEN_52521 = 6'h23 == _T_6589 ? _T_5936_35_fp_val : _GEN_52431;
  assign _GEN_52581 = 6'h24 == _T_6589 ? _T_5936_36_pdst : _GEN_52491;
  assign _GEN_52588 = 6'h24 == _T_6589 ? _T_5936_36_stale_pdst : _GEN_52498;
  assign _GEN_52595 = 6'h24 == _T_6589 ? _T_5936_36_is_fencei : _GEN_52505;
  assign _GEN_52596 = 6'h24 == _T_6589 ? _T_5936_36_is_store : _GEN_52506;
  assign _GEN_52598 = 6'h24 == _T_6589 ? _T_5936_36_is_load : _GEN_52508;
  assign _GEN_52599 = 6'h24 == _T_6589 ? _T_5936_36_is_sys_pc2epc : _GEN_52509;
  assign _GEN_52601 = 6'h24 == _T_6589 ? _T_5936_36_flush_on_commit : _GEN_52511;
  assign _GEN_52602 = 6'h24 == _T_6589 ? _T_5936_36_ldst : _GEN_52512;
  assign _GEN_52607 = 6'h24 == _T_6589 ? _T_5936_36_dst_rtype : _GEN_52517;
  assign _GEN_52611 = 6'h24 == _T_6589 ? _T_5936_36_fp_val : _GEN_52521;
  assign _GEN_52671 = 6'h25 == _T_6589 ? _T_5936_37_pdst : _GEN_52581;
  assign _GEN_52678 = 6'h25 == _T_6589 ? _T_5936_37_stale_pdst : _GEN_52588;
  assign _GEN_52685 = 6'h25 == _T_6589 ? _T_5936_37_is_fencei : _GEN_52595;
  assign _GEN_52686 = 6'h25 == _T_6589 ? _T_5936_37_is_store : _GEN_52596;
  assign _GEN_52688 = 6'h25 == _T_6589 ? _T_5936_37_is_load : _GEN_52598;
  assign _GEN_52689 = 6'h25 == _T_6589 ? _T_5936_37_is_sys_pc2epc : _GEN_52599;
  assign _GEN_52691 = 6'h25 == _T_6589 ? _T_5936_37_flush_on_commit : _GEN_52601;
  assign _GEN_52692 = 6'h25 == _T_6589 ? _T_5936_37_ldst : _GEN_52602;
  assign _GEN_52697 = 6'h25 == _T_6589 ? _T_5936_37_dst_rtype : _GEN_52607;
  assign _GEN_52701 = 6'h25 == _T_6589 ? _T_5936_37_fp_val : _GEN_52611;
  assign _GEN_52761 = 6'h26 == _T_6589 ? _T_5936_38_pdst : _GEN_52671;
  assign _GEN_52768 = 6'h26 == _T_6589 ? _T_5936_38_stale_pdst : _GEN_52678;
  assign _GEN_52775 = 6'h26 == _T_6589 ? _T_5936_38_is_fencei : _GEN_52685;
  assign _GEN_52776 = 6'h26 == _T_6589 ? _T_5936_38_is_store : _GEN_52686;
  assign _GEN_52778 = 6'h26 == _T_6589 ? _T_5936_38_is_load : _GEN_52688;
  assign _GEN_52779 = 6'h26 == _T_6589 ? _T_5936_38_is_sys_pc2epc : _GEN_52689;
  assign _GEN_52781 = 6'h26 == _T_6589 ? _T_5936_38_flush_on_commit : _GEN_52691;
  assign _GEN_52782 = 6'h26 == _T_6589 ? _T_5936_38_ldst : _GEN_52692;
  assign _GEN_52787 = 6'h26 == _T_6589 ? _T_5936_38_dst_rtype : _GEN_52697;
  assign _GEN_52791 = 6'h26 == _T_6589 ? _T_5936_38_fp_val : _GEN_52701;
  assign _GEN_52851 = 6'h27 == _T_6589 ? _T_5936_39_pdst : _GEN_52761;
  assign _GEN_52858 = 6'h27 == _T_6589 ? _T_5936_39_stale_pdst : _GEN_52768;
  assign _GEN_52865 = 6'h27 == _T_6589 ? _T_5936_39_is_fencei : _GEN_52775;
  assign _GEN_52866 = 6'h27 == _T_6589 ? _T_5936_39_is_store : _GEN_52776;
  assign _GEN_52868 = 6'h27 == _T_6589 ? _T_5936_39_is_load : _GEN_52778;
  assign _GEN_52869 = 6'h27 == _T_6589 ? _T_5936_39_is_sys_pc2epc : _GEN_52779;
  assign _GEN_52871 = 6'h27 == _T_6589 ? _T_5936_39_flush_on_commit : _GEN_52781;
  assign _GEN_52872 = 6'h27 == _T_6589 ? _T_5936_39_ldst : _GEN_52782;
  assign _GEN_52877 = 6'h27 == _T_6589 ? _T_5936_39_dst_rtype : _GEN_52787;
  assign _GEN_52881 = 6'h27 == _T_6589 ? _T_5936_39_fp_val : _GEN_52791;
  assign _GEN_52889 = 6'h1 == _T_6589 ? _T_5637_1 : _T_5637_0;
  assign _GEN_52890 = 6'h2 == _T_6589 ? _T_5637_2 : _GEN_52889;
  assign _GEN_52891 = 6'h3 == _T_6589 ? _T_5637_3 : _GEN_52890;
  assign _GEN_52892 = 6'h4 == _T_6589 ? _T_5637_4 : _GEN_52891;
  assign _GEN_52893 = 6'h5 == _T_6589 ? _T_5637_5 : _GEN_52892;
  assign _GEN_52894 = 6'h6 == _T_6589 ? _T_5637_6 : _GEN_52893;
  assign _GEN_52895 = 6'h7 == _T_6589 ? _T_5637_7 : _GEN_52894;
  assign _GEN_52896 = 6'h8 == _T_6589 ? _T_5637_8 : _GEN_52895;
  assign _GEN_52897 = 6'h9 == _T_6589 ? _T_5637_9 : _GEN_52896;
  assign _GEN_52898 = 6'ha == _T_6589 ? _T_5637_10 : _GEN_52897;
  assign _GEN_52899 = 6'hb == _T_6589 ? _T_5637_11 : _GEN_52898;
  assign _GEN_52900 = 6'hc == _T_6589 ? _T_5637_12 : _GEN_52899;
  assign _GEN_52901 = 6'hd == _T_6589 ? _T_5637_13 : _GEN_52900;
  assign _GEN_52902 = 6'he == _T_6589 ? _T_5637_14 : _GEN_52901;
  assign _GEN_52903 = 6'hf == _T_6589 ? _T_5637_15 : _GEN_52902;
  assign _GEN_52904 = 6'h10 == _T_6589 ? _T_5637_16 : _GEN_52903;
  assign _GEN_52905 = 6'h11 == _T_6589 ? _T_5637_17 : _GEN_52904;
  assign _GEN_52906 = 6'h12 == _T_6589 ? _T_5637_18 : _GEN_52905;
  assign _GEN_52907 = 6'h13 == _T_6589 ? _T_5637_19 : _GEN_52906;
  assign _GEN_52908 = 6'h14 == _T_6589 ? _T_5637_20 : _GEN_52907;
  assign _GEN_52909 = 6'h15 == _T_6589 ? _T_5637_21 : _GEN_52908;
  assign _GEN_52910 = 6'h16 == _T_6589 ? _T_5637_22 : _GEN_52909;
  assign _GEN_52911 = 6'h17 == _T_6589 ? _T_5637_23 : _GEN_52910;
  assign _GEN_52912 = 6'h18 == _T_6589 ? _T_5637_24 : _GEN_52911;
  assign _GEN_52913 = 6'h19 == _T_6589 ? _T_5637_25 : _GEN_52912;
  assign _GEN_52914 = 6'h1a == _T_6589 ? _T_5637_26 : _GEN_52913;
  assign _GEN_52915 = 6'h1b == _T_6589 ? _T_5637_27 : _GEN_52914;
  assign _GEN_52916 = 6'h1c == _T_6589 ? _T_5637_28 : _GEN_52915;
  assign _GEN_52917 = 6'h1d == _T_6589 ? _T_5637_29 : _GEN_52916;
  assign _GEN_52918 = 6'h1e == _T_6589 ? _T_5637_30 : _GEN_52917;
  assign _GEN_52919 = 6'h1f == _T_6589 ? _T_5637_31 : _GEN_52918;
  assign _GEN_52920 = 6'h20 == _T_6589 ? _T_5637_32 : _GEN_52919;
  assign _GEN_52921 = 6'h21 == _T_6589 ? _T_5637_33 : _GEN_52920;
  assign _GEN_52922 = 6'h22 == _T_6589 ? _T_5637_34 : _GEN_52921;
  assign _GEN_52923 = 6'h23 == _T_6589 ? _T_5637_35 : _GEN_52922;
  assign _GEN_52924 = 6'h24 == _T_6589 ? _T_5637_36 : _GEN_52923;
  assign _GEN_52925 = 6'h25 == _T_6589 ? _T_5637_37 : _GEN_52924;
  assign _GEN_52926 = 6'h26 == _T_6589 ? _T_5637_38 : _GEN_52925;
  assign _GEN_52927 = 6'h27 == _T_6589 ? _T_5637_39 : _GEN_52926;
  assign _T_6610 = _T_4026 & _GEN_422;
  assign _T_6623 = _GEN_423_dst_rtype == 2'h0;
  assign _T_6636 = _GEN_424_dst_rtype == 2'h1;
  assign _T_6637 = _T_6623 | _T_6636;
  assign _T_6638 = _T_6610 & _T_6637;
  assign _T_6641 = rob_state == 2'h2;
  assign _GEN_59948 = 6'h0 == _T_6589 ? 1'h0 : _GEN_45169;
  assign _GEN_59949 = 6'h1 == _T_6589 ? 1'h0 : _GEN_45170;
  assign _GEN_59950 = 6'h2 == _T_6589 ? 1'h0 : _GEN_45171;
  assign _GEN_59951 = 6'h3 == _T_6589 ? 1'h0 : _GEN_45172;
  assign _GEN_59952 = 6'h4 == _T_6589 ? 1'h0 : _GEN_45173;
  assign _GEN_59953 = 6'h5 == _T_6589 ? 1'h0 : _GEN_45174;
  assign _GEN_59954 = 6'h6 == _T_6589 ? 1'h0 : _GEN_45175;
  assign _GEN_59955 = 6'h7 == _T_6589 ? 1'h0 : _GEN_45176;
  assign _GEN_59956 = 6'h8 == _T_6589 ? 1'h0 : _GEN_45177;
  assign _GEN_59957 = 6'h9 == _T_6589 ? 1'h0 : _GEN_45178;
  assign _GEN_59958 = 6'ha == _T_6589 ? 1'h0 : _GEN_45179;
  assign _GEN_59959 = 6'hb == _T_6589 ? 1'h0 : _GEN_45180;
  assign _GEN_59960 = 6'hc == _T_6589 ? 1'h0 : _GEN_45181;
  assign _GEN_59961 = 6'hd == _T_6589 ? 1'h0 : _GEN_45182;
  assign _GEN_59962 = 6'he == _T_6589 ? 1'h0 : _GEN_45183;
  assign _GEN_59963 = 6'hf == _T_6589 ? 1'h0 : _GEN_45184;
  assign _GEN_59964 = 6'h10 == _T_6589 ? 1'h0 : _GEN_45185;
  assign _GEN_59965 = 6'h11 == _T_6589 ? 1'h0 : _GEN_45186;
  assign _GEN_59966 = 6'h12 == _T_6589 ? 1'h0 : _GEN_45187;
  assign _GEN_59967 = 6'h13 == _T_6589 ? 1'h0 : _GEN_45188;
  assign _GEN_59968 = 6'h14 == _T_6589 ? 1'h0 : _GEN_45189;
  assign _GEN_59969 = 6'h15 == _T_6589 ? 1'h0 : _GEN_45190;
  assign _GEN_59970 = 6'h16 == _T_6589 ? 1'h0 : _GEN_45191;
  assign _GEN_59971 = 6'h17 == _T_6589 ? 1'h0 : _GEN_45192;
  assign _GEN_59972 = 6'h18 == _T_6589 ? 1'h0 : _GEN_45193;
  assign _GEN_59973 = 6'h19 == _T_6589 ? 1'h0 : _GEN_45194;
  assign _GEN_59974 = 6'h1a == _T_6589 ? 1'h0 : _GEN_45195;
  assign _GEN_59975 = 6'h1b == _T_6589 ? 1'h0 : _GEN_45196;
  assign _GEN_59976 = 6'h1c == _T_6589 ? 1'h0 : _GEN_45197;
  assign _GEN_59977 = 6'h1d == _T_6589 ? 1'h0 : _GEN_45198;
  assign _GEN_59978 = 6'h1e == _T_6589 ? 1'h0 : _GEN_45199;
  assign _GEN_59979 = 6'h1f == _T_6589 ? 1'h0 : _GEN_45200;
  assign _GEN_59980 = 6'h20 == _T_6589 ? 1'h0 : _GEN_45201;
  assign _GEN_59981 = 6'h21 == _T_6589 ? 1'h0 : _GEN_45202;
  assign _GEN_59982 = 6'h22 == _T_6589 ? 1'h0 : _GEN_45203;
  assign _GEN_59983 = 6'h23 == _T_6589 ? 1'h0 : _GEN_45204;
  assign _GEN_59984 = 6'h24 == _T_6589 ? 1'h0 : _GEN_45205;
  assign _GEN_59985 = 6'h25 == _T_6589 ? 1'h0 : _GEN_45206;
  assign _GEN_59986 = 6'h26 == _T_6589 ? 1'h0 : _GEN_45207;
  assign _GEN_59987 = 6'h27 == _T_6589 ? 1'h0 : _GEN_45208;
  assign _GEN_59988 = _T_4026 ? _GEN_59948 : _GEN_45169;
  assign _GEN_59989 = _T_4026 ? _GEN_59949 : _GEN_45170;
  assign _GEN_59990 = _T_4026 ? _GEN_59950 : _GEN_45171;
  assign _GEN_59991 = _T_4026 ? _GEN_59951 : _GEN_45172;
  assign _GEN_59992 = _T_4026 ? _GEN_59952 : _GEN_45173;
  assign _GEN_59993 = _T_4026 ? _GEN_59953 : _GEN_45174;
  assign _GEN_59994 = _T_4026 ? _GEN_59954 : _GEN_45175;
  assign _GEN_59995 = _T_4026 ? _GEN_59955 : _GEN_45176;
  assign _GEN_59996 = _T_4026 ? _GEN_59956 : _GEN_45177;
  assign _GEN_59997 = _T_4026 ? _GEN_59957 : _GEN_45178;
  assign _GEN_59998 = _T_4026 ? _GEN_59958 : _GEN_45179;
  assign _GEN_59999 = _T_4026 ? _GEN_59959 : _GEN_45180;
  assign _GEN_60000 = _T_4026 ? _GEN_59960 : _GEN_45181;
  assign _GEN_60001 = _T_4026 ? _GEN_59961 : _GEN_45182;
  assign _GEN_60002 = _T_4026 ? _GEN_59962 : _GEN_45183;
  assign _GEN_60003 = _T_4026 ? _GEN_59963 : _GEN_45184;
  assign _GEN_60004 = _T_4026 ? _GEN_59964 : _GEN_45185;
  assign _GEN_60005 = _T_4026 ? _GEN_59965 : _GEN_45186;
  assign _GEN_60006 = _T_4026 ? _GEN_59966 : _GEN_45187;
  assign _GEN_60007 = _T_4026 ? _GEN_59967 : _GEN_45188;
  assign _GEN_60008 = _T_4026 ? _GEN_59968 : _GEN_45189;
  assign _GEN_60009 = _T_4026 ? _GEN_59969 : _GEN_45190;
  assign _GEN_60010 = _T_4026 ? _GEN_59970 : _GEN_45191;
  assign _GEN_60011 = _T_4026 ? _GEN_59971 : _GEN_45192;
  assign _GEN_60012 = _T_4026 ? _GEN_59972 : _GEN_45193;
  assign _GEN_60013 = _T_4026 ? _GEN_59973 : _GEN_45194;
  assign _GEN_60014 = _T_4026 ? _GEN_59974 : _GEN_45195;
  assign _GEN_60015 = _T_4026 ? _GEN_59975 : _GEN_45196;
  assign _GEN_60016 = _T_4026 ? _GEN_59976 : _GEN_45197;
  assign _GEN_60017 = _T_4026 ? _GEN_59977 : _GEN_45198;
  assign _GEN_60018 = _T_4026 ? _GEN_59978 : _GEN_45199;
  assign _GEN_60019 = _T_4026 ? _GEN_59979 : _GEN_45200;
  assign _GEN_60020 = _T_4026 ? _GEN_59980 : _GEN_45201;
  assign _GEN_60021 = _T_4026 ? _GEN_59981 : _GEN_45202;
  assign _GEN_60022 = _T_4026 ? _GEN_59982 : _GEN_45203;
  assign _GEN_60023 = _T_4026 ? _GEN_59983 : _GEN_45204;
  assign _GEN_60024 = _T_4026 ? _GEN_59984 : _GEN_45205;
  assign _GEN_60025 = _T_4026 ? _GEN_59985 : _GEN_45206;
  assign _GEN_60026 = _T_4026 ? _GEN_59986 : _GEN_45207;
  assign _GEN_60027 = _T_4026 ? _GEN_59987 : _GEN_45208;
  assign _T_6654 = io_brinfo_mask & _T_5936_0_br_mask;
  assign _T_6656 = _T_6654 != 8'h0;
  assign _T_6657 = _T_5637_0 & _T_6656;
  assign _T_6659 = _T_4094 & _T_6657;
  assign _T_6674 = _T_4109 & _T_6657;
  assign _T_6676 = _T_5936_0_br_mask & _T_4111;
  assign _GEN_60032 = _T_6674 ? _T_6676 : _GEN_46173;
  assign _GEN_60033 = _T_6659 ? 1'h0 : _GEN_59988;
  assign _GEN_60035 = _T_6659 ? _GEN_46173 : _GEN_60032;
  assign _T_6677 = io_brinfo_mask & _T_5936_1_br_mask;
  assign _T_6679 = _T_6677 != 8'h0;
  assign _T_6680 = _T_5637_1 & _T_6679;
  assign _T_6682 = _T_4094 & _T_6680;
  assign _T_6697 = _T_4109 & _T_6680;
  assign _T_6699 = _T_5936_1_br_mask & _T_4111;
  assign _GEN_60036 = _T_6697 ? _T_6699 : _GEN_46174;
  assign _GEN_60037 = _T_6682 ? 1'h0 : _GEN_59989;
  assign _GEN_60039 = _T_6682 ? _GEN_46174 : _GEN_60036;
  assign _T_6700 = io_brinfo_mask & _T_5936_2_br_mask;
  assign _T_6702 = _T_6700 != 8'h0;
  assign _T_6703 = _T_5637_2 & _T_6702;
  assign _T_6705 = _T_4094 & _T_6703;
  assign _T_6720 = _T_4109 & _T_6703;
  assign _T_6722 = _T_5936_2_br_mask & _T_4111;
  assign _GEN_60040 = _T_6720 ? _T_6722 : _GEN_46175;
  assign _GEN_60041 = _T_6705 ? 1'h0 : _GEN_59990;
  assign _GEN_60043 = _T_6705 ? _GEN_46175 : _GEN_60040;
  assign _T_6723 = io_brinfo_mask & _T_5936_3_br_mask;
  assign _T_6725 = _T_6723 != 8'h0;
  assign _T_6726 = _T_5637_3 & _T_6725;
  assign _T_6728 = _T_4094 & _T_6726;
  assign _T_6743 = _T_4109 & _T_6726;
  assign _T_6745 = _T_5936_3_br_mask & _T_4111;
  assign _GEN_60044 = _T_6743 ? _T_6745 : _GEN_46176;
  assign _GEN_60045 = _T_6728 ? 1'h0 : _GEN_59991;
  assign _GEN_60047 = _T_6728 ? _GEN_46176 : _GEN_60044;
  assign _T_6746 = io_brinfo_mask & _T_5936_4_br_mask;
  assign _T_6748 = _T_6746 != 8'h0;
  assign _T_6749 = _T_5637_4 & _T_6748;
  assign _T_6751 = _T_4094 & _T_6749;
  assign _T_6766 = _T_4109 & _T_6749;
  assign _T_6768 = _T_5936_4_br_mask & _T_4111;
  assign _GEN_60048 = _T_6766 ? _T_6768 : _GEN_46177;
  assign _GEN_60049 = _T_6751 ? 1'h0 : _GEN_59992;
  assign _GEN_60051 = _T_6751 ? _GEN_46177 : _GEN_60048;
  assign _T_6769 = io_brinfo_mask & _T_5936_5_br_mask;
  assign _T_6771 = _T_6769 != 8'h0;
  assign _T_6772 = _T_5637_5 & _T_6771;
  assign _T_6774 = _T_4094 & _T_6772;
  assign _T_6789 = _T_4109 & _T_6772;
  assign _T_6791 = _T_5936_5_br_mask & _T_4111;
  assign _GEN_60052 = _T_6789 ? _T_6791 : _GEN_46178;
  assign _GEN_60053 = _T_6774 ? 1'h0 : _GEN_59993;
  assign _GEN_60055 = _T_6774 ? _GEN_46178 : _GEN_60052;
  assign _T_6792 = io_brinfo_mask & _T_5936_6_br_mask;
  assign _T_6794 = _T_6792 != 8'h0;
  assign _T_6795 = _T_5637_6 & _T_6794;
  assign _T_6797 = _T_4094 & _T_6795;
  assign _T_6812 = _T_4109 & _T_6795;
  assign _T_6814 = _T_5936_6_br_mask & _T_4111;
  assign _GEN_60056 = _T_6812 ? _T_6814 : _GEN_46179;
  assign _GEN_60057 = _T_6797 ? 1'h0 : _GEN_59994;
  assign _GEN_60059 = _T_6797 ? _GEN_46179 : _GEN_60056;
  assign _T_6815 = io_brinfo_mask & _T_5936_7_br_mask;
  assign _T_6817 = _T_6815 != 8'h0;
  assign _T_6818 = _T_5637_7 & _T_6817;
  assign _T_6820 = _T_4094 & _T_6818;
  assign _T_6835 = _T_4109 & _T_6818;
  assign _T_6837 = _T_5936_7_br_mask & _T_4111;
  assign _GEN_60060 = _T_6835 ? _T_6837 : _GEN_46180;
  assign _GEN_60061 = _T_6820 ? 1'h0 : _GEN_59995;
  assign _GEN_60063 = _T_6820 ? _GEN_46180 : _GEN_60060;
  assign _T_6838 = io_brinfo_mask & _T_5936_8_br_mask;
  assign _T_6840 = _T_6838 != 8'h0;
  assign _T_6841 = _T_5637_8 & _T_6840;
  assign _T_6843 = _T_4094 & _T_6841;
  assign _T_6858 = _T_4109 & _T_6841;
  assign _T_6860 = _T_5936_8_br_mask & _T_4111;
  assign _GEN_60064 = _T_6858 ? _T_6860 : _GEN_46181;
  assign _GEN_60065 = _T_6843 ? 1'h0 : _GEN_59996;
  assign _GEN_60067 = _T_6843 ? _GEN_46181 : _GEN_60064;
  assign _T_6861 = io_brinfo_mask & _T_5936_9_br_mask;
  assign _T_6863 = _T_6861 != 8'h0;
  assign _T_6864 = _T_5637_9 & _T_6863;
  assign _T_6866 = _T_4094 & _T_6864;
  assign _T_6881 = _T_4109 & _T_6864;
  assign _T_6883 = _T_5936_9_br_mask & _T_4111;
  assign _GEN_60068 = _T_6881 ? _T_6883 : _GEN_46182;
  assign _GEN_60069 = _T_6866 ? 1'h0 : _GEN_59997;
  assign _GEN_60071 = _T_6866 ? _GEN_46182 : _GEN_60068;
  assign _T_6884 = io_brinfo_mask & _T_5936_10_br_mask;
  assign _T_6886 = _T_6884 != 8'h0;
  assign _T_6887 = _T_5637_10 & _T_6886;
  assign _T_6889 = _T_4094 & _T_6887;
  assign _T_6904 = _T_4109 & _T_6887;
  assign _T_6906 = _T_5936_10_br_mask & _T_4111;
  assign _GEN_60072 = _T_6904 ? _T_6906 : _GEN_46183;
  assign _GEN_60073 = _T_6889 ? 1'h0 : _GEN_59998;
  assign _GEN_60075 = _T_6889 ? _GEN_46183 : _GEN_60072;
  assign _T_6907 = io_brinfo_mask & _T_5936_11_br_mask;
  assign _T_6909 = _T_6907 != 8'h0;
  assign _T_6910 = _T_5637_11 & _T_6909;
  assign _T_6912 = _T_4094 & _T_6910;
  assign _T_6927 = _T_4109 & _T_6910;
  assign _T_6929 = _T_5936_11_br_mask & _T_4111;
  assign _GEN_60076 = _T_6927 ? _T_6929 : _GEN_46184;
  assign _GEN_60077 = _T_6912 ? 1'h0 : _GEN_59999;
  assign _GEN_60079 = _T_6912 ? _GEN_46184 : _GEN_60076;
  assign _T_6930 = io_brinfo_mask & _T_5936_12_br_mask;
  assign _T_6932 = _T_6930 != 8'h0;
  assign _T_6933 = _T_5637_12 & _T_6932;
  assign _T_6935 = _T_4094 & _T_6933;
  assign _T_6950 = _T_4109 & _T_6933;
  assign _T_6952 = _T_5936_12_br_mask & _T_4111;
  assign _GEN_60080 = _T_6950 ? _T_6952 : _GEN_46185;
  assign _GEN_60081 = _T_6935 ? 1'h0 : _GEN_60000;
  assign _GEN_60083 = _T_6935 ? _GEN_46185 : _GEN_60080;
  assign _T_6953 = io_brinfo_mask & _T_5936_13_br_mask;
  assign _T_6955 = _T_6953 != 8'h0;
  assign _T_6956 = _T_5637_13 & _T_6955;
  assign _T_6958 = _T_4094 & _T_6956;
  assign _T_6973 = _T_4109 & _T_6956;
  assign _T_6975 = _T_5936_13_br_mask & _T_4111;
  assign _GEN_60084 = _T_6973 ? _T_6975 : _GEN_46186;
  assign _GEN_60085 = _T_6958 ? 1'h0 : _GEN_60001;
  assign _GEN_60087 = _T_6958 ? _GEN_46186 : _GEN_60084;
  assign _T_6976 = io_brinfo_mask & _T_5936_14_br_mask;
  assign _T_6978 = _T_6976 != 8'h0;
  assign _T_6979 = _T_5637_14 & _T_6978;
  assign _T_6981 = _T_4094 & _T_6979;
  assign _T_6996 = _T_4109 & _T_6979;
  assign _T_6998 = _T_5936_14_br_mask & _T_4111;
  assign _GEN_60088 = _T_6996 ? _T_6998 : _GEN_46187;
  assign _GEN_60089 = _T_6981 ? 1'h0 : _GEN_60002;
  assign _GEN_60091 = _T_6981 ? _GEN_46187 : _GEN_60088;
  assign _T_6999 = io_brinfo_mask & _T_5936_15_br_mask;
  assign _T_7001 = _T_6999 != 8'h0;
  assign _T_7002 = _T_5637_15 & _T_7001;
  assign _T_7004 = _T_4094 & _T_7002;
  assign _T_7019 = _T_4109 & _T_7002;
  assign _T_7021 = _T_5936_15_br_mask & _T_4111;
  assign _GEN_60092 = _T_7019 ? _T_7021 : _GEN_46188;
  assign _GEN_60093 = _T_7004 ? 1'h0 : _GEN_60003;
  assign _GEN_60095 = _T_7004 ? _GEN_46188 : _GEN_60092;
  assign _T_7022 = io_brinfo_mask & _T_5936_16_br_mask;
  assign _T_7024 = _T_7022 != 8'h0;
  assign _T_7025 = _T_5637_16 & _T_7024;
  assign _T_7027 = _T_4094 & _T_7025;
  assign _T_7042 = _T_4109 & _T_7025;
  assign _T_7044 = _T_5936_16_br_mask & _T_4111;
  assign _GEN_60096 = _T_7042 ? _T_7044 : _GEN_46189;
  assign _GEN_60097 = _T_7027 ? 1'h0 : _GEN_60004;
  assign _GEN_60099 = _T_7027 ? _GEN_46189 : _GEN_60096;
  assign _T_7045 = io_brinfo_mask & _T_5936_17_br_mask;
  assign _T_7047 = _T_7045 != 8'h0;
  assign _T_7048 = _T_5637_17 & _T_7047;
  assign _T_7050 = _T_4094 & _T_7048;
  assign _T_7065 = _T_4109 & _T_7048;
  assign _T_7067 = _T_5936_17_br_mask & _T_4111;
  assign _GEN_60100 = _T_7065 ? _T_7067 : _GEN_46190;
  assign _GEN_60101 = _T_7050 ? 1'h0 : _GEN_60005;
  assign _GEN_60103 = _T_7050 ? _GEN_46190 : _GEN_60100;
  assign _T_7068 = io_brinfo_mask & _T_5936_18_br_mask;
  assign _T_7070 = _T_7068 != 8'h0;
  assign _T_7071 = _T_5637_18 & _T_7070;
  assign _T_7073 = _T_4094 & _T_7071;
  assign _T_7088 = _T_4109 & _T_7071;
  assign _T_7090 = _T_5936_18_br_mask & _T_4111;
  assign _GEN_60104 = _T_7088 ? _T_7090 : _GEN_46191;
  assign _GEN_60105 = _T_7073 ? 1'h0 : _GEN_60006;
  assign _GEN_60107 = _T_7073 ? _GEN_46191 : _GEN_60104;
  assign _T_7091 = io_brinfo_mask & _T_5936_19_br_mask;
  assign _T_7093 = _T_7091 != 8'h0;
  assign _T_7094 = _T_5637_19 & _T_7093;
  assign _T_7096 = _T_4094 & _T_7094;
  assign _T_7111 = _T_4109 & _T_7094;
  assign _T_7113 = _T_5936_19_br_mask & _T_4111;
  assign _GEN_60108 = _T_7111 ? _T_7113 : _GEN_46192;
  assign _GEN_60109 = _T_7096 ? 1'h0 : _GEN_60007;
  assign _GEN_60111 = _T_7096 ? _GEN_46192 : _GEN_60108;
  assign _T_7114 = io_brinfo_mask & _T_5936_20_br_mask;
  assign _T_7116 = _T_7114 != 8'h0;
  assign _T_7117 = _T_5637_20 & _T_7116;
  assign _T_7119 = _T_4094 & _T_7117;
  assign _T_7134 = _T_4109 & _T_7117;
  assign _T_7136 = _T_5936_20_br_mask & _T_4111;
  assign _GEN_60112 = _T_7134 ? _T_7136 : _GEN_46193;
  assign _GEN_60113 = _T_7119 ? 1'h0 : _GEN_60008;
  assign _GEN_60115 = _T_7119 ? _GEN_46193 : _GEN_60112;
  assign _T_7137 = io_brinfo_mask & _T_5936_21_br_mask;
  assign _T_7139 = _T_7137 != 8'h0;
  assign _T_7140 = _T_5637_21 & _T_7139;
  assign _T_7142 = _T_4094 & _T_7140;
  assign _T_7157 = _T_4109 & _T_7140;
  assign _T_7159 = _T_5936_21_br_mask & _T_4111;
  assign _GEN_60116 = _T_7157 ? _T_7159 : _GEN_46194;
  assign _GEN_60117 = _T_7142 ? 1'h0 : _GEN_60009;
  assign _GEN_60119 = _T_7142 ? _GEN_46194 : _GEN_60116;
  assign _T_7160 = io_brinfo_mask & _T_5936_22_br_mask;
  assign _T_7162 = _T_7160 != 8'h0;
  assign _T_7163 = _T_5637_22 & _T_7162;
  assign _T_7165 = _T_4094 & _T_7163;
  assign _T_7180 = _T_4109 & _T_7163;
  assign _T_7182 = _T_5936_22_br_mask & _T_4111;
  assign _GEN_60120 = _T_7180 ? _T_7182 : _GEN_46195;
  assign _GEN_60121 = _T_7165 ? 1'h0 : _GEN_60010;
  assign _GEN_60123 = _T_7165 ? _GEN_46195 : _GEN_60120;
  assign _T_7183 = io_brinfo_mask & _T_5936_23_br_mask;
  assign _T_7185 = _T_7183 != 8'h0;
  assign _T_7186 = _T_5637_23 & _T_7185;
  assign _T_7188 = _T_4094 & _T_7186;
  assign _T_7203 = _T_4109 & _T_7186;
  assign _T_7205 = _T_5936_23_br_mask & _T_4111;
  assign _GEN_60124 = _T_7203 ? _T_7205 : _GEN_46196;
  assign _GEN_60125 = _T_7188 ? 1'h0 : _GEN_60011;
  assign _GEN_60127 = _T_7188 ? _GEN_46196 : _GEN_60124;
  assign _T_7206 = io_brinfo_mask & _T_5936_24_br_mask;
  assign _T_7208 = _T_7206 != 8'h0;
  assign _T_7209 = _T_5637_24 & _T_7208;
  assign _T_7211 = _T_4094 & _T_7209;
  assign _T_7226 = _T_4109 & _T_7209;
  assign _T_7228 = _T_5936_24_br_mask & _T_4111;
  assign _GEN_60128 = _T_7226 ? _T_7228 : _GEN_46197;
  assign _GEN_60129 = _T_7211 ? 1'h0 : _GEN_60012;
  assign _GEN_60131 = _T_7211 ? _GEN_46197 : _GEN_60128;
  assign _T_7229 = io_brinfo_mask & _T_5936_25_br_mask;
  assign _T_7231 = _T_7229 != 8'h0;
  assign _T_7232 = _T_5637_25 & _T_7231;
  assign _T_7234 = _T_4094 & _T_7232;
  assign _T_7249 = _T_4109 & _T_7232;
  assign _T_7251 = _T_5936_25_br_mask & _T_4111;
  assign _GEN_60132 = _T_7249 ? _T_7251 : _GEN_46198;
  assign _GEN_60133 = _T_7234 ? 1'h0 : _GEN_60013;
  assign _GEN_60135 = _T_7234 ? _GEN_46198 : _GEN_60132;
  assign _T_7252 = io_brinfo_mask & _T_5936_26_br_mask;
  assign _T_7254 = _T_7252 != 8'h0;
  assign _T_7255 = _T_5637_26 & _T_7254;
  assign _T_7257 = _T_4094 & _T_7255;
  assign _T_7272 = _T_4109 & _T_7255;
  assign _T_7274 = _T_5936_26_br_mask & _T_4111;
  assign _GEN_60136 = _T_7272 ? _T_7274 : _GEN_46199;
  assign _GEN_60137 = _T_7257 ? 1'h0 : _GEN_60014;
  assign _GEN_60139 = _T_7257 ? _GEN_46199 : _GEN_60136;
  assign _T_7275 = io_brinfo_mask & _T_5936_27_br_mask;
  assign _T_7277 = _T_7275 != 8'h0;
  assign _T_7278 = _T_5637_27 & _T_7277;
  assign _T_7280 = _T_4094 & _T_7278;
  assign _T_7295 = _T_4109 & _T_7278;
  assign _T_7297 = _T_5936_27_br_mask & _T_4111;
  assign _GEN_60140 = _T_7295 ? _T_7297 : _GEN_46200;
  assign _GEN_60141 = _T_7280 ? 1'h0 : _GEN_60015;
  assign _GEN_60143 = _T_7280 ? _GEN_46200 : _GEN_60140;
  assign _T_7298 = io_brinfo_mask & _T_5936_28_br_mask;
  assign _T_7300 = _T_7298 != 8'h0;
  assign _T_7301 = _T_5637_28 & _T_7300;
  assign _T_7303 = _T_4094 & _T_7301;
  assign _T_7318 = _T_4109 & _T_7301;
  assign _T_7320 = _T_5936_28_br_mask & _T_4111;
  assign _GEN_60144 = _T_7318 ? _T_7320 : _GEN_46201;
  assign _GEN_60145 = _T_7303 ? 1'h0 : _GEN_60016;
  assign _GEN_60147 = _T_7303 ? _GEN_46201 : _GEN_60144;
  assign _T_7321 = io_brinfo_mask & _T_5936_29_br_mask;
  assign _T_7323 = _T_7321 != 8'h0;
  assign _T_7324 = _T_5637_29 & _T_7323;
  assign _T_7326 = _T_4094 & _T_7324;
  assign _T_7341 = _T_4109 & _T_7324;
  assign _T_7343 = _T_5936_29_br_mask & _T_4111;
  assign _GEN_60148 = _T_7341 ? _T_7343 : _GEN_46202;
  assign _GEN_60149 = _T_7326 ? 1'h0 : _GEN_60017;
  assign _GEN_60151 = _T_7326 ? _GEN_46202 : _GEN_60148;
  assign _T_7344 = io_brinfo_mask & _T_5936_30_br_mask;
  assign _T_7346 = _T_7344 != 8'h0;
  assign _T_7347 = _T_5637_30 & _T_7346;
  assign _T_7349 = _T_4094 & _T_7347;
  assign _T_7364 = _T_4109 & _T_7347;
  assign _T_7366 = _T_5936_30_br_mask & _T_4111;
  assign _GEN_60152 = _T_7364 ? _T_7366 : _GEN_46203;
  assign _GEN_60153 = _T_7349 ? 1'h0 : _GEN_60018;
  assign _GEN_60155 = _T_7349 ? _GEN_46203 : _GEN_60152;
  assign _T_7367 = io_brinfo_mask & _T_5936_31_br_mask;
  assign _T_7369 = _T_7367 != 8'h0;
  assign _T_7370 = _T_5637_31 & _T_7369;
  assign _T_7372 = _T_4094 & _T_7370;
  assign _T_7387 = _T_4109 & _T_7370;
  assign _T_7389 = _T_5936_31_br_mask & _T_4111;
  assign _GEN_60156 = _T_7387 ? _T_7389 : _GEN_46204;
  assign _GEN_60157 = _T_7372 ? 1'h0 : _GEN_60019;
  assign _GEN_60159 = _T_7372 ? _GEN_46204 : _GEN_60156;
  assign _T_7390 = io_brinfo_mask & _T_5936_32_br_mask;
  assign _T_7392 = _T_7390 != 8'h0;
  assign _T_7393 = _T_5637_32 & _T_7392;
  assign _T_7395 = _T_4094 & _T_7393;
  assign _T_7410 = _T_4109 & _T_7393;
  assign _T_7412 = _T_5936_32_br_mask & _T_4111;
  assign _GEN_60160 = _T_7410 ? _T_7412 : _GEN_46205;
  assign _GEN_60161 = _T_7395 ? 1'h0 : _GEN_60020;
  assign _GEN_60163 = _T_7395 ? _GEN_46205 : _GEN_60160;
  assign _T_7413 = io_brinfo_mask & _T_5936_33_br_mask;
  assign _T_7415 = _T_7413 != 8'h0;
  assign _T_7416 = _T_5637_33 & _T_7415;
  assign _T_7418 = _T_4094 & _T_7416;
  assign _T_7433 = _T_4109 & _T_7416;
  assign _T_7435 = _T_5936_33_br_mask & _T_4111;
  assign _GEN_60164 = _T_7433 ? _T_7435 : _GEN_46206;
  assign _GEN_60165 = _T_7418 ? 1'h0 : _GEN_60021;
  assign _GEN_60167 = _T_7418 ? _GEN_46206 : _GEN_60164;
  assign _T_7436 = io_brinfo_mask & _T_5936_34_br_mask;
  assign _T_7438 = _T_7436 != 8'h0;
  assign _T_7439 = _T_5637_34 & _T_7438;
  assign _T_7441 = _T_4094 & _T_7439;
  assign _T_7456 = _T_4109 & _T_7439;
  assign _T_7458 = _T_5936_34_br_mask & _T_4111;
  assign _GEN_60168 = _T_7456 ? _T_7458 : _GEN_46207;
  assign _GEN_60169 = _T_7441 ? 1'h0 : _GEN_60022;
  assign _GEN_60171 = _T_7441 ? _GEN_46207 : _GEN_60168;
  assign _T_7459 = io_brinfo_mask & _T_5936_35_br_mask;
  assign _T_7461 = _T_7459 != 8'h0;
  assign _T_7462 = _T_5637_35 & _T_7461;
  assign _T_7464 = _T_4094 & _T_7462;
  assign _T_7479 = _T_4109 & _T_7462;
  assign _T_7481 = _T_5936_35_br_mask & _T_4111;
  assign _GEN_60172 = _T_7479 ? _T_7481 : _GEN_46208;
  assign _GEN_60173 = _T_7464 ? 1'h0 : _GEN_60023;
  assign _GEN_60175 = _T_7464 ? _GEN_46208 : _GEN_60172;
  assign _T_7482 = io_brinfo_mask & _T_5936_36_br_mask;
  assign _T_7484 = _T_7482 != 8'h0;
  assign _T_7485 = _T_5637_36 & _T_7484;
  assign _T_7487 = _T_4094 & _T_7485;
  assign _T_7502 = _T_4109 & _T_7485;
  assign _T_7504 = _T_5936_36_br_mask & _T_4111;
  assign _GEN_60176 = _T_7502 ? _T_7504 : _GEN_46209;
  assign _GEN_60177 = _T_7487 ? 1'h0 : _GEN_60024;
  assign _GEN_60179 = _T_7487 ? _GEN_46209 : _GEN_60176;
  assign _T_7505 = io_brinfo_mask & _T_5936_37_br_mask;
  assign _T_7507 = _T_7505 != 8'h0;
  assign _T_7508 = _T_5637_37 & _T_7507;
  assign _T_7510 = _T_4094 & _T_7508;
  assign _T_7525 = _T_4109 & _T_7508;
  assign _T_7527 = _T_5936_37_br_mask & _T_4111;
  assign _GEN_60180 = _T_7525 ? _T_7527 : _GEN_46210;
  assign _GEN_60181 = _T_7510 ? 1'h0 : _GEN_60025;
  assign _GEN_60183 = _T_7510 ? _GEN_46210 : _GEN_60180;
  assign _T_7528 = io_brinfo_mask & _T_5936_38_br_mask;
  assign _T_7530 = _T_7528 != 8'h0;
  assign _T_7531 = _T_5637_38 & _T_7530;
  assign _T_7533 = _T_4094 & _T_7531;
  assign _T_7548 = _T_4109 & _T_7531;
  assign _T_7550 = _T_5936_38_br_mask & _T_4111;
  assign _GEN_60184 = _T_7548 ? _T_7550 : _GEN_46211;
  assign _GEN_60185 = _T_7533 ? 1'h0 : _GEN_60026;
  assign _GEN_60187 = _T_7533 ? _GEN_46211 : _GEN_60184;
  assign _T_7551 = io_brinfo_mask & _T_5936_39_br_mask;
  assign _T_7553 = _T_7551 != 8'h0;
  assign _T_7554 = _T_5637_39 & _T_7553;
  assign _T_7556 = _T_4094 & _T_7554;
  assign _T_7571 = _T_4109 & _T_7554;
  assign _T_7573 = _T_5936_39_br_mask & _T_4111;
  assign _GEN_60188 = _T_7571 ? _T_7573 : _GEN_46212;
  assign _GEN_60189 = _T_7556 ? 1'h0 : _GEN_60027;
  assign _GEN_60191 = _T_7556 ? _GEN_46212 : _GEN_60188;
  assign _GEN_60192 = 6'h0 == rob_head ? 1'h0 : _GEN_60033;
  assign _GEN_60193 = 6'h1 == rob_head ? 1'h0 : _GEN_60037;
  assign _GEN_60194 = 6'h2 == rob_head ? 1'h0 : _GEN_60041;
  assign _GEN_60195 = 6'h3 == rob_head ? 1'h0 : _GEN_60045;
  assign _GEN_60196 = 6'h4 == rob_head ? 1'h0 : _GEN_60049;
  assign _GEN_60197 = 6'h5 == rob_head ? 1'h0 : _GEN_60053;
  assign _GEN_60198 = 6'h6 == rob_head ? 1'h0 : _GEN_60057;
  assign _GEN_60199 = 6'h7 == rob_head ? 1'h0 : _GEN_60061;
  assign _GEN_60200 = 6'h8 == rob_head ? 1'h0 : _GEN_60065;
  assign _GEN_60201 = 6'h9 == rob_head ? 1'h0 : _GEN_60069;
  assign _GEN_60202 = 6'ha == rob_head ? 1'h0 : _GEN_60073;
  assign _GEN_60203 = 6'hb == rob_head ? 1'h0 : _GEN_60077;
  assign _GEN_60204 = 6'hc == rob_head ? 1'h0 : _GEN_60081;
  assign _GEN_60205 = 6'hd == rob_head ? 1'h0 : _GEN_60085;
  assign _GEN_60206 = 6'he == rob_head ? 1'h0 : _GEN_60089;
  assign _GEN_60207 = 6'hf == rob_head ? 1'h0 : _GEN_60093;
  assign _GEN_60208 = 6'h10 == rob_head ? 1'h0 : _GEN_60097;
  assign _GEN_60209 = 6'h11 == rob_head ? 1'h0 : _GEN_60101;
  assign _GEN_60210 = 6'h12 == rob_head ? 1'h0 : _GEN_60105;
  assign _GEN_60211 = 6'h13 == rob_head ? 1'h0 : _GEN_60109;
  assign _GEN_60212 = 6'h14 == rob_head ? 1'h0 : _GEN_60113;
  assign _GEN_60213 = 6'h15 == rob_head ? 1'h0 : _GEN_60117;
  assign _GEN_60214 = 6'h16 == rob_head ? 1'h0 : _GEN_60121;
  assign _GEN_60215 = 6'h17 == rob_head ? 1'h0 : _GEN_60125;
  assign _GEN_60216 = 6'h18 == rob_head ? 1'h0 : _GEN_60129;
  assign _GEN_60217 = 6'h19 == rob_head ? 1'h0 : _GEN_60133;
  assign _GEN_60218 = 6'h1a == rob_head ? 1'h0 : _GEN_60137;
  assign _GEN_60219 = 6'h1b == rob_head ? 1'h0 : _GEN_60141;
  assign _GEN_60220 = 6'h1c == rob_head ? 1'h0 : _GEN_60145;
  assign _GEN_60221 = 6'h1d == rob_head ? 1'h0 : _GEN_60149;
  assign _GEN_60222 = 6'h1e == rob_head ? 1'h0 : _GEN_60153;
  assign _GEN_60223 = 6'h1f == rob_head ? 1'h0 : _GEN_60157;
  assign _GEN_60224 = 6'h20 == rob_head ? 1'h0 : _GEN_60161;
  assign _GEN_60225 = 6'h21 == rob_head ? 1'h0 : _GEN_60165;
  assign _GEN_60226 = 6'h22 == rob_head ? 1'h0 : _GEN_60169;
  assign _GEN_60227 = 6'h23 == rob_head ? 1'h0 : _GEN_60173;
  assign _GEN_60228 = 6'h24 == rob_head ? 1'h0 : _GEN_60177;
  assign _GEN_60229 = 6'h25 == rob_head ? 1'h0 : _GEN_60181;
  assign _GEN_60230 = 6'h26 == rob_head ? 1'h0 : _GEN_60185;
  assign _GEN_60231 = 6'h27 == rob_head ? 1'h0 : _GEN_60189;
  assign _GEN_60232 = will_commit_1 ? _GEN_60192 : _GEN_60033;
  assign _GEN_60233 = will_commit_1 ? _GEN_60193 : _GEN_60037;
  assign _GEN_60234 = will_commit_1 ? _GEN_60194 : _GEN_60041;
  assign _GEN_60235 = will_commit_1 ? _GEN_60195 : _GEN_60045;
  assign _GEN_60236 = will_commit_1 ? _GEN_60196 : _GEN_60049;
  assign _GEN_60237 = will_commit_1 ? _GEN_60197 : _GEN_60053;
  assign _GEN_60238 = will_commit_1 ? _GEN_60198 : _GEN_60057;
  assign _GEN_60239 = will_commit_1 ? _GEN_60199 : _GEN_60061;
  assign _GEN_60240 = will_commit_1 ? _GEN_60200 : _GEN_60065;
  assign _GEN_60241 = will_commit_1 ? _GEN_60201 : _GEN_60069;
  assign _GEN_60242 = will_commit_1 ? _GEN_60202 : _GEN_60073;
  assign _GEN_60243 = will_commit_1 ? _GEN_60203 : _GEN_60077;
  assign _GEN_60244 = will_commit_1 ? _GEN_60204 : _GEN_60081;
  assign _GEN_60245 = will_commit_1 ? _GEN_60205 : _GEN_60085;
  assign _GEN_60246 = will_commit_1 ? _GEN_60206 : _GEN_60089;
  assign _GEN_60247 = will_commit_1 ? _GEN_60207 : _GEN_60093;
  assign _GEN_60248 = will_commit_1 ? _GEN_60208 : _GEN_60097;
  assign _GEN_60249 = will_commit_1 ? _GEN_60209 : _GEN_60101;
  assign _GEN_60250 = will_commit_1 ? _GEN_60210 : _GEN_60105;
  assign _GEN_60251 = will_commit_1 ? _GEN_60211 : _GEN_60109;
  assign _GEN_60252 = will_commit_1 ? _GEN_60212 : _GEN_60113;
  assign _GEN_60253 = will_commit_1 ? _GEN_60213 : _GEN_60117;
  assign _GEN_60254 = will_commit_1 ? _GEN_60214 : _GEN_60121;
  assign _GEN_60255 = will_commit_1 ? _GEN_60215 : _GEN_60125;
  assign _GEN_60256 = will_commit_1 ? _GEN_60216 : _GEN_60129;
  assign _GEN_60257 = will_commit_1 ? _GEN_60217 : _GEN_60133;
  assign _GEN_60258 = will_commit_1 ? _GEN_60218 : _GEN_60137;
  assign _GEN_60259 = will_commit_1 ? _GEN_60219 : _GEN_60141;
  assign _GEN_60260 = will_commit_1 ? _GEN_60220 : _GEN_60145;
  assign _GEN_60261 = will_commit_1 ? _GEN_60221 : _GEN_60149;
  assign _GEN_60262 = will_commit_1 ? _GEN_60222 : _GEN_60153;
  assign _GEN_60263 = will_commit_1 ? _GEN_60223 : _GEN_60157;
  assign _GEN_60264 = will_commit_1 ? _GEN_60224 : _GEN_60161;
  assign _GEN_60265 = will_commit_1 ? _GEN_60225 : _GEN_60165;
  assign _GEN_60266 = will_commit_1 ? _GEN_60226 : _GEN_60169;
  assign _GEN_60267 = will_commit_1 ? _GEN_60227 : _GEN_60173;
  assign _GEN_60268 = will_commit_1 ? _GEN_60228 : _GEN_60177;
  assign _GEN_60269 = will_commit_1 ? _GEN_60229 : _GEN_60181;
  assign _GEN_60270 = will_commit_1 ? _GEN_60230 : _GEN_60185;
  assign _GEN_60271 = will_commit_1 ? _GEN_60231 : _GEN_60189;
  assign _GEN_60339 = 6'h1 == rob_head ? _T_5936_1_is_store : _T_5936_0_is_store;
  assign _GEN_60341 = 6'h1 == rob_head ? _T_5936_1_is_load : _T_5936_0_is_load;
  assign _GEN_60429 = 6'h2 == rob_head ? _T_5936_2_is_store : _GEN_60339;
  assign _GEN_60431 = 6'h2 == rob_head ? _T_5936_2_is_load : _GEN_60341;
  assign _GEN_60519 = 6'h3 == rob_head ? _T_5936_3_is_store : _GEN_60429;
  assign _GEN_60521 = 6'h3 == rob_head ? _T_5936_3_is_load : _GEN_60431;
  assign _GEN_60609 = 6'h4 == rob_head ? _T_5936_4_is_store : _GEN_60519;
  assign _GEN_60611 = 6'h4 == rob_head ? _T_5936_4_is_load : _GEN_60521;
  assign _GEN_60699 = 6'h5 == rob_head ? _T_5936_5_is_store : _GEN_60609;
  assign _GEN_60701 = 6'h5 == rob_head ? _T_5936_5_is_load : _GEN_60611;
  assign _GEN_60789 = 6'h6 == rob_head ? _T_5936_6_is_store : _GEN_60699;
  assign _GEN_60791 = 6'h6 == rob_head ? _T_5936_6_is_load : _GEN_60701;
  assign _GEN_60879 = 6'h7 == rob_head ? _T_5936_7_is_store : _GEN_60789;
  assign _GEN_60881 = 6'h7 == rob_head ? _T_5936_7_is_load : _GEN_60791;
  assign _GEN_60969 = 6'h8 == rob_head ? _T_5936_8_is_store : _GEN_60879;
  assign _GEN_60971 = 6'h8 == rob_head ? _T_5936_8_is_load : _GEN_60881;
  assign _GEN_61059 = 6'h9 == rob_head ? _T_5936_9_is_store : _GEN_60969;
  assign _GEN_61061 = 6'h9 == rob_head ? _T_5936_9_is_load : _GEN_60971;
  assign _GEN_61149 = 6'ha == rob_head ? _T_5936_10_is_store : _GEN_61059;
  assign _GEN_61151 = 6'ha == rob_head ? _T_5936_10_is_load : _GEN_61061;
  assign _GEN_61239 = 6'hb == rob_head ? _T_5936_11_is_store : _GEN_61149;
  assign _GEN_61241 = 6'hb == rob_head ? _T_5936_11_is_load : _GEN_61151;
  assign _GEN_61329 = 6'hc == rob_head ? _T_5936_12_is_store : _GEN_61239;
  assign _GEN_61331 = 6'hc == rob_head ? _T_5936_12_is_load : _GEN_61241;
  assign _GEN_61419 = 6'hd == rob_head ? _T_5936_13_is_store : _GEN_61329;
  assign _GEN_61421 = 6'hd == rob_head ? _T_5936_13_is_load : _GEN_61331;
  assign _GEN_61509 = 6'he == rob_head ? _T_5936_14_is_store : _GEN_61419;
  assign _GEN_61511 = 6'he == rob_head ? _T_5936_14_is_load : _GEN_61421;
  assign _GEN_61599 = 6'hf == rob_head ? _T_5936_15_is_store : _GEN_61509;
  assign _GEN_61601 = 6'hf == rob_head ? _T_5936_15_is_load : _GEN_61511;
  assign _GEN_61689 = 6'h10 == rob_head ? _T_5936_16_is_store : _GEN_61599;
  assign _GEN_61691 = 6'h10 == rob_head ? _T_5936_16_is_load : _GEN_61601;
  assign _GEN_61779 = 6'h11 == rob_head ? _T_5936_17_is_store : _GEN_61689;
  assign _GEN_61781 = 6'h11 == rob_head ? _T_5936_17_is_load : _GEN_61691;
  assign _GEN_61869 = 6'h12 == rob_head ? _T_5936_18_is_store : _GEN_61779;
  assign _GEN_61871 = 6'h12 == rob_head ? _T_5936_18_is_load : _GEN_61781;
  assign _GEN_61959 = 6'h13 == rob_head ? _T_5936_19_is_store : _GEN_61869;
  assign _GEN_61961 = 6'h13 == rob_head ? _T_5936_19_is_load : _GEN_61871;
  assign _GEN_62049 = 6'h14 == rob_head ? _T_5936_20_is_store : _GEN_61959;
  assign _GEN_62051 = 6'h14 == rob_head ? _T_5936_20_is_load : _GEN_61961;
  assign _GEN_62139 = 6'h15 == rob_head ? _T_5936_21_is_store : _GEN_62049;
  assign _GEN_62141 = 6'h15 == rob_head ? _T_5936_21_is_load : _GEN_62051;
  assign _GEN_62229 = 6'h16 == rob_head ? _T_5936_22_is_store : _GEN_62139;
  assign _GEN_62231 = 6'h16 == rob_head ? _T_5936_22_is_load : _GEN_62141;
  assign _GEN_62319 = 6'h17 == rob_head ? _T_5936_23_is_store : _GEN_62229;
  assign _GEN_62321 = 6'h17 == rob_head ? _T_5936_23_is_load : _GEN_62231;
  assign _GEN_62409 = 6'h18 == rob_head ? _T_5936_24_is_store : _GEN_62319;
  assign _GEN_62411 = 6'h18 == rob_head ? _T_5936_24_is_load : _GEN_62321;
  assign _GEN_62499 = 6'h19 == rob_head ? _T_5936_25_is_store : _GEN_62409;
  assign _GEN_62501 = 6'h19 == rob_head ? _T_5936_25_is_load : _GEN_62411;
  assign _GEN_62589 = 6'h1a == rob_head ? _T_5936_26_is_store : _GEN_62499;
  assign _GEN_62591 = 6'h1a == rob_head ? _T_5936_26_is_load : _GEN_62501;
  assign _GEN_62679 = 6'h1b == rob_head ? _T_5936_27_is_store : _GEN_62589;
  assign _GEN_62681 = 6'h1b == rob_head ? _T_5936_27_is_load : _GEN_62591;
  assign _GEN_62769 = 6'h1c == rob_head ? _T_5936_28_is_store : _GEN_62679;
  assign _GEN_62771 = 6'h1c == rob_head ? _T_5936_28_is_load : _GEN_62681;
  assign _GEN_62859 = 6'h1d == rob_head ? _T_5936_29_is_store : _GEN_62769;
  assign _GEN_62861 = 6'h1d == rob_head ? _T_5936_29_is_load : _GEN_62771;
  assign _GEN_62949 = 6'h1e == rob_head ? _T_5936_30_is_store : _GEN_62859;
  assign _GEN_62951 = 6'h1e == rob_head ? _T_5936_30_is_load : _GEN_62861;
  assign _GEN_63039 = 6'h1f == rob_head ? _T_5936_31_is_store : _GEN_62949;
  assign _GEN_63041 = 6'h1f == rob_head ? _T_5936_31_is_load : _GEN_62951;
  assign _GEN_63129 = 6'h20 == rob_head ? _T_5936_32_is_store : _GEN_63039;
  assign _GEN_63131 = 6'h20 == rob_head ? _T_5936_32_is_load : _GEN_63041;
  assign _GEN_63219 = 6'h21 == rob_head ? _T_5936_33_is_store : _GEN_63129;
  assign _GEN_63221 = 6'h21 == rob_head ? _T_5936_33_is_load : _GEN_63131;
  assign _GEN_63309 = 6'h22 == rob_head ? _T_5936_34_is_store : _GEN_63219;
  assign _GEN_63311 = 6'h22 == rob_head ? _T_5936_34_is_load : _GEN_63221;
  assign _GEN_63399 = 6'h23 == rob_head ? _T_5936_35_is_store : _GEN_63309;
  assign _GEN_63401 = 6'h23 == rob_head ? _T_5936_35_is_load : _GEN_63311;
  assign _GEN_63489 = 6'h24 == rob_head ? _T_5936_36_is_store : _GEN_63399;
  assign _GEN_63491 = 6'h24 == rob_head ? _T_5936_36_is_load : _GEN_63401;
  assign _GEN_63579 = 6'h25 == rob_head ? _T_5936_37_is_store : _GEN_63489;
  assign _GEN_63581 = 6'h25 == rob_head ? _T_5936_37_is_load : _GEN_63491;
  assign _GEN_63669 = 6'h26 == rob_head ? _T_5936_38_is_store : _GEN_63579;
  assign _GEN_63671 = 6'h26 == rob_head ? _T_5936_38_is_load : _GEN_63581;
  assign _GEN_63759 = 6'h27 == rob_head ? _T_5936_39_is_store : _GEN_63669;
  assign _GEN_63761 = 6'h27 == rob_head ? _T_5936_39_is_load : _GEN_63671;
  assign _GEN_63782 = 6'h1 == _T_2899 ? _T_5637_1 : _T_5637_0;
  assign _GEN_63783 = 6'h2 == _T_2899 ? _T_5637_2 : _GEN_63782;
  assign _GEN_63784 = 6'h3 == _T_2899 ? _T_5637_3 : _GEN_63783;
  assign _GEN_63785 = 6'h4 == _T_2899 ? _T_5637_4 : _GEN_63784;
  assign _GEN_63786 = 6'h5 == _T_2899 ? _T_5637_5 : _GEN_63785;
  assign _GEN_63787 = 6'h6 == _T_2899 ? _T_5637_6 : _GEN_63786;
  assign _GEN_63788 = 6'h7 == _T_2899 ? _T_5637_7 : _GEN_63787;
  assign _GEN_63789 = 6'h8 == _T_2899 ? _T_5637_8 : _GEN_63788;
  assign _GEN_63790 = 6'h9 == _T_2899 ? _T_5637_9 : _GEN_63789;
  assign _GEN_63791 = 6'ha == _T_2899 ? _T_5637_10 : _GEN_63790;
  assign _GEN_63792 = 6'hb == _T_2899 ? _T_5637_11 : _GEN_63791;
  assign _GEN_63793 = 6'hc == _T_2899 ? _T_5637_12 : _GEN_63792;
  assign _GEN_63794 = 6'hd == _T_2899 ? _T_5637_13 : _GEN_63793;
  assign _GEN_63795 = 6'he == _T_2899 ? _T_5637_14 : _GEN_63794;
  assign _GEN_63796 = 6'hf == _T_2899 ? _T_5637_15 : _GEN_63795;
  assign _GEN_63797 = 6'h10 == _T_2899 ? _T_5637_16 : _GEN_63796;
  assign _GEN_63798 = 6'h11 == _T_2899 ? _T_5637_17 : _GEN_63797;
  assign _GEN_63799 = 6'h12 == _T_2899 ? _T_5637_18 : _GEN_63798;
  assign _GEN_63800 = 6'h13 == _T_2899 ? _T_5637_19 : _GEN_63799;
  assign _GEN_63801 = 6'h14 == _T_2899 ? _T_5637_20 : _GEN_63800;
  assign _GEN_63802 = 6'h15 == _T_2899 ? _T_5637_21 : _GEN_63801;
  assign _GEN_63803 = 6'h16 == _T_2899 ? _T_5637_22 : _GEN_63802;
  assign _GEN_63804 = 6'h17 == _T_2899 ? _T_5637_23 : _GEN_63803;
  assign _GEN_63805 = 6'h18 == _T_2899 ? _T_5637_24 : _GEN_63804;
  assign _GEN_63806 = 6'h19 == _T_2899 ? _T_5637_25 : _GEN_63805;
  assign _GEN_63807 = 6'h1a == _T_2899 ? _T_5637_26 : _GEN_63806;
  assign _GEN_63808 = 6'h1b == _T_2899 ? _T_5637_27 : _GEN_63807;
  assign _GEN_63809 = 6'h1c == _T_2899 ? _T_5637_28 : _GEN_63808;
  assign _GEN_63810 = 6'h1d == _T_2899 ? _T_5637_29 : _GEN_63809;
  assign _GEN_63811 = 6'h1e == _T_2899 ? _T_5637_30 : _GEN_63810;
  assign _GEN_63812 = 6'h1f == _T_2899 ? _T_5637_31 : _GEN_63811;
  assign _GEN_63813 = 6'h20 == _T_2899 ? _T_5637_32 : _GEN_63812;
  assign _GEN_63814 = 6'h21 == _T_2899 ? _T_5637_33 : _GEN_63813;
  assign _GEN_63815 = 6'h22 == _T_2899 ? _T_5637_34 : _GEN_63814;
  assign _GEN_63816 = 6'h23 == _T_2899 ? _T_5637_35 : _GEN_63815;
  assign _GEN_63817 = 6'h24 == _T_2899 ? _T_5637_36 : _GEN_63816;
  assign _GEN_63818 = 6'h25 == _T_2899 ? _T_5637_37 : _GEN_63817;
  assign _GEN_63819 = 6'h26 == _T_2899 ? _T_5637_38 : _GEN_63818;
  assign _GEN_63820 = 6'h27 == _T_2899 ? _T_5637_39 : _GEN_63819;
  assign _GEN_63821 = 6'h1 == _T_5054 ? _T_5637_1 : _T_5637_0;
  assign _GEN_63822 = 6'h2 == _T_5054 ? _T_5637_2 : _GEN_63821;
  assign _GEN_63823 = 6'h3 == _T_5054 ? _T_5637_3 : _GEN_63822;
  assign _GEN_63824 = 6'h4 == _T_5054 ? _T_5637_4 : _GEN_63823;
  assign _GEN_63825 = 6'h5 == _T_5054 ? _T_5637_5 : _GEN_63824;
  assign _GEN_63826 = 6'h6 == _T_5054 ? _T_5637_6 : _GEN_63825;
  assign _GEN_63827 = 6'h7 == _T_5054 ? _T_5637_7 : _GEN_63826;
  assign _GEN_63828 = 6'h8 == _T_5054 ? _T_5637_8 : _GEN_63827;
  assign _GEN_63829 = 6'h9 == _T_5054 ? _T_5637_9 : _GEN_63828;
  assign _GEN_63830 = 6'ha == _T_5054 ? _T_5637_10 : _GEN_63829;
  assign _GEN_63831 = 6'hb == _T_5054 ? _T_5637_11 : _GEN_63830;
  assign _GEN_63832 = 6'hc == _T_5054 ? _T_5637_12 : _GEN_63831;
  assign _GEN_63833 = 6'hd == _T_5054 ? _T_5637_13 : _GEN_63832;
  assign _GEN_63834 = 6'he == _T_5054 ? _T_5637_14 : _GEN_63833;
  assign _GEN_63835 = 6'hf == _T_5054 ? _T_5637_15 : _GEN_63834;
  assign _GEN_63836 = 6'h10 == _T_5054 ? _T_5637_16 : _GEN_63835;
  assign _GEN_63837 = 6'h11 == _T_5054 ? _T_5637_17 : _GEN_63836;
  assign _GEN_63838 = 6'h12 == _T_5054 ? _T_5637_18 : _GEN_63837;
  assign _GEN_63839 = 6'h13 == _T_5054 ? _T_5637_19 : _GEN_63838;
  assign _GEN_63840 = 6'h14 == _T_5054 ? _T_5637_20 : _GEN_63839;
  assign _GEN_63841 = 6'h15 == _T_5054 ? _T_5637_21 : _GEN_63840;
  assign _GEN_63842 = 6'h16 == _T_5054 ? _T_5637_22 : _GEN_63841;
  assign _GEN_63843 = 6'h17 == _T_5054 ? _T_5637_23 : _GEN_63842;
  assign _GEN_63844 = 6'h18 == _T_5054 ? _T_5637_24 : _GEN_63843;
  assign _GEN_63845 = 6'h19 == _T_5054 ? _T_5637_25 : _GEN_63844;
  assign _GEN_63846 = 6'h1a == _T_5054 ? _T_5637_26 : _GEN_63845;
  assign _GEN_63847 = 6'h1b == _T_5054 ? _T_5637_27 : _GEN_63846;
  assign _GEN_63848 = 6'h1c == _T_5054 ? _T_5637_28 : _GEN_63847;
  assign _GEN_63849 = 6'h1d == _T_5054 ? _T_5637_29 : _GEN_63848;
  assign _GEN_63850 = 6'h1e == _T_5054 ? _T_5637_30 : _GEN_63849;
  assign _GEN_63851 = 6'h1f == _T_5054 ? _T_5637_31 : _GEN_63850;
  assign _GEN_63852 = 6'h20 == _T_5054 ? _T_5637_32 : _GEN_63851;
  assign _GEN_63853 = 6'h21 == _T_5054 ? _T_5637_33 : _GEN_63852;
  assign _GEN_63854 = 6'h22 == _T_5054 ? _T_5637_34 : _GEN_63853;
  assign _GEN_63855 = 6'h23 == _T_5054 ? _T_5637_35 : _GEN_63854;
  assign _GEN_63856 = 6'h24 == _T_5054 ? _T_5637_36 : _GEN_63855;
  assign _GEN_63857 = 6'h25 == _T_5054 ? _T_5637_37 : _GEN_63856;
  assign _GEN_63858 = 6'h26 == _T_5054 ? _T_5637_38 : _GEN_63857;
  assign _GEN_63859 = 6'h27 == _T_5054 ? _T_5637_39 : _GEN_63858;
  assign _GEN_64100 = 6'h1 == _T_3818 ? _T_5637_1 : _T_5637_0;
  assign _GEN_64101 = 6'h2 == _T_3818 ? _T_5637_2 : _GEN_64100;
  assign _GEN_64102 = 6'h3 == _T_3818 ? _T_5637_3 : _GEN_64101;
  assign _GEN_64103 = 6'h4 == _T_3818 ? _T_5637_4 : _GEN_64102;
  assign _GEN_64104 = 6'h5 == _T_3818 ? _T_5637_5 : _GEN_64103;
  assign _GEN_64105 = 6'h6 == _T_3818 ? _T_5637_6 : _GEN_64104;
  assign _GEN_64106 = 6'h7 == _T_3818 ? _T_5637_7 : _GEN_64105;
  assign _GEN_64107 = 6'h8 == _T_3818 ? _T_5637_8 : _GEN_64106;
  assign _GEN_64108 = 6'h9 == _T_3818 ? _T_5637_9 : _GEN_64107;
  assign _GEN_64109 = 6'ha == _T_3818 ? _T_5637_10 : _GEN_64108;
  assign _GEN_64110 = 6'hb == _T_3818 ? _T_5637_11 : _GEN_64109;
  assign _GEN_64111 = 6'hc == _T_3818 ? _T_5637_12 : _GEN_64110;
  assign _GEN_64112 = 6'hd == _T_3818 ? _T_5637_13 : _GEN_64111;
  assign _GEN_64113 = 6'he == _T_3818 ? _T_5637_14 : _GEN_64112;
  assign _GEN_64114 = 6'hf == _T_3818 ? _T_5637_15 : _GEN_64113;
  assign _GEN_64115 = 6'h10 == _T_3818 ? _T_5637_16 : _GEN_64114;
  assign _GEN_64116 = 6'h11 == _T_3818 ? _T_5637_17 : _GEN_64115;
  assign _GEN_64117 = 6'h12 == _T_3818 ? _T_5637_18 : _GEN_64116;
  assign _GEN_64118 = 6'h13 == _T_3818 ? _T_5637_19 : _GEN_64117;
  assign _GEN_64119 = 6'h14 == _T_3818 ? _T_5637_20 : _GEN_64118;
  assign _GEN_64120 = 6'h15 == _T_3818 ? _T_5637_21 : _GEN_64119;
  assign _GEN_64121 = 6'h16 == _T_3818 ? _T_5637_22 : _GEN_64120;
  assign _GEN_64122 = 6'h17 == _T_3818 ? _T_5637_23 : _GEN_64121;
  assign _GEN_64123 = 6'h18 == _T_3818 ? _T_5637_24 : _GEN_64122;
  assign _GEN_64124 = 6'h19 == _T_3818 ? _T_5637_25 : _GEN_64123;
  assign _GEN_64125 = 6'h1a == _T_3818 ? _T_5637_26 : _GEN_64124;
  assign _GEN_64126 = 6'h1b == _T_3818 ? _T_5637_27 : _GEN_64125;
  assign _GEN_64127 = 6'h1c == _T_3818 ? _T_5637_28 : _GEN_64126;
  assign _GEN_64128 = 6'h1d == _T_3818 ? _T_5637_29 : _GEN_64127;
  assign _GEN_64129 = 6'h1e == _T_3818 ? _T_5637_30 : _GEN_64128;
  assign _GEN_64130 = 6'h1f == _T_3818 ? _T_5637_31 : _GEN_64129;
  assign _GEN_64131 = 6'h20 == _T_3818 ? _T_5637_32 : _GEN_64130;
  assign _GEN_64132 = 6'h21 == _T_3818 ? _T_5637_33 : _GEN_64131;
  assign _GEN_64133 = 6'h22 == _T_3818 ? _T_5637_34 : _GEN_64132;
  assign _GEN_64134 = 6'h23 == _T_3818 ? _T_5637_35 : _GEN_64133;
  assign _GEN_64135 = 6'h24 == _T_3818 ? _T_5637_36 : _GEN_64134;
  assign _GEN_64136 = 6'h25 == _T_3818 ? _T_5637_37 : _GEN_64135;
  assign _GEN_64137 = 6'h26 == _T_3818 ? _T_5637_38 : _GEN_64136;
  assign _GEN_64138 = 6'h27 == _T_3818 ? _T_5637_39 : _GEN_64137;
  assign _T_7677 = _GEN_435 == 1'h0;
  assign _T_7678 = _T_6381 & _T_7677;
  assign _T_7680 = _T_7678 == 1'h0;
  assign _T_7682 = _T_7680 | reset;
  assign _T_7684 = _T_7682 == 1'h0;
  assign _T_7691 = _T_3813[5:0];
  assign _T_7694 = _T_5764__T_7692_data == 1'h0;
  assign _T_7695 = _T_6381 & _T_7694;
  assign _T_7697 = _T_7695 == 1'h0;
  assign _T_7699 = _T_7697 | reset;
  assign _T_7701 = _T_7699 == 1'h0;
  assign _GEN_64191 = 6'h1 == _T_3818 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_64216 = 6'h1 == _T_3818 ? _T_5936_1_ldst_val : _T_5936_0_ldst_val;
  assign _GEN_64281 = 6'h2 == _T_3818 ? _T_5936_2_pdst : _GEN_64191;
  assign _GEN_64306 = 6'h2 == _T_3818 ? _T_5936_2_ldst_val : _GEN_64216;
  assign _GEN_64371 = 6'h3 == _T_3818 ? _T_5936_3_pdst : _GEN_64281;
  assign _GEN_64396 = 6'h3 == _T_3818 ? _T_5936_3_ldst_val : _GEN_64306;
  assign _GEN_64461 = 6'h4 == _T_3818 ? _T_5936_4_pdst : _GEN_64371;
  assign _GEN_64486 = 6'h4 == _T_3818 ? _T_5936_4_ldst_val : _GEN_64396;
  assign _GEN_64551 = 6'h5 == _T_3818 ? _T_5936_5_pdst : _GEN_64461;
  assign _GEN_64576 = 6'h5 == _T_3818 ? _T_5936_5_ldst_val : _GEN_64486;
  assign _GEN_64641 = 6'h6 == _T_3818 ? _T_5936_6_pdst : _GEN_64551;
  assign _GEN_64666 = 6'h6 == _T_3818 ? _T_5936_6_ldst_val : _GEN_64576;
  assign _GEN_64731 = 6'h7 == _T_3818 ? _T_5936_7_pdst : _GEN_64641;
  assign _GEN_64756 = 6'h7 == _T_3818 ? _T_5936_7_ldst_val : _GEN_64666;
  assign _GEN_64821 = 6'h8 == _T_3818 ? _T_5936_8_pdst : _GEN_64731;
  assign _GEN_64846 = 6'h8 == _T_3818 ? _T_5936_8_ldst_val : _GEN_64756;
  assign _GEN_64911 = 6'h9 == _T_3818 ? _T_5936_9_pdst : _GEN_64821;
  assign _GEN_64936 = 6'h9 == _T_3818 ? _T_5936_9_ldst_val : _GEN_64846;
  assign _GEN_65001 = 6'ha == _T_3818 ? _T_5936_10_pdst : _GEN_64911;
  assign _GEN_65026 = 6'ha == _T_3818 ? _T_5936_10_ldst_val : _GEN_64936;
  assign _GEN_65091 = 6'hb == _T_3818 ? _T_5936_11_pdst : _GEN_65001;
  assign _GEN_65116 = 6'hb == _T_3818 ? _T_5936_11_ldst_val : _GEN_65026;
  assign _GEN_65181 = 6'hc == _T_3818 ? _T_5936_12_pdst : _GEN_65091;
  assign _GEN_65206 = 6'hc == _T_3818 ? _T_5936_12_ldst_val : _GEN_65116;
  assign _GEN_65271 = 6'hd == _T_3818 ? _T_5936_13_pdst : _GEN_65181;
  assign _GEN_65296 = 6'hd == _T_3818 ? _T_5936_13_ldst_val : _GEN_65206;
  assign _GEN_65361 = 6'he == _T_3818 ? _T_5936_14_pdst : _GEN_65271;
  assign _GEN_65386 = 6'he == _T_3818 ? _T_5936_14_ldst_val : _GEN_65296;
  assign _GEN_65451 = 6'hf == _T_3818 ? _T_5936_15_pdst : _GEN_65361;
  assign _GEN_65476 = 6'hf == _T_3818 ? _T_5936_15_ldst_val : _GEN_65386;
  assign _GEN_65541 = 6'h10 == _T_3818 ? _T_5936_16_pdst : _GEN_65451;
  assign _GEN_65566 = 6'h10 == _T_3818 ? _T_5936_16_ldst_val : _GEN_65476;
  assign _GEN_65631 = 6'h11 == _T_3818 ? _T_5936_17_pdst : _GEN_65541;
  assign _GEN_65656 = 6'h11 == _T_3818 ? _T_5936_17_ldst_val : _GEN_65566;
  assign _GEN_65721 = 6'h12 == _T_3818 ? _T_5936_18_pdst : _GEN_65631;
  assign _GEN_65746 = 6'h12 == _T_3818 ? _T_5936_18_ldst_val : _GEN_65656;
  assign _GEN_65811 = 6'h13 == _T_3818 ? _T_5936_19_pdst : _GEN_65721;
  assign _GEN_65836 = 6'h13 == _T_3818 ? _T_5936_19_ldst_val : _GEN_65746;
  assign _GEN_65901 = 6'h14 == _T_3818 ? _T_5936_20_pdst : _GEN_65811;
  assign _GEN_65926 = 6'h14 == _T_3818 ? _T_5936_20_ldst_val : _GEN_65836;
  assign _GEN_65991 = 6'h15 == _T_3818 ? _T_5936_21_pdst : _GEN_65901;
  assign _GEN_66016 = 6'h15 == _T_3818 ? _T_5936_21_ldst_val : _GEN_65926;
  assign _GEN_66081 = 6'h16 == _T_3818 ? _T_5936_22_pdst : _GEN_65991;
  assign _GEN_66106 = 6'h16 == _T_3818 ? _T_5936_22_ldst_val : _GEN_66016;
  assign _GEN_66171 = 6'h17 == _T_3818 ? _T_5936_23_pdst : _GEN_66081;
  assign _GEN_66196 = 6'h17 == _T_3818 ? _T_5936_23_ldst_val : _GEN_66106;
  assign _GEN_66261 = 6'h18 == _T_3818 ? _T_5936_24_pdst : _GEN_66171;
  assign _GEN_66286 = 6'h18 == _T_3818 ? _T_5936_24_ldst_val : _GEN_66196;
  assign _GEN_66351 = 6'h19 == _T_3818 ? _T_5936_25_pdst : _GEN_66261;
  assign _GEN_66376 = 6'h19 == _T_3818 ? _T_5936_25_ldst_val : _GEN_66286;
  assign _GEN_66441 = 6'h1a == _T_3818 ? _T_5936_26_pdst : _GEN_66351;
  assign _GEN_66466 = 6'h1a == _T_3818 ? _T_5936_26_ldst_val : _GEN_66376;
  assign _GEN_66531 = 6'h1b == _T_3818 ? _T_5936_27_pdst : _GEN_66441;
  assign _GEN_66556 = 6'h1b == _T_3818 ? _T_5936_27_ldst_val : _GEN_66466;
  assign _GEN_66621 = 6'h1c == _T_3818 ? _T_5936_28_pdst : _GEN_66531;
  assign _GEN_66646 = 6'h1c == _T_3818 ? _T_5936_28_ldst_val : _GEN_66556;
  assign _GEN_66711 = 6'h1d == _T_3818 ? _T_5936_29_pdst : _GEN_66621;
  assign _GEN_66736 = 6'h1d == _T_3818 ? _T_5936_29_ldst_val : _GEN_66646;
  assign _GEN_66801 = 6'h1e == _T_3818 ? _T_5936_30_pdst : _GEN_66711;
  assign _GEN_66826 = 6'h1e == _T_3818 ? _T_5936_30_ldst_val : _GEN_66736;
  assign _GEN_66891 = 6'h1f == _T_3818 ? _T_5936_31_pdst : _GEN_66801;
  assign _GEN_66916 = 6'h1f == _T_3818 ? _T_5936_31_ldst_val : _GEN_66826;
  assign _GEN_66981 = 6'h20 == _T_3818 ? _T_5936_32_pdst : _GEN_66891;
  assign _GEN_67006 = 6'h20 == _T_3818 ? _T_5936_32_ldst_val : _GEN_66916;
  assign _GEN_67071 = 6'h21 == _T_3818 ? _T_5936_33_pdst : _GEN_66981;
  assign _GEN_67096 = 6'h21 == _T_3818 ? _T_5936_33_ldst_val : _GEN_67006;
  assign _GEN_67161 = 6'h22 == _T_3818 ? _T_5936_34_pdst : _GEN_67071;
  assign _GEN_67186 = 6'h22 == _T_3818 ? _T_5936_34_ldst_val : _GEN_67096;
  assign _GEN_67251 = 6'h23 == _T_3818 ? _T_5936_35_pdst : _GEN_67161;
  assign _GEN_67276 = 6'h23 == _T_3818 ? _T_5936_35_ldst_val : _GEN_67186;
  assign _GEN_67341 = 6'h24 == _T_3818 ? _T_5936_36_pdst : _GEN_67251;
  assign _GEN_67366 = 6'h24 == _T_3818 ? _T_5936_36_ldst_val : _GEN_67276;
  assign _GEN_67431 = 6'h25 == _T_3818 ? _T_5936_37_pdst : _GEN_67341;
  assign _GEN_67456 = 6'h25 == _T_3818 ? _T_5936_37_ldst_val : _GEN_67366;
  assign _GEN_67521 = 6'h26 == _T_3818 ? _T_5936_38_pdst : _GEN_67431;
  assign _GEN_67546 = 6'h26 == _T_3818 ? _T_5936_38_ldst_val : _GEN_67456;
  assign _GEN_67611 = 6'h27 == _T_3818 ? _T_5936_39_pdst : _GEN_67521;
  assign _GEN_67636 = 6'h27 == _T_3818 ? _T_5936_39_ldst_val : _GEN_67546;
  assign _T_7706 = _T_6381 & _GEN_436_ldst_val;
  assign _T_7707 = _GEN_437_pdst != io_wb_resps_0_bits_uop_pdst;
  assign _T_7708 = _T_7706 & _T_7707;
  assign _T_7710 = _T_7708 == 1'h0;
  assign _T_7712 = _T_7710 | reset;
  assign _T_7714 = _T_7712 == 1'h0;
  assign _GEN_67729 = 6'h1 == _T_3827 ? _T_5637_1 : _T_5637_0;
  assign _GEN_67730 = 6'h2 == _T_3827 ? _T_5637_2 : _GEN_67729;
  assign _GEN_67731 = 6'h3 == _T_3827 ? _T_5637_3 : _GEN_67730;
  assign _GEN_67732 = 6'h4 == _T_3827 ? _T_5637_4 : _GEN_67731;
  assign _GEN_67733 = 6'h5 == _T_3827 ? _T_5637_5 : _GEN_67732;
  assign _GEN_67734 = 6'h6 == _T_3827 ? _T_5637_6 : _GEN_67733;
  assign _GEN_67735 = 6'h7 == _T_3827 ? _T_5637_7 : _GEN_67734;
  assign _GEN_67736 = 6'h8 == _T_3827 ? _T_5637_8 : _GEN_67735;
  assign _GEN_67737 = 6'h9 == _T_3827 ? _T_5637_9 : _GEN_67736;
  assign _GEN_67738 = 6'ha == _T_3827 ? _T_5637_10 : _GEN_67737;
  assign _GEN_67739 = 6'hb == _T_3827 ? _T_5637_11 : _GEN_67738;
  assign _GEN_67740 = 6'hc == _T_3827 ? _T_5637_12 : _GEN_67739;
  assign _GEN_67741 = 6'hd == _T_3827 ? _T_5637_13 : _GEN_67740;
  assign _GEN_67742 = 6'he == _T_3827 ? _T_5637_14 : _GEN_67741;
  assign _GEN_67743 = 6'hf == _T_3827 ? _T_5637_15 : _GEN_67742;
  assign _GEN_67744 = 6'h10 == _T_3827 ? _T_5637_16 : _GEN_67743;
  assign _GEN_67745 = 6'h11 == _T_3827 ? _T_5637_17 : _GEN_67744;
  assign _GEN_67746 = 6'h12 == _T_3827 ? _T_5637_18 : _GEN_67745;
  assign _GEN_67747 = 6'h13 == _T_3827 ? _T_5637_19 : _GEN_67746;
  assign _GEN_67748 = 6'h14 == _T_3827 ? _T_5637_20 : _GEN_67747;
  assign _GEN_67749 = 6'h15 == _T_3827 ? _T_5637_21 : _GEN_67748;
  assign _GEN_67750 = 6'h16 == _T_3827 ? _T_5637_22 : _GEN_67749;
  assign _GEN_67751 = 6'h17 == _T_3827 ? _T_5637_23 : _GEN_67750;
  assign _GEN_67752 = 6'h18 == _T_3827 ? _T_5637_24 : _GEN_67751;
  assign _GEN_67753 = 6'h19 == _T_3827 ? _T_5637_25 : _GEN_67752;
  assign _GEN_67754 = 6'h1a == _T_3827 ? _T_5637_26 : _GEN_67753;
  assign _GEN_67755 = 6'h1b == _T_3827 ? _T_5637_27 : _GEN_67754;
  assign _GEN_67756 = 6'h1c == _T_3827 ? _T_5637_28 : _GEN_67755;
  assign _GEN_67757 = 6'h1d == _T_3827 ? _T_5637_29 : _GEN_67756;
  assign _GEN_67758 = 6'h1e == _T_3827 ? _T_5637_30 : _GEN_67757;
  assign _GEN_67759 = 6'h1f == _T_3827 ? _T_5637_31 : _GEN_67758;
  assign _GEN_67760 = 6'h20 == _T_3827 ? _T_5637_32 : _GEN_67759;
  assign _GEN_67761 = 6'h21 == _T_3827 ? _T_5637_33 : _GEN_67760;
  assign _GEN_67762 = 6'h22 == _T_3827 ? _T_5637_34 : _GEN_67761;
  assign _GEN_67763 = 6'h23 == _T_3827 ? _T_5637_35 : _GEN_67762;
  assign _GEN_67764 = 6'h24 == _T_3827 ? _T_5637_36 : _GEN_67763;
  assign _GEN_67765 = 6'h25 == _T_3827 ? _T_5637_37 : _GEN_67764;
  assign _GEN_67766 = 6'h26 == _T_3827 ? _T_5637_38 : _GEN_67765;
  assign _GEN_67767 = 6'h27 == _T_3827 ? _T_5637_39 : _GEN_67766;
  assign _T_7754 = _GEN_439 == 1'h0;
  assign _T_7755 = _T_6390 & _T_7754;
  assign _T_7757 = _T_7755 == 1'h0;
  assign _T_7759 = _T_7757 | reset;
  assign _T_7761 = _T_7759 == 1'h0;
  assign _T_7768 = _T_3822[5:0];
  assign _T_7771 = _T_5764__T_7769_data == 1'h0;
  assign _T_7772 = _T_6390 & _T_7771;
  assign _T_7774 = _T_7772 == 1'h0;
  assign _T_7776 = _T_7774 | reset;
  assign _T_7778 = _T_7776 == 1'h0;
  assign _GEN_67820 = 6'h1 == _T_3827 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_67845 = 6'h1 == _T_3827 ? _T_5936_1_ldst_val : _T_5936_0_ldst_val;
  assign _GEN_67910 = 6'h2 == _T_3827 ? _T_5936_2_pdst : _GEN_67820;
  assign _GEN_67935 = 6'h2 == _T_3827 ? _T_5936_2_ldst_val : _GEN_67845;
  assign _GEN_68000 = 6'h3 == _T_3827 ? _T_5936_3_pdst : _GEN_67910;
  assign _GEN_68025 = 6'h3 == _T_3827 ? _T_5936_3_ldst_val : _GEN_67935;
  assign _GEN_68090 = 6'h4 == _T_3827 ? _T_5936_4_pdst : _GEN_68000;
  assign _GEN_68115 = 6'h4 == _T_3827 ? _T_5936_4_ldst_val : _GEN_68025;
  assign _GEN_68180 = 6'h5 == _T_3827 ? _T_5936_5_pdst : _GEN_68090;
  assign _GEN_68205 = 6'h5 == _T_3827 ? _T_5936_5_ldst_val : _GEN_68115;
  assign _GEN_68270 = 6'h6 == _T_3827 ? _T_5936_6_pdst : _GEN_68180;
  assign _GEN_68295 = 6'h6 == _T_3827 ? _T_5936_6_ldst_val : _GEN_68205;
  assign _GEN_68360 = 6'h7 == _T_3827 ? _T_5936_7_pdst : _GEN_68270;
  assign _GEN_68385 = 6'h7 == _T_3827 ? _T_5936_7_ldst_val : _GEN_68295;
  assign _GEN_68450 = 6'h8 == _T_3827 ? _T_5936_8_pdst : _GEN_68360;
  assign _GEN_68475 = 6'h8 == _T_3827 ? _T_5936_8_ldst_val : _GEN_68385;
  assign _GEN_68540 = 6'h9 == _T_3827 ? _T_5936_9_pdst : _GEN_68450;
  assign _GEN_68565 = 6'h9 == _T_3827 ? _T_5936_9_ldst_val : _GEN_68475;
  assign _GEN_68630 = 6'ha == _T_3827 ? _T_5936_10_pdst : _GEN_68540;
  assign _GEN_68655 = 6'ha == _T_3827 ? _T_5936_10_ldst_val : _GEN_68565;
  assign _GEN_68720 = 6'hb == _T_3827 ? _T_5936_11_pdst : _GEN_68630;
  assign _GEN_68745 = 6'hb == _T_3827 ? _T_5936_11_ldst_val : _GEN_68655;
  assign _GEN_68810 = 6'hc == _T_3827 ? _T_5936_12_pdst : _GEN_68720;
  assign _GEN_68835 = 6'hc == _T_3827 ? _T_5936_12_ldst_val : _GEN_68745;
  assign _GEN_68900 = 6'hd == _T_3827 ? _T_5936_13_pdst : _GEN_68810;
  assign _GEN_68925 = 6'hd == _T_3827 ? _T_5936_13_ldst_val : _GEN_68835;
  assign _GEN_68990 = 6'he == _T_3827 ? _T_5936_14_pdst : _GEN_68900;
  assign _GEN_69015 = 6'he == _T_3827 ? _T_5936_14_ldst_val : _GEN_68925;
  assign _GEN_69080 = 6'hf == _T_3827 ? _T_5936_15_pdst : _GEN_68990;
  assign _GEN_69105 = 6'hf == _T_3827 ? _T_5936_15_ldst_val : _GEN_69015;
  assign _GEN_69170 = 6'h10 == _T_3827 ? _T_5936_16_pdst : _GEN_69080;
  assign _GEN_69195 = 6'h10 == _T_3827 ? _T_5936_16_ldst_val : _GEN_69105;
  assign _GEN_69260 = 6'h11 == _T_3827 ? _T_5936_17_pdst : _GEN_69170;
  assign _GEN_69285 = 6'h11 == _T_3827 ? _T_5936_17_ldst_val : _GEN_69195;
  assign _GEN_69350 = 6'h12 == _T_3827 ? _T_5936_18_pdst : _GEN_69260;
  assign _GEN_69375 = 6'h12 == _T_3827 ? _T_5936_18_ldst_val : _GEN_69285;
  assign _GEN_69440 = 6'h13 == _T_3827 ? _T_5936_19_pdst : _GEN_69350;
  assign _GEN_69465 = 6'h13 == _T_3827 ? _T_5936_19_ldst_val : _GEN_69375;
  assign _GEN_69530 = 6'h14 == _T_3827 ? _T_5936_20_pdst : _GEN_69440;
  assign _GEN_69555 = 6'h14 == _T_3827 ? _T_5936_20_ldst_val : _GEN_69465;
  assign _GEN_69620 = 6'h15 == _T_3827 ? _T_5936_21_pdst : _GEN_69530;
  assign _GEN_69645 = 6'h15 == _T_3827 ? _T_5936_21_ldst_val : _GEN_69555;
  assign _GEN_69710 = 6'h16 == _T_3827 ? _T_5936_22_pdst : _GEN_69620;
  assign _GEN_69735 = 6'h16 == _T_3827 ? _T_5936_22_ldst_val : _GEN_69645;
  assign _GEN_69800 = 6'h17 == _T_3827 ? _T_5936_23_pdst : _GEN_69710;
  assign _GEN_69825 = 6'h17 == _T_3827 ? _T_5936_23_ldst_val : _GEN_69735;
  assign _GEN_69890 = 6'h18 == _T_3827 ? _T_5936_24_pdst : _GEN_69800;
  assign _GEN_69915 = 6'h18 == _T_3827 ? _T_5936_24_ldst_val : _GEN_69825;
  assign _GEN_69980 = 6'h19 == _T_3827 ? _T_5936_25_pdst : _GEN_69890;
  assign _GEN_70005 = 6'h19 == _T_3827 ? _T_5936_25_ldst_val : _GEN_69915;
  assign _GEN_70070 = 6'h1a == _T_3827 ? _T_5936_26_pdst : _GEN_69980;
  assign _GEN_70095 = 6'h1a == _T_3827 ? _T_5936_26_ldst_val : _GEN_70005;
  assign _GEN_70160 = 6'h1b == _T_3827 ? _T_5936_27_pdst : _GEN_70070;
  assign _GEN_70185 = 6'h1b == _T_3827 ? _T_5936_27_ldst_val : _GEN_70095;
  assign _GEN_70250 = 6'h1c == _T_3827 ? _T_5936_28_pdst : _GEN_70160;
  assign _GEN_70275 = 6'h1c == _T_3827 ? _T_5936_28_ldst_val : _GEN_70185;
  assign _GEN_70340 = 6'h1d == _T_3827 ? _T_5936_29_pdst : _GEN_70250;
  assign _GEN_70365 = 6'h1d == _T_3827 ? _T_5936_29_ldst_val : _GEN_70275;
  assign _GEN_70430 = 6'h1e == _T_3827 ? _T_5936_30_pdst : _GEN_70340;
  assign _GEN_70455 = 6'h1e == _T_3827 ? _T_5936_30_ldst_val : _GEN_70365;
  assign _GEN_70520 = 6'h1f == _T_3827 ? _T_5936_31_pdst : _GEN_70430;
  assign _GEN_70545 = 6'h1f == _T_3827 ? _T_5936_31_ldst_val : _GEN_70455;
  assign _GEN_70610 = 6'h20 == _T_3827 ? _T_5936_32_pdst : _GEN_70520;
  assign _GEN_70635 = 6'h20 == _T_3827 ? _T_5936_32_ldst_val : _GEN_70545;
  assign _GEN_70700 = 6'h21 == _T_3827 ? _T_5936_33_pdst : _GEN_70610;
  assign _GEN_70725 = 6'h21 == _T_3827 ? _T_5936_33_ldst_val : _GEN_70635;
  assign _GEN_70790 = 6'h22 == _T_3827 ? _T_5936_34_pdst : _GEN_70700;
  assign _GEN_70815 = 6'h22 == _T_3827 ? _T_5936_34_ldst_val : _GEN_70725;
  assign _GEN_70880 = 6'h23 == _T_3827 ? _T_5936_35_pdst : _GEN_70790;
  assign _GEN_70905 = 6'h23 == _T_3827 ? _T_5936_35_ldst_val : _GEN_70815;
  assign _GEN_70970 = 6'h24 == _T_3827 ? _T_5936_36_pdst : _GEN_70880;
  assign _GEN_70995 = 6'h24 == _T_3827 ? _T_5936_36_ldst_val : _GEN_70905;
  assign _GEN_71060 = 6'h25 == _T_3827 ? _T_5936_37_pdst : _GEN_70970;
  assign _GEN_71085 = 6'h25 == _T_3827 ? _T_5936_37_ldst_val : _GEN_70995;
  assign _GEN_71150 = 6'h26 == _T_3827 ? _T_5936_38_pdst : _GEN_71060;
  assign _GEN_71175 = 6'h26 == _T_3827 ? _T_5936_38_ldst_val : _GEN_71085;
  assign _GEN_71240 = 6'h27 == _T_3827 ? _T_5936_39_pdst : _GEN_71150;
  assign _GEN_71265 = 6'h27 == _T_3827 ? _T_5936_39_ldst_val : _GEN_71175;
  assign _T_7783 = _T_6390 & _GEN_440_ldst_val;
  assign _T_7784 = _GEN_441_pdst != io_wb_resps_1_bits_uop_pdst;
  assign _T_7785 = _T_7783 & _T_7784;
  assign _T_7787 = _T_7785 == 1'h0;
  assign _T_7789 = _T_7787 | reset;
  assign _T_7791 = _T_7789 == 1'h0;
  assign _GEN_71358 = 6'h1 == _T_3836 ? _T_5637_1 : _T_5637_0;
  assign _GEN_71359 = 6'h2 == _T_3836 ? _T_5637_2 : _GEN_71358;
  assign _GEN_71360 = 6'h3 == _T_3836 ? _T_5637_3 : _GEN_71359;
  assign _GEN_71361 = 6'h4 == _T_3836 ? _T_5637_4 : _GEN_71360;
  assign _GEN_71362 = 6'h5 == _T_3836 ? _T_5637_5 : _GEN_71361;
  assign _GEN_71363 = 6'h6 == _T_3836 ? _T_5637_6 : _GEN_71362;
  assign _GEN_71364 = 6'h7 == _T_3836 ? _T_5637_7 : _GEN_71363;
  assign _GEN_71365 = 6'h8 == _T_3836 ? _T_5637_8 : _GEN_71364;
  assign _GEN_71366 = 6'h9 == _T_3836 ? _T_5637_9 : _GEN_71365;
  assign _GEN_71367 = 6'ha == _T_3836 ? _T_5637_10 : _GEN_71366;
  assign _GEN_71368 = 6'hb == _T_3836 ? _T_5637_11 : _GEN_71367;
  assign _GEN_71369 = 6'hc == _T_3836 ? _T_5637_12 : _GEN_71368;
  assign _GEN_71370 = 6'hd == _T_3836 ? _T_5637_13 : _GEN_71369;
  assign _GEN_71371 = 6'he == _T_3836 ? _T_5637_14 : _GEN_71370;
  assign _GEN_71372 = 6'hf == _T_3836 ? _T_5637_15 : _GEN_71371;
  assign _GEN_71373 = 6'h10 == _T_3836 ? _T_5637_16 : _GEN_71372;
  assign _GEN_71374 = 6'h11 == _T_3836 ? _T_5637_17 : _GEN_71373;
  assign _GEN_71375 = 6'h12 == _T_3836 ? _T_5637_18 : _GEN_71374;
  assign _GEN_71376 = 6'h13 == _T_3836 ? _T_5637_19 : _GEN_71375;
  assign _GEN_71377 = 6'h14 == _T_3836 ? _T_5637_20 : _GEN_71376;
  assign _GEN_71378 = 6'h15 == _T_3836 ? _T_5637_21 : _GEN_71377;
  assign _GEN_71379 = 6'h16 == _T_3836 ? _T_5637_22 : _GEN_71378;
  assign _GEN_71380 = 6'h17 == _T_3836 ? _T_5637_23 : _GEN_71379;
  assign _GEN_71381 = 6'h18 == _T_3836 ? _T_5637_24 : _GEN_71380;
  assign _GEN_71382 = 6'h19 == _T_3836 ? _T_5637_25 : _GEN_71381;
  assign _GEN_71383 = 6'h1a == _T_3836 ? _T_5637_26 : _GEN_71382;
  assign _GEN_71384 = 6'h1b == _T_3836 ? _T_5637_27 : _GEN_71383;
  assign _GEN_71385 = 6'h1c == _T_3836 ? _T_5637_28 : _GEN_71384;
  assign _GEN_71386 = 6'h1d == _T_3836 ? _T_5637_29 : _GEN_71385;
  assign _GEN_71387 = 6'h1e == _T_3836 ? _T_5637_30 : _GEN_71386;
  assign _GEN_71388 = 6'h1f == _T_3836 ? _T_5637_31 : _GEN_71387;
  assign _GEN_71389 = 6'h20 == _T_3836 ? _T_5637_32 : _GEN_71388;
  assign _GEN_71390 = 6'h21 == _T_3836 ? _T_5637_33 : _GEN_71389;
  assign _GEN_71391 = 6'h22 == _T_3836 ? _T_5637_34 : _GEN_71390;
  assign _GEN_71392 = 6'h23 == _T_3836 ? _T_5637_35 : _GEN_71391;
  assign _GEN_71393 = 6'h24 == _T_3836 ? _T_5637_36 : _GEN_71392;
  assign _GEN_71394 = 6'h25 == _T_3836 ? _T_5637_37 : _GEN_71393;
  assign _GEN_71395 = 6'h26 == _T_3836 ? _T_5637_38 : _GEN_71394;
  assign _GEN_71396 = 6'h27 == _T_3836 ? _T_5637_39 : _GEN_71395;
  assign _T_7831 = _GEN_443 == 1'h0;
  assign _T_7832 = _T_6399 & _T_7831;
  assign _T_7834 = _T_7832 == 1'h0;
  assign _T_7836 = _T_7834 | reset;
  assign _T_7838 = _T_7836 == 1'h0;
  assign _T_7845 = _T_3831[5:0];
  assign _T_7848 = _T_5764__T_7846_data == 1'h0;
  assign _T_7849 = _T_6399 & _T_7848;
  assign _T_7851 = _T_7849 == 1'h0;
  assign _T_7853 = _T_7851 | reset;
  assign _T_7855 = _T_7853 == 1'h0;
  assign _GEN_71449 = 6'h1 == _T_3836 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_71474 = 6'h1 == _T_3836 ? _T_5936_1_ldst_val : _T_5936_0_ldst_val;
  assign _GEN_71539 = 6'h2 == _T_3836 ? _T_5936_2_pdst : _GEN_71449;
  assign _GEN_71564 = 6'h2 == _T_3836 ? _T_5936_2_ldst_val : _GEN_71474;
  assign _GEN_71629 = 6'h3 == _T_3836 ? _T_5936_3_pdst : _GEN_71539;
  assign _GEN_71654 = 6'h3 == _T_3836 ? _T_5936_3_ldst_val : _GEN_71564;
  assign _GEN_71719 = 6'h4 == _T_3836 ? _T_5936_4_pdst : _GEN_71629;
  assign _GEN_71744 = 6'h4 == _T_3836 ? _T_5936_4_ldst_val : _GEN_71654;
  assign _GEN_71809 = 6'h5 == _T_3836 ? _T_5936_5_pdst : _GEN_71719;
  assign _GEN_71834 = 6'h5 == _T_3836 ? _T_5936_5_ldst_val : _GEN_71744;
  assign _GEN_71899 = 6'h6 == _T_3836 ? _T_5936_6_pdst : _GEN_71809;
  assign _GEN_71924 = 6'h6 == _T_3836 ? _T_5936_6_ldst_val : _GEN_71834;
  assign _GEN_71989 = 6'h7 == _T_3836 ? _T_5936_7_pdst : _GEN_71899;
  assign _GEN_72014 = 6'h7 == _T_3836 ? _T_5936_7_ldst_val : _GEN_71924;
  assign _GEN_72079 = 6'h8 == _T_3836 ? _T_5936_8_pdst : _GEN_71989;
  assign _GEN_72104 = 6'h8 == _T_3836 ? _T_5936_8_ldst_val : _GEN_72014;
  assign _GEN_72169 = 6'h9 == _T_3836 ? _T_5936_9_pdst : _GEN_72079;
  assign _GEN_72194 = 6'h9 == _T_3836 ? _T_5936_9_ldst_val : _GEN_72104;
  assign _GEN_72259 = 6'ha == _T_3836 ? _T_5936_10_pdst : _GEN_72169;
  assign _GEN_72284 = 6'ha == _T_3836 ? _T_5936_10_ldst_val : _GEN_72194;
  assign _GEN_72349 = 6'hb == _T_3836 ? _T_5936_11_pdst : _GEN_72259;
  assign _GEN_72374 = 6'hb == _T_3836 ? _T_5936_11_ldst_val : _GEN_72284;
  assign _GEN_72439 = 6'hc == _T_3836 ? _T_5936_12_pdst : _GEN_72349;
  assign _GEN_72464 = 6'hc == _T_3836 ? _T_5936_12_ldst_val : _GEN_72374;
  assign _GEN_72529 = 6'hd == _T_3836 ? _T_5936_13_pdst : _GEN_72439;
  assign _GEN_72554 = 6'hd == _T_3836 ? _T_5936_13_ldst_val : _GEN_72464;
  assign _GEN_72619 = 6'he == _T_3836 ? _T_5936_14_pdst : _GEN_72529;
  assign _GEN_72644 = 6'he == _T_3836 ? _T_5936_14_ldst_val : _GEN_72554;
  assign _GEN_72709 = 6'hf == _T_3836 ? _T_5936_15_pdst : _GEN_72619;
  assign _GEN_72734 = 6'hf == _T_3836 ? _T_5936_15_ldst_val : _GEN_72644;
  assign _GEN_72799 = 6'h10 == _T_3836 ? _T_5936_16_pdst : _GEN_72709;
  assign _GEN_72824 = 6'h10 == _T_3836 ? _T_5936_16_ldst_val : _GEN_72734;
  assign _GEN_72889 = 6'h11 == _T_3836 ? _T_5936_17_pdst : _GEN_72799;
  assign _GEN_72914 = 6'h11 == _T_3836 ? _T_5936_17_ldst_val : _GEN_72824;
  assign _GEN_72979 = 6'h12 == _T_3836 ? _T_5936_18_pdst : _GEN_72889;
  assign _GEN_73004 = 6'h12 == _T_3836 ? _T_5936_18_ldst_val : _GEN_72914;
  assign _GEN_73069 = 6'h13 == _T_3836 ? _T_5936_19_pdst : _GEN_72979;
  assign _GEN_73094 = 6'h13 == _T_3836 ? _T_5936_19_ldst_val : _GEN_73004;
  assign _GEN_73159 = 6'h14 == _T_3836 ? _T_5936_20_pdst : _GEN_73069;
  assign _GEN_73184 = 6'h14 == _T_3836 ? _T_5936_20_ldst_val : _GEN_73094;
  assign _GEN_73249 = 6'h15 == _T_3836 ? _T_5936_21_pdst : _GEN_73159;
  assign _GEN_73274 = 6'h15 == _T_3836 ? _T_5936_21_ldst_val : _GEN_73184;
  assign _GEN_73339 = 6'h16 == _T_3836 ? _T_5936_22_pdst : _GEN_73249;
  assign _GEN_73364 = 6'h16 == _T_3836 ? _T_5936_22_ldst_val : _GEN_73274;
  assign _GEN_73429 = 6'h17 == _T_3836 ? _T_5936_23_pdst : _GEN_73339;
  assign _GEN_73454 = 6'h17 == _T_3836 ? _T_5936_23_ldst_val : _GEN_73364;
  assign _GEN_73519 = 6'h18 == _T_3836 ? _T_5936_24_pdst : _GEN_73429;
  assign _GEN_73544 = 6'h18 == _T_3836 ? _T_5936_24_ldst_val : _GEN_73454;
  assign _GEN_73609 = 6'h19 == _T_3836 ? _T_5936_25_pdst : _GEN_73519;
  assign _GEN_73634 = 6'h19 == _T_3836 ? _T_5936_25_ldst_val : _GEN_73544;
  assign _GEN_73699 = 6'h1a == _T_3836 ? _T_5936_26_pdst : _GEN_73609;
  assign _GEN_73724 = 6'h1a == _T_3836 ? _T_5936_26_ldst_val : _GEN_73634;
  assign _GEN_73789 = 6'h1b == _T_3836 ? _T_5936_27_pdst : _GEN_73699;
  assign _GEN_73814 = 6'h1b == _T_3836 ? _T_5936_27_ldst_val : _GEN_73724;
  assign _GEN_73879 = 6'h1c == _T_3836 ? _T_5936_28_pdst : _GEN_73789;
  assign _GEN_73904 = 6'h1c == _T_3836 ? _T_5936_28_ldst_val : _GEN_73814;
  assign _GEN_73969 = 6'h1d == _T_3836 ? _T_5936_29_pdst : _GEN_73879;
  assign _GEN_73994 = 6'h1d == _T_3836 ? _T_5936_29_ldst_val : _GEN_73904;
  assign _GEN_74059 = 6'h1e == _T_3836 ? _T_5936_30_pdst : _GEN_73969;
  assign _GEN_74084 = 6'h1e == _T_3836 ? _T_5936_30_ldst_val : _GEN_73994;
  assign _GEN_74149 = 6'h1f == _T_3836 ? _T_5936_31_pdst : _GEN_74059;
  assign _GEN_74174 = 6'h1f == _T_3836 ? _T_5936_31_ldst_val : _GEN_74084;
  assign _GEN_74239 = 6'h20 == _T_3836 ? _T_5936_32_pdst : _GEN_74149;
  assign _GEN_74264 = 6'h20 == _T_3836 ? _T_5936_32_ldst_val : _GEN_74174;
  assign _GEN_74329 = 6'h21 == _T_3836 ? _T_5936_33_pdst : _GEN_74239;
  assign _GEN_74354 = 6'h21 == _T_3836 ? _T_5936_33_ldst_val : _GEN_74264;
  assign _GEN_74419 = 6'h22 == _T_3836 ? _T_5936_34_pdst : _GEN_74329;
  assign _GEN_74444 = 6'h22 == _T_3836 ? _T_5936_34_ldst_val : _GEN_74354;
  assign _GEN_74509 = 6'h23 == _T_3836 ? _T_5936_35_pdst : _GEN_74419;
  assign _GEN_74534 = 6'h23 == _T_3836 ? _T_5936_35_ldst_val : _GEN_74444;
  assign _GEN_74599 = 6'h24 == _T_3836 ? _T_5936_36_pdst : _GEN_74509;
  assign _GEN_74624 = 6'h24 == _T_3836 ? _T_5936_36_ldst_val : _GEN_74534;
  assign _GEN_74689 = 6'h25 == _T_3836 ? _T_5936_37_pdst : _GEN_74599;
  assign _GEN_74714 = 6'h25 == _T_3836 ? _T_5936_37_ldst_val : _GEN_74624;
  assign _GEN_74779 = 6'h26 == _T_3836 ? _T_5936_38_pdst : _GEN_74689;
  assign _GEN_74804 = 6'h26 == _T_3836 ? _T_5936_38_ldst_val : _GEN_74714;
  assign _GEN_74869 = 6'h27 == _T_3836 ? _T_5936_39_pdst : _GEN_74779;
  assign _GEN_74894 = 6'h27 == _T_3836 ? _T_5936_39_ldst_val : _GEN_74804;
  assign _T_7860 = _T_6399 & _GEN_444_ldst_val;
  assign _T_7861 = _GEN_445_pdst != io_wb_resps_2_bits_uop_pdst;
  assign _T_7862 = _T_7860 & _T_7861;
  assign _T_7864 = _T_7862 == 1'h0;
  assign _T_7866 = _T_7864 | reset;
  assign _T_7868 = _T_7866 == 1'h0;
  assign _GEN_74987 = 6'h1 == _T_3845 ? _T_5637_1 : _T_5637_0;
  assign _GEN_74988 = 6'h2 == _T_3845 ? _T_5637_2 : _GEN_74987;
  assign _GEN_74989 = 6'h3 == _T_3845 ? _T_5637_3 : _GEN_74988;
  assign _GEN_74990 = 6'h4 == _T_3845 ? _T_5637_4 : _GEN_74989;
  assign _GEN_74991 = 6'h5 == _T_3845 ? _T_5637_5 : _GEN_74990;
  assign _GEN_74992 = 6'h6 == _T_3845 ? _T_5637_6 : _GEN_74991;
  assign _GEN_74993 = 6'h7 == _T_3845 ? _T_5637_7 : _GEN_74992;
  assign _GEN_74994 = 6'h8 == _T_3845 ? _T_5637_8 : _GEN_74993;
  assign _GEN_74995 = 6'h9 == _T_3845 ? _T_5637_9 : _GEN_74994;
  assign _GEN_74996 = 6'ha == _T_3845 ? _T_5637_10 : _GEN_74995;
  assign _GEN_74997 = 6'hb == _T_3845 ? _T_5637_11 : _GEN_74996;
  assign _GEN_74998 = 6'hc == _T_3845 ? _T_5637_12 : _GEN_74997;
  assign _GEN_74999 = 6'hd == _T_3845 ? _T_5637_13 : _GEN_74998;
  assign _GEN_75000 = 6'he == _T_3845 ? _T_5637_14 : _GEN_74999;
  assign _GEN_75001 = 6'hf == _T_3845 ? _T_5637_15 : _GEN_75000;
  assign _GEN_75002 = 6'h10 == _T_3845 ? _T_5637_16 : _GEN_75001;
  assign _GEN_75003 = 6'h11 == _T_3845 ? _T_5637_17 : _GEN_75002;
  assign _GEN_75004 = 6'h12 == _T_3845 ? _T_5637_18 : _GEN_75003;
  assign _GEN_75005 = 6'h13 == _T_3845 ? _T_5637_19 : _GEN_75004;
  assign _GEN_75006 = 6'h14 == _T_3845 ? _T_5637_20 : _GEN_75005;
  assign _GEN_75007 = 6'h15 == _T_3845 ? _T_5637_21 : _GEN_75006;
  assign _GEN_75008 = 6'h16 == _T_3845 ? _T_5637_22 : _GEN_75007;
  assign _GEN_75009 = 6'h17 == _T_3845 ? _T_5637_23 : _GEN_75008;
  assign _GEN_75010 = 6'h18 == _T_3845 ? _T_5637_24 : _GEN_75009;
  assign _GEN_75011 = 6'h19 == _T_3845 ? _T_5637_25 : _GEN_75010;
  assign _GEN_75012 = 6'h1a == _T_3845 ? _T_5637_26 : _GEN_75011;
  assign _GEN_75013 = 6'h1b == _T_3845 ? _T_5637_27 : _GEN_75012;
  assign _GEN_75014 = 6'h1c == _T_3845 ? _T_5637_28 : _GEN_75013;
  assign _GEN_75015 = 6'h1d == _T_3845 ? _T_5637_29 : _GEN_75014;
  assign _GEN_75016 = 6'h1e == _T_3845 ? _T_5637_30 : _GEN_75015;
  assign _GEN_75017 = 6'h1f == _T_3845 ? _T_5637_31 : _GEN_75016;
  assign _GEN_75018 = 6'h20 == _T_3845 ? _T_5637_32 : _GEN_75017;
  assign _GEN_75019 = 6'h21 == _T_3845 ? _T_5637_33 : _GEN_75018;
  assign _GEN_75020 = 6'h22 == _T_3845 ? _T_5637_34 : _GEN_75019;
  assign _GEN_75021 = 6'h23 == _T_3845 ? _T_5637_35 : _GEN_75020;
  assign _GEN_75022 = 6'h24 == _T_3845 ? _T_5637_36 : _GEN_75021;
  assign _GEN_75023 = 6'h25 == _T_3845 ? _T_5637_37 : _GEN_75022;
  assign _GEN_75024 = 6'h26 == _T_3845 ? _T_5637_38 : _GEN_75023;
  assign _GEN_75025 = 6'h27 == _T_3845 ? _T_5637_39 : _GEN_75024;
  assign _T_7908 = _GEN_447 == 1'h0;
  assign _T_7909 = _T_6408 & _T_7908;
  assign _T_7911 = _T_7909 == 1'h0;
  assign _T_7913 = _T_7911 | reset;
  assign _T_7915 = _T_7913 == 1'h0;
  assign _T_7922 = _T_3840[5:0];
  assign _T_7925 = _T_5764__T_7923_data == 1'h0;
  assign _T_7926 = _T_6408 & _T_7925;
  assign _T_7928 = _T_7926 == 1'h0;
  assign _T_7930 = _T_7928 | reset;
  assign _T_7932 = _T_7930 == 1'h0;
  assign _GEN_75078 = 6'h1 == _T_3845 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_75103 = 6'h1 == _T_3845 ? _T_5936_1_ldst_val : _T_5936_0_ldst_val;
  assign _GEN_75168 = 6'h2 == _T_3845 ? _T_5936_2_pdst : _GEN_75078;
  assign _GEN_75193 = 6'h2 == _T_3845 ? _T_5936_2_ldst_val : _GEN_75103;
  assign _GEN_75258 = 6'h3 == _T_3845 ? _T_5936_3_pdst : _GEN_75168;
  assign _GEN_75283 = 6'h3 == _T_3845 ? _T_5936_3_ldst_val : _GEN_75193;
  assign _GEN_75348 = 6'h4 == _T_3845 ? _T_5936_4_pdst : _GEN_75258;
  assign _GEN_75373 = 6'h4 == _T_3845 ? _T_5936_4_ldst_val : _GEN_75283;
  assign _GEN_75438 = 6'h5 == _T_3845 ? _T_5936_5_pdst : _GEN_75348;
  assign _GEN_75463 = 6'h5 == _T_3845 ? _T_5936_5_ldst_val : _GEN_75373;
  assign _GEN_75528 = 6'h6 == _T_3845 ? _T_5936_6_pdst : _GEN_75438;
  assign _GEN_75553 = 6'h6 == _T_3845 ? _T_5936_6_ldst_val : _GEN_75463;
  assign _GEN_75618 = 6'h7 == _T_3845 ? _T_5936_7_pdst : _GEN_75528;
  assign _GEN_75643 = 6'h7 == _T_3845 ? _T_5936_7_ldst_val : _GEN_75553;
  assign _GEN_75708 = 6'h8 == _T_3845 ? _T_5936_8_pdst : _GEN_75618;
  assign _GEN_75733 = 6'h8 == _T_3845 ? _T_5936_8_ldst_val : _GEN_75643;
  assign _GEN_75798 = 6'h9 == _T_3845 ? _T_5936_9_pdst : _GEN_75708;
  assign _GEN_75823 = 6'h9 == _T_3845 ? _T_5936_9_ldst_val : _GEN_75733;
  assign _GEN_75888 = 6'ha == _T_3845 ? _T_5936_10_pdst : _GEN_75798;
  assign _GEN_75913 = 6'ha == _T_3845 ? _T_5936_10_ldst_val : _GEN_75823;
  assign _GEN_75978 = 6'hb == _T_3845 ? _T_5936_11_pdst : _GEN_75888;
  assign _GEN_76003 = 6'hb == _T_3845 ? _T_5936_11_ldst_val : _GEN_75913;
  assign _GEN_76068 = 6'hc == _T_3845 ? _T_5936_12_pdst : _GEN_75978;
  assign _GEN_76093 = 6'hc == _T_3845 ? _T_5936_12_ldst_val : _GEN_76003;
  assign _GEN_76158 = 6'hd == _T_3845 ? _T_5936_13_pdst : _GEN_76068;
  assign _GEN_76183 = 6'hd == _T_3845 ? _T_5936_13_ldst_val : _GEN_76093;
  assign _GEN_76248 = 6'he == _T_3845 ? _T_5936_14_pdst : _GEN_76158;
  assign _GEN_76273 = 6'he == _T_3845 ? _T_5936_14_ldst_val : _GEN_76183;
  assign _GEN_76338 = 6'hf == _T_3845 ? _T_5936_15_pdst : _GEN_76248;
  assign _GEN_76363 = 6'hf == _T_3845 ? _T_5936_15_ldst_val : _GEN_76273;
  assign _GEN_76428 = 6'h10 == _T_3845 ? _T_5936_16_pdst : _GEN_76338;
  assign _GEN_76453 = 6'h10 == _T_3845 ? _T_5936_16_ldst_val : _GEN_76363;
  assign _GEN_76518 = 6'h11 == _T_3845 ? _T_5936_17_pdst : _GEN_76428;
  assign _GEN_76543 = 6'h11 == _T_3845 ? _T_5936_17_ldst_val : _GEN_76453;
  assign _GEN_76608 = 6'h12 == _T_3845 ? _T_5936_18_pdst : _GEN_76518;
  assign _GEN_76633 = 6'h12 == _T_3845 ? _T_5936_18_ldst_val : _GEN_76543;
  assign _GEN_76698 = 6'h13 == _T_3845 ? _T_5936_19_pdst : _GEN_76608;
  assign _GEN_76723 = 6'h13 == _T_3845 ? _T_5936_19_ldst_val : _GEN_76633;
  assign _GEN_76788 = 6'h14 == _T_3845 ? _T_5936_20_pdst : _GEN_76698;
  assign _GEN_76813 = 6'h14 == _T_3845 ? _T_5936_20_ldst_val : _GEN_76723;
  assign _GEN_76878 = 6'h15 == _T_3845 ? _T_5936_21_pdst : _GEN_76788;
  assign _GEN_76903 = 6'h15 == _T_3845 ? _T_5936_21_ldst_val : _GEN_76813;
  assign _GEN_76968 = 6'h16 == _T_3845 ? _T_5936_22_pdst : _GEN_76878;
  assign _GEN_76993 = 6'h16 == _T_3845 ? _T_5936_22_ldst_val : _GEN_76903;
  assign _GEN_77058 = 6'h17 == _T_3845 ? _T_5936_23_pdst : _GEN_76968;
  assign _GEN_77083 = 6'h17 == _T_3845 ? _T_5936_23_ldst_val : _GEN_76993;
  assign _GEN_77148 = 6'h18 == _T_3845 ? _T_5936_24_pdst : _GEN_77058;
  assign _GEN_77173 = 6'h18 == _T_3845 ? _T_5936_24_ldst_val : _GEN_77083;
  assign _GEN_77238 = 6'h19 == _T_3845 ? _T_5936_25_pdst : _GEN_77148;
  assign _GEN_77263 = 6'h19 == _T_3845 ? _T_5936_25_ldst_val : _GEN_77173;
  assign _GEN_77328 = 6'h1a == _T_3845 ? _T_5936_26_pdst : _GEN_77238;
  assign _GEN_77353 = 6'h1a == _T_3845 ? _T_5936_26_ldst_val : _GEN_77263;
  assign _GEN_77418 = 6'h1b == _T_3845 ? _T_5936_27_pdst : _GEN_77328;
  assign _GEN_77443 = 6'h1b == _T_3845 ? _T_5936_27_ldst_val : _GEN_77353;
  assign _GEN_77508 = 6'h1c == _T_3845 ? _T_5936_28_pdst : _GEN_77418;
  assign _GEN_77533 = 6'h1c == _T_3845 ? _T_5936_28_ldst_val : _GEN_77443;
  assign _GEN_77598 = 6'h1d == _T_3845 ? _T_5936_29_pdst : _GEN_77508;
  assign _GEN_77623 = 6'h1d == _T_3845 ? _T_5936_29_ldst_val : _GEN_77533;
  assign _GEN_77688 = 6'h1e == _T_3845 ? _T_5936_30_pdst : _GEN_77598;
  assign _GEN_77713 = 6'h1e == _T_3845 ? _T_5936_30_ldst_val : _GEN_77623;
  assign _GEN_77778 = 6'h1f == _T_3845 ? _T_5936_31_pdst : _GEN_77688;
  assign _GEN_77803 = 6'h1f == _T_3845 ? _T_5936_31_ldst_val : _GEN_77713;
  assign _GEN_77868 = 6'h20 == _T_3845 ? _T_5936_32_pdst : _GEN_77778;
  assign _GEN_77893 = 6'h20 == _T_3845 ? _T_5936_32_ldst_val : _GEN_77803;
  assign _GEN_77958 = 6'h21 == _T_3845 ? _T_5936_33_pdst : _GEN_77868;
  assign _GEN_77983 = 6'h21 == _T_3845 ? _T_5936_33_ldst_val : _GEN_77893;
  assign _GEN_78048 = 6'h22 == _T_3845 ? _T_5936_34_pdst : _GEN_77958;
  assign _GEN_78073 = 6'h22 == _T_3845 ? _T_5936_34_ldst_val : _GEN_77983;
  assign _GEN_78138 = 6'h23 == _T_3845 ? _T_5936_35_pdst : _GEN_78048;
  assign _GEN_78163 = 6'h23 == _T_3845 ? _T_5936_35_ldst_val : _GEN_78073;
  assign _GEN_78228 = 6'h24 == _T_3845 ? _T_5936_36_pdst : _GEN_78138;
  assign _GEN_78253 = 6'h24 == _T_3845 ? _T_5936_36_ldst_val : _GEN_78163;
  assign _GEN_78318 = 6'h25 == _T_3845 ? _T_5936_37_pdst : _GEN_78228;
  assign _GEN_78343 = 6'h25 == _T_3845 ? _T_5936_37_ldst_val : _GEN_78253;
  assign _GEN_78408 = 6'h26 == _T_3845 ? _T_5936_38_pdst : _GEN_78318;
  assign _GEN_78433 = 6'h26 == _T_3845 ? _T_5936_38_ldst_val : _GEN_78343;
  assign _GEN_78498 = 6'h27 == _T_3845 ? _T_5936_39_pdst : _GEN_78408;
  assign _GEN_78523 = 6'h27 == _T_3845 ? _T_5936_39_ldst_val : _GEN_78433;
  assign _T_7937 = _T_6408 & _GEN_448_ldst_val;
  assign _T_7938 = _GEN_449_pdst != io_wb_resps_3_bits_uop_pdst;
  assign _T_7939 = _T_7937 & _T_7938;
  assign _T_7941 = _T_7939 == 1'h0;
  assign _T_7943 = _T_7941 | reset;
  assign _T_7945 = _T_7943 == 1'h0;
  assign _GEN_78616 = 6'h1 == _T_3854 ? _T_5637_1 : _T_5637_0;
  assign _GEN_78617 = 6'h2 == _T_3854 ? _T_5637_2 : _GEN_78616;
  assign _GEN_78618 = 6'h3 == _T_3854 ? _T_5637_3 : _GEN_78617;
  assign _GEN_78619 = 6'h4 == _T_3854 ? _T_5637_4 : _GEN_78618;
  assign _GEN_78620 = 6'h5 == _T_3854 ? _T_5637_5 : _GEN_78619;
  assign _GEN_78621 = 6'h6 == _T_3854 ? _T_5637_6 : _GEN_78620;
  assign _GEN_78622 = 6'h7 == _T_3854 ? _T_5637_7 : _GEN_78621;
  assign _GEN_78623 = 6'h8 == _T_3854 ? _T_5637_8 : _GEN_78622;
  assign _GEN_78624 = 6'h9 == _T_3854 ? _T_5637_9 : _GEN_78623;
  assign _GEN_78625 = 6'ha == _T_3854 ? _T_5637_10 : _GEN_78624;
  assign _GEN_78626 = 6'hb == _T_3854 ? _T_5637_11 : _GEN_78625;
  assign _GEN_78627 = 6'hc == _T_3854 ? _T_5637_12 : _GEN_78626;
  assign _GEN_78628 = 6'hd == _T_3854 ? _T_5637_13 : _GEN_78627;
  assign _GEN_78629 = 6'he == _T_3854 ? _T_5637_14 : _GEN_78628;
  assign _GEN_78630 = 6'hf == _T_3854 ? _T_5637_15 : _GEN_78629;
  assign _GEN_78631 = 6'h10 == _T_3854 ? _T_5637_16 : _GEN_78630;
  assign _GEN_78632 = 6'h11 == _T_3854 ? _T_5637_17 : _GEN_78631;
  assign _GEN_78633 = 6'h12 == _T_3854 ? _T_5637_18 : _GEN_78632;
  assign _GEN_78634 = 6'h13 == _T_3854 ? _T_5637_19 : _GEN_78633;
  assign _GEN_78635 = 6'h14 == _T_3854 ? _T_5637_20 : _GEN_78634;
  assign _GEN_78636 = 6'h15 == _T_3854 ? _T_5637_21 : _GEN_78635;
  assign _GEN_78637 = 6'h16 == _T_3854 ? _T_5637_22 : _GEN_78636;
  assign _GEN_78638 = 6'h17 == _T_3854 ? _T_5637_23 : _GEN_78637;
  assign _GEN_78639 = 6'h18 == _T_3854 ? _T_5637_24 : _GEN_78638;
  assign _GEN_78640 = 6'h19 == _T_3854 ? _T_5637_25 : _GEN_78639;
  assign _GEN_78641 = 6'h1a == _T_3854 ? _T_5637_26 : _GEN_78640;
  assign _GEN_78642 = 6'h1b == _T_3854 ? _T_5637_27 : _GEN_78641;
  assign _GEN_78643 = 6'h1c == _T_3854 ? _T_5637_28 : _GEN_78642;
  assign _GEN_78644 = 6'h1d == _T_3854 ? _T_5637_29 : _GEN_78643;
  assign _GEN_78645 = 6'h1e == _T_3854 ? _T_5637_30 : _GEN_78644;
  assign _GEN_78646 = 6'h1f == _T_3854 ? _T_5637_31 : _GEN_78645;
  assign _GEN_78647 = 6'h20 == _T_3854 ? _T_5637_32 : _GEN_78646;
  assign _GEN_78648 = 6'h21 == _T_3854 ? _T_5637_33 : _GEN_78647;
  assign _GEN_78649 = 6'h22 == _T_3854 ? _T_5637_34 : _GEN_78648;
  assign _GEN_78650 = 6'h23 == _T_3854 ? _T_5637_35 : _GEN_78649;
  assign _GEN_78651 = 6'h24 == _T_3854 ? _T_5637_36 : _GEN_78650;
  assign _GEN_78652 = 6'h25 == _T_3854 ? _T_5637_37 : _GEN_78651;
  assign _GEN_78653 = 6'h26 == _T_3854 ? _T_5637_38 : _GEN_78652;
  assign _GEN_78654 = 6'h27 == _T_3854 ? _T_5637_39 : _GEN_78653;
  assign _T_7985 = _GEN_451 == 1'h0;
  assign _T_7986 = _T_6417 & _T_7985;
  assign _T_7988 = _T_7986 == 1'h0;
  assign _T_7990 = _T_7988 | reset;
  assign _T_7992 = _T_7990 == 1'h0;
  assign _T_7999 = _T_3849[5:0];
  assign _T_8002 = _T_5764__T_8000_data == 1'h0;
  assign _T_8003 = _T_6417 & _T_8002;
  assign _T_8005 = _T_8003 == 1'h0;
  assign _T_8007 = _T_8005 | reset;
  assign _T_8009 = _T_8007 == 1'h0;
  assign _GEN_78707 = 6'h1 == _T_3854 ? _T_5936_1_pdst : _T_5936_0_pdst;
  assign _GEN_78732 = 6'h1 == _T_3854 ? _T_5936_1_ldst_val : _T_5936_0_ldst_val;
  assign _GEN_78797 = 6'h2 == _T_3854 ? _T_5936_2_pdst : _GEN_78707;
  assign _GEN_78822 = 6'h2 == _T_3854 ? _T_5936_2_ldst_val : _GEN_78732;
  assign _GEN_78887 = 6'h3 == _T_3854 ? _T_5936_3_pdst : _GEN_78797;
  assign _GEN_78912 = 6'h3 == _T_3854 ? _T_5936_3_ldst_val : _GEN_78822;
  assign _GEN_78977 = 6'h4 == _T_3854 ? _T_5936_4_pdst : _GEN_78887;
  assign _GEN_79002 = 6'h4 == _T_3854 ? _T_5936_4_ldst_val : _GEN_78912;
  assign _GEN_79067 = 6'h5 == _T_3854 ? _T_5936_5_pdst : _GEN_78977;
  assign _GEN_79092 = 6'h5 == _T_3854 ? _T_5936_5_ldst_val : _GEN_79002;
  assign _GEN_79157 = 6'h6 == _T_3854 ? _T_5936_6_pdst : _GEN_79067;
  assign _GEN_79182 = 6'h6 == _T_3854 ? _T_5936_6_ldst_val : _GEN_79092;
  assign _GEN_79247 = 6'h7 == _T_3854 ? _T_5936_7_pdst : _GEN_79157;
  assign _GEN_79272 = 6'h7 == _T_3854 ? _T_5936_7_ldst_val : _GEN_79182;
  assign _GEN_79337 = 6'h8 == _T_3854 ? _T_5936_8_pdst : _GEN_79247;
  assign _GEN_79362 = 6'h8 == _T_3854 ? _T_5936_8_ldst_val : _GEN_79272;
  assign _GEN_79427 = 6'h9 == _T_3854 ? _T_5936_9_pdst : _GEN_79337;
  assign _GEN_79452 = 6'h9 == _T_3854 ? _T_5936_9_ldst_val : _GEN_79362;
  assign _GEN_79517 = 6'ha == _T_3854 ? _T_5936_10_pdst : _GEN_79427;
  assign _GEN_79542 = 6'ha == _T_3854 ? _T_5936_10_ldst_val : _GEN_79452;
  assign _GEN_79607 = 6'hb == _T_3854 ? _T_5936_11_pdst : _GEN_79517;
  assign _GEN_79632 = 6'hb == _T_3854 ? _T_5936_11_ldst_val : _GEN_79542;
  assign _GEN_79697 = 6'hc == _T_3854 ? _T_5936_12_pdst : _GEN_79607;
  assign _GEN_79722 = 6'hc == _T_3854 ? _T_5936_12_ldst_val : _GEN_79632;
  assign _GEN_79787 = 6'hd == _T_3854 ? _T_5936_13_pdst : _GEN_79697;
  assign _GEN_79812 = 6'hd == _T_3854 ? _T_5936_13_ldst_val : _GEN_79722;
  assign _GEN_79877 = 6'he == _T_3854 ? _T_5936_14_pdst : _GEN_79787;
  assign _GEN_79902 = 6'he == _T_3854 ? _T_5936_14_ldst_val : _GEN_79812;
  assign _GEN_79967 = 6'hf == _T_3854 ? _T_5936_15_pdst : _GEN_79877;
  assign _GEN_79992 = 6'hf == _T_3854 ? _T_5936_15_ldst_val : _GEN_79902;
  assign _GEN_80057 = 6'h10 == _T_3854 ? _T_5936_16_pdst : _GEN_79967;
  assign _GEN_80082 = 6'h10 == _T_3854 ? _T_5936_16_ldst_val : _GEN_79992;
  assign _GEN_80147 = 6'h11 == _T_3854 ? _T_5936_17_pdst : _GEN_80057;
  assign _GEN_80172 = 6'h11 == _T_3854 ? _T_5936_17_ldst_val : _GEN_80082;
  assign _GEN_80237 = 6'h12 == _T_3854 ? _T_5936_18_pdst : _GEN_80147;
  assign _GEN_80262 = 6'h12 == _T_3854 ? _T_5936_18_ldst_val : _GEN_80172;
  assign _GEN_80327 = 6'h13 == _T_3854 ? _T_5936_19_pdst : _GEN_80237;
  assign _GEN_80352 = 6'h13 == _T_3854 ? _T_5936_19_ldst_val : _GEN_80262;
  assign _GEN_80417 = 6'h14 == _T_3854 ? _T_5936_20_pdst : _GEN_80327;
  assign _GEN_80442 = 6'h14 == _T_3854 ? _T_5936_20_ldst_val : _GEN_80352;
  assign _GEN_80507 = 6'h15 == _T_3854 ? _T_5936_21_pdst : _GEN_80417;
  assign _GEN_80532 = 6'h15 == _T_3854 ? _T_5936_21_ldst_val : _GEN_80442;
  assign _GEN_80597 = 6'h16 == _T_3854 ? _T_5936_22_pdst : _GEN_80507;
  assign _GEN_80622 = 6'h16 == _T_3854 ? _T_5936_22_ldst_val : _GEN_80532;
  assign _GEN_80687 = 6'h17 == _T_3854 ? _T_5936_23_pdst : _GEN_80597;
  assign _GEN_80712 = 6'h17 == _T_3854 ? _T_5936_23_ldst_val : _GEN_80622;
  assign _GEN_80777 = 6'h18 == _T_3854 ? _T_5936_24_pdst : _GEN_80687;
  assign _GEN_80802 = 6'h18 == _T_3854 ? _T_5936_24_ldst_val : _GEN_80712;
  assign _GEN_80867 = 6'h19 == _T_3854 ? _T_5936_25_pdst : _GEN_80777;
  assign _GEN_80892 = 6'h19 == _T_3854 ? _T_5936_25_ldst_val : _GEN_80802;
  assign _GEN_80957 = 6'h1a == _T_3854 ? _T_5936_26_pdst : _GEN_80867;
  assign _GEN_80982 = 6'h1a == _T_3854 ? _T_5936_26_ldst_val : _GEN_80892;
  assign _GEN_81047 = 6'h1b == _T_3854 ? _T_5936_27_pdst : _GEN_80957;
  assign _GEN_81072 = 6'h1b == _T_3854 ? _T_5936_27_ldst_val : _GEN_80982;
  assign _GEN_81137 = 6'h1c == _T_3854 ? _T_5936_28_pdst : _GEN_81047;
  assign _GEN_81162 = 6'h1c == _T_3854 ? _T_5936_28_ldst_val : _GEN_81072;
  assign _GEN_81227 = 6'h1d == _T_3854 ? _T_5936_29_pdst : _GEN_81137;
  assign _GEN_81252 = 6'h1d == _T_3854 ? _T_5936_29_ldst_val : _GEN_81162;
  assign _GEN_81317 = 6'h1e == _T_3854 ? _T_5936_30_pdst : _GEN_81227;
  assign _GEN_81342 = 6'h1e == _T_3854 ? _T_5936_30_ldst_val : _GEN_81252;
  assign _GEN_81407 = 6'h1f == _T_3854 ? _T_5936_31_pdst : _GEN_81317;
  assign _GEN_81432 = 6'h1f == _T_3854 ? _T_5936_31_ldst_val : _GEN_81342;
  assign _GEN_81497 = 6'h20 == _T_3854 ? _T_5936_32_pdst : _GEN_81407;
  assign _GEN_81522 = 6'h20 == _T_3854 ? _T_5936_32_ldst_val : _GEN_81432;
  assign _GEN_81587 = 6'h21 == _T_3854 ? _T_5936_33_pdst : _GEN_81497;
  assign _GEN_81612 = 6'h21 == _T_3854 ? _T_5936_33_ldst_val : _GEN_81522;
  assign _GEN_81677 = 6'h22 == _T_3854 ? _T_5936_34_pdst : _GEN_81587;
  assign _GEN_81702 = 6'h22 == _T_3854 ? _T_5936_34_ldst_val : _GEN_81612;
  assign _GEN_81767 = 6'h23 == _T_3854 ? _T_5936_35_pdst : _GEN_81677;
  assign _GEN_81792 = 6'h23 == _T_3854 ? _T_5936_35_ldst_val : _GEN_81702;
  assign _GEN_81857 = 6'h24 == _T_3854 ? _T_5936_36_pdst : _GEN_81767;
  assign _GEN_81882 = 6'h24 == _T_3854 ? _T_5936_36_ldst_val : _GEN_81792;
  assign _GEN_81947 = 6'h25 == _T_3854 ? _T_5936_37_pdst : _GEN_81857;
  assign _GEN_81972 = 6'h25 == _T_3854 ? _T_5936_37_ldst_val : _GEN_81882;
  assign _GEN_82037 = 6'h26 == _T_3854 ? _T_5936_38_pdst : _GEN_81947;
  assign _GEN_82062 = 6'h26 == _T_3854 ? _T_5936_38_ldst_val : _GEN_81972;
  assign _GEN_82127 = 6'h27 == _T_3854 ? _T_5936_39_pdst : _GEN_82037;
  assign _GEN_82152 = 6'h27 == _T_3854 ? _T_5936_39_ldst_val : _GEN_82062;
  assign _T_8014 = _T_6417 & _GEN_452_ldst_val;
  assign _T_8015 = _GEN_453_pdst != io_wb_resps_4_bits_uop_pdst;
  assign _T_8016 = _T_8014 & _T_8015;
  assign _T_8018 = _T_8016 == 1'h0;
  assign _T_8020 = _T_8018 | reset;
  assign _T_8022 = _T_8020 == 1'h0;
  assign _T_8032 = rob_state != 2'h1;
  assign _T_8033 = rob_state != 2'h3;
  assign _T_8034 = _T_8032 & _T_8033;
  assign _T_8038 = _T_8034 == 1'h0;
  assign _T_8039 = can_throw_exception_0 & _T_8038;
  assign _T_8045 = can_throw_exception_0 == 1'h0;
  assign _T_8046 = can_commit_0 & _T_8045;
  assign _T_8049 = _T_8046 & _T_8038;
  assign _T_8051 = can_commit_0 == 1'h0;
  assign _T_8052 = _T_8051 | can_throw_exception_0;
  assign _T_8053 = rob_head_vals_0 & _T_8052;
  assign _T_8054 = _T_8053 | _T_8034;
  assign _T_8056 = _T_8054 == 1'h0;
  assign _T_8057 = can_throw_exception_1 & _T_8056;
  assign _T_8059 = will_commit_0 == 1'h0;
  assign _T_8060 = _T_8057 & _T_8059;
  assign will_throw_exception = _T_8060 | _T_8039;
  assign _T_8062 = can_throw_exception_1 == 1'h0;
  assign _T_8063 = can_commit_1 & _T_8062;
  assign _T_8066 = _T_8063 & _T_8056;
  assign _T_8072 = io_com_xcpt_bits_cause == 64'h10;
  assign _T_8073 = io_com_xcpt_bits_cause == 64'h11;
  assign is_mini_exception = _T_8072 | _T_8073;
  assign _T_8075 = is_mini_exception == 1'h0;
  assign _T_8076 = exception_thrown & _T_8075;
  assign _T_8077 = rob_head_vals_0 | rob_head_vals_1;
  assign _T_8078 = rob_head_vals_0 ? io_commit_uops_0_is_sys_pc2epc : io_commit_uops_1_is_sys_pc2epc;
  assign insn_sys_pc2epc = _T_8077 & _T_8078;
  assign refetch_inst = exception_thrown | insn_sys_pc2epc;
  assign _T_8082 = rob_head >> 1'h1;
  assign _T_8083 = _T_8082[4:0];
  assign _GEN_440 = {{3'd0}, _T_2772__T_8084_data};
  assign _T_8086 = _GEN_440 << 2'h3;
  assign _T_8087 = rob_head[0];
  assign _T_8090 = _T_8082[4:0];
  assign _GEN_441 = {{3'd0}, _T_2775__T_8091_data};
  assign _T_8093 = _GEN_441 << 2'h3;
  assign _GEN_82168 = _T_8087 ? _T_8093 : _T_8086;
  assign _T_8094 = _T_8080[39:0];
  assign _T_8095 = _T_8094[39];
  assign _T_8099 = _T_8095 ? 24'hffffff : 24'h0;
  assign _T_8100 = {_T_8099,_T_8094};
  assign _T_8103 = rob_head_vals_0 ? 3'h0 : 3'h4;
  assign _GEN_444 = {{61'd0}, _T_8103};
  assign _T_8104 = _T_8100 + _GEN_444;
  assign _T_8105 = _T_8104[63:0];
  assign _T_8108 = refetch_inst ? 3'h0 : 3'h4;
  assign _GEN_445 = {{61'd0}, _T_8108};
  assign _T_8109 = _T_8105 + _GEN_445;
  assign flush_pc = _T_8109[63:0];
  assign _T_8110 = exception_thrown | io_csr_eret;
  assign _T_8111 = io_commit_valids_0 & io_commit_uops_0_flush_on_commit;
  assign _T_8112 = io_commit_valids_1 & io_commit_uops_1_flush_on_commit;
  assign _T_8113 = _T_8111 | _T_8112;
  assign flush_val = _T_8110 | _T_8113;
  assign _T_8117 = io_com_xcpt_valid | io_csr_eret;
  assign _T_8118 = _T_8117 ? {{24'd0}, io_csr_evec} : flush_pc;
  assign _T_8122 = exception_thrown & _T_8072;
  assign _T_8125 = io_flush_valid == 1'h0;
  assign _T_8126 = com_lsu_misspec & _T_8125;
  assign _T_8128 = _T_8126 == 1'h0;
  assign _T_8130 = _T_8128 | reset;
  assign _T_8132 = _T_8130 == 1'h0;
  assign _T_8147 = io_commit_valids_0 & io_commit_uops_0_fp_val;
  assign _T_8148 = io_commit_uops_0_is_load | io_commit_uops_0_is_store;
  assign _T_8150 = _T_8148 == 1'h0;
  assign _T_8151 = _T_8147 & _T_8150;
  assign _T_8153 = fflags_val_0 ? rob_head_fflags_0 : 5'h0;
  assign _T_8155 = io_commit_uops_0_fp_val == 1'h0;
  assign _T_8156 = io_commit_valids_0 & _T_8155;
  assign _T_8158 = rob_head_fflags_0 != 5'h0;
  assign _T_8159 = _T_8156 & _T_8158;
  assign _T_8161 = _T_8159 == 1'h0;
  assign _T_8163 = _T_8161 | reset;
  assign _T_8165 = _T_8163 == 1'h0;
  assign _T_8168 = _T_8147 & _T_8148;
  assign _T_8171 = _T_8168 & _T_8158;
  assign _T_8173 = _T_8171 == 1'h0;
  assign _T_8175 = _T_8173 | reset;
  assign _T_8177 = _T_8175 == 1'h0;
  assign _T_8178 = io_commit_valids_1 & io_commit_uops_1_fp_val;
  assign _T_8179 = io_commit_uops_1_is_load | io_commit_uops_1_is_store;
  assign _T_8181 = _T_8179 == 1'h0;
  assign _T_8182 = _T_8178 & _T_8181;
  assign _T_8184 = fflags_val_1 ? rob_head_fflags_1 : 5'h0;
  assign _T_8186 = io_commit_uops_1_fp_val == 1'h0;
  assign _T_8187 = io_commit_valids_1 & _T_8186;
  assign _T_8189 = rob_head_fflags_1 != 5'h0;
  assign _T_8190 = _T_8187 & _T_8189;
  assign _T_8192 = _T_8190 == 1'h0;
  assign _T_8194 = _T_8192 | reset;
  assign _T_8196 = _T_8194 == 1'h0;
  assign _T_8199 = _T_8178 & _T_8179;
  assign _T_8202 = _T_8199 & _T_8189;
  assign _T_8204 = _T_8202 == 1'h0;
  assign _T_8206 = _T_8204 | reset;
  assign _T_8208 = _T_8206 == 1'h0;
  assign _T_8209 = fflags_val_0 | fflags_val_1;
  assign _T_8210 = fflags_0 | fflags_1;
  assign _T_8227 = io_enq_valids_0 & io_enq_uops_0_exception;
  assign _T_8228 = io_enq_valids_1 & io_enq_uops_1_exception;
  assign _T_8229 = io_flush_valid | exception_thrown;
  assign _T_8231 = _T_8229 == 1'h0;
  assign _T_8232 = rob_state != 2'h2;
  assign _T_8233 = _T_8231 & _T_8232;
  assign _T_8234 = io_lxcpt_valid | io_bxcpt_valid;
  assign _T_8236 = io_bxcpt_valid == 1'h0;
  assign _T_8237 = io_lxcpt_valid & _T_8236;
  assign _T_8238 = io_lxcpt_valid & io_bxcpt_valid;
  assign _T_8239 = io_lxcpt_bits_uop_rob_idx <= rob_tail_idx;
  assign _T_8240 = {_T_8239,io_lxcpt_bits_uop_rob_idx};
  assign _T_8241 = io_bxcpt_bits_uop_rob_idx <= rob_tail_idx;
  assign _T_8242 = {_T_8241,io_bxcpt_bits_uop_rob_idx};
  assign _T_8243 = _T_8240 < _T_8242;
  assign _T_8244 = _T_8238 & _T_8243;
  assign _T_8245 = _T_8237 | _T_8244;
  assign _T_8246_br_mask = _T_8245 ? io_lxcpt_bits_uop_br_mask : io_bxcpt_bits_uop_br_mask;
  assign _T_8246_rob_idx = _T_8245 ? io_lxcpt_bits_uop_rob_idx : io_bxcpt_bits_uop_rob_idx;
  assign _T_8252 = r_xcpt_val == 1'h0;
  assign _T_8253 = _T_8246_rob_idx <= rob_tail_idx;
  assign _T_8254 = {_T_8253,_T_8246_rob_idx};
  assign _T_8255 = r_xcpt_uop_rob_idx <= rob_tail_idx;
  assign _T_8256 = {_T_8255,r_xcpt_uop_rob_idx};
  assign _T_8257 = _T_8254 < _T_8256;
  assign _T_8258 = _T_8252 | _T_8257;
  assign _T_8260 = io_lxcpt_valid ? io_lxcpt_bits_cause : 5'h0;
  assign _T_8261 = io_lxcpt_valid ? io_lxcpt_bits_badvaddr : io_bxcpt_bits_badvaddr;
  assign _GEN_82169 = _T_8258 ? 1'h1 : r_xcpt_val;
  assign _GEN_82194 = _T_8258 ? _T_8246_br_mask : r_xcpt_uop_br_mask;
  assign _GEN_82218 = _T_8258 ? _T_8246_rob_idx : r_xcpt_uop_rob_idx;
  assign _GEN_82231 = _T_8258 ? {{59'd0}, _T_8260} : r_xcpt_uop_exc_cause;
  assign _GEN_82260 = _T_8258 ? {{24'd0}, _T_8261} : r_xcpt_badvaddr;
  assign _T_8264 = enq_xcpts_0 | enq_xcpts_1;
  assign _T_8265 = _T_8252 & _T_8264;
  assign _T_8268 = enq_xcpts_0 ? 1'h0 : 1'h1;
  assign _GEN_82285 = _T_8268 ? io_enq_uops_1_br_mask : io_enq_uops_0_br_mask;
  assign _GEN_82309 = _T_8268 ? io_enq_uops_1_rob_idx : io_enq_uops_0_rob_idx;
  assign _GEN_82322 = _T_8268 ? io_enq_uops_1_exc_cause : io_enq_uops_0_exc_cause;
  assign _T_8289 = _GEN_545_exc_cause == 64'h2;
  assign _GEN_448 = {{3'd0}, _T_8268};
  assign _T_8292 = _GEN_448 << 2'h2;
  assign _GEN_449 = {{36'd0}, _T_8292};
  assign _T_8293 = io_enq_uops_0_pc + _GEN_449;
  assign _T_8294 = _T_8293[39:0];
  assign _T_8295 = _T_8289 ? 40'h0 : _T_8294;
  assign _GEN_82351 = _T_8265 ? 1'h1 : r_xcpt_val;
  assign _GEN_82376 = _T_8265 ? _GEN_479_br_mask : r_xcpt_uop_br_mask;
  assign _GEN_82400 = _T_8265 ? _GEN_503_rob_idx : r_xcpt_uop_rob_idx;
  assign _GEN_82413 = _T_8265 ? _GEN_516_exc_cause : r_xcpt_uop_exc_cause;
  assign _GEN_82442 = _T_8265 ? {{24'd0}, _T_8295} : r_xcpt_badvaddr;
  assign _GEN_82443 = _T_8234 ? _GEN_82169 : _GEN_82351;
  assign _GEN_82468 = _T_8234 ? _GEN_82194 : _GEN_82376;
  assign _GEN_82492 = _T_8234 ? _GEN_82218 : _GEN_82400;
  assign _GEN_82505 = _T_8234 ? _GEN_82231 : _GEN_82413;
  assign _GEN_82534 = _T_8234 ? _GEN_82260 : _GEN_82442;
  assign _GEN_82535 = _T_8233 ? _GEN_82443 : r_xcpt_val;
  assign _GEN_82560 = _T_8233 ? _GEN_82468 : r_xcpt_uop_br_mask;
  assign _GEN_82584 = _T_8233 ? _GEN_82492 : r_xcpt_uop_rob_idx;
  assign _GEN_82597 = _T_8233 ? _GEN_82505 : r_xcpt_uop_exc_cause;
  assign _GEN_82626 = _T_8233 ? _GEN_82534 : r_xcpt_badvaddr;
  assign _T_8297 = next_xcpt_uop_br_mask & _T_4111;
  assign _T_8298 = io_brinfo_valid ? _T_8297 : next_xcpt_uop_br_mask;
  assign _T_8300 = io_brinfo_mask & next_xcpt_uop_br_mask;
  assign _T_8302 = _T_8300 != 8'h0;
  assign _T_8303 = _T_4094 & _T_8302;
  assign _T_8304 = io_flush_valid | _T_8303;
  assign _GEN_82627 = _T_8304 ? 1'h0 : _GEN_82535;
  assign _T_8311 = exception_thrown & _T_8252;
  assign _T_8313 = _T_8311 == 1'h0;
  assign _T_8315 = _T_8313 | reset;
  assign _T_8317 = _T_8315 == 1'h0;
  assign _T_8318 = io_empty & r_xcpt_val;
  assign _T_8320 = _T_8318 == 1'h0;
  assign _T_8322 = _T_8320 | reset;
  assign _T_8324 = _T_8322 == 1'h0;
  assign _T_8326 = r_xcpt_uop_rob_idx >> 1'h1;
  assign _GEN_452 = {{1'd0}, rob_head};
  assign _T_8327 = _T_8326 != _GEN_452;
  assign _T_8328 = will_throw_exception & _T_8327;
  assign _T_8330 = _T_8328 == 1'h0;
  assign _T_8332 = _T_8330 | reset;
  assign _T_8334 = _T_8332 == 1'h0;
  assign _T_8335 = {io_commit_valids_1,io_commit_valids_0};
  assign _T_8337 = _T_8335 != 2'h0;
  assign _T_8338 = {will_commit_1,will_commit_0};
  assign _T_8339 = {rob_head_vals_1,rob_head_vals_0};
  assign _T_8340 = _T_8338 ^ _T_8339;
  assign _T_8342 = _T_8340 == 2'h0;
  assign _T_8343 = _T_8337 & _T_8342;
  assign _T_8344 = rob_head == rob_tail;
  assign _T_8345 = r_partial_row & _T_8344;
  assign _T_8347 = _T_8345 == 1'h0;
  assign _T_8348 = _T_8343 & _T_8347;
  assign _T_8350 = rob_head == 6'h27;
  assign _T_8353 = rob_head + 6'h1;
  assign _T_8354 = _T_8353[5:0];
  assign _T_8355 = _T_8350 ? 6'h0 : _T_8354;
  assign _GEN_82628 = finished_committing_row ? _T_8355 : rob_head;
  assign _T_8357 = rob_tail != rob_head;
  assign _T_8358 = _T_4026 & _T_8357;
  assign _T_8360 = rob_tail == 6'h0;
  assign _T_8363 = rob_tail - 6'h1;
  assign _T_8364 = $unsigned(_T_8363);
  assign _T_8365 = _T_8364[5:0];
  assign _T_8366 = _T_8360 ? 6'h27 : _T_8365;
  assign _T_8371 = _T_3916 == 7'h27;
  assign _T_8374 = _T_3916 + 7'h1;
  assign _T_8375 = _T_8374[6:0];
  assign _T_8376 = _T_8371 ? 7'h0 : _T_8375;
  assign _T_8379 = _T_2855 != 2'h0;
  assign _T_8381 = io_enq_partial_stall == 1'h0;
  assign _T_8382 = _T_8379 & _T_8381;
  assign _T_8384 = rob_tail == 6'h27;
  assign _T_8387 = rob_tail + 6'h1;
  assign _T_8388 = _T_8387[5:0];
  assign _T_8389 = _T_8384 ? 6'h0 : _T_8388;
  assign _GEN_82629 = _T_8382 ? _T_8389 : rob_tail;
  assign _GEN_82630 = _T_4094 ? _T_8376 : {{1'd0}, _GEN_82629};
  assign _GEN_82631 = _T_8358 ? {{1'd0}, _T_8366} : _GEN_82630;
  assign full = _T_8389 == rob_head;
  assign _T_8400 = _T_8339 == 2'h0;
  assign _T_8401 = _T_8344 & _T_8400;
  assign _T_8402 = rob_state == 2'h1;
  assign _T_8404 = full == 1'h0;
  assign _T_8405 = _T_8402 & _T_8404;
  assign _T_8406 = 2'h0 == rob_state;
  assign _GEN_82632 = _T_8406 ? 2'h1 : rob_state;
  assign _T_8407 = 2'h1 == rob_state;
  assign _GEN_82633 = _T_2901 ? 2'h3 : _GEN_82632;
  assign _GEN_82634 = _T_2902 ? 2'h3 : _GEN_82633;
  assign _GEN_82635 = exception_thrown ? 2'h2 : _GEN_82634;
  assign _GEN_82636 = _T_8407 ? _GEN_82635 : _GEN_82632;
  assign _T_8410 = 2'h2 == rob_state;
  assign _GEN_82637 = io_empty ? 2'h1 : _GEN_82636;
  assign _GEN_82638 = _T_8410 ? _GEN_82637 : _GEN_82636;
  assign _T_8411 = 2'h3 == rob_state;
  assign _GEN_82639 = io_empty ? 2'h1 : _GEN_82638;
  assign _GEN_82640 = exception_thrown ? 2'h2 : _GEN_82639;
  assign _GEN_82641 = _T_8411 ? _GEN_82640 : _GEN_82638;
  assign _T_8412 = io_commit_valids_0 & rob_head_is_store_0;
  assign _T_8413 = io_commit_valids_0 & rob_head_is_load_0;
  assign _T_8414 = io_commit_valids_1 & rob_head_is_store_1;
  assign _T_8415 = io_commit_valids_1 & rob_head_is_load_1;
  assign _T_8417 = _T_8339[0];
  assign _T_8421 = _T_8417 ? 1'h0 : 1'h1;
  assign _GEN_82642 = _T_8421 ? rob_head_is_load_1 : rob_head_is_load_0;
  assign io_curr_rob_tail = {{1'd0}, rob_tail};
  assign io_get_pc_curr_pc = _T_2838[39:0];
  assign io_get_pc_curr_brob_idx = row_metadata_brob_idx__T_2900_data;
  assign io_get_pc_next_val = _T_2870;
  assign io_get_pc_next_pc = _T_2876[39:0];
  assign io_commit_valids_0 = will_commit_0;
  assign io_commit_valids_1 = will_commit_1;
  assign io_commit_uops_0_pdst = _GEN_157_pdst;
  assign io_commit_uops_0_stale_pdst = _GEN_164_stale_pdst;
  assign io_commit_uops_0_is_fencei = _GEN_171_is_fencei;
  assign io_commit_uops_0_is_store = _GEN_172_is_store;
  assign io_commit_uops_0_is_load = _GEN_174_is_load;
  assign io_commit_uops_0_is_sys_pc2epc = _GEN_175_is_sys_pc2epc;
  assign io_commit_uops_0_flush_on_commit = _GEN_177_flush_on_commit;
  assign io_commit_uops_0_ldst = _GEN_178_ldst;
  assign io_commit_uops_0_dst_rtype = _GEN_183_dst_rtype;
  assign io_commit_uops_0_fp_val = _GEN_187_fp_val;
  assign io_commit_uops_1_pdst = _GEN_384_pdst;
  assign io_commit_uops_1_stale_pdst = _GEN_391_stale_pdst;
  assign io_commit_uops_1_is_fencei = _GEN_398_is_fencei;
  assign io_commit_uops_1_is_store = _GEN_399_is_store;
  assign io_commit_uops_1_is_load = _GEN_401_is_load;
  assign io_commit_uops_1_is_sys_pc2epc = _GEN_402_is_sys_pc2epc;
  assign io_commit_uops_1_flush_on_commit = _GEN_404_flush_on_commit;
  assign io_commit_uops_1_ldst = _GEN_405_ldst;
  assign io_commit_uops_1_dst_rtype = _GEN_410_dst_rtype;
  assign io_commit_uops_1_fp_val = _GEN_414_fp_val;
  assign io_commit_fflags_valid = _T_8209;
  assign io_commit_fflags_bits = _T_8210;
  assign io_commit_rbk_valids_0 = _T_4074;
  assign io_commit_rbk_valids_1 = _T_6638;
  assign io_commit_st_mask_0 = _T_8412;
  assign io_commit_st_mask_1 = _T_8414;
  assign io_commit_ld_mask_0 = _T_8413;
  assign io_commit_ld_mask_1 = _T_8415;
  assign io_com_load_is_at_rob_head = _GEN_546;
  assign io_com_xcpt_valid = _T_8076;
  assign io_com_xcpt_bits_pc = flush_pc;
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause;
  assign io_com_xcpt_bits_badvaddr = r_xcpt_badvaddr;
  assign io_flush_valid = _T_8115;
  assign io_flush_bits_pc = _T_8120;
  assign io_clear_brob = _T_2903;
  assign io_empty = _T_8401;
  assign io_ready = _T_8405;
  assign io_brob_deallocate_valid = _T_2895;
  assign io_brob_deallocate_bits_brob_idx = row_metadata_brob_idx__T_2896_data;
  assign will_commit_0 = _T_8049;
  assign will_commit_1 = _T_8066;
  assign can_commit_0 = _T_4023;
  assign can_commit_1 = _T_6587;
  assign can_throw_exception_0 = _T_4013;
  assign can_throw_exception_1 = _T_6577;
  assign rob_head_vals_0 = _GEN_200;
  assign rob_head_vals_1 = _GEN_427;
  assign rob_head_is_store_0 = _GEN_201_is_store;
  assign rob_head_is_store_1 = _GEN_428_is_store;
  assign rob_head_is_load_0 = _GEN_202_is_load;
  assign rob_head_is_load_1 = _GEN_429_is_load;
  assign rob_head_fflags_0 = _T_3748__T_5017_data;
  assign rob_head_fflags_1 = _T_6312__T_7581_data;
  assign rob_getpc_next_vals_0 = _GEN_204;
  assign rob_getpc_next_vals_1 = _GEN_431;
  assign rob_getpc_curr_vals_0 = _GEN_203;
  assign rob_getpc_curr_vals_1 = _GEN_430;
  assign exception_thrown = will_throw_exception;
  assign _T_2815 = {{24'd0}, _T_2819};
  assign _T_2817 = {{24'd0}, _T_2821};
  assign curr_row_next_pc_val = _T_2846;
  assign _GEN_0 = _GEN_563;
  assign finished_committing_row = _T_8348;
  assign _GEN_26 = io_enq_uops_0_br_mask;
  assign _GEN_54 = io_enq_uops_0_pdst;
  assign _GEN_61 = io_enq_uops_0_stale_pdst;
  assign _GEN_68 = io_enq_uops_0_is_fencei;
  assign _GEN_69 = io_enq_uops_0_is_store;
  assign _GEN_71 = io_enq_uops_0_is_load;
  assign _GEN_72 = io_enq_uops_0_is_sys_pc2epc;
  assign _GEN_74 = io_enq_uops_0_flush_on_commit;
  assign _GEN_75 = io_enq_uops_0_ldst;
  assign _GEN_79 = io_enq_uops_0_ldst_val;
  assign _GEN_80 = io_enq_uops_0_dst_rtype;
  assign _GEN_84 = io_enq_uops_0_fp_val;
  assign _GEN_93 = _GEN_4293;
  assign _GEN_96 = _GEN_8078;
  assign _GEN_97 = _GEN_8122;
  assign _GEN_103 = _GEN_8582;
  assign _GEN_104 = _GEN_8582;
  assign _T_4025 = _GEN_8583;
  assign _GEN_157_pdst = _GEN_12056;
  assign _GEN_164_stale_pdst = _GEN_12063;
  assign _GEN_171_is_fencei = _GEN_12070;
  assign _GEN_172_is_store = _GEN_12071;
  assign _GEN_174_is_load = _GEN_12073;
  assign _GEN_175_is_sys_pc2epc = _GEN_12074;
  assign _GEN_177_flush_on_commit = _GEN_12076;
  assign _GEN_178_ldst = _GEN_12077;
  assign _GEN_183_dst_rtype = _GEN_12082;
  assign _GEN_187_fp_val = _GEN_12086;
  assign _GEN_195 = _GEN_12132;
  assign _GEN_196_dst_rtype = _GEN_12082;
  assign _GEN_197_dst_rtype = _GEN_12082;
  assign _GEN_200 = _GEN_8582;
  assign _GEN_201_is_store = _GEN_22964;
  assign _GEN_202_is_load = _GEN_22966;
  assign _GEN_203 = _GEN_23025;
  assign _GEN_204 = _GEN_23064;
  assign _GEN_208 = _GEN_23343;
  assign _GEN_209_ldst_val = _GEN_26841;
  assign _GEN_210_pdst = _GEN_26816;
  assign _GEN_212 = _GEN_26972;
  assign _GEN_213_ldst_val = _GEN_30470;
  assign _GEN_214_pdst = _GEN_30445;
  assign _GEN_216 = _GEN_30601;
  assign _GEN_217_ldst_val = _GEN_34099;
  assign _GEN_218_pdst = _GEN_34074;
  assign _GEN_220 = _GEN_34230;
  assign _GEN_221_ldst_val = _GEN_37728;
  assign _GEN_222_pdst = _GEN_37703;
  assign _GEN_224 = _GEN_37859;
  assign _GEN_225_ldst_val = _GEN_41357;
  assign _GEN_226_pdst = _GEN_41332;
  assign _GEN_253 = io_enq_uops_1_br_mask;
  assign _GEN_281 = io_enq_uops_1_pdst;
  assign _GEN_288 = io_enq_uops_1_stale_pdst;
  assign _GEN_295 = io_enq_uops_1_is_fencei;
  assign _GEN_296 = io_enq_uops_1_is_store;
  assign _GEN_298 = io_enq_uops_1_is_load;
  assign _GEN_299 = io_enq_uops_1_is_sys_pc2epc;
  assign _GEN_301 = io_enq_uops_1_flush_on_commit;
  assign _GEN_302 = io_enq_uops_1_ldst;
  assign _GEN_306 = io_enq_uops_1_ldst_val;
  assign _GEN_307 = io_enq_uops_1_dst_rtype;
  assign _GEN_311 = io_enq_uops_1_fp_val;
  assign _GEN_320 = _GEN_45088;
  assign _GEN_323 = _GEN_48873;
  assign _GEN_324 = _GEN_48917;
  assign _GEN_330 = _GEN_49377;
  assign _GEN_331 = _GEN_49377;
  assign _T_6589 = _GEN_8583;
  assign _GEN_384_pdst = _GEN_52851;
  assign _GEN_391_stale_pdst = _GEN_52858;
  assign _GEN_398_is_fencei = _GEN_52865;
  assign _GEN_399_is_store = _GEN_52866;
  assign _GEN_401_is_load = _GEN_52868;
  assign _GEN_402_is_sys_pc2epc = _GEN_52869;
  assign _GEN_404_flush_on_commit = _GEN_52871;
  assign _GEN_405_ldst = _GEN_52872;
  assign _GEN_410_dst_rtype = _GEN_52877;
  assign _GEN_414_fp_val = _GEN_52881;
  assign _GEN_422 = _GEN_52927;
  assign _GEN_423_dst_rtype = _GEN_52877;
  assign _GEN_424_dst_rtype = _GEN_52877;
  assign _GEN_427 = _GEN_49377;
  assign _GEN_428_is_store = _GEN_63759;
  assign _GEN_429_is_load = _GEN_63761;
  assign _GEN_430 = _GEN_63820;
  assign _GEN_431 = _GEN_63859;
  assign _GEN_435 = _GEN_64138;
  assign _GEN_436_ldst_val = _GEN_67636;
  assign _GEN_437_pdst = _GEN_67611;
  assign _GEN_439 = _GEN_67767;
  assign _GEN_440_ldst_val = _GEN_71265;
  assign _GEN_441_pdst = _GEN_71240;
  assign _GEN_443 = _GEN_71396;
  assign _GEN_444_ldst_val = _GEN_74894;
  assign _GEN_445_pdst = _GEN_74869;
  assign _GEN_447 = _GEN_75025;
  assign _GEN_448_ldst_val = _GEN_78523;
  assign _GEN_449_pdst = _GEN_78498;
  assign _GEN_451 = _GEN_78654;
  assign _GEN_452_ldst_val = _GEN_82152;
  assign _GEN_453_pdst = _GEN_82127;
  assign _T_8080 = {{24'd0}, _GEN_82168};
  assign fflags_val_0 = _T_8151;
  assign fflags_val_1 = _T_8182;
  assign fflags_0 = _T_8153;
  assign fflags_1 = _T_8184;
  assign next_xcpt_uop_br_mask = _GEN_82560;
  assign next_xcpt_uop_rob_idx = _GEN_82584;
  assign next_xcpt_uop_exc_cause = _GEN_82597;
  assign enq_xcpts_0 = _T_8227;
  assign enq_xcpts_1 = _T_8228;
  assign _GEN_479_br_mask = _GEN_82285;
  assign _GEN_503_rob_idx = _GEN_82309;
  assign _GEN_516_exc_cause = _GEN_82322;
  assign _GEN_545_exc_cause = _GEN_82322;
  assign _GEN_546 = _GEN_82642;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  rob_state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  rob_head = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  rob_tail = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  r_xcpt_val = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  r_xcpt_uop_br_mask = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  r_xcpt_uop_rob_idx = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{$random}};
  r_xcpt_uop_exc_cause = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  r_xcpt_badvaddr = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    _T_2772[initvar] = _RAND_8[36:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {2{$random}};
  _RAND_10 = {2{$random}};
  _RAND_11 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    _T_2775[initvar] = _RAND_11[36:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {2{$random}};
  _RAND_13 = {2{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  r_partial_row = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    row_metadata_brob_idx[initvar] = _RAND_15[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {1{$random}};
  _RAND_17 = {1{$random}};
  _RAND_18 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    row_metadata_has_brorjalr[initvar] = _RAND_18[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_3073_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_3073_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_3073_2 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_3073_3 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_3073_4 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_3073_5 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_3073_6 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_3073_7 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_3073_8 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_3073_9 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_3073_10 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_3073_11 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_3073_12 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_3073_13 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_3073_14 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_3073_15 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_3073_16 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_3073_17 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_3073_18 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_3073_19 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_3073_20 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_3073_21 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_3073_22 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_3073_23 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_3073_24 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_3073_25 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_3073_26 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_3073_27 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_3073_28 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_3073_29 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_3073_30 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_3073_31 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_3073_32 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_3073_33 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_3073_34 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_3073_35 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_3073_36 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_3073_37 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_3073_38 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_3073_39 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_3200[initvar] = _RAND_60[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{$random}};
  _RAND_62 = {1{$random}};
  _RAND_63 = {1{$random}};
  _RAND_64 = {1{$random}};
  _RAND_65 = {1{$random}};
  _RAND_66 = {1{$random}};
  _RAND_67 = {1{$random}};
  _RAND_68 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_3372_0_br_mask = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_3372_0_pdst = _RAND_70[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_3372_0_stale_pdst = _RAND_71[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_3372_0_is_fencei = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_3372_0_is_store = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_3372_0_is_load = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_3372_0_is_sys_pc2epc = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_3372_0_flush_on_commit = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_3372_0_ldst = _RAND_77[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_3372_0_ldst_val = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_3372_0_dst_rtype = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_3372_0_fp_val = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_3372_1_br_mask = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_3372_1_pdst = _RAND_82[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_3372_1_stale_pdst = _RAND_83[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_3372_1_is_fencei = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_3372_1_is_store = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_3372_1_is_load = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_3372_1_is_sys_pc2epc = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_3372_1_flush_on_commit = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_3372_1_ldst = _RAND_89[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_3372_1_ldst_val = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_3372_1_dst_rtype = _RAND_91[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_3372_1_fp_val = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_3372_2_br_mask = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_3372_2_pdst = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_3372_2_stale_pdst = _RAND_95[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_3372_2_is_fencei = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_3372_2_is_store = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_3372_2_is_load = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_3372_2_is_sys_pc2epc = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_3372_2_flush_on_commit = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_3372_2_ldst = _RAND_101[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_3372_2_ldst_val = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_3372_2_dst_rtype = _RAND_103[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_3372_2_fp_val = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_3372_3_br_mask = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_3372_3_pdst = _RAND_106[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_3372_3_stale_pdst = _RAND_107[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_3372_3_is_fencei = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_3372_3_is_store = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_3372_3_is_load = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_3372_3_is_sys_pc2epc = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_3372_3_flush_on_commit = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_3372_3_ldst = _RAND_113[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_3372_3_ldst_val = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_3372_3_dst_rtype = _RAND_115[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_3372_3_fp_val = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_3372_4_br_mask = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_3372_4_pdst = _RAND_118[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_3372_4_stale_pdst = _RAND_119[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_3372_4_is_fencei = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_3372_4_is_store = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_3372_4_is_load = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_3372_4_is_sys_pc2epc = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_3372_4_flush_on_commit = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_3372_4_ldst = _RAND_125[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_3372_4_ldst_val = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_3372_4_dst_rtype = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_3372_4_fp_val = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_3372_5_br_mask = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_3372_5_pdst = _RAND_130[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_3372_5_stale_pdst = _RAND_131[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_3372_5_is_fencei = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_3372_5_is_store = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_3372_5_is_load = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_3372_5_is_sys_pc2epc = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_3372_5_flush_on_commit = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_3372_5_ldst = _RAND_137[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_3372_5_ldst_val = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_3372_5_dst_rtype = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_3372_5_fp_val = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_3372_6_br_mask = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_3372_6_pdst = _RAND_142[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_3372_6_stale_pdst = _RAND_143[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_3372_6_is_fencei = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_3372_6_is_store = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_3372_6_is_load = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_3372_6_is_sys_pc2epc = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_3372_6_flush_on_commit = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_3372_6_ldst = _RAND_149[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_3372_6_ldst_val = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_3372_6_dst_rtype = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_3372_6_fp_val = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_3372_7_br_mask = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_3372_7_pdst = _RAND_154[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_3372_7_stale_pdst = _RAND_155[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_3372_7_is_fencei = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_3372_7_is_store = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_3372_7_is_load = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_3372_7_is_sys_pc2epc = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_3372_7_flush_on_commit = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_3372_7_ldst = _RAND_161[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_3372_7_ldst_val = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_3372_7_dst_rtype = _RAND_163[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_3372_7_fp_val = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_3372_8_br_mask = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_3372_8_pdst = _RAND_166[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_3372_8_stale_pdst = _RAND_167[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_3372_8_is_fencei = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_3372_8_is_store = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_3372_8_is_load = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_3372_8_is_sys_pc2epc = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_3372_8_flush_on_commit = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_3372_8_ldst = _RAND_173[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _T_3372_8_ldst_val = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _T_3372_8_dst_rtype = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _T_3372_8_fp_val = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _T_3372_9_br_mask = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _T_3372_9_pdst = _RAND_178[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _T_3372_9_stale_pdst = _RAND_179[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  _T_3372_9_is_fencei = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  _T_3372_9_is_store = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  _T_3372_9_is_load = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  _T_3372_9_is_sys_pc2epc = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  _T_3372_9_flush_on_commit = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  _T_3372_9_ldst = _RAND_185[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  _T_3372_9_ldst_val = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  _T_3372_9_dst_rtype = _RAND_187[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  _T_3372_9_fp_val = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  _T_3372_10_br_mask = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  _T_3372_10_pdst = _RAND_190[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  _T_3372_10_stale_pdst = _RAND_191[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  _T_3372_10_is_fencei = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  _T_3372_10_is_store = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  _T_3372_10_is_load = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  _T_3372_10_is_sys_pc2epc = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  _T_3372_10_flush_on_commit = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  _T_3372_10_ldst = _RAND_197[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  _T_3372_10_ldst_val = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  _T_3372_10_dst_rtype = _RAND_199[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  _T_3372_10_fp_val = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  _T_3372_11_br_mask = _RAND_201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  _T_3372_11_pdst = _RAND_202[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  _T_3372_11_stale_pdst = _RAND_203[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  _T_3372_11_is_fencei = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  _T_3372_11_is_store = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  _T_3372_11_is_load = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  _T_3372_11_is_sys_pc2epc = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  _T_3372_11_flush_on_commit = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  _T_3372_11_ldst = _RAND_209[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  _T_3372_11_ldst_val = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  _T_3372_11_dst_rtype = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  _T_3372_11_fp_val = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  _T_3372_12_br_mask = _RAND_213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  _T_3372_12_pdst = _RAND_214[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  _T_3372_12_stale_pdst = _RAND_215[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  _T_3372_12_is_fencei = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  _T_3372_12_is_store = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  _T_3372_12_is_load = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  _T_3372_12_is_sys_pc2epc = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  _T_3372_12_flush_on_commit = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  _T_3372_12_ldst = _RAND_221[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  _T_3372_12_ldst_val = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  _T_3372_12_dst_rtype = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  _T_3372_12_fp_val = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  _T_3372_13_br_mask = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  _T_3372_13_pdst = _RAND_226[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  _T_3372_13_stale_pdst = _RAND_227[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  _T_3372_13_is_fencei = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  _T_3372_13_is_store = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  _T_3372_13_is_load = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  _T_3372_13_is_sys_pc2epc = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  _T_3372_13_flush_on_commit = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  _T_3372_13_ldst = _RAND_233[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  _T_3372_13_ldst_val = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  _T_3372_13_dst_rtype = _RAND_235[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  _T_3372_13_fp_val = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  _T_3372_14_br_mask = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  _T_3372_14_pdst = _RAND_238[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  _T_3372_14_stale_pdst = _RAND_239[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  _T_3372_14_is_fencei = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  _T_3372_14_is_store = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  _T_3372_14_is_load = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  _T_3372_14_is_sys_pc2epc = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  _T_3372_14_flush_on_commit = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  _T_3372_14_ldst = _RAND_245[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  _T_3372_14_ldst_val = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  _T_3372_14_dst_rtype = _RAND_247[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  _T_3372_14_fp_val = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  _T_3372_15_br_mask = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  _T_3372_15_pdst = _RAND_250[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  _T_3372_15_stale_pdst = _RAND_251[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  _T_3372_15_is_fencei = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  _T_3372_15_is_store = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  _T_3372_15_is_load = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  _T_3372_15_is_sys_pc2epc = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  _T_3372_15_flush_on_commit = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  _T_3372_15_ldst = _RAND_257[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  _T_3372_15_ldst_val = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  _T_3372_15_dst_rtype = _RAND_259[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  _T_3372_15_fp_val = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  _T_3372_16_br_mask = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  _T_3372_16_pdst = _RAND_262[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  _T_3372_16_stale_pdst = _RAND_263[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  _T_3372_16_is_fencei = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  _T_3372_16_is_store = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  _T_3372_16_is_load = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  _T_3372_16_is_sys_pc2epc = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  _T_3372_16_flush_on_commit = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  _T_3372_16_ldst = _RAND_269[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  _T_3372_16_ldst_val = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  _T_3372_16_dst_rtype = _RAND_271[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  _T_3372_16_fp_val = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  _T_3372_17_br_mask = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  _T_3372_17_pdst = _RAND_274[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  _T_3372_17_stale_pdst = _RAND_275[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  _T_3372_17_is_fencei = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  _T_3372_17_is_store = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  _T_3372_17_is_load = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  _T_3372_17_is_sys_pc2epc = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  _T_3372_17_flush_on_commit = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  _T_3372_17_ldst = _RAND_281[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  _T_3372_17_ldst_val = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  _T_3372_17_dst_rtype = _RAND_283[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  _T_3372_17_fp_val = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  _T_3372_18_br_mask = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  _T_3372_18_pdst = _RAND_286[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  _T_3372_18_stale_pdst = _RAND_287[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  _T_3372_18_is_fencei = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  _T_3372_18_is_store = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  _T_3372_18_is_load = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  _T_3372_18_is_sys_pc2epc = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  _T_3372_18_flush_on_commit = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  _T_3372_18_ldst = _RAND_293[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  _T_3372_18_ldst_val = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  _T_3372_18_dst_rtype = _RAND_295[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  _T_3372_18_fp_val = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  _T_3372_19_br_mask = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  _T_3372_19_pdst = _RAND_298[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  _T_3372_19_stale_pdst = _RAND_299[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  _T_3372_19_is_fencei = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  _T_3372_19_is_store = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  _T_3372_19_is_load = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  _T_3372_19_is_sys_pc2epc = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  _T_3372_19_flush_on_commit = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  _T_3372_19_ldst = _RAND_305[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  _T_3372_19_ldst_val = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  _T_3372_19_dst_rtype = _RAND_307[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  _T_3372_19_fp_val = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  _T_3372_20_br_mask = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  _T_3372_20_pdst = _RAND_310[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  _T_3372_20_stale_pdst = _RAND_311[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  _T_3372_20_is_fencei = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  _T_3372_20_is_store = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  _T_3372_20_is_load = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  _T_3372_20_is_sys_pc2epc = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  _T_3372_20_flush_on_commit = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  _T_3372_20_ldst = _RAND_317[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  _T_3372_20_ldst_val = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  _T_3372_20_dst_rtype = _RAND_319[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  _T_3372_20_fp_val = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  _T_3372_21_br_mask = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  _T_3372_21_pdst = _RAND_322[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  _T_3372_21_stale_pdst = _RAND_323[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  _T_3372_21_is_fencei = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  _T_3372_21_is_store = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  _T_3372_21_is_load = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  _T_3372_21_is_sys_pc2epc = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  _T_3372_21_flush_on_commit = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  _T_3372_21_ldst = _RAND_329[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  _T_3372_21_ldst_val = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  _T_3372_21_dst_rtype = _RAND_331[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{$random}};
  _T_3372_21_fp_val = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{$random}};
  _T_3372_22_br_mask = _RAND_333[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{$random}};
  _T_3372_22_pdst = _RAND_334[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{$random}};
  _T_3372_22_stale_pdst = _RAND_335[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{$random}};
  _T_3372_22_is_fencei = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{$random}};
  _T_3372_22_is_store = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{$random}};
  _T_3372_22_is_load = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{$random}};
  _T_3372_22_is_sys_pc2epc = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{$random}};
  _T_3372_22_flush_on_commit = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{$random}};
  _T_3372_22_ldst = _RAND_341[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{$random}};
  _T_3372_22_ldst_val = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{$random}};
  _T_3372_22_dst_rtype = _RAND_343[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{$random}};
  _T_3372_22_fp_val = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{$random}};
  _T_3372_23_br_mask = _RAND_345[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{$random}};
  _T_3372_23_pdst = _RAND_346[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{$random}};
  _T_3372_23_stale_pdst = _RAND_347[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{$random}};
  _T_3372_23_is_fencei = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{$random}};
  _T_3372_23_is_store = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{$random}};
  _T_3372_23_is_load = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{$random}};
  _T_3372_23_is_sys_pc2epc = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{$random}};
  _T_3372_23_flush_on_commit = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{$random}};
  _T_3372_23_ldst = _RAND_353[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{$random}};
  _T_3372_23_ldst_val = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{$random}};
  _T_3372_23_dst_rtype = _RAND_355[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{$random}};
  _T_3372_23_fp_val = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{$random}};
  _T_3372_24_br_mask = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{$random}};
  _T_3372_24_pdst = _RAND_358[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{$random}};
  _T_3372_24_stale_pdst = _RAND_359[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{$random}};
  _T_3372_24_is_fencei = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{$random}};
  _T_3372_24_is_store = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{$random}};
  _T_3372_24_is_load = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{$random}};
  _T_3372_24_is_sys_pc2epc = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{$random}};
  _T_3372_24_flush_on_commit = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{$random}};
  _T_3372_24_ldst = _RAND_365[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{$random}};
  _T_3372_24_ldst_val = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{$random}};
  _T_3372_24_dst_rtype = _RAND_367[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{$random}};
  _T_3372_24_fp_val = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{$random}};
  _T_3372_25_br_mask = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{$random}};
  _T_3372_25_pdst = _RAND_370[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{$random}};
  _T_3372_25_stale_pdst = _RAND_371[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{$random}};
  _T_3372_25_is_fencei = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{$random}};
  _T_3372_25_is_store = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{$random}};
  _T_3372_25_is_load = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{$random}};
  _T_3372_25_is_sys_pc2epc = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{$random}};
  _T_3372_25_flush_on_commit = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{$random}};
  _T_3372_25_ldst = _RAND_377[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{$random}};
  _T_3372_25_ldst_val = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{$random}};
  _T_3372_25_dst_rtype = _RAND_379[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{$random}};
  _T_3372_25_fp_val = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{$random}};
  _T_3372_26_br_mask = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{$random}};
  _T_3372_26_pdst = _RAND_382[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{$random}};
  _T_3372_26_stale_pdst = _RAND_383[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{$random}};
  _T_3372_26_is_fencei = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{$random}};
  _T_3372_26_is_store = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{$random}};
  _T_3372_26_is_load = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{$random}};
  _T_3372_26_is_sys_pc2epc = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{$random}};
  _T_3372_26_flush_on_commit = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{$random}};
  _T_3372_26_ldst = _RAND_389[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{$random}};
  _T_3372_26_ldst_val = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{$random}};
  _T_3372_26_dst_rtype = _RAND_391[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{$random}};
  _T_3372_26_fp_val = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{$random}};
  _T_3372_27_br_mask = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{$random}};
  _T_3372_27_pdst = _RAND_394[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{$random}};
  _T_3372_27_stale_pdst = _RAND_395[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{$random}};
  _T_3372_27_is_fencei = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{$random}};
  _T_3372_27_is_store = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{$random}};
  _T_3372_27_is_load = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{$random}};
  _T_3372_27_is_sys_pc2epc = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{$random}};
  _T_3372_27_flush_on_commit = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{$random}};
  _T_3372_27_ldst = _RAND_401[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{$random}};
  _T_3372_27_ldst_val = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{$random}};
  _T_3372_27_dst_rtype = _RAND_403[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{$random}};
  _T_3372_27_fp_val = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{$random}};
  _T_3372_28_br_mask = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{$random}};
  _T_3372_28_pdst = _RAND_406[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{$random}};
  _T_3372_28_stale_pdst = _RAND_407[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{$random}};
  _T_3372_28_is_fencei = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{$random}};
  _T_3372_28_is_store = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{$random}};
  _T_3372_28_is_load = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{$random}};
  _T_3372_28_is_sys_pc2epc = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{$random}};
  _T_3372_28_flush_on_commit = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{$random}};
  _T_3372_28_ldst = _RAND_413[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{$random}};
  _T_3372_28_ldst_val = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{$random}};
  _T_3372_28_dst_rtype = _RAND_415[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{$random}};
  _T_3372_28_fp_val = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{$random}};
  _T_3372_29_br_mask = _RAND_417[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{$random}};
  _T_3372_29_pdst = _RAND_418[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{$random}};
  _T_3372_29_stale_pdst = _RAND_419[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{$random}};
  _T_3372_29_is_fencei = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{$random}};
  _T_3372_29_is_store = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{$random}};
  _T_3372_29_is_load = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{$random}};
  _T_3372_29_is_sys_pc2epc = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{$random}};
  _T_3372_29_flush_on_commit = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{$random}};
  _T_3372_29_ldst = _RAND_425[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{$random}};
  _T_3372_29_ldst_val = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{$random}};
  _T_3372_29_dst_rtype = _RAND_427[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{$random}};
  _T_3372_29_fp_val = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{$random}};
  _T_3372_30_br_mask = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{$random}};
  _T_3372_30_pdst = _RAND_430[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{$random}};
  _T_3372_30_stale_pdst = _RAND_431[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{$random}};
  _T_3372_30_is_fencei = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{$random}};
  _T_3372_30_is_store = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{$random}};
  _T_3372_30_is_load = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{$random}};
  _T_3372_30_is_sys_pc2epc = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{$random}};
  _T_3372_30_flush_on_commit = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{$random}};
  _T_3372_30_ldst = _RAND_437[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{$random}};
  _T_3372_30_ldst_val = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{$random}};
  _T_3372_30_dst_rtype = _RAND_439[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{$random}};
  _T_3372_30_fp_val = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{$random}};
  _T_3372_31_br_mask = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{$random}};
  _T_3372_31_pdst = _RAND_442[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{$random}};
  _T_3372_31_stale_pdst = _RAND_443[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{$random}};
  _T_3372_31_is_fencei = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{$random}};
  _T_3372_31_is_store = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{$random}};
  _T_3372_31_is_load = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{$random}};
  _T_3372_31_is_sys_pc2epc = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{$random}};
  _T_3372_31_flush_on_commit = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{$random}};
  _T_3372_31_ldst = _RAND_449[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{$random}};
  _T_3372_31_ldst_val = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{$random}};
  _T_3372_31_dst_rtype = _RAND_451[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{$random}};
  _T_3372_31_fp_val = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{$random}};
  _T_3372_32_br_mask = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{$random}};
  _T_3372_32_pdst = _RAND_454[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{$random}};
  _T_3372_32_stale_pdst = _RAND_455[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{$random}};
  _T_3372_32_is_fencei = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{$random}};
  _T_3372_32_is_store = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{$random}};
  _T_3372_32_is_load = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{$random}};
  _T_3372_32_is_sys_pc2epc = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{$random}};
  _T_3372_32_flush_on_commit = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{$random}};
  _T_3372_32_ldst = _RAND_461[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{$random}};
  _T_3372_32_ldst_val = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{$random}};
  _T_3372_32_dst_rtype = _RAND_463[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{$random}};
  _T_3372_32_fp_val = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{$random}};
  _T_3372_33_br_mask = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{$random}};
  _T_3372_33_pdst = _RAND_466[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{$random}};
  _T_3372_33_stale_pdst = _RAND_467[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{$random}};
  _T_3372_33_is_fencei = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{$random}};
  _T_3372_33_is_store = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{$random}};
  _T_3372_33_is_load = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{$random}};
  _T_3372_33_is_sys_pc2epc = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{$random}};
  _T_3372_33_flush_on_commit = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{$random}};
  _T_3372_33_ldst = _RAND_473[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{$random}};
  _T_3372_33_ldst_val = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{$random}};
  _T_3372_33_dst_rtype = _RAND_475[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{$random}};
  _T_3372_33_fp_val = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{$random}};
  _T_3372_34_br_mask = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{$random}};
  _T_3372_34_pdst = _RAND_478[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{$random}};
  _T_3372_34_stale_pdst = _RAND_479[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{$random}};
  _T_3372_34_is_fencei = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{$random}};
  _T_3372_34_is_store = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{$random}};
  _T_3372_34_is_load = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{$random}};
  _T_3372_34_is_sys_pc2epc = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{$random}};
  _T_3372_34_flush_on_commit = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{$random}};
  _T_3372_34_ldst = _RAND_485[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{$random}};
  _T_3372_34_ldst_val = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{$random}};
  _T_3372_34_dst_rtype = _RAND_487[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{$random}};
  _T_3372_34_fp_val = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{$random}};
  _T_3372_35_br_mask = _RAND_489[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{$random}};
  _T_3372_35_pdst = _RAND_490[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{$random}};
  _T_3372_35_stale_pdst = _RAND_491[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{$random}};
  _T_3372_35_is_fencei = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{$random}};
  _T_3372_35_is_store = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{$random}};
  _T_3372_35_is_load = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{$random}};
  _T_3372_35_is_sys_pc2epc = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{$random}};
  _T_3372_35_flush_on_commit = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{$random}};
  _T_3372_35_ldst = _RAND_497[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{$random}};
  _T_3372_35_ldst_val = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{$random}};
  _T_3372_35_dst_rtype = _RAND_499[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{$random}};
  _T_3372_35_fp_val = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{$random}};
  _T_3372_36_br_mask = _RAND_501[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{$random}};
  _T_3372_36_pdst = _RAND_502[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{$random}};
  _T_3372_36_stale_pdst = _RAND_503[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{$random}};
  _T_3372_36_is_fencei = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{$random}};
  _T_3372_36_is_store = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{$random}};
  _T_3372_36_is_load = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{$random}};
  _T_3372_36_is_sys_pc2epc = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{$random}};
  _T_3372_36_flush_on_commit = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{$random}};
  _T_3372_36_ldst = _RAND_509[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{$random}};
  _T_3372_36_ldst_val = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{$random}};
  _T_3372_36_dst_rtype = _RAND_511[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{$random}};
  _T_3372_36_fp_val = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{$random}};
  _T_3372_37_br_mask = _RAND_513[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{$random}};
  _T_3372_37_pdst = _RAND_514[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{$random}};
  _T_3372_37_stale_pdst = _RAND_515[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{$random}};
  _T_3372_37_is_fencei = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{$random}};
  _T_3372_37_is_store = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{$random}};
  _T_3372_37_is_load = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{$random}};
  _T_3372_37_is_sys_pc2epc = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{$random}};
  _T_3372_37_flush_on_commit = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{$random}};
  _T_3372_37_ldst = _RAND_521[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{$random}};
  _T_3372_37_ldst_val = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{$random}};
  _T_3372_37_dst_rtype = _RAND_523[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{$random}};
  _T_3372_37_fp_val = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{$random}};
  _T_3372_38_br_mask = _RAND_525[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{$random}};
  _T_3372_38_pdst = _RAND_526[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{$random}};
  _T_3372_38_stale_pdst = _RAND_527[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{$random}};
  _T_3372_38_is_fencei = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{$random}};
  _T_3372_38_is_store = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{$random}};
  _T_3372_38_is_load = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{$random}};
  _T_3372_38_is_sys_pc2epc = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{$random}};
  _T_3372_38_flush_on_commit = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{$random}};
  _T_3372_38_ldst = _RAND_533[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{$random}};
  _T_3372_38_ldst_val = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{$random}};
  _T_3372_38_dst_rtype = _RAND_535[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{$random}};
  _T_3372_38_fp_val = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{$random}};
  _T_3372_39_br_mask = _RAND_537[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{$random}};
  _T_3372_39_pdst = _RAND_538[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{$random}};
  _T_3372_39_stale_pdst = _RAND_539[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{$random}};
  _T_3372_39_is_fencei = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{$random}};
  _T_3372_39_is_store = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{$random}};
  _T_3372_39_is_load = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{$random}};
  _T_3372_39_is_sys_pc2epc = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{$random}};
  _T_3372_39_flush_on_commit = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{$random}};
  _T_3372_39_ldst = _RAND_545[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{$random}};
  _T_3372_39_ldst_val = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{$random}};
  _T_3372_39_dst_rtype = _RAND_547[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{$random}};
  _T_3372_39_fp_val = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_549 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_3745[initvar] = _RAND_549[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_550 = {1{$random}};
  _RAND_551 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_3748[initvar] = _RAND_551[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_552 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{$random}};
  _T_5637_0 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{$random}};
  _T_5637_1 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{$random}};
  _T_5637_2 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{$random}};
  _T_5637_3 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{$random}};
  _T_5637_4 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{$random}};
  _T_5637_5 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{$random}};
  _T_5637_6 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{$random}};
  _T_5637_7 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{$random}};
  _T_5637_8 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{$random}};
  _T_5637_9 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{$random}};
  _T_5637_10 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{$random}};
  _T_5637_11 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{$random}};
  _T_5637_12 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{$random}};
  _T_5637_13 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{$random}};
  _T_5637_14 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{$random}};
  _T_5637_15 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{$random}};
  _T_5637_16 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{$random}};
  _T_5637_17 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{$random}};
  _T_5637_18 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{$random}};
  _T_5637_19 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{$random}};
  _T_5637_20 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{$random}};
  _T_5637_21 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{$random}};
  _T_5637_22 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{$random}};
  _T_5637_23 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{$random}};
  _T_5637_24 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{$random}};
  _T_5637_25 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{$random}};
  _T_5637_26 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{$random}};
  _T_5637_27 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{$random}};
  _T_5637_28 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{$random}};
  _T_5637_29 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{$random}};
  _T_5637_30 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{$random}};
  _T_5637_31 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{$random}};
  _T_5637_32 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{$random}};
  _T_5637_33 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{$random}};
  _T_5637_34 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{$random}};
  _T_5637_35 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{$random}};
  _T_5637_36 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{$random}};
  _T_5637_37 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{$random}};
  _T_5637_38 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{$random}};
  _T_5637_39 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_593 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_5764[initvar] = _RAND_593[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_594 = {1{$random}};
  _RAND_595 = {1{$random}};
  _RAND_596 = {1{$random}};
  _RAND_597 = {1{$random}};
  _RAND_598 = {1{$random}};
  _RAND_599 = {1{$random}};
  _RAND_600 = {1{$random}};
  _RAND_601 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{$random}};
  _T_5936_0_br_mask = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{$random}};
  _T_5936_0_pdst = _RAND_603[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{$random}};
  _T_5936_0_stale_pdst = _RAND_604[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{$random}};
  _T_5936_0_is_fencei = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{$random}};
  _T_5936_0_is_store = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{$random}};
  _T_5936_0_is_load = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{$random}};
  _T_5936_0_is_sys_pc2epc = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{$random}};
  _T_5936_0_flush_on_commit = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{$random}};
  _T_5936_0_ldst = _RAND_610[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{$random}};
  _T_5936_0_ldst_val = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{$random}};
  _T_5936_0_dst_rtype = _RAND_612[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{$random}};
  _T_5936_0_fp_val = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{$random}};
  _T_5936_1_br_mask = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{$random}};
  _T_5936_1_pdst = _RAND_615[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{$random}};
  _T_5936_1_stale_pdst = _RAND_616[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{$random}};
  _T_5936_1_is_fencei = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{$random}};
  _T_5936_1_is_store = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{$random}};
  _T_5936_1_is_load = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{$random}};
  _T_5936_1_is_sys_pc2epc = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{$random}};
  _T_5936_1_flush_on_commit = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{$random}};
  _T_5936_1_ldst = _RAND_622[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{$random}};
  _T_5936_1_ldst_val = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{$random}};
  _T_5936_1_dst_rtype = _RAND_624[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{$random}};
  _T_5936_1_fp_val = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{$random}};
  _T_5936_2_br_mask = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{$random}};
  _T_5936_2_pdst = _RAND_627[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{$random}};
  _T_5936_2_stale_pdst = _RAND_628[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{$random}};
  _T_5936_2_is_fencei = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{$random}};
  _T_5936_2_is_store = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{$random}};
  _T_5936_2_is_load = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{$random}};
  _T_5936_2_is_sys_pc2epc = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{$random}};
  _T_5936_2_flush_on_commit = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{$random}};
  _T_5936_2_ldst = _RAND_634[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{$random}};
  _T_5936_2_ldst_val = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{$random}};
  _T_5936_2_dst_rtype = _RAND_636[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{$random}};
  _T_5936_2_fp_val = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{$random}};
  _T_5936_3_br_mask = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{$random}};
  _T_5936_3_pdst = _RAND_639[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{$random}};
  _T_5936_3_stale_pdst = _RAND_640[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{$random}};
  _T_5936_3_is_fencei = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{$random}};
  _T_5936_3_is_store = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{$random}};
  _T_5936_3_is_load = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{$random}};
  _T_5936_3_is_sys_pc2epc = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{$random}};
  _T_5936_3_flush_on_commit = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{$random}};
  _T_5936_3_ldst = _RAND_646[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{$random}};
  _T_5936_3_ldst_val = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{$random}};
  _T_5936_3_dst_rtype = _RAND_648[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{$random}};
  _T_5936_3_fp_val = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{$random}};
  _T_5936_4_br_mask = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{$random}};
  _T_5936_4_pdst = _RAND_651[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{$random}};
  _T_5936_4_stale_pdst = _RAND_652[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{$random}};
  _T_5936_4_is_fencei = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{$random}};
  _T_5936_4_is_store = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{$random}};
  _T_5936_4_is_load = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{$random}};
  _T_5936_4_is_sys_pc2epc = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{$random}};
  _T_5936_4_flush_on_commit = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{$random}};
  _T_5936_4_ldst = _RAND_658[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{$random}};
  _T_5936_4_ldst_val = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{$random}};
  _T_5936_4_dst_rtype = _RAND_660[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{$random}};
  _T_5936_4_fp_val = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{$random}};
  _T_5936_5_br_mask = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{$random}};
  _T_5936_5_pdst = _RAND_663[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{$random}};
  _T_5936_5_stale_pdst = _RAND_664[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{$random}};
  _T_5936_5_is_fencei = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{$random}};
  _T_5936_5_is_store = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{$random}};
  _T_5936_5_is_load = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{$random}};
  _T_5936_5_is_sys_pc2epc = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{$random}};
  _T_5936_5_flush_on_commit = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{$random}};
  _T_5936_5_ldst = _RAND_670[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{$random}};
  _T_5936_5_ldst_val = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{$random}};
  _T_5936_5_dst_rtype = _RAND_672[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{$random}};
  _T_5936_5_fp_val = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{$random}};
  _T_5936_6_br_mask = _RAND_674[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{$random}};
  _T_5936_6_pdst = _RAND_675[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{$random}};
  _T_5936_6_stale_pdst = _RAND_676[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{$random}};
  _T_5936_6_is_fencei = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{$random}};
  _T_5936_6_is_store = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{$random}};
  _T_5936_6_is_load = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{$random}};
  _T_5936_6_is_sys_pc2epc = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{$random}};
  _T_5936_6_flush_on_commit = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{$random}};
  _T_5936_6_ldst = _RAND_682[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{$random}};
  _T_5936_6_ldst_val = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{$random}};
  _T_5936_6_dst_rtype = _RAND_684[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{$random}};
  _T_5936_6_fp_val = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{$random}};
  _T_5936_7_br_mask = _RAND_686[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{$random}};
  _T_5936_7_pdst = _RAND_687[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{$random}};
  _T_5936_7_stale_pdst = _RAND_688[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{$random}};
  _T_5936_7_is_fencei = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{$random}};
  _T_5936_7_is_store = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{$random}};
  _T_5936_7_is_load = _RAND_691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{$random}};
  _T_5936_7_is_sys_pc2epc = _RAND_692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{$random}};
  _T_5936_7_flush_on_commit = _RAND_693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{$random}};
  _T_5936_7_ldst = _RAND_694[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{$random}};
  _T_5936_7_ldst_val = _RAND_695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{$random}};
  _T_5936_7_dst_rtype = _RAND_696[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{$random}};
  _T_5936_7_fp_val = _RAND_697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{$random}};
  _T_5936_8_br_mask = _RAND_698[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{$random}};
  _T_5936_8_pdst = _RAND_699[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{$random}};
  _T_5936_8_stale_pdst = _RAND_700[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{$random}};
  _T_5936_8_is_fencei = _RAND_701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{$random}};
  _T_5936_8_is_store = _RAND_702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{$random}};
  _T_5936_8_is_load = _RAND_703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{$random}};
  _T_5936_8_is_sys_pc2epc = _RAND_704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{$random}};
  _T_5936_8_flush_on_commit = _RAND_705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{$random}};
  _T_5936_8_ldst = _RAND_706[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{$random}};
  _T_5936_8_ldst_val = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{$random}};
  _T_5936_8_dst_rtype = _RAND_708[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{$random}};
  _T_5936_8_fp_val = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{$random}};
  _T_5936_9_br_mask = _RAND_710[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{$random}};
  _T_5936_9_pdst = _RAND_711[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{$random}};
  _T_5936_9_stale_pdst = _RAND_712[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{$random}};
  _T_5936_9_is_fencei = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{$random}};
  _T_5936_9_is_store = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{$random}};
  _T_5936_9_is_load = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{$random}};
  _T_5936_9_is_sys_pc2epc = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{$random}};
  _T_5936_9_flush_on_commit = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{$random}};
  _T_5936_9_ldst = _RAND_718[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{$random}};
  _T_5936_9_ldst_val = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{$random}};
  _T_5936_9_dst_rtype = _RAND_720[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{$random}};
  _T_5936_9_fp_val = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{$random}};
  _T_5936_10_br_mask = _RAND_722[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{$random}};
  _T_5936_10_pdst = _RAND_723[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{$random}};
  _T_5936_10_stale_pdst = _RAND_724[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{$random}};
  _T_5936_10_is_fencei = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{$random}};
  _T_5936_10_is_store = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{$random}};
  _T_5936_10_is_load = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{$random}};
  _T_5936_10_is_sys_pc2epc = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{$random}};
  _T_5936_10_flush_on_commit = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{$random}};
  _T_5936_10_ldst = _RAND_730[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{$random}};
  _T_5936_10_ldst_val = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{$random}};
  _T_5936_10_dst_rtype = _RAND_732[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{$random}};
  _T_5936_10_fp_val = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{$random}};
  _T_5936_11_br_mask = _RAND_734[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{$random}};
  _T_5936_11_pdst = _RAND_735[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{$random}};
  _T_5936_11_stale_pdst = _RAND_736[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{$random}};
  _T_5936_11_is_fencei = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{$random}};
  _T_5936_11_is_store = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{$random}};
  _T_5936_11_is_load = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{$random}};
  _T_5936_11_is_sys_pc2epc = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{$random}};
  _T_5936_11_flush_on_commit = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{$random}};
  _T_5936_11_ldst = _RAND_742[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{$random}};
  _T_5936_11_ldst_val = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{$random}};
  _T_5936_11_dst_rtype = _RAND_744[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{$random}};
  _T_5936_11_fp_val = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{$random}};
  _T_5936_12_br_mask = _RAND_746[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{$random}};
  _T_5936_12_pdst = _RAND_747[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{$random}};
  _T_5936_12_stale_pdst = _RAND_748[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{$random}};
  _T_5936_12_is_fencei = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{$random}};
  _T_5936_12_is_store = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{$random}};
  _T_5936_12_is_load = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{$random}};
  _T_5936_12_is_sys_pc2epc = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{$random}};
  _T_5936_12_flush_on_commit = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{$random}};
  _T_5936_12_ldst = _RAND_754[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{$random}};
  _T_5936_12_ldst_val = _RAND_755[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{$random}};
  _T_5936_12_dst_rtype = _RAND_756[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{$random}};
  _T_5936_12_fp_val = _RAND_757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{$random}};
  _T_5936_13_br_mask = _RAND_758[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{$random}};
  _T_5936_13_pdst = _RAND_759[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{$random}};
  _T_5936_13_stale_pdst = _RAND_760[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{$random}};
  _T_5936_13_is_fencei = _RAND_761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{$random}};
  _T_5936_13_is_store = _RAND_762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{$random}};
  _T_5936_13_is_load = _RAND_763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{$random}};
  _T_5936_13_is_sys_pc2epc = _RAND_764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{$random}};
  _T_5936_13_flush_on_commit = _RAND_765[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{$random}};
  _T_5936_13_ldst = _RAND_766[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{$random}};
  _T_5936_13_ldst_val = _RAND_767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{$random}};
  _T_5936_13_dst_rtype = _RAND_768[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{$random}};
  _T_5936_13_fp_val = _RAND_769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{$random}};
  _T_5936_14_br_mask = _RAND_770[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{$random}};
  _T_5936_14_pdst = _RAND_771[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{$random}};
  _T_5936_14_stale_pdst = _RAND_772[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{$random}};
  _T_5936_14_is_fencei = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{$random}};
  _T_5936_14_is_store = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{$random}};
  _T_5936_14_is_load = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{$random}};
  _T_5936_14_is_sys_pc2epc = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{$random}};
  _T_5936_14_flush_on_commit = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{$random}};
  _T_5936_14_ldst = _RAND_778[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{$random}};
  _T_5936_14_ldst_val = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{$random}};
  _T_5936_14_dst_rtype = _RAND_780[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{$random}};
  _T_5936_14_fp_val = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{$random}};
  _T_5936_15_br_mask = _RAND_782[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{$random}};
  _T_5936_15_pdst = _RAND_783[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{$random}};
  _T_5936_15_stale_pdst = _RAND_784[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{$random}};
  _T_5936_15_is_fencei = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{$random}};
  _T_5936_15_is_store = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{$random}};
  _T_5936_15_is_load = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{$random}};
  _T_5936_15_is_sys_pc2epc = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{$random}};
  _T_5936_15_flush_on_commit = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{$random}};
  _T_5936_15_ldst = _RAND_790[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{$random}};
  _T_5936_15_ldst_val = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{$random}};
  _T_5936_15_dst_rtype = _RAND_792[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{$random}};
  _T_5936_15_fp_val = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{$random}};
  _T_5936_16_br_mask = _RAND_794[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{$random}};
  _T_5936_16_pdst = _RAND_795[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{$random}};
  _T_5936_16_stale_pdst = _RAND_796[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{$random}};
  _T_5936_16_is_fencei = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{$random}};
  _T_5936_16_is_store = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{$random}};
  _T_5936_16_is_load = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{$random}};
  _T_5936_16_is_sys_pc2epc = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{$random}};
  _T_5936_16_flush_on_commit = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{$random}};
  _T_5936_16_ldst = _RAND_802[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{$random}};
  _T_5936_16_ldst_val = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{$random}};
  _T_5936_16_dst_rtype = _RAND_804[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{$random}};
  _T_5936_16_fp_val = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{$random}};
  _T_5936_17_br_mask = _RAND_806[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{$random}};
  _T_5936_17_pdst = _RAND_807[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{$random}};
  _T_5936_17_stale_pdst = _RAND_808[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{$random}};
  _T_5936_17_is_fencei = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{$random}};
  _T_5936_17_is_store = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{$random}};
  _T_5936_17_is_load = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{$random}};
  _T_5936_17_is_sys_pc2epc = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{$random}};
  _T_5936_17_flush_on_commit = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{$random}};
  _T_5936_17_ldst = _RAND_814[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{$random}};
  _T_5936_17_ldst_val = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{$random}};
  _T_5936_17_dst_rtype = _RAND_816[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{$random}};
  _T_5936_17_fp_val = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{$random}};
  _T_5936_18_br_mask = _RAND_818[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{$random}};
  _T_5936_18_pdst = _RAND_819[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{$random}};
  _T_5936_18_stale_pdst = _RAND_820[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{$random}};
  _T_5936_18_is_fencei = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{$random}};
  _T_5936_18_is_store = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{$random}};
  _T_5936_18_is_load = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{$random}};
  _T_5936_18_is_sys_pc2epc = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{$random}};
  _T_5936_18_flush_on_commit = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{$random}};
  _T_5936_18_ldst = _RAND_826[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{$random}};
  _T_5936_18_ldst_val = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{$random}};
  _T_5936_18_dst_rtype = _RAND_828[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{$random}};
  _T_5936_18_fp_val = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{$random}};
  _T_5936_19_br_mask = _RAND_830[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{$random}};
  _T_5936_19_pdst = _RAND_831[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{$random}};
  _T_5936_19_stale_pdst = _RAND_832[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{$random}};
  _T_5936_19_is_fencei = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{$random}};
  _T_5936_19_is_store = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{$random}};
  _T_5936_19_is_load = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{$random}};
  _T_5936_19_is_sys_pc2epc = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{$random}};
  _T_5936_19_flush_on_commit = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{$random}};
  _T_5936_19_ldst = _RAND_838[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{$random}};
  _T_5936_19_ldst_val = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{$random}};
  _T_5936_19_dst_rtype = _RAND_840[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{$random}};
  _T_5936_19_fp_val = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{$random}};
  _T_5936_20_br_mask = _RAND_842[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{$random}};
  _T_5936_20_pdst = _RAND_843[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{$random}};
  _T_5936_20_stale_pdst = _RAND_844[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{$random}};
  _T_5936_20_is_fencei = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{$random}};
  _T_5936_20_is_store = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{$random}};
  _T_5936_20_is_load = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{$random}};
  _T_5936_20_is_sys_pc2epc = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{$random}};
  _T_5936_20_flush_on_commit = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{$random}};
  _T_5936_20_ldst = _RAND_850[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{$random}};
  _T_5936_20_ldst_val = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{$random}};
  _T_5936_20_dst_rtype = _RAND_852[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{$random}};
  _T_5936_20_fp_val = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{$random}};
  _T_5936_21_br_mask = _RAND_854[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{$random}};
  _T_5936_21_pdst = _RAND_855[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{$random}};
  _T_5936_21_stale_pdst = _RAND_856[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{$random}};
  _T_5936_21_is_fencei = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{$random}};
  _T_5936_21_is_store = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{$random}};
  _T_5936_21_is_load = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{$random}};
  _T_5936_21_is_sys_pc2epc = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{$random}};
  _T_5936_21_flush_on_commit = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{$random}};
  _T_5936_21_ldst = _RAND_862[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{$random}};
  _T_5936_21_ldst_val = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{$random}};
  _T_5936_21_dst_rtype = _RAND_864[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{$random}};
  _T_5936_21_fp_val = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{$random}};
  _T_5936_22_br_mask = _RAND_866[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{$random}};
  _T_5936_22_pdst = _RAND_867[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{$random}};
  _T_5936_22_stale_pdst = _RAND_868[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{$random}};
  _T_5936_22_is_fencei = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{$random}};
  _T_5936_22_is_store = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{$random}};
  _T_5936_22_is_load = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{$random}};
  _T_5936_22_is_sys_pc2epc = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{$random}};
  _T_5936_22_flush_on_commit = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{$random}};
  _T_5936_22_ldst = _RAND_874[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{$random}};
  _T_5936_22_ldst_val = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{$random}};
  _T_5936_22_dst_rtype = _RAND_876[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{$random}};
  _T_5936_22_fp_val = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{$random}};
  _T_5936_23_br_mask = _RAND_878[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{$random}};
  _T_5936_23_pdst = _RAND_879[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{$random}};
  _T_5936_23_stale_pdst = _RAND_880[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{$random}};
  _T_5936_23_is_fencei = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{$random}};
  _T_5936_23_is_store = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{$random}};
  _T_5936_23_is_load = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{$random}};
  _T_5936_23_is_sys_pc2epc = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{$random}};
  _T_5936_23_flush_on_commit = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{$random}};
  _T_5936_23_ldst = _RAND_886[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{$random}};
  _T_5936_23_ldst_val = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{$random}};
  _T_5936_23_dst_rtype = _RAND_888[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{$random}};
  _T_5936_23_fp_val = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{$random}};
  _T_5936_24_br_mask = _RAND_890[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{$random}};
  _T_5936_24_pdst = _RAND_891[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{$random}};
  _T_5936_24_stale_pdst = _RAND_892[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{$random}};
  _T_5936_24_is_fencei = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{$random}};
  _T_5936_24_is_store = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{$random}};
  _T_5936_24_is_load = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{$random}};
  _T_5936_24_is_sys_pc2epc = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{$random}};
  _T_5936_24_flush_on_commit = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{$random}};
  _T_5936_24_ldst = _RAND_898[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{$random}};
  _T_5936_24_ldst_val = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{$random}};
  _T_5936_24_dst_rtype = _RAND_900[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{$random}};
  _T_5936_24_fp_val = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{$random}};
  _T_5936_25_br_mask = _RAND_902[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{$random}};
  _T_5936_25_pdst = _RAND_903[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{$random}};
  _T_5936_25_stale_pdst = _RAND_904[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{$random}};
  _T_5936_25_is_fencei = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{$random}};
  _T_5936_25_is_store = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{$random}};
  _T_5936_25_is_load = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{$random}};
  _T_5936_25_is_sys_pc2epc = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{$random}};
  _T_5936_25_flush_on_commit = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{$random}};
  _T_5936_25_ldst = _RAND_910[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{$random}};
  _T_5936_25_ldst_val = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{$random}};
  _T_5936_25_dst_rtype = _RAND_912[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{$random}};
  _T_5936_25_fp_val = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{$random}};
  _T_5936_26_br_mask = _RAND_914[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{$random}};
  _T_5936_26_pdst = _RAND_915[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{$random}};
  _T_5936_26_stale_pdst = _RAND_916[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{$random}};
  _T_5936_26_is_fencei = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{$random}};
  _T_5936_26_is_store = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{$random}};
  _T_5936_26_is_load = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{$random}};
  _T_5936_26_is_sys_pc2epc = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{$random}};
  _T_5936_26_flush_on_commit = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{$random}};
  _T_5936_26_ldst = _RAND_922[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{$random}};
  _T_5936_26_ldst_val = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{$random}};
  _T_5936_26_dst_rtype = _RAND_924[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{$random}};
  _T_5936_26_fp_val = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{$random}};
  _T_5936_27_br_mask = _RAND_926[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{$random}};
  _T_5936_27_pdst = _RAND_927[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{$random}};
  _T_5936_27_stale_pdst = _RAND_928[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{$random}};
  _T_5936_27_is_fencei = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{$random}};
  _T_5936_27_is_store = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{$random}};
  _T_5936_27_is_load = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{$random}};
  _T_5936_27_is_sys_pc2epc = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{$random}};
  _T_5936_27_flush_on_commit = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{$random}};
  _T_5936_27_ldst = _RAND_934[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{$random}};
  _T_5936_27_ldst_val = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{$random}};
  _T_5936_27_dst_rtype = _RAND_936[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{$random}};
  _T_5936_27_fp_val = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{$random}};
  _T_5936_28_br_mask = _RAND_938[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{$random}};
  _T_5936_28_pdst = _RAND_939[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{$random}};
  _T_5936_28_stale_pdst = _RAND_940[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{$random}};
  _T_5936_28_is_fencei = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{$random}};
  _T_5936_28_is_store = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{$random}};
  _T_5936_28_is_load = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{$random}};
  _T_5936_28_is_sys_pc2epc = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{$random}};
  _T_5936_28_flush_on_commit = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{$random}};
  _T_5936_28_ldst = _RAND_946[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{$random}};
  _T_5936_28_ldst_val = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{$random}};
  _T_5936_28_dst_rtype = _RAND_948[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{$random}};
  _T_5936_28_fp_val = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{$random}};
  _T_5936_29_br_mask = _RAND_950[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{$random}};
  _T_5936_29_pdst = _RAND_951[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{$random}};
  _T_5936_29_stale_pdst = _RAND_952[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{$random}};
  _T_5936_29_is_fencei = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{$random}};
  _T_5936_29_is_store = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{$random}};
  _T_5936_29_is_load = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{$random}};
  _T_5936_29_is_sys_pc2epc = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{$random}};
  _T_5936_29_flush_on_commit = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{$random}};
  _T_5936_29_ldst = _RAND_958[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{$random}};
  _T_5936_29_ldst_val = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{$random}};
  _T_5936_29_dst_rtype = _RAND_960[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{$random}};
  _T_5936_29_fp_val = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{$random}};
  _T_5936_30_br_mask = _RAND_962[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{$random}};
  _T_5936_30_pdst = _RAND_963[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{$random}};
  _T_5936_30_stale_pdst = _RAND_964[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{$random}};
  _T_5936_30_is_fencei = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{$random}};
  _T_5936_30_is_store = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{$random}};
  _T_5936_30_is_load = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{$random}};
  _T_5936_30_is_sys_pc2epc = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{$random}};
  _T_5936_30_flush_on_commit = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{$random}};
  _T_5936_30_ldst = _RAND_970[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{$random}};
  _T_5936_30_ldst_val = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{$random}};
  _T_5936_30_dst_rtype = _RAND_972[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{$random}};
  _T_5936_30_fp_val = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{$random}};
  _T_5936_31_br_mask = _RAND_974[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{$random}};
  _T_5936_31_pdst = _RAND_975[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{$random}};
  _T_5936_31_stale_pdst = _RAND_976[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{$random}};
  _T_5936_31_is_fencei = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{$random}};
  _T_5936_31_is_store = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{$random}};
  _T_5936_31_is_load = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{$random}};
  _T_5936_31_is_sys_pc2epc = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{$random}};
  _T_5936_31_flush_on_commit = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{$random}};
  _T_5936_31_ldst = _RAND_982[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{$random}};
  _T_5936_31_ldst_val = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{$random}};
  _T_5936_31_dst_rtype = _RAND_984[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{$random}};
  _T_5936_31_fp_val = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{$random}};
  _T_5936_32_br_mask = _RAND_986[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{$random}};
  _T_5936_32_pdst = _RAND_987[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{$random}};
  _T_5936_32_stale_pdst = _RAND_988[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{$random}};
  _T_5936_32_is_fencei = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{$random}};
  _T_5936_32_is_store = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{$random}};
  _T_5936_32_is_load = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{$random}};
  _T_5936_32_is_sys_pc2epc = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{$random}};
  _T_5936_32_flush_on_commit = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{$random}};
  _T_5936_32_ldst = _RAND_994[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{$random}};
  _T_5936_32_ldst_val = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{$random}};
  _T_5936_32_dst_rtype = _RAND_996[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{$random}};
  _T_5936_32_fp_val = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{$random}};
  _T_5936_33_br_mask = _RAND_998[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{$random}};
  _T_5936_33_pdst = _RAND_999[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{$random}};
  _T_5936_33_stale_pdst = _RAND_1000[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{$random}};
  _T_5936_33_is_fencei = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{$random}};
  _T_5936_33_is_store = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{$random}};
  _T_5936_33_is_load = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{$random}};
  _T_5936_33_is_sys_pc2epc = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{$random}};
  _T_5936_33_flush_on_commit = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{$random}};
  _T_5936_33_ldst = _RAND_1006[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{$random}};
  _T_5936_33_ldst_val = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{$random}};
  _T_5936_33_dst_rtype = _RAND_1008[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{$random}};
  _T_5936_33_fp_val = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{$random}};
  _T_5936_34_br_mask = _RAND_1010[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{$random}};
  _T_5936_34_pdst = _RAND_1011[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{$random}};
  _T_5936_34_stale_pdst = _RAND_1012[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{$random}};
  _T_5936_34_is_fencei = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{$random}};
  _T_5936_34_is_store = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{$random}};
  _T_5936_34_is_load = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{$random}};
  _T_5936_34_is_sys_pc2epc = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{$random}};
  _T_5936_34_flush_on_commit = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{$random}};
  _T_5936_34_ldst = _RAND_1018[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{$random}};
  _T_5936_34_ldst_val = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{$random}};
  _T_5936_34_dst_rtype = _RAND_1020[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{$random}};
  _T_5936_34_fp_val = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{$random}};
  _T_5936_35_br_mask = _RAND_1022[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{$random}};
  _T_5936_35_pdst = _RAND_1023[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{$random}};
  _T_5936_35_stale_pdst = _RAND_1024[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{$random}};
  _T_5936_35_is_fencei = _RAND_1025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{$random}};
  _T_5936_35_is_store = _RAND_1026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{$random}};
  _T_5936_35_is_load = _RAND_1027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{$random}};
  _T_5936_35_is_sys_pc2epc = _RAND_1028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{$random}};
  _T_5936_35_flush_on_commit = _RAND_1029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{$random}};
  _T_5936_35_ldst = _RAND_1030[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{$random}};
  _T_5936_35_ldst_val = _RAND_1031[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{$random}};
  _T_5936_35_dst_rtype = _RAND_1032[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{$random}};
  _T_5936_35_fp_val = _RAND_1033[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{$random}};
  _T_5936_36_br_mask = _RAND_1034[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{$random}};
  _T_5936_36_pdst = _RAND_1035[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{$random}};
  _T_5936_36_stale_pdst = _RAND_1036[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{$random}};
  _T_5936_36_is_fencei = _RAND_1037[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{$random}};
  _T_5936_36_is_store = _RAND_1038[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{$random}};
  _T_5936_36_is_load = _RAND_1039[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{$random}};
  _T_5936_36_is_sys_pc2epc = _RAND_1040[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{$random}};
  _T_5936_36_flush_on_commit = _RAND_1041[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{$random}};
  _T_5936_36_ldst = _RAND_1042[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{$random}};
  _T_5936_36_ldst_val = _RAND_1043[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{$random}};
  _T_5936_36_dst_rtype = _RAND_1044[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{$random}};
  _T_5936_36_fp_val = _RAND_1045[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{$random}};
  _T_5936_37_br_mask = _RAND_1046[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{$random}};
  _T_5936_37_pdst = _RAND_1047[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{$random}};
  _T_5936_37_stale_pdst = _RAND_1048[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{$random}};
  _T_5936_37_is_fencei = _RAND_1049[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{$random}};
  _T_5936_37_is_store = _RAND_1050[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{$random}};
  _T_5936_37_is_load = _RAND_1051[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{$random}};
  _T_5936_37_is_sys_pc2epc = _RAND_1052[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{$random}};
  _T_5936_37_flush_on_commit = _RAND_1053[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{$random}};
  _T_5936_37_ldst = _RAND_1054[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{$random}};
  _T_5936_37_ldst_val = _RAND_1055[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{$random}};
  _T_5936_37_dst_rtype = _RAND_1056[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{$random}};
  _T_5936_37_fp_val = _RAND_1057[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{$random}};
  _T_5936_38_br_mask = _RAND_1058[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{$random}};
  _T_5936_38_pdst = _RAND_1059[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{$random}};
  _T_5936_38_stale_pdst = _RAND_1060[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{$random}};
  _T_5936_38_is_fencei = _RAND_1061[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{$random}};
  _T_5936_38_is_store = _RAND_1062[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{$random}};
  _T_5936_38_is_load = _RAND_1063[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{$random}};
  _T_5936_38_is_sys_pc2epc = _RAND_1064[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{$random}};
  _T_5936_38_flush_on_commit = _RAND_1065[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{$random}};
  _T_5936_38_ldst = _RAND_1066[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{$random}};
  _T_5936_38_ldst_val = _RAND_1067[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{$random}};
  _T_5936_38_dst_rtype = _RAND_1068[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{$random}};
  _T_5936_38_fp_val = _RAND_1069[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{$random}};
  _T_5936_39_br_mask = _RAND_1070[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{$random}};
  _T_5936_39_pdst = _RAND_1071[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{$random}};
  _T_5936_39_stale_pdst = _RAND_1072[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{$random}};
  _T_5936_39_is_fencei = _RAND_1073[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{$random}};
  _T_5936_39_is_store = _RAND_1074[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{$random}};
  _T_5936_39_is_load = _RAND_1075[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{$random}};
  _T_5936_39_is_sys_pc2epc = _RAND_1076[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{$random}};
  _T_5936_39_flush_on_commit = _RAND_1077[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{$random}};
  _T_5936_39_ldst = _RAND_1078[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{$random}};
  _T_5936_39_ldst_val = _RAND_1079[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{$random}};
  _T_5936_39_dst_rtype = _RAND_1080[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{$random}};
  _T_5936_39_fp_val = _RAND_1081[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_1082 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_6309[initvar] = _RAND_1082[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1083 = {1{$random}};
  _RAND_1084 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 40; initvar = initvar+1)
    _T_6312[initvar] = _RAND_1084[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1085 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{$random}};
  _T_8115 = _RAND_1086[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {2{$random}};
  _T_8120 = _RAND_1087[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{$random}};
  com_lsu_misspec = _RAND_1088[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      rob_state <= 2'h0;
    end else begin
      if (_T_8411) begin
        if (exception_thrown) begin
          rob_state <= 2'h2;
        end else begin
          if (io_empty) begin
            rob_state <= 2'h1;
          end else begin
            if (_T_8410) begin
              if (io_empty) begin
                rob_state <= 2'h1;
              end else begin
                if (_T_8407) begin
                  if (exception_thrown) begin
                    rob_state <= 2'h2;
                  end else begin
                    if (_T_2902) begin
                      rob_state <= 2'h3;
                    end else begin
                      if (_T_2901) begin
                        rob_state <= 2'h3;
                      end else begin
                        if (_T_8406) begin
                          rob_state <= 2'h1;
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_8406) begin
                    rob_state <= 2'h1;
                  end
                end
              end
            end else begin
              if (_T_8407) begin
                if (exception_thrown) begin
                  rob_state <= 2'h2;
                end else begin
                  if (_T_2902) begin
                    rob_state <= 2'h3;
                  end else begin
                    if (_T_2901) begin
                      rob_state <= 2'h3;
                    end else begin
                      if (_T_8406) begin
                        rob_state <= 2'h1;
                      end
                    end
                  end
                end
              end else begin
                if (_T_8406) begin
                  rob_state <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_8410) begin
          if (io_empty) begin
            rob_state <= 2'h1;
          end else begin
            if (_T_8407) begin
              if (exception_thrown) begin
                rob_state <= 2'h2;
              end else begin
                if (_T_2902) begin
                  rob_state <= 2'h3;
                end else begin
                  if (_T_2901) begin
                    rob_state <= 2'h3;
                  end else begin
                    rob_state <= _GEN_82632;
                  end
                end
              end
            end else begin
              rob_state <= _GEN_82632;
            end
          end
        end else begin
          if (_T_8407) begin
            if (exception_thrown) begin
              rob_state <= 2'h2;
            end else begin
              if (_T_2902) begin
                rob_state <= 2'h3;
              end else begin
                if (_T_2901) begin
                  rob_state <= 2'h3;
                end else begin
                  rob_state <= _GEN_82632;
                end
              end
            end
          end else begin
            rob_state <= _GEN_82632;
          end
        end
      end
    end
    if (reset) begin
      rob_head <= 6'h0;
    end else begin
      if (finished_committing_row) begin
        if (_T_8350) begin
          rob_head <= 6'h0;
        end else begin
          rob_head <= _T_8354;
        end
      end
    end
    if (reset) begin
      rob_tail <= 6'h0;
    end else begin
      rob_tail <= _GEN_82631[5:0];
    end
    if (reset) begin
      r_xcpt_val <= 1'h0;
    end else begin
      if (_T_8304) begin
        r_xcpt_val <= 1'h0;
      end else begin
        if (_T_8233) begin
          if (_T_8234) begin
            if (_T_8258) begin
              r_xcpt_val <= 1'h1;
            end
          end else begin
            if (_T_8265) begin
              r_xcpt_val <= 1'h1;
            end
          end
        end
      end
    end
    if (io_brinfo_valid) begin
      r_xcpt_uop_br_mask <= _T_8297;
    end else begin
      r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask;
    end
    r_xcpt_uop_rob_idx <= next_xcpt_uop_rob_idx;
    r_xcpt_uop_exc_cause <= next_xcpt_uop_exc_cause;
    if (_T_8233) begin
      if (_T_8234) begin
        if (_T_8258) begin
          r_xcpt_badvaddr <= {{24'd0}, _T_8261};
        end
      end else begin
        if (_T_8265) begin
          r_xcpt_badvaddr <= {{24'd0}, _T_8295};
        end
      end
    end
    if(_T_2772__T_2788_en & _T_2772__T_2788_mask) begin
      _T_2772[_T_2772__T_2788_addr] <= _T_2772__T_2788_data;
    end
    if(_T_2775__T_2784_en & _T_2775__T_2784_mask) begin
      _T_2775[_T_2775__T_2784_addr] <= _T_2775__T_2784_data;
    end
    if (reset) begin
      r_partial_row <= 1'h0;
    end else begin
      if (_T_2885) begin
        r_partial_row <= io_enq_partial_stall;
      end else begin
        if (_T_2891) begin
          r_partial_row <= io_enq_partial_stall;
        end
      end
    end
    if(row_metadata_brob_idx__T_2886_en & row_metadata_brob_idx__T_2886_mask) begin
      row_metadata_brob_idx[row_metadata_brob_idx__T_2886_addr] <= row_metadata_brob_idx__T_2886_data;
    end
    if(row_metadata_has_brorjalr__T_2887_en & row_metadata_has_brorjalr__T_2887_mask) begin
      row_metadata_has_brorjalr[row_metadata_has_brorjalr__T_2887_addr] <= row_metadata_has_brorjalr__T_2887_data;
    end
    if(row_metadata_has_brorjalr__T_2892_en & row_metadata_has_brorjalr__T_2892_mask) begin
      row_metadata_has_brorjalr[row_metadata_has_brorjalr__T_2892_addr] <= row_metadata_has_brorjalr__T_2892_data;
    end
    if (reset) begin
      _T_3073_0 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h0 == rob_head) begin
          _T_3073_0 <= 1'h0;
        end else begin
          if (_T_4095) begin
            _T_3073_0 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h0 == _T_4025) begin
                _T_3073_0 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h0 == rob_tail) begin
                    _T_3073_0 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h0 == rob_tail) begin
                  _T_3073_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4095) begin
          _T_3073_0 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h0 == _T_4025) begin
              _T_3073_0 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h0 == rob_tail) begin
                  _T_3073_0 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h0 == rob_tail) begin
                _T_3073_0 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_1 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1 == rob_head) begin
          _T_3073_1 <= 1'h0;
        end else begin
          if (_T_4118) begin
            _T_3073_1 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1 == _T_4025) begin
                _T_3073_1 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1 == rob_tail) begin
                    _T_3073_1 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1 == rob_tail) begin
                  _T_3073_1 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4118) begin
          _T_3073_1 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1 == _T_4025) begin
              _T_3073_1 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1 == rob_tail) begin
                  _T_3073_1 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1 == rob_tail) begin
                _T_3073_1 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_2 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h2 == rob_head) begin
          _T_3073_2 <= 1'h0;
        end else begin
          if (_T_4141) begin
            _T_3073_2 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h2 == _T_4025) begin
                _T_3073_2 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h2 == rob_tail) begin
                    _T_3073_2 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h2 == rob_tail) begin
                  _T_3073_2 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4141) begin
          _T_3073_2 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h2 == _T_4025) begin
              _T_3073_2 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h2 == rob_tail) begin
                  _T_3073_2 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h2 == rob_tail) begin
                _T_3073_2 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_3 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h3 == rob_head) begin
          _T_3073_3 <= 1'h0;
        end else begin
          if (_T_4164) begin
            _T_3073_3 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h3 == _T_4025) begin
                _T_3073_3 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h3 == rob_tail) begin
                    _T_3073_3 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h3 == rob_tail) begin
                  _T_3073_3 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4164) begin
          _T_3073_3 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h3 == _T_4025) begin
              _T_3073_3 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h3 == rob_tail) begin
                  _T_3073_3 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h3 == rob_tail) begin
                _T_3073_3 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_4 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h4 == rob_head) begin
          _T_3073_4 <= 1'h0;
        end else begin
          if (_T_4187) begin
            _T_3073_4 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h4 == _T_4025) begin
                _T_3073_4 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h4 == rob_tail) begin
                    _T_3073_4 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h4 == rob_tail) begin
                  _T_3073_4 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4187) begin
          _T_3073_4 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h4 == _T_4025) begin
              _T_3073_4 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h4 == rob_tail) begin
                  _T_3073_4 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h4 == rob_tail) begin
                _T_3073_4 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_5 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h5 == rob_head) begin
          _T_3073_5 <= 1'h0;
        end else begin
          if (_T_4210) begin
            _T_3073_5 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h5 == _T_4025) begin
                _T_3073_5 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h5 == rob_tail) begin
                    _T_3073_5 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h5 == rob_tail) begin
                  _T_3073_5 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4210) begin
          _T_3073_5 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h5 == _T_4025) begin
              _T_3073_5 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h5 == rob_tail) begin
                  _T_3073_5 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h5 == rob_tail) begin
                _T_3073_5 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_6 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h6 == rob_head) begin
          _T_3073_6 <= 1'h0;
        end else begin
          if (_T_4233) begin
            _T_3073_6 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h6 == _T_4025) begin
                _T_3073_6 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h6 == rob_tail) begin
                    _T_3073_6 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h6 == rob_tail) begin
                  _T_3073_6 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4233) begin
          _T_3073_6 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h6 == _T_4025) begin
              _T_3073_6 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h6 == rob_tail) begin
                  _T_3073_6 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h6 == rob_tail) begin
                _T_3073_6 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_7 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h7 == rob_head) begin
          _T_3073_7 <= 1'h0;
        end else begin
          if (_T_4256) begin
            _T_3073_7 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h7 == _T_4025) begin
                _T_3073_7 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h7 == rob_tail) begin
                    _T_3073_7 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h7 == rob_tail) begin
                  _T_3073_7 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4256) begin
          _T_3073_7 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h7 == _T_4025) begin
              _T_3073_7 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h7 == rob_tail) begin
                  _T_3073_7 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h7 == rob_tail) begin
                _T_3073_7 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_8 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h8 == rob_head) begin
          _T_3073_8 <= 1'h0;
        end else begin
          if (_T_4279) begin
            _T_3073_8 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h8 == _T_4025) begin
                _T_3073_8 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h8 == rob_tail) begin
                    _T_3073_8 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h8 == rob_tail) begin
                  _T_3073_8 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4279) begin
          _T_3073_8 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h8 == _T_4025) begin
              _T_3073_8 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h8 == rob_tail) begin
                  _T_3073_8 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h8 == rob_tail) begin
                _T_3073_8 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_9 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h9 == rob_head) begin
          _T_3073_9 <= 1'h0;
        end else begin
          if (_T_4302) begin
            _T_3073_9 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h9 == _T_4025) begin
                _T_3073_9 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h9 == rob_tail) begin
                    _T_3073_9 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h9 == rob_tail) begin
                  _T_3073_9 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4302) begin
          _T_3073_9 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h9 == _T_4025) begin
              _T_3073_9 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h9 == rob_tail) begin
                  _T_3073_9 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h9 == rob_tail) begin
                _T_3073_9 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_10 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'ha == rob_head) begin
          _T_3073_10 <= 1'h0;
        end else begin
          if (_T_4325) begin
            _T_3073_10 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'ha == _T_4025) begin
                _T_3073_10 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'ha == rob_tail) begin
                    _T_3073_10 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'ha == rob_tail) begin
                  _T_3073_10 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4325) begin
          _T_3073_10 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'ha == _T_4025) begin
              _T_3073_10 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'ha == rob_tail) begin
                  _T_3073_10 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'ha == rob_tail) begin
                _T_3073_10 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_11 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'hb == rob_head) begin
          _T_3073_11 <= 1'h0;
        end else begin
          if (_T_4348) begin
            _T_3073_11 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hb == _T_4025) begin
                _T_3073_11 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'hb == rob_tail) begin
                    _T_3073_11 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'hb == rob_tail) begin
                  _T_3073_11 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4348) begin
          _T_3073_11 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hb == _T_4025) begin
              _T_3073_11 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'hb == rob_tail) begin
                  _T_3073_11 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'hb == rob_tail) begin
                _T_3073_11 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_12 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'hc == rob_head) begin
          _T_3073_12 <= 1'h0;
        end else begin
          if (_T_4371) begin
            _T_3073_12 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hc == _T_4025) begin
                _T_3073_12 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'hc == rob_tail) begin
                    _T_3073_12 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'hc == rob_tail) begin
                  _T_3073_12 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4371) begin
          _T_3073_12 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hc == _T_4025) begin
              _T_3073_12 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'hc == rob_tail) begin
                  _T_3073_12 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'hc == rob_tail) begin
                _T_3073_12 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_13 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'hd == rob_head) begin
          _T_3073_13 <= 1'h0;
        end else begin
          if (_T_4394) begin
            _T_3073_13 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hd == _T_4025) begin
                _T_3073_13 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'hd == rob_tail) begin
                    _T_3073_13 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'hd == rob_tail) begin
                  _T_3073_13 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4394) begin
          _T_3073_13 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hd == _T_4025) begin
              _T_3073_13 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'hd == rob_tail) begin
                  _T_3073_13 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'hd == rob_tail) begin
                _T_3073_13 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_14 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'he == rob_head) begin
          _T_3073_14 <= 1'h0;
        end else begin
          if (_T_4417) begin
            _T_3073_14 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'he == _T_4025) begin
                _T_3073_14 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'he == rob_tail) begin
                    _T_3073_14 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'he == rob_tail) begin
                  _T_3073_14 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4417) begin
          _T_3073_14 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'he == _T_4025) begin
              _T_3073_14 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'he == rob_tail) begin
                  _T_3073_14 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'he == rob_tail) begin
                _T_3073_14 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_15 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'hf == rob_head) begin
          _T_3073_15 <= 1'h0;
        end else begin
          if (_T_4440) begin
            _T_3073_15 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hf == _T_4025) begin
                _T_3073_15 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'hf == rob_tail) begin
                    _T_3073_15 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'hf == rob_tail) begin
                  _T_3073_15 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4440) begin
          _T_3073_15 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hf == _T_4025) begin
              _T_3073_15 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'hf == rob_tail) begin
                  _T_3073_15 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'hf == rob_tail) begin
                _T_3073_15 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_16 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h10 == rob_head) begin
          _T_3073_16 <= 1'h0;
        end else begin
          if (_T_4463) begin
            _T_3073_16 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h10 == _T_4025) begin
                _T_3073_16 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h10 == rob_tail) begin
                    _T_3073_16 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h10 == rob_tail) begin
                  _T_3073_16 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4463) begin
          _T_3073_16 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h10 == _T_4025) begin
              _T_3073_16 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h10 == rob_tail) begin
                  _T_3073_16 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h10 == rob_tail) begin
                _T_3073_16 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_17 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h11 == rob_head) begin
          _T_3073_17 <= 1'h0;
        end else begin
          if (_T_4486) begin
            _T_3073_17 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h11 == _T_4025) begin
                _T_3073_17 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h11 == rob_tail) begin
                    _T_3073_17 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h11 == rob_tail) begin
                  _T_3073_17 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4486) begin
          _T_3073_17 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h11 == _T_4025) begin
              _T_3073_17 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h11 == rob_tail) begin
                  _T_3073_17 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h11 == rob_tail) begin
                _T_3073_17 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_18 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h12 == rob_head) begin
          _T_3073_18 <= 1'h0;
        end else begin
          if (_T_4509) begin
            _T_3073_18 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h12 == _T_4025) begin
                _T_3073_18 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h12 == rob_tail) begin
                    _T_3073_18 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h12 == rob_tail) begin
                  _T_3073_18 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4509) begin
          _T_3073_18 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h12 == _T_4025) begin
              _T_3073_18 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h12 == rob_tail) begin
                  _T_3073_18 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h12 == rob_tail) begin
                _T_3073_18 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_19 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h13 == rob_head) begin
          _T_3073_19 <= 1'h0;
        end else begin
          if (_T_4532) begin
            _T_3073_19 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h13 == _T_4025) begin
                _T_3073_19 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h13 == rob_tail) begin
                    _T_3073_19 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h13 == rob_tail) begin
                  _T_3073_19 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4532) begin
          _T_3073_19 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h13 == _T_4025) begin
              _T_3073_19 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h13 == rob_tail) begin
                  _T_3073_19 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h13 == rob_tail) begin
                _T_3073_19 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_20 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h14 == rob_head) begin
          _T_3073_20 <= 1'h0;
        end else begin
          if (_T_4555) begin
            _T_3073_20 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h14 == _T_4025) begin
                _T_3073_20 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h14 == rob_tail) begin
                    _T_3073_20 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h14 == rob_tail) begin
                  _T_3073_20 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4555) begin
          _T_3073_20 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h14 == _T_4025) begin
              _T_3073_20 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h14 == rob_tail) begin
                  _T_3073_20 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h14 == rob_tail) begin
                _T_3073_20 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_21 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h15 == rob_head) begin
          _T_3073_21 <= 1'h0;
        end else begin
          if (_T_4578) begin
            _T_3073_21 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h15 == _T_4025) begin
                _T_3073_21 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h15 == rob_tail) begin
                    _T_3073_21 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h15 == rob_tail) begin
                  _T_3073_21 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4578) begin
          _T_3073_21 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h15 == _T_4025) begin
              _T_3073_21 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h15 == rob_tail) begin
                  _T_3073_21 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h15 == rob_tail) begin
                _T_3073_21 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_22 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h16 == rob_head) begin
          _T_3073_22 <= 1'h0;
        end else begin
          if (_T_4601) begin
            _T_3073_22 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h16 == _T_4025) begin
                _T_3073_22 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h16 == rob_tail) begin
                    _T_3073_22 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h16 == rob_tail) begin
                  _T_3073_22 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4601) begin
          _T_3073_22 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h16 == _T_4025) begin
              _T_3073_22 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h16 == rob_tail) begin
                  _T_3073_22 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h16 == rob_tail) begin
                _T_3073_22 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_23 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h17 == rob_head) begin
          _T_3073_23 <= 1'h0;
        end else begin
          if (_T_4624) begin
            _T_3073_23 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h17 == _T_4025) begin
                _T_3073_23 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h17 == rob_tail) begin
                    _T_3073_23 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h17 == rob_tail) begin
                  _T_3073_23 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4624) begin
          _T_3073_23 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h17 == _T_4025) begin
              _T_3073_23 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h17 == rob_tail) begin
                  _T_3073_23 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h17 == rob_tail) begin
                _T_3073_23 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_24 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h18 == rob_head) begin
          _T_3073_24 <= 1'h0;
        end else begin
          if (_T_4647) begin
            _T_3073_24 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h18 == _T_4025) begin
                _T_3073_24 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h18 == rob_tail) begin
                    _T_3073_24 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h18 == rob_tail) begin
                  _T_3073_24 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4647) begin
          _T_3073_24 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h18 == _T_4025) begin
              _T_3073_24 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h18 == rob_tail) begin
                  _T_3073_24 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h18 == rob_tail) begin
                _T_3073_24 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_25 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h19 == rob_head) begin
          _T_3073_25 <= 1'h0;
        end else begin
          if (_T_4670) begin
            _T_3073_25 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h19 == _T_4025) begin
                _T_3073_25 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h19 == rob_tail) begin
                    _T_3073_25 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h19 == rob_tail) begin
                  _T_3073_25 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4670) begin
          _T_3073_25 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h19 == _T_4025) begin
              _T_3073_25 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h19 == rob_tail) begin
                  _T_3073_25 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h19 == rob_tail) begin
                _T_3073_25 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_26 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1a == rob_head) begin
          _T_3073_26 <= 1'h0;
        end else begin
          if (_T_4693) begin
            _T_3073_26 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1a == _T_4025) begin
                _T_3073_26 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1a == rob_tail) begin
                    _T_3073_26 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1a == rob_tail) begin
                  _T_3073_26 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4693) begin
          _T_3073_26 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1a == _T_4025) begin
              _T_3073_26 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1a == rob_tail) begin
                  _T_3073_26 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1a == rob_tail) begin
                _T_3073_26 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_27 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1b == rob_head) begin
          _T_3073_27 <= 1'h0;
        end else begin
          if (_T_4716) begin
            _T_3073_27 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1b == _T_4025) begin
                _T_3073_27 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1b == rob_tail) begin
                    _T_3073_27 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1b == rob_tail) begin
                  _T_3073_27 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4716) begin
          _T_3073_27 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1b == _T_4025) begin
              _T_3073_27 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1b == rob_tail) begin
                  _T_3073_27 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1b == rob_tail) begin
                _T_3073_27 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_28 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1c == rob_head) begin
          _T_3073_28 <= 1'h0;
        end else begin
          if (_T_4739) begin
            _T_3073_28 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1c == _T_4025) begin
                _T_3073_28 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1c == rob_tail) begin
                    _T_3073_28 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1c == rob_tail) begin
                  _T_3073_28 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4739) begin
          _T_3073_28 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1c == _T_4025) begin
              _T_3073_28 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1c == rob_tail) begin
                  _T_3073_28 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1c == rob_tail) begin
                _T_3073_28 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_29 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1d == rob_head) begin
          _T_3073_29 <= 1'h0;
        end else begin
          if (_T_4762) begin
            _T_3073_29 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1d == _T_4025) begin
                _T_3073_29 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1d == rob_tail) begin
                    _T_3073_29 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1d == rob_tail) begin
                  _T_3073_29 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4762) begin
          _T_3073_29 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1d == _T_4025) begin
              _T_3073_29 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1d == rob_tail) begin
                  _T_3073_29 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1d == rob_tail) begin
                _T_3073_29 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_30 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1e == rob_head) begin
          _T_3073_30 <= 1'h0;
        end else begin
          if (_T_4785) begin
            _T_3073_30 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1e == _T_4025) begin
                _T_3073_30 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1e == rob_tail) begin
                    _T_3073_30 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1e == rob_tail) begin
                  _T_3073_30 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4785) begin
          _T_3073_30 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1e == _T_4025) begin
              _T_3073_30 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1e == rob_tail) begin
                  _T_3073_30 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1e == rob_tail) begin
                _T_3073_30 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_31 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h1f == rob_head) begin
          _T_3073_31 <= 1'h0;
        end else begin
          if (_T_4808) begin
            _T_3073_31 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1f == _T_4025) begin
                _T_3073_31 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h1f == rob_tail) begin
                    _T_3073_31 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1f == rob_tail) begin
                  _T_3073_31 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4808) begin
          _T_3073_31 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1f == _T_4025) begin
              _T_3073_31 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h1f == rob_tail) begin
                  _T_3073_31 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h1f == rob_tail) begin
                _T_3073_31 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_32 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h20 == rob_head) begin
          _T_3073_32 <= 1'h0;
        end else begin
          if (_T_4831) begin
            _T_3073_32 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h20 == _T_4025) begin
                _T_3073_32 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h20 == rob_tail) begin
                    _T_3073_32 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h20 == rob_tail) begin
                  _T_3073_32 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4831) begin
          _T_3073_32 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h20 == _T_4025) begin
              _T_3073_32 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h20 == rob_tail) begin
                  _T_3073_32 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h20 == rob_tail) begin
                _T_3073_32 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_33 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h21 == rob_head) begin
          _T_3073_33 <= 1'h0;
        end else begin
          if (_T_4854) begin
            _T_3073_33 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h21 == _T_4025) begin
                _T_3073_33 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h21 == rob_tail) begin
                    _T_3073_33 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h21 == rob_tail) begin
                  _T_3073_33 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4854) begin
          _T_3073_33 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h21 == _T_4025) begin
              _T_3073_33 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h21 == rob_tail) begin
                  _T_3073_33 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h21 == rob_tail) begin
                _T_3073_33 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_34 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h22 == rob_head) begin
          _T_3073_34 <= 1'h0;
        end else begin
          if (_T_4877) begin
            _T_3073_34 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h22 == _T_4025) begin
                _T_3073_34 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h22 == rob_tail) begin
                    _T_3073_34 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h22 == rob_tail) begin
                  _T_3073_34 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4877) begin
          _T_3073_34 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h22 == _T_4025) begin
              _T_3073_34 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h22 == rob_tail) begin
                  _T_3073_34 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h22 == rob_tail) begin
                _T_3073_34 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_35 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h23 == rob_head) begin
          _T_3073_35 <= 1'h0;
        end else begin
          if (_T_4900) begin
            _T_3073_35 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h23 == _T_4025) begin
                _T_3073_35 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h23 == rob_tail) begin
                    _T_3073_35 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h23 == rob_tail) begin
                  _T_3073_35 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4900) begin
          _T_3073_35 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h23 == _T_4025) begin
              _T_3073_35 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h23 == rob_tail) begin
                  _T_3073_35 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h23 == rob_tail) begin
                _T_3073_35 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_36 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h24 == rob_head) begin
          _T_3073_36 <= 1'h0;
        end else begin
          if (_T_4923) begin
            _T_3073_36 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h24 == _T_4025) begin
                _T_3073_36 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h24 == rob_tail) begin
                    _T_3073_36 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h24 == rob_tail) begin
                  _T_3073_36 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4923) begin
          _T_3073_36 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h24 == _T_4025) begin
              _T_3073_36 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h24 == rob_tail) begin
                  _T_3073_36 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h24 == rob_tail) begin
                _T_3073_36 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_37 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h25 == rob_head) begin
          _T_3073_37 <= 1'h0;
        end else begin
          if (_T_4946) begin
            _T_3073_37 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h25 == _T_4025) begin
                _T_3073_37 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h25 == rob_tail) begin
                    _T_3073_37 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h25 == rob_tail) begin
                  _T_3073_37 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4946) begin
          _T_3073_37 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h25 == _T_4025) begin
              _T_3073_37 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h25 == rob_tail) begin
                  _T_3073_37 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h25 == rob_tail) begin
                _T_3073_37 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_38 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h26 == rob_head) begin
          _T_3073_38 <= 1'h0;
        end else begin
          if (_T_4969) begin
            _T_3073_38 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h26 == _T_4025) begin
                _T_3073_38 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h26 == rob_tail) begin
                    _T_3073_38 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h26 == rob_tail) begin
                  _T_3073_38 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4969) begin
          _T_3073_38 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h26 == _T_4025) begin
              _T_3073_38 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h26 == rob_tail) begin
                  _T_3073_38 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h26 == rob_tail) begin
                _T_3073_38 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_3073_39 <= 1'h0;
    end else begin
      if (will_commit_0) begin
        if (6'h27 == rob_head) begin
          _T_3073_39 <= 1'h0;
        end else begin
          if (_T_4992) begin
            _T_3073_39 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h27 == _T_4025) begin
                _T_3073_39 <= 1'h0;
              end else begin
                if (io_enq_valids_0) begin
                  if (6'h27 == rob_tail) begin
                    _T_3073_39 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_0) begin
                if (6'h27 == rob_tail) begin
                  _T_3073_39 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_4992) begin
          _T_3073_39 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h27 == _T_4025) begin
              _T_3073_39 <= 1'h0;
            end else begin
              if (io_enq_valids_0) begin
                if (6'h27 == rob_tail) begin
                  _T_3073_39 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_0) begin
              if (6'h27 == rob_tail) begin
                _T_3073_39 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if(_T_3200__T_3753_en & _T_3200__T_3753_mask) begin
      _T_3200[_T_3200__T_3753_addr] <= _T_3200__T_3753_data;
    end
    if(_T_3200__T_3819_en & _T_3200__T_3819_mask) begin
      _T_3200[_T_3200__T_3819_addr] <= _T_3200__T_3819_data;
    end
    if(_T_3200__T_3828_en & _T_3200__T_3828_mask) begin
      _T_3200[_T_3200__T_3828_addr] <= _T_3200__T_3828_data;
    end
    if(_T_3200__T_3837_en & _T_3200__T_3837_mask) begin
      _T_3200[_T_3200__T_3837_addr] <= _T_3200__T_3837_data;
    end
    if(_T_3200__T_3846_en & _T_3200__T_3846_mask) begin
      _T_3200[_T_3200__T_3846_addr] <= _T_3200__T_3846_data;
    end
    if(_T_3200__T_3855_en & _T_3200__T_3855_mask) begin
      _T_3200[_T_3200__T_3855_addr] <= _T_3200__T_3855_data;
    end
    if(_T_3200__T_3864_en & _T_3200__T_3864_mask) begin
      _T_3200[_T_3200__T_3864_addr] <= _T_3200__T_3864_data;
    end
    if(_T_3200__T_3891_en & _T_3200__T_3891_mask) begin
      _T_3200[_T_3200__T_3891_addr] <= _T_3200__T_3891_data;
    end
    if (_T_4095) begin
      if (io_enq_valids_0) begin
        if (6'h0 == rob_tail) begin
          _T_3372_0_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4110) begin
        _T_3372_0_br_mask <= _T_4112;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h0 == rob_tail) begin
            _T_3372_0_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h0 == rob_tail) begin
        _T_3372_0_fp_val <= _GEN_84;
      end
    end
    if (_T_4118) begin
      if (io_enq_valids_0) begin
        if (6'h1 == rob_tail) begin
          _T_3372_1_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4133) begin
        _T_3372_1_br_mask <= _T_4135;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1 == rob_tail) begin
            _T_3372_1_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1 == rob_tail) begin
        _T_3372_1_fp_val <= _GEN_84;
      end
    end
    if (_T_4141) begin
      if (io_enq_valids_0) begin
        if (6'h2 == rob_tail) begin
          _T_3372_2_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4156) begin
        _T_3372_2_br_mask <= _T_4158;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h2 == rob_tail) begin
            _T_3372_2_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h2 == rob_tail) begin
        _T_3372_2_fp_val <= _GEN_84;
      end
    end
    if (_T_4164) begin
      if (io_enq_valids_0) begin
        if (6'h3 == rob_tail) begin
          _T_3372_3_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4179) begin
        _T_3372_3_br_mask <= _T_4181;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h3 == rob_tail) begin
            _T_3372_3_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h3 == rob_tail) begin
        _T_3372_3_fp_val <= _GEN_84;
      end
    end
    if (_T_4187) begin
      if (io_enq_valids_0) begin
        if (6'h4 == rob_tail) begin
          _T_3372_4_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4202) begin
        _T_3372_4_br_mask <= _T_4204;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h4 == rob_tail) begin
            _T_3372_4_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h4 == rob_tail) begin
        _T_3372_4_fp_val <= _GEN_84;
      end
    end
    if (_T_4210) begin
      if (io_enq_valids_0) begin
        if (6'h5 == rob_tail) begin
          _T_3372_5_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4225) begin
        _T_3372_5_br_mask <= _T_4227;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h5 == rob_tail) begin
            _T_3372_5_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h5 == rob_tail) begin
        _T_3372_5_fp_val <= _GEN_84;
      end
    end
    if (_T_4233) begin
      if (io_enq_valids_0) begin
        if (6'h6 == rob_tail) begin
          _T_3372_6_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4248) begin
        _T_3372_6_br_mask <= _T_4250;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h6 == rob_tail) begin
            _T_3372_6_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h6 == rob_tail) begin
        _T_3372_6_fp_val <= _GEN_84;
      end
    end
    if (_T_4256) begin
      if (io_enq_valids_0) begin
        if (6'h7 == rob_tail) begin
          _T_3372_7_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4271) begin
        _T_3372_7_br_mask <= _T_4273;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h7 == rob_tail) begin
            _T_3372_7_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h7 == rob_tail) begin
        _T_3372_7_fp_val <= _GEN_84;
      end
    end
    if (_T_4279) begin
      if (io_enq_valids_0) begin
        if (6'h8 == rob_tail) begin
          _T_3372_8_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4294) begin
        _T_3372_8_br_mask <= _T_4296;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h8 == rob_tail) begin
            _T_3372_8_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h8 == rob_tail) begin
        _T_3372_8_fp_val <= _GEN_84;
      end
    end
    if (_T_4302) begin
      if (io_enq_valids_0) begin
        if (6'h9 == rob_tail) begin
          _T_3372_9_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4317) begin
        _T_3372_9_br_mask <= _T_4319;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h9 == rob_tail) begin
            _T_3372_9_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h9 == rob_tail) begin
        _T_3372_9_fp_val <= _GEN_84;
      end
    end
    if (_T_4325) begin
      if (io_enq_valids_0) begin
        if (6'ha == rob_tail) begin
          _T_3372_10_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4340) begin
        _T_3372_10_br_mask <= _T_4342;
      end else begin
        if (io_enq_valids_0) begin
          if (6'ha == rob_tail) begin
            _T_3372_10_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'ha == rob_tail) begin
        _T_3372_10_fp_val <= _GEN_84;
      end
    end
    if (_T_4348) begin
      if (io_enq_valids_0) begin
        if (6'hb == rob_tail) begin
          _T_3372_11_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4363) begin
        _T_3372_11_br_mask <= _T_4365;
      end else begin
        if (io_enq_valids_0) begin
          if (6'hb == rob_tail) begin
            _T_3372_11_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hb == rob_tail) begin
        _T_3372_11_fp_val <= _GEN_84;
      end
    end
    if (_T_4371) begin
      if (io_enq_valids_0) begin
        if (6'hc == rob_tail) begin
          _T_3372_12_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4386) begin
        _T_3372_12_br_mask <= _T_4388;
      end else begin
        if (io_enq_valids_0) begin
          if (6'hc == rob_tail) begin
            _T_3372_12_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hc == rob_tail) begin
        _T_3372_12_fp_val <= _GEN_84;
      end
    end
    if (_T_4394) begin
      if (io_enq_valids_0) begin
        if (6'hd == rob_tail) begin
          _T_3372_13_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4409) begin
        _T_3372_13_br_mask <= _T_4411;
      end else begin
        if (io_enq_valids_0) begin
          if (6'hd == rob_tail) begin
            _T_3372_13_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hd == rob_tail) begin
        _T_3372_13_fp_val <= _GEN_84;
      end
    end
    if (_T_4417) begin
      if (io_enq_valids_0) begin
        if (6'he == rob_tail) begin
          _T_3372_14_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4432) begin
        _T_3372_14_br_mask <= _T_4434;
      end else begin
        if (io_enq_valids_0) begin
          if (6'he == rob_tail) begin
            _T_3372_14_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'he == rob_tail) begin
        _T_3372_14_fp_val <= _GEN_84;
      end
    end
    if (_T_4440) begin
      if (io_enq_valids_0) begin
        if (6'hf == rob_tail) begin
          _T_3372_15_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4455) begin
        _T_3372_15_br_mask <= _T_4457;
      end else begin
        if (io_enq_valids_0) begin
          if (6'hf == rob_tail) begin
            _T_3372_15_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'hf == rob_tail) begin
        _T_3372_15_fp_val <= _GEN_84;
      end
    end
    if (_T_4463) begin
      if (io_enq_valids_0) begin
        if (6'h10 == rob_tail) begin
          _T_3372_16_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4478) begin
        _T_3372_16_br_mask <= _T_4480;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h10 == rob_tail) begin
            _T_3372_16_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h10 == rob_tail) begin
        _T_3372_16_fp_val <= _GEN_84;
      end
    end
    if (_T_4486) begin
      if (io_enq_valids_0) begin
        if (6'h11 == rob_tail) begin
          _T_3372_17_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4501) begin
        _T_3372_17_br_mask <= _T_4503;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h11 == rob_tail) begin
            _T_3372_17_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h11 == rob_tail) begin
        _T_3372_17_fp_val <= _GEN_84;
      end
    end
    if (_T_4509) begin
      if (io_enq_valids_0) begin
        if (6'h12 == rob_tail) begin
          _T_3372_18_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4524) begin
        _T_3372_18_br_mask <= _T_4526;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h12 == rob_tail) begin
            _T_3372_18_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h12 == rob_tail) begin
        _T_3372_18_fp_val <= _GEN_84;
      end
    end
    if (_T_4532) begin
      if (io_enq_valids_0) begin
        if (6'h13 == rob_tail) begin
          _T_3372_19_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4547) begin
        _T_3372_19_br_mask <= _T_4549;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h13 == rob_tail) begin
            _T_3372_19_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h13 == rob_tail) begin
        _T_3372_19_fp_val <= _GEN_84;
      end
    end
    if (_T_4555) begin
      if (io_enq_valids_0) begin
        if (6'h14 == rob_tail) begin
          _T_3372_20_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4570) begin
        _T_3372_20_br_mask <= _T_4572;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h14 == rob_tail) begin
            _T_3372_20_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h14 == rob_tail) begin
        _T_3372_20_fp_val <= _GEN_84;
      end
    end
    if (_T_4578) begin
      if (io_enq_valids_0) begin
        if (6'h15 == rob_tail) begin
          _T_3372_21_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4593) begin
        _T_3372_21_br_mask <= _T_4595;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h15 == rob_tail) begin
            _T_3372_21_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h15 == rob_tail) begin
        _T_3372_21_fp_val <= _GEN_84;
      end
    end
    if (_T_4601) begin
      if (io_enq_valids_0) begin
        if (6'h16 == rob_tail) begin
          _T_3372_22_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4616) begin
        _T_3372_22_br_mask <= _T_4618;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h16 == rob_tail) begin
            _T_3372_22_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h16 == rob_tail) begin
        _T_3372_22_fp_val <= _GEN_84;
      end
    end
    if (_T_4624) begin
      if (io_enq_valids_0) begin
        if (6'h17 == rob_tail) begin
          _T_3372_23_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4639) begin
        _T_3372_23_br_mask <= _T_4641;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h17 == rob_tail) begin
            _T_3372_23_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h17 == rob_tail) begin
        _T_3372_23_fp_val <= _GEN_84;
      end
    end
    if (_T_4647) begin
      if (io_enq_valids_0) begin
        if (6'h18 == rob_tail) begin
          _T_3372_24_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4662) begin
        _T_3372_24_br_mask <= _T_4664;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h18 == rob_tail) begin
            _T_3372_24_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h18 == rob_tail) begin
        _T_3372_24_fp_val <= _GEN_84;
      end
    end
    if (_T_4670) begin
      if (io_enq_valids_0) begin
        if (6'h19 == rob_tail) begin
          _T_3372_25_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4685) begin
        _T_3372_25_br_mask <= _T_4687;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h19 == rob_tail) begin
            _T_3372_25_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h19 == rob_tail) begin
        _T_3372_25_fp_val <= _GEN_84;
      end
    end
    if (_T_4693) begin
      if (io_enq_valids_0) begin
        if (6'h1a == rob_tail) begin
          _T_3372_26_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4708) begin
        _T_3372_26_br_mask <= _T_4710;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1a == rob_tail) begin
            _T_3372_26_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1a == rob_tail) begin
        _T_3372_26_fp_val <= _GEN_84;
      end
    end
    if (_T_4716) begin
      if (io_enq_valids_0) begin
        if (6'h1b == rob_tail) begin
          _T_3372_27_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4731) begin
        _T_3372_27_br_mask <= _T_4733;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1b == rob_tail) begin
            _T_3372_27_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1b == rob_tail) begin
        _T_3372_27_fp_val <= _GEN_84;
      end
    end
    if (_T_4739) begin
      if (io_enq_valids_0) begin
        if (6'h1c == rob_tail) begin
          _T_3372_28_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4754) begin
        _T_3372_28_br_mask <= _T_4756;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1c == rob_tail) begin
            _T_3372_28_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1c == rob_tail) begin
        _T_3372_28_fp_val <= _GEN_84;
      end
    end
    if (_T_4762) begin
      if (io_enq_valids_0) begin
        if (6'h1d == rob_tail) begin
          _T_3372_29_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4777) begin
        _T_3372_29_br_mask <= _T_4779;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1d == rob_tail) begin
            _T_3372_29_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1d == rob_tail) begin
        _T_3372_29_fp_val <= _GEN_84;
      end
    end
    if (_T_4785) begin
      if (io_enq_valids_0) begin
        if (6'h1e == rob_tail) begin
          _T_3372_30_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4800) begin
        _T_3372_30_br_mask <= _T_4802;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1e == rob_tail) begin
            _T_3372_30_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1e == rob_tail) begin
        _T_3372_30_fp_val <= _GEN_84;
      end
    end
    if (_T_4808) begin
      if (io_enq_valids_0) begin
        if (6'h1f == rob_tail) begin
          _T_3372_31_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4823) begin
        _T_3372_31_br_mask <= _T_4825;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h1f == rob_tail) begin
            _T_3372_31_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h1f == rob_tail) begin
        _T_3372_31_fp_val <= _GEN_84;
      end
    end
    if (_T_4831) begin
      if (io_enq_valids_0) begin
        if (6'h20 == rob_tail) begin
          _T_3372_32_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4846) begin
        _T_3372_32_br_mask <= _T_4848;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h20 == rob_tail) begin
            _T_3372_32_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h20 == rob_tail) begin
        _T_3372_32_fp_val <= _GEN_84;
      end
    end
    if (_T_4854) begin
      if (io_enq_valids_0) begin
        if (6'h21 == rob_tail) begin
          _T_3372_33_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4869) begin
        _T_3372_33_br_mask <= _T_4871;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h21 == rob_tail) begin
            _T_3372_33_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h21 == rob_tail) begin
        _T_3372_33_fp_val <= _GEN_84;
      end
    end
    if (_T_4877) begin
      if (io_enq_valids_0) begin
        if (6'h22 == rob_tail) begin
          _T_3372_34_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4892) begin
        _T_3372_34_br_mask <= _T_4894;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h22 == rob_tail) begin
            _T_3372_34_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h22 == rob_tail) begin
        _T_3372_34_fp_val <= _GEN_84;
      end
    end
    if (_T_4900) begin
      if (io_enq_valids_0) begin
        if (6'h23 == rob_tail) begin
          _T_3372_35_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4915) begin
        _T_3372_35_br_mask <= _T_4917;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h23 == rob_tail) begin
            _T_3372_35_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h23 == rob_tail) begin
        _T_3372_35_fp_val <= _GEN_84;
      end
    end
    if (_T_4923) begin
      if (io_enq_valids_0) begin
        if (6'h24 == rob_tail) begin
          _T_3372_36_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4938) begin
        _T_3372_36_br_mask <= _T_4940;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h24 == rob_tail) begin
            _T_3372_36_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h24 == rob_tail) begin
        _T_3372_36_fp_val <= _GEN_84;
      end
    end
    if (_T_4946) begin
      if (io_enq_valids_0) begin
        if (6'h25 == rob_tail) begin
          _T_3372_37_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4961) begin
        _T_3372_37_br_mask <= _T_4963;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h25 == rob_tail) begin
            _T_3372_37_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h25 == rob_tail) begin
        _T_3372_37_fp_val <= _GEN_84;
      end
    end
    if (_T_4969) begin
      if (io_enq_valids_0) begin
        if (6'h26 == rob_tail) begin
          _T_3372_38_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_4984) begin
        _T_3372_38_br_mask <= _T_4986;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h26 == rob_tail) begin
            _T_3372_38_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h26 == rob_tail) begin
        _T_3372_38_fp_val <= _GEN_84;
      end
    end
    if (_T_4992) begin
      if (io_enq_valids_0) begin
        if (6'h27 == rob_tail) begin
          _T_3372_39_br_mask <= _GEN_26;
        end
      end
    end else begin
      if (_T_5007) begin
        _T_3372_39_br_mask <= _T_5009;
      end else begin
        if (io_enq_valids_0) begin
          if (6'h27 == rob_tail) begin
            _T_3372_39_br_mask <= _GEN_26;
          end
        end
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_pdst <= _GEN_54;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_stale_pdst <= _GEN_61;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_is_fencei <= _GEN_68;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_is_store <= _GEN_69;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_is_load <= _GEN_71;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_is_sys_pc2epc <= _GEN_72;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_flush_on_commit <= _GEN_74;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_ldst <= _GEN_75;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_ldst_val <= _GEN_79;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_dst_rtype <= _GEN_80;
      end
    end
    if (io_enq_valids_0) begin
      if (6'h27 == rob_tail) begin
        _T_3372_39_fp_val <= _GEN_84;
      end
    end
    if(_T_3745__T_3768_en & _T_3745__T_3768_mask) begin
      _T_3745[_T_3745__T_3768_addr] <= _T_3745__T_3768_data;
    end
    if(_T_3745__T_3998_en & _T_3745__T_3998_mask) begin
      _T_3745[_T_3745__T_3998_addr] <= _T_3745__T_3998_data;
    end
    if(_T_3745__T_4007_en & _T_3745__T_4007_mask) begin
      _T_3745[_T_3745__T_4007_addr] <= _T_3745__T_4007_data;
    end
    if(_T_3745__T_4088_en & _T_3745__T_4088_mask) begin
      _T_3745[_T_3745__T_4088_addr] <= _T_3745__T_4088_data;
    end
    if(_T_3748__T_3769_en & _T_3748__T_3769_mask) begin
      _T_3748[_T_3748__T_3769_addr] <= _T_3748__T_3769_data;
    end
    if(_T_3748__T_3982_en & _T_3748__T_3982_mask) begin
      _T_3748[_T_3748__T_3982_addr] <= _T_3748__T_3982_data;
    end
    if(_T_3748__T_3990_en & _T_3748__T_3990_mask) begin
      _T_3748[_T_3748__T_3990_addr] <= _T_3748__T_3990_data;
    end
    if (reset) begin
      _T_5637_0 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h0 == rob_head) begin
          _T_5637_0 <= 1'h0;
        end else begin
          if (_T_6659) begin
            _T_5637_0 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h0 == _T_6589) begin
                _T_5637_0 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h0 == rob_tail) begin
                    _T_5637_0 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h0 == rob_tail) begin
                  _T_5637_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6659) begin
          _T_5637_0 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h0 == _T_6589) begin
              _T_5637_0 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h0 == rob_tail) begin
                  _T_5637_0 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h0 == rob_tail) begin
                _T_5637_0 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_1 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1 == rob_head) begin
          _T_5637_1 <= 1'h0;
        end else begin
          if (_T_6682) begin
            _T_5637_1 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1 == _T_6589) begin
                _T_5637_1 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1 == rob_tail) begin
                    _T_5637_1 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1 == rob_tail) begin
                  _T_5637_1 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6682) begin
          _T_5637_1 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1 == _T_6589) begin
              _T_5637_1 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1 == rob_tail) begin
                  _T_5637_1 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1 == rob_tail) begin
                _T_5637_1 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_2 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h2 == rob_head) begin
          _T_5637_2 <= 1'h0;
        end else begin
          if (_T_6705) begin
            _T_5637_2 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h2 == _T_6589) begin
                _T_5637_2 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h2 == rob_tail) begin
                    _T_5637_2 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h2 == rob_tail) begin
                  _T_5637_2 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6705) begin
          _T_5637_2 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h2 == _T_6589) begin
              _T_5637_2 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h2 == rob_tail) begin
                  _T_5637_2 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h2 == rob_tail) begin
                _T_5637_2 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_3 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h3 == rob_head) begin
          _T_5637_3 <= 1'h0;
        end else begin
          if (_T_6728) begin
            _T_5637_3 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h3 == _T_6589) begin
                _T_5637_3 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h3 == rob_tail) begin
                    _T_5637_3 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h3 == rob_tail) begin
                  _T_5637_3 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6728) begin
          _T_5637_3 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h3 == _T_6589) begin
              _T_5637_3 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h3 == rob_tail) begin
                  _T_5637_3 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h3 == rob_tail) begin
                _T_5637_3 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_4 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h4 == rob_head) begin
          _T_5637_4 <= 1'h0;
        end else begin
          if (_T_6751) begin
            _T_5637_4 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h4 == _T_6589) begin
                _T_5637_4 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h4 == rob_tail) begin
                    _T_5637_4 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h4 == rob_tail) begin
                  _T_5637_4 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6751) begin
          _T_5637_4 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h4 == _T_6589) begin
              _T_5637_4 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h4 == rob_tail) begin
                  _T_5637_4 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h4 == rob_tail) begin
                _T_5637_4 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_5 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h5 == rob_head) begin
          _T_5637_5 <= 1'h0;
        end else begin
          if (_T_6774) begin
            _T_5637_5 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h5 == _T_6589) begin
                _T_5637_5 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h5 == rob_tail) begin
                    _T_5637_5 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h5 == rob_tail) begin
                  _T_5637_5 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6774) begin
          _T_5637_5 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h5 == _T_6589) begin
              _T_5637_5 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h5 == rob_tail) begin
                  _T_5637_5 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h5 == rob_tail) begin
                _T_5637_5 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_6 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h6 == rob_head) begin
          _T_5637_6 <= 1'h0;
        end else begin
          if (_T_6797) begin
            _T_5637_6 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h6 == _T_6589) begin
                _T_5637_6 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h6 == rob_tail) begin
                    _T_5637_6 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h6 == rob_tail) begin
                  _T_5637_6 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6797) begin
          _T_5637_6 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h6 == _T_6589) begin
              _T_5637_6 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h6 == rob_tail) begin
                  _T_5637_6 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h6 == rob_tail) begin
                _T_5637_6 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_7 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h7 == rob_head) begin
          _T_5637_7 <= 1'h0;
        end else begin
          if (_T_6820) begin
            _T_5637_7 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h7 == _T_6589) begin
                _T_5637_7 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h7 == rob_tail) begin
                    _T_5637_7 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h7 == rob_tail) begin
                  _T_5637_7 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6820) begin
          _T_5637_7 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h7 == _T_6589) begin
              _T_5637_7 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h7 == rob_tail) begin
                  _T_5637_7 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h7 == rob_tail) begin
                _T_5637_7 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_8 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h8 == rob_head) begin
          _T_5637_8 <= 1'h0;
        end else begin
          if (_T_6843) begin
            _T_5637_8 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h8 == _T_6589) begin
                _T_5637_8 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h8 == rob_tail) begin
                    _T_5637_8 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h8 == rob_tail) begin
                  _T_5637_8 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6843) begin
          _T_5637_8 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h8 == _T_6589) begin
              _T_5637_8 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h8 == rob_tail) begin
                  _T_5637_8 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h8 == rob_tail) begin
                _T_5637_8 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_9 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h9 == rob_head) begin
          _T_5637_9 <= 1'h0;
        end else begin
          if (_T_6866) begin
            _T_5637_9 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h9 == _T_6589) begin
                _T_5637_9 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h9 == rob_tail) begin
                    _T_5637_9 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h9 == rob_tail) begin
                  _T_5637_9 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6866) begin
          _T_5637_9 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h9 == _T_6589) begin
              _T_5637_9 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h9 == rob_tail) begin
                  _T_5637_9 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h9 == rob_tail) begin
                _T_5637_9 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_10 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'ha == rob_head) begin
          _T_5637_10 <= 1'h0;
        end else begin
          if (_T_6889) begin
            _T_5637_10 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'ha == _T_6589) begin
                _T_5637_10 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'ha == rob_tail) begin
                    _T_5637_10 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'ha == rob_tail) begin
                  _T_5637_10 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6889) begin
          _T_5637_10 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'ha == _T_6589) begin
              _T_5637_10 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'ha == rob_tail) begin
                  _T_5637_10 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'ha == rob_tail) begin
                _T_5637_10 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_11 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'hb == rob_head) begin
          _T_5637_11 <= 1'h0;
        end else begin
          if (_T_6912) begin
            _T_5637_11 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hb == _T_6589) begin
                _T_5637_11 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'hb == rob_tail) begin
                    _T_5637_11 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'hb == rob_tail) begin
                  _T_5637_11 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6912) begin
          _T_5637_11 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hb == _T_6589) begin
              _T_5637_11 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'hb == rob_tail) begin
                  _T_5637_11 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'hb == rob_tail) begin
                _T_5637_11 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_12 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'hc == rob_head) begin
          _T_5637_12 <= 1'h0;
        end else begin
          if (_T_6935) begin
            _T_5637_12 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hc == _T_6589) begin
                _T_5637_12 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'hc == rob_tail) begin
                    _T_5637_12 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'hc == rob_tail) begin
                  _T_5637_12 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6935) begin
          _T_5637_12 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hc == _T_6589) begin
              _T_5637_12 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'hc == rob_tail) begin
                  _T_5637_12 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'hc == rob_tail) begin
                _T_5637_12 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_13 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'hd == rob_head) begin
          _T_5637_13 <= 1'h0;
        end else begin
          if (_T_6958) begin
            _T_5637_13 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hd == _T_6589) begin
                _T_5637_13 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'hd == rob_tail) begin
                    _T_5637_13 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'hd == rob_tail) begin
                  _T_5637_13 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6958) begin
          _T_5637_13 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hd == _T_6589) begin
              _T_5637_13 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'hd == rob_tail) begin
                  _T_5637_13 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'hd == rob_tail) begin
                _T_5637_13 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_14 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'he == rob_head) begin
          _T_5637_14 <= 1'h0;
        end else begin
          if (_T_6981) begin
            _T_5637_14 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'he == _T_6589) begin
                _T_5637_14 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'he == rob_tail) begin
                    _T_5637_14 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'he == rob_tail) begin
                  _T_5637_14 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_6981) begin
          _T_5637_14 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'he == _T_6589) begin
              _T_5637_14 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'he == rob_tail) begin
                  _T_5637_14 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'he == rob_tail) begin
                _T_5637_14 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_15 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'hf == rob_head) begin
          _T_5637_15 <= 1'h0;
        end else begin
          if (_T_7004) begin
            _T_5637_15 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'hf == _T_6589) begin
                _T_5637_15 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'hf == rob_tail) begin
                    _T_5637_15 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'hf == rob_tail) begin
                  _T_5637_15 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7004) begin
          _T_5637_15 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'hf == _T_6589) begin
              _T_5637_15 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'hf == rob_tail) begin
                  _T_5637_15 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'hf == rob_tail) begin
                _T_5637_15 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_16 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h10 == rob_head) begin
          _T_5637_16 <= 1'h0;
        end else begin
          if (_T_7027) begin
            _T_5637_16 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h10 == _T_6589) begin
                _T_5637_16 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h10 == rob_tail) begin
                    _T_5637_16 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h10 == rob_tail) begin
                  _T_5637_16 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7027) begin
          _T_5637_16 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h10 == _T_6589) begin
              _T_5637_16 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h10 == rob_tail) begin
                  _T_5637_16 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h10 == rob_tail) begin
                _T_5637_16 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_17 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h11 == rob_head) begin
          _T_5637_17 <= 1'h0;
        end else begin
          if (_T_7050) begin
            _T_5637_17 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h11 == _T_6589) begin
                _T_5637_17 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h11 == rob_tail) begin
                    _T_5637_17 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h11 == rob_tail) begin
                  _T_5637_17 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7050) begin
          _T_5637_17 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h11 == _T_6589) begin
              _T_5637_17 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h11 == rob_tail) begin
                  _T_5637_17 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h11 == rob_tail) begin
                _T_5637_17 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_18 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h12 == rob_head) begin
          _T_5637_18 <= 1'h0;
        end else begin
          if (_T_7073) begin
            _T_5637_18 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h12 == _T_6589) begin
                _T_5637_18 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h12 == rob_tail) begin
                    _T_5637_18 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h12 == rob_tail) begin
                  _T_5637_18 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7073) begin
          _T_5637_18 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h12 == _T_6589) begin
              _T_5637_18 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h12 == rob_tail) begin
                  _T_5637_18 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h12 == rob_tail) begin
                _T_5637_18 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_19 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h13 == rob_head) begin
          _T_5637_19 <= 1'h0;
        end else begin
          if (_T_7096) begin
            _T_5637_19 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h13 == _T_6589) begin
                _T_5637_19 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h13 == rob_tail) begin
                    _T_5637_19 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h13 == rob_tail) begin
                  _T_5637_19 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7096) begin
          _T_5637_19 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h13 == _T_6589) begin
              _T_5637_19 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h13 == rob_tail) begin
                  _T_5637_19 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h13 == rob_tail) begin
                _T_5637_19 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_20 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h14 == rob_head) begin
          _T_5637_20 <= 1'h0;
        end else begin
          if (_T_7119) begin
            _T_5637_20 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h14 == _T_6589) begin
                _T_5637_20 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h14 == rob_tail) begin
                    _T_5637_20 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h14 == rob_tail) begin
                  _T_5637_20 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7119) begin
          _T_5637_20 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h14 == _T_6589) begin
              _T_5637_20 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h14 == rob_tail) begin
                  _T_5637_20 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h14 == rob_tail) begin
                _T_5637_20 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_21 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h15 == rob_head) begin
          _T_5637_21 <= 1'h0;
        end else begin
          if (_T_7142) begin
            _T_5637_21 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h15 == _T_6589) begin
                _T_5637_21 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h15 == rob_tail) begin
                    _T_5637_21 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h15 == rob_tail) begin
                  _T_5637_21 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7142) begin
          _T_5637_21 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h15 == _T_6589) begin
              _T_5637_21 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h15 == rob_tail) begin
                  _T_5637_21 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h15 == rob_tail) begin
                _T_5637_21 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_22 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h16 == rob_head) begin
          _T_5637_22 <= 1'h0;
        end else begin
          if (_T_7165) begin
            _T_5637_22 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h16 == _T_6589) begin
                _T_5637_22 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h16 == rob_tail) begin
                    _T_5637_22 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h16 == rob_tail) begin
                  _T_5637_22 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7165) begin
          _T_5637_22 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h16 == _T_6589) begin
              _T_5637_22 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h16 == rob_tail) begin
                  _T_5637_22 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h16 == rob_tail) begin
                _T_5637_22 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_23 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h17 == rob_head) begin
          _T_5637_23 <= 1'h0;
        end else begin
          if (_T_7188) begin
            _T_5637_23 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h17 == _T_6589) begin
                _T_5637_23 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h17 == rob_tail) begin
                    _T_5637_23 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h17 == rob_tail) begin
                  _T_5637_23 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7188) begin
          _T_5637_23 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h17 == _T_6589) begin
              _T_5637_23 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h17 == rob_tail) begin
                  _T_5637_23 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h17 == rob_tail) begin
                _T_5637_23 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_24 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h18 == rob_head) begin
          _T_5637_24 <= 1'h0;
        end else begin
          if (_T_7211) begin
            _T_5637_24 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h18 == _T_6589) begin
                _T_5637_24 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h18 == rob_tail) begin
                    _T_5637_24 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h18 == rob_tail) begin
                  _T_5637_24 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7211) begin
          _T_5637_24 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h18 == _T_6589) begin
              _T_5637_24 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h18 == rob_tail) begin
                  _T_5637_24 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h18 == rob_tail) begin
                _T_5637_24 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_25 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h19 == rob_head) begin
          _T_5637_25 <= 1'h0;
        end else begin
          if (_T_7234) begin
            _T_5637_25 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h19 == _T_6589) begin
                _T_5637_25 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h19 == rob_tail) begin
                    _T_5637_25 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h19 == rob_tail) begin
                  _T_5637_25 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7234) begin
          _T_5637_25 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h19 == _T_6589) begin
              _T_5637_25 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h19 == rob_tail) begin
                  _T_5637_25 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h19 == rob_tail) begin
                _T_5637_25 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_26 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1a == rob_head) begin
          _T_5637_26 <= 1'h0;
        end else begin
          if (_T_7257) begin
            _T_5637_26 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1a == _T_6589) begin
                _T_5637_26 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1a == rob_tail) begin
                    _T_5637_26 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1a == rob_tail) begin
                  _T_5637_26 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7257) begin
          _T_5637_26 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1a == _T_6589) begin
              _T_5637_26 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1a == rob_tail) begin
                  _T_5637_26 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1a == rob_tail) begin
                _T_5637_26 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_27 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1b == rob_head) begin
          _T_5637_27 <= 1'h0;
        end else begin
          if (_T_7280) begin
            _T_5637_27 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1b == _T_6589) begin
                _T_5637_27 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1b == rob_tail) begin
                    _T_5637_27 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1b == rob_tail) begin
                  _T_5637_27 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7280) begin
          _T_5637_27 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1b == _T_6589) begin
              _T_5637_27 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1b == rob_tail) begin
                  _T_5637_27 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1b == rob_tail) begin
                _T_5637_27 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_28 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1c == rob_head) begin
          _T_5637_28 <= 1'h0;
        end else begin
          if (_T_7303) begin
            _T_5637_28 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1c == _T_6589) begin
                _T_5637_28 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1c == rob_tail) begin
                    _T_5637_28 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1c == rob_tail) begin
                  _T_5637_28 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7303) begin
          _T_5637_28 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1c == _T_6589) begin
              _T_5637_28 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1c == rob_tail) begin
                  _T_5637_28 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1c == rob_tail) begin
                _T_5637_28 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_29 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1d == rob_head) begin
          _T_5637_29 <= 1'h0;
        end else begin
          if (_T_7326) begin
            _T_5637_29 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1d == _T_6589) begin
                _T_5637_29 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1d == rob_tail) begin
                    _T_5637_29 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1d == rob_tail) begin
                  _T_5637_29 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7326) begin
          _T_5637_29 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1d == _T_6589) begin
              _T_5637_29 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1d == rob_tail) begin
                  _T_5637_29 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1d == rob_tail) begin
                _T_5637_29 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_30 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1e == rob_head) begin
          _T_5637_30 <= 1'h0;
        end else begin
          if (_T_7349) begin
            _T_5637_30 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1e == _T_6589) begin
                _T_5637_30 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1e == rob_tail) begin
                    _T_5637_30 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1e == rob_tail) begin
                  _T_5637_30 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7349) begin
          _T_5637_30 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1e == _T_6589) begin
              _T_5637_30 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1e == rob_tail) begin
                  _T_5637_30 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1e == rob_tail) begin
                _T_5637_30 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_31 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h1f == rob_head) begin
          _T_5637_31 <= 1'h0;
        end else begin
          if (_T_7372) begin
            _T_5637_31 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h1f == _T_6589) begin
                _T_5637_31 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h1f == rob_tail) begin
                    _T_5637_31 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1f == rob_tail) begin
                  _T_5637_31 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7372) begin
          _T_5637_31 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h1f == _T_6589) begin
              _T_5637_31 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h1f == rob_tail) begin
                  _T_5637_31 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h1f == rob_tail) begin
                _T_5637_31 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_32 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h20 == rob_head) begin
          _T_5637_32 <= 1'h0;
        end else begin
          if (_T_7395) begin
            _T_5637_32 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h20 == _T_6589) begin
                _T_5637_32 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h20 == rob_tail) begin
                    _T_5637_32 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h20 == rob_tail) begin
                  _T_5637_32 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7395) begin
          _T_5637_32 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h20 == _T_6589) begin
              _T_5637_32 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h20 == rob_tail) begin
                  _T_5637_32 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h20 == rob_tail) begin
                _T_5637_32 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_33 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h21 == rob_head) begin
          _T_5637_33 <= 1'h0;
        end else begin
          if (_T_7418) begin
            _T_5637_33 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h21 == _T_6589) begin
                _T_5637_33 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h21 == rob_tail) begin
                    _T_5637_33 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h21 == rob_tail) begin
                  _T_5637_33 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7418) begin
          _T_5637_33 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h21 == _T_6589) begin
              _T_5637_33 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h21 == rob_tail) begin
                  _T_5637_33 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h21 == rob_tail) begin
                _T_5637_33 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_34 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h22 == rob_head) begin
          _T_5637_34 <= 1'h0;
        end else begin
          if (_T_7441) begin
            _T_5637_34 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h22 == _T_6589) begin
                _T_5637_34 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h22 == rob_tail) begin
                    _T_5637_34 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h22 == rob_tail) begin
                  _T_5637_34 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7441) begin
          _T_5637_34 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h22 == _T_6589) begin
              _T_5637_34 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h22 == rob_tail) begin
                  _T_5637_34 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h22 == rob_tail) begin
                _T_5637_34 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_35 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h23 == rob_head) begin
          _T_5637_35 <= 1'h0;
        end else begin
          if (_T_7464) begin
            _T_5637_35 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h23 == _T_6589) begin
                _T_5637_35 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h23 == rob_tail) begin
                    _T_5637_35 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h23 == rob_tail) begin
                  _T_5637_35 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7464) begin
          _T_5637_35 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h23 == _T_6589) begin
              _T_5637_35 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h23 == rob_tail) begin
                  _T_5637_35 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h23 == rob_tail) begin
                _T_5637_35 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_36 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h24 == rob_head) begin
          _T_5637_36 <= 1'h0;
        end else begin
          if (_T_7487) begin
            _T_5637_36 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h24 == _T_6589) begin
                _T_5637_36 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h24 == rob_tail) begin
                    _T_5637_36 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h24 == rob_tail) begin
                  _T_5637_36 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7487) begin
          _T_5637_36 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h24 == _T_6589) begin
              _T_5637_36 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h24 == rob_tail) begin
                  _T_5637_36 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h24 == rob_tail) begin
                _T_5637_36 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_37 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h25 == rob_head) begin
          _T_5637_37 <= 1'h0;
        end else begin
          if (_T_7510) begin
            _T_5637_37 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h25 == _T_6589) begin
                _T_5637_37 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h25 == rob_tail) begin
                    _T_5637_37 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h25 == rob_tail) begin
                  _T_5637_37 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7510) begin
          _T_5637_37 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h25 == _T_6589) begin
              _T_5637_37 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h25 == rob_tail) begin
                  _T_5637_37 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h25 == rob_tail) begin
                _T_5637_37 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_38 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h26 == rob_head) begin
          _T_5637_38 <= 1'h0;
        end else begin
          if (_T_7533) begin
            _T_5637_38 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h26 == _T_6589) begin
                _T_5637_38 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h26 == rob_tail) begin
                    _T_5637_38 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h26 == rob_tail) begin
                  _T_5637_38 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7533) begin
          _T_5637_38 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h26 == _T_6589) begin
              _T_5637_38 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h26 == rob_tail) begin
                  _T_5637_38 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h26 == rob_tail) begin
                _T_5637_38 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5637_39 <= 1'h0;
    end else begin
      if (will_commit_1) begin
        if (6'h27 == rob_head) begin
          _T_5637_39 <= 1'h0;
        end else begin
          if (_T_7556) begin
            _T_5637_39 <= 1'h0;
          end else begin
            if (_T_4026) begin
              if (6'h27 == _T_6589) begin
                _T_5637_39 <= 1'h0;
              end else begin
                if (io_enq_valids_1) begin
                  if (6'h27 == rob_tail) begin
                    _T_5637_39 <= 1'h1;
                  end
                end
              end
            end else begin
              if (io_enq_valids_1) begin
                if (6'h27 == rob_tail) begin
                  _T_5637_39 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_7556) begin
          _T_5637_39 <= 1'h0;
        end else begin
          if (_T_4026) begin
            if (6'h27 == _T_6589) begin
              _T_5637_39 <= 1'h0;
            end else begin
              if (io_enq_valids_1) begin
                if (6'h27 == rob_tail) begin
                  _T_5637_39 <= 1'h1;
                end
              end
            end
          end else begin
            if (io_enq_valids_1) begin
              if (6'h27 == rob_tail) begin
                _T_5637_39 <= 1'h1;
              end
            end
          end
        end
      end
    end
    if(_T_5764__T_6317_en & _T_5764__T_6317_mask) begin
      _T_5764[_T_5764__T_6317_addr] <= _T_5764__T_6317_data;
    end
    if(_T_5764__T_6383_en & _T_5764__T_6383_mask) begin
      _T_5764[_T_5764__T_6383_addr] <= _T_5764__T_6383_data;
    end
    if(_T_5764__T_6392_en & _T_5764__T_6392_mask) begin
      _T_5764[_T_5764__T_6392_addr] <= _T_5764__T_6392_data;
    end
    if(_T_5764__T_6401_en & _T_5764__T_6401_mask) begin
      _T_5764[_T_5764__T_6401_addr] <= _T_5764__T_6401_data;
    end
    if(_T_5764__T_6410_en & _T_5764__T_6410_mask) begin
      _T_5764[_T_5764__T_6410_addr] <= _T_5764__T_6410_data;
    end
    if(_T_5764__T_6419_en & _T_5764__T_6419_mask) begin
      _T_5764[_T_5764__T_6419_addr] <= _T_5764__T_6419_data;
    end
    if(_T_5764__T_6428_en & _T_5764__T_6428_mask) begin
      _T_5764[_T_5764__T_6428_addr] <= _T_5764__T_6428_data;
    end
    if(_T_5764__T_6455_en & _T_5764__T_6455_mask) begin
      _T_5764[_T_5764__T_6455_addr] <= _T_5764__T_6455_data;
    end
    if (_T_6659) begin
      if (io_enq_valids_1) begin
        if (6'h0 == rob_tail) begin
          _T_5936_0_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6674) begin
        _T_5936_0_br_mask <= _T_6676;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h0 == rob_tail) begin
            _T_5936_0_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h0 == rob_tail) begin
        _T_5936_0_fp_val <= _GEN_311;
      end
    end
    if (_T_6682) begin
      if (io_enq_valids_1) begin
        if (6'h1 == rob_tail) begin
          _T_5936_1_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6697) begin
        _T_5936_1_br_mask <= _T_6699;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1 == rob_tail) begin
            _T_5936_1_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1 == rob_tail) begin
        _T_5936_1_fp_val <= _GEN_311;
      end
    end
    if (_T_6705) begin
      if (io_enq_valids_1) begin
        if (6'h2 == rob_tail) begin
          _T_5936_2_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6720) begin
        _T_5936_2_br_mask <= _T_6722;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h2 == rob_tail) begin
            _T_5936_2_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h2 == rob_tail) begin
        _T_5936_2_fp_val <= _GEN_311;
      end
    end
    if (_T_6728) begin
      if (io_enq_valids_1) begin
        if (6'h3 == rob_tail) begin
          _T_5936_3_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6743) begin
        _T_5936_3_br_mask <= _T_6745;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h3 == rob_tail) begin
            _T_5936_3_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h3 == rob_tail) begin
        _T_5936_3_fp_val <= _GEN_311;
      end
    end
    if (_T_6751) begin
      if (io_enq_valids_1) begin
        if (6'h4 == rob_tail) begin
          _T_5936_4_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6766) begin
        _T_5936_4_br_mask <= _T_6768;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h4 == rob_tail) begin
            _T_5936_4_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h4 == rob_tail) begin
        _T_5936_4_fp_val <= _GEN_311;
      end
    end
    if (_T_6774) begin
      if (io_enq_valids_1) begin
        if (6'h5 == rob_tail) begin
          _T_5936_5_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6789) begin
        _T_5936_5_br_mask <= _T_6791;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h5 == rob_tail) begin
            _T_5936_5_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h5 == rob_tail) begin
        _T_5936_5_fp_val <= _GEN_311;
      end
    end
    if (_T_6797) begin
      if (io_enq_valids_1) begin
        if (6'h6 == rob_tail) begin
          _T_5936_6_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6812) begin
        _T_5936_6_br_mask <= _T_6814;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h6 == rob_tail) begin
            _T_5936_6_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h6 == rob_tail) begin
        _T_5936_6_fp_val <= _GEN_311;
      end
    end
    if (_T_6820) begin
      if (io_enq_valids_1) begin
        if (6'h7 == rob_tail) begin
          _T_5936_7_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6835) begin
        _T_5936_7_br_mask <= _T_6837;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h7 == rob_tail) begin
            _T_5936_7_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h7 == rob_tail) begin
        _T_5936_7_fp_val <= _GEN_311;
      end
    end
    if (_T_6843) begin
      if (io_enq_valids_1) begin
        if (6'h8 == rob_tail) begin
          _T_5936_8_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6858) begin
        _T_5936_8_br_mask <= _T_6860;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h8 == rob_tail) begin
            _T_5936_8_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h8 == rob_tail) begin
        _T_5936_8_fp_val <= _GEN_311;
      end
    end
    if (_T_6866) begin
      if (io_enq_valids_1) begin
        if (6'h9 == rob_tail) begin
          _T_5936_9_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6881) begin
        _T_5936_9_br_mask <= _T_6883;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h9 == rob_tail) begin
            _T_5936_9_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h9 == rob_tail) begin
        _T_5936_9_fp_val <= _GEN_311;
      end
    end
    if (_T_6889) begin
      if (io_enq_valids_1) begin
        if (6'ha == rob_tail) begin
          _T_5936_10_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6904) begin
        _T_5936_10_br_mask <= _T_6906;
      end else begin
        if (io_enq_valids_1) begin
          if (6'ha == rob_tail) begin
            _T_5936_10_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'ha == rob_tail) begin
        _T_5936_10_fp_val <= _GEN_311;
      end
    end
    if (_T_6912) begin
      if (io_enq_valids_1) begin
        if (6'hb == rob_tail) begin
          _T_5936_11_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6927) begin
        _T_5936_11_br_mask <= _T_6929;
      end else begin
        if (io_enq_valids_1) begin
          if (6'hb == rob_tail) begin
            _T_5936_11_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hb == rob_tail) begin
        _T_5936_11_fp_val <= _GEN_311;
      end
    end
    if (_T_6935) begin
      if (io_enq_valids_1) begin
        if (6'hc == rob_tail) begin
          _T_5936_12_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6950) begin
        _T_5936_12_br_mask <= _T_6952;
      end else begin
        if (io_enq_valids_1) begin
          if (6'hc == rob_tail) begin
            _T_5936_12_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hc == rob_tail) begin
        _T_5936_12_fp_val <= _GEN_311;
      end
    end
    if (_T_6958) begin
      if (io_enq_valids_1) begin
        if (6'hd == rob_tail) begin
          _T_5936_13_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6973) begin
        _T_5936_13_br_mask <= _T_6975;
      end else begin
        if (io_enq_valids_1) begin
          if (6'hd == rob_tail) begin
            _T_5936_13_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hd == rob_tail) begin
        _T_5936_13_fp_val <= _GEN_311;
      end
    end
    if (_T_6981) begin
      if (io_enq_valids_1) begin
        if (6'he == rob_tail) begin
          _T_5936_14_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_6996) begin
        _T_5936_14_br_mask <= _T_6998;
      end else begin
        if (io_enq_valids_1) begin
          if (6'he == rob_tail) begin
            _T_5936_14_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'he == rob_tail) begin
        _T_5936_14_fp_val <= _GEN_311;
      end
    end
    if (_T_7004) begin
      if (io_enq_valids_1) begin
        if (6'hf == rob_tail) begin
          _T_5936_15_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7019) begin
        _T_5936_15_br_mask <= _T_7021;
      end else begin
        if (io_enq_valids_1) begin
          if (6'hf == rob_tail) begin
            _T_5936_15_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'hf == rob_tail) begin
        _T_5936_15_fp_val <= _GEN_311;
      end
    end
    if (_T_7027) begin
      if (io_enq_valids_1) begin
        if (6'h10 == rob_tail) begin
          _T_5936_16_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7042) begin
        _T_5936_16_br_mask <= _T_7044;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h10 == rob_tail) begin
            _T_5936_16_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h10 == rob_tail) begin
        _T_5936_16_fp_val <= _GEN_311;
      end
    end
    if (_T_7050) begin
      if (io_enq_valids_1) begin
        if (6'h11 == rob_tail) begin
          _T_5936_17_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7065) begin
        _T_5936_17_br_mask <= _T_7067;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h11 == rob_tail) begin
            _T_5936_17_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h11 == rob_tail) begin
        _T_5936_17_fp_val <= _GEN_311;
      end
    end
    if (_T_7073) begin
      if (io_enq_valids_1) begin
        if (6'h12 == rob_tail) begin
          _T_5936_18_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7088) begin
        _T_5936_18_br_mask <= _T_7090;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h12 == rob_tail) begin
            _T_5936_18_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h12 == rob_tail) begin
        _T_5936_18_fp_val <= _GEN_311;
      end
    end
    if (_T_7096) begin
      if (io_enq_valids_1) begin
        if (6'h13 == rob_tail) begin
          _T_5936_19_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7111) begin
        _T_5936_19_br_mask <= _T_7113;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h13 == rob_tail) begin
            _T_5936_19_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h13 == rob_tail) begin
        _T_5936_19_fp_val <= _GEN_311;
      end
    end
    if (_T_7119) begin
      if (io_enq_valids_1) begin
        if (6'h14 == rob_tail) begin
          _T_5936_20_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7134) begin
        _T_5936_20_br_mask <= _T_7136;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h14 == rob_tail) begin
            _T_5936_20_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h14 == rob_tail) begin
        _T_5936_20_fp_val <= _GEN_311;
      end
    end
    if (_T_7142) begin
      if (io_enq_valids_1) begin
        if (6'h15 == rob_tail) begin
          _T_5936_21_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7157) begin
        _T_5936_21_br_mask <= _T_7159;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h15 == rob_tail) begin
            _T_5936_21_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h15 == rob_tail) begin
        _T_5936_21_fp_val <= _GEN_311;
      end
    end
    if (_T_7165) begin
      if (io_enq_valids_1) begin
        if (6'h16 == rob_tail) begin
          _T_5936_22_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7180) begin
        _T_5936_22_br_mask <= _T_7182;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h16 == rob_tail) begin
            _T_5936_22_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h16 == rob_tail) begin
        _T_5936_22_fp_val <= _GEN_311;
      end
    end
    if (_T_7188) begin
      if (io_enq_valids_1) begin
        if (6'h17 == rob_tail) begin
          _T_5936_23_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7203) begin
        _T_5936_23_br_mask <= _T_7205;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h17 == rob_tail) begin
            _T_5936_23_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h17 == rob_tail) begin
        _T_5936_23_fp_val <= _GEN_311;
      end
    end
    if (_T_7211) begin
      if (io_enq_valids_1) begin
        if (6'h18 == rob_tail) begin
          _T_5936_24_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7226) begin
        _T_5936_24_br_mask <= _T_7228;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h18 == rob_tail) begin
            _T_5936_24_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h18 == rob_tail) begin
        _T_5936_24_fp_val <= _GEN_311;
      end
    end
    if (_T_7234) begin
      if (io_enq_valids_1) begin
        if (6'h19 == rob_tail) begin
          _T_5936_25_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7249) begin
        _T_5936_25_br_mask <= _T_7251;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h19 == rob_tail) begin
            _T_5936_25_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h19 == rob_tail) begin
        _T_5936_25_fp_val <= _GEN_311;
      end
    end
    if (_T_7257) begin
      if (io_enq_valids_1) begin
        if (6'h1a == rob_tail) begin
          _T_5936_26_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7272) begin
        _T_5936_26_br_mask <= _T_7274;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1a == rob_tail) begin
            _T_5936_26_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1a == rob_tail) begin
        _T_5936_26_fp_val <= _GEN_311;
      end
    end
    if (_T_7280) begin
      if (io_enq_valids_1) begin
        if (6'h1b == rob_tail) begin
          _T_5936_27_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7295) begin
        _T_5936_27_br_mask <= _T_7297;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1b == rob_tail) begin
            _T_5936_27_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1b == rob_tail) begin
        _T_5936_27_fp_val <= _GEN_311;
      end
    end
    if (_T_7303) begin
      if (io_enq_valids_1) begin
        if (6'h1c == rob_tail) begin
          _T_5936_28_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7318) begin
        _T_5936_28_br_mask <= _T_7320;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1c == rob_tail) begin
            _T_5936_28_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1c == rob_tail) begin
        _T_5936_28_fp_val <= _GEN_311;
      end
    end
    if (_T_7326) begin
      if (io_enq_valids_1) begin
        if (6'h1d == rob_tail) begin
          _T_5936_29_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7341) begin
        _T_5936_29_br_mask <= _T_7343;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1d == rob_tail) begin
            _T_5936_29_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1d == rob_tail) begin
        _T_5936_29_fp_val <= _GEN_311;
      end
    end
    if (_T_7349) begin
      if (io_enq_valids_1) begin
        if (6'h1e == rob_tail) begin
          _T_5936_30_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7364) begin
        _T_5936_30_br_mask <= _T_7366;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1e == rob_tail) begin
            _T_5936_30_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1e == rob_tail) begin
        _T_5936_30_fp_val <= _GEN_311;
      end
    end
    if (_T_7372) begin
      if (io_enq_valids_1) begin
        if (6'h1f == rob_tail) begin
          _T_5936_31_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7387) begin
        _T_5936_31_br_mask <= _T_7389;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h1f == rob_tail) begin
            _T_5936_31_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h1f == rob_tail) begin
        _T_5936_31_fp_val <= _GEN_311;
      end
    end
    if (_T_7395) begin
      if (io_enq_valids_1) begin
        if (6'h20 == rob_tail) begin
          _T_5936_32_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7410) begin
        _T_5936_32_br_mask <= _T_7412;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h20 == rob_tail) begin
            _T_5936_32_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h20 == rob_tail) begin
        _T_5936_32_fp_val <= _GEN_311;
      end
    end
    if (_T_7418) begin
      if (io_enq_valids_1) begin
        if (6'h21 == rob_tail) begin
          _T_5936_33_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7433) begin
        _T_5936_33_br_mask <= _T_7435;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h21 == rob_tail) begin
            _T_5936_33_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h21 == rob_tail) begin
        _T_5936_33_fp_val <= _GEN_311;
      end
    end
    if (_T_7441) begin
      if (io_enq_valids_1) begin
        if (6'h22 == rob_tail) begin
          _T_5936_34_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7456) begin
        _T_5936_34_br_mask <= _T_7458;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h22 == rob_tail) begin
            _T_5936_34_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h22 == rob_tail) begin
        _T_5936_34_fp_val <= _GEN_311;
      end
    end
    if (_T_7464) begin
      if (io_enq_valids_1) begin
        if (6'h23 == rob_tail) begin
          _T_5936_35_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7479) begin
        _T_5936_35_br_mask <= _T_7481;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h23 == rob_tail) begin
            _T_5936_35_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h23 == rob_tail) begin
        _T_5936_35_fp_val <= _GEN_311;
      end
    end
    if (_T_7487) begin
      if (io_enq_valids_1) begin
        if (6'h24 == rob_tail) begin
          _T_5936_36_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7502) begin
        _T_5936_36_br_mask <= _T_7504;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h24 == rob_tail) begin
            _T_5936_36_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h24 == rob_tail) begin
        _T_5936_36_fp_val <= _GEN_311;
      end
    end
    if (_T_7510) begin
      if (io_enq_valids_1) begin
        if (6'h25 == rob_tail) begin
          _T_5936_37_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7525) begin
        _T_5936_37_br_mask <= _T_7527;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h25 == rob_tail) begin
            _T_5936_37_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h25 == rob_tail) begin
        _T_5936_37_fp_val <= _GEN_311;
      end
    end
    if (_T_7533) begin
      if (io_enq_valids_1) begin
        if (6'h26 == rob_tail) begin
          _T_5936_38_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7548) begin
        _T_5936_38_br_mask <= _T_7550;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h26 == rob_tail) begin
            _T_5936_38_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h26 == rob_tail) begin
        _T_5936_38_fp_val <= _GEN_311;
      end
    end
    if (_T_7556) begin
      if (io_enq_valids_1) begin
        if (6'h27 == rob_tail) begin
          _T_5936_39_br_mask <= _GEN_253;
        end
      end
    end else begin
      if (_T_7571) begin
        _T_5936_39_br_mask <= _T_7573;
      end else begin
        if (io_enq_valids_1) begin
          if (6'h27 == rob_tail) begin
            _T_5936_39_br_mask <= _GEN_253;
          end
        end
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_pdst <= _GEN_281;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_stale_pdst <= _GEN_288;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_is_fencei <= _GEN_295;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_is_store <= _GEN_296;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_is_load <= _GEN_298;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_is_sys_pc2epc <= _GEN_299;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_flush_on_commit <= _GEN_301;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_ldst <= _GEN_302;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_ldst_val <= _GEN_306;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_dst_rtype <= _GEN_307;
      end
    end
    if (io_enq_valids_1) begin
      if (6'h27 == rob_tail) begin
        _T_5936_39_fp_val <= _GEN_311;
      end
    end
    if(_T_6309__T_6332_en & _T_6309__T_6332_mask) begin
      _T_6309[_T_6309__T_6332_addr] <= _T_6309__T_6332_data;
    end
    if(_T_6309__T_6562_en & _T_6309__T_6562_mask) begin
      _T_6309[_T_6309__T_6562_addr] <= _T_6309__T_6562_data;
    end
    if(_T_6309__T_6571_en & _T_6309__T_6571_mask) begin
      _T_6309[_T_6309__T_6571_addr] <= _T_6309__T_6571_data;
    end
    if(_T_6309__T_6652_en & _T_6309__T_6652_mask) begin
      _T_6309[_T_6309__T_6652_addr] <= _T_6309__T_6652_data;
    end
    if(_T_6312__T_6333_en & _T_6312__T_6333_mask) begin
      _T_6312[_T_6312__T_6333_addr] <= _T_6312__T_6333_data;
    end
    if(_T_6312__T_6546_en & _T_6312__T_6546_mask) begin
      _T_6312[_T_6312__T_6546_addr] <= _T_6312__T_6546_data;
    end
    if(_T_6312__T_6554_en & _T_6312__T_6554_mask) begin
      _T_6312[_T_6312__T_6554_addr] <= _T_6312__T_6554_data;
    end
    _T_8115 <= flush_val;
    if (_T_8117) begin
      _T_8120 <= {{24'd0}, io_csr_evec};
    end else begin
      _T_8120 <= flush_pc;
    end
    com_lsu_misspec <= _T_8122;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_0 & _T_3789) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:388 assert (rob_val(rob_tail) === Bool(false),\"[rob] overwriting a valid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_0 & _T_3789) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_0 & _T_3795) begin
          $fwrite(32'h80000002,"Assertion failed\n    at rob.scala:389 assert ((io.enq_uops(w).rob_idx >> log2Ceil(width)) === rob_tail)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_0 & _T_3795) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3860 & _T_3875) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:431 assert (rob_val(cidx) === Bool(true), \"[rob] store writing back to invalid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3860 & _T_3875) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3860 & _T_3883) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:432 assert (rob_bsy(cidx) === Bool(true), \"[rob] store writing back to a not-busy entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3860 & _T_3883) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3887 & _T_3902) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:431 assert (rob_val(cidx) === Bool(true), \"[rob] store writing back to invalid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3887 & _T_3902) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3887 & _T_3910) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:432 assert (rob_bsy(cidx) === Bool(true), \"[rob] store writing back to a not-busy entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3887 & _T_3910) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5120) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5137) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5150) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5197) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5214) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5227) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5274) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5274) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5291) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5304) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5351) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5351) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5368) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5368) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5381) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5381) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5428) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5428) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5445) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5445) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5458) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5458) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_1 & _T_6353) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:388 assert (rob_val(rob_tail) === Bool(false),\"[rob] overwriting a valid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_1 & _T_6353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_enq_valids_1 & _T_6359) begin
          $fwrite(32'h80000002,"Assertion failed\n    at rob.scala:389 assert ((io.enq_uops(w).rob_idx >> log2Ceil(width)) === rob_tail)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_enq_valids_1 & _T_6359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6424 & _T_6439) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:431 assert (rob_val(cidx) === Bool(true), \"[rob] store writing back to invalid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6424 & _T_6439) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6424 & _T_6447) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:432 assert (rob_bsy(cidx) === Bool(true), \"[rob] store writing back to a not-busy entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6424 & _T_6447) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6451 & _T_6466) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:431 assert (rob_val(cidx) === Bool(true), \"[rob] store writing back to invalid entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6451 & _T_6466) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6451 & _T_6474) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:432 assert (rob_bsy(cidx) === Bool(true), \"[rob] store writing back to a not-busy entry.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6451 & _T_6474) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7684) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7684) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7701) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7701) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7714) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7714) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7761) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7761) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7778) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7778) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7791) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7791) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7838) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7838) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7855) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7855) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7868) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7868) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7915) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7915) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7932) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7932) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7945) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7945) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7992) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:580 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7992) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8009) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:583 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8009) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8022) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:586 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8022) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8132) begin
          $fwrite(32'h80000002,"Assertion failed: [rob] pipeline flush not be excercised during a LSU misspeculation\n    at rob.scala:668 assert (!(com_lsu_misspec && !io.flush.valid), \"[rob] pipeline flush not be excercised during a LSU misspeculation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8165) begin
          $fwrite(32'h80000002,"Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:686 assert (!(io.commit.valids(w) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8177) begin
          $fwrite(32'h80000002,"Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:690 assert (!(io.commit.valids(w) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8196) begin
          $fwrite(32'h80000002,"Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:686 assert (!(io.commit.valids(w) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8208) begin
          $fwrite(32'h80000002,"Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:690 assert (!(io.commit.valids(w) &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8317) begin
          $fwrite(32'h80000002,"Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:753 assert (!(exception_thrown && !io.cxcpt.valid && !r_xcpt_val),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8324) begin
          $fwrite(32'h80000002,"Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:756 assert (!(io.empty && r_xcpt_val),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8324) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8334) begin
          $fwrite(32'h80000002,"Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:759 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_8334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  input  [11:0] io_decode_0_csr,
  output        io_decode_0_fp_illegal,
  output        io_decode_0_read_illegal,
  output        io_decode_0_write_illegal,
  output        io_decode_0_write_flush,
  output        io_decode_0_system_illegal,
  input  [11:0] io_decode_1_csr,
  output        io_decode_1_fp_illegal,
  output        io_decode_1_read_illegal,
  output        io_decode_1_write_illegal,
  output        io_decode_1_write_flush,
  output        io_decode_1_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_hpp,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [3:0]  io_ptbr_mode,
  output [43:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input         io_exception,
  input  [1:0]  io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_badaddr,
  output [2:0]  io_fcsr_rm,
  input         io_fcsr_flags_valid,
  input  [4:0]  io_fcsr_flags_bits,
  output        io_interrupt,
  output [63:0] io_interrupt_cause,
  output [63:0] io_counters_0_eventSel,
  input  [1:0]  io_counters_0_inc,
  output [63:0] io_counters_1_eventSel,
  input  [1:0]  io_counters_1_inc,
  output [63:0] io_counters_2_eventSel,
  input  [1:0]  io_counters_2_inc,
  output [63:0] io_counters_3_eventSel,
  input  [1:0]  io_counters_3_inc,
  output [63:0] io_counters_4_eventSel,
  input  [1:0]  io_counters_4_inc,
  output [63:0] io_counters_5_eventSel,
  input  [1:0]  io_counters_5_inc,
  output [63:0] io_counters_6_eventSel,
  input  [1:0]  io_counters_6_inc,
  output [63:0] io_counters_7_eventSel,
  input  [1:0]  io_counters_7_inc,
  output [63:0] io_counters_8_eventSel,
  input  [1:0]  io_counters_8_inc,
  output [63:0] io_counters_9_eventSel,
  input  [1:0]  io_counters_9_inc,
  output [63:0] io_counters_10_eventSel,
  input  [1:0]  io_counters_10_inc,
  output [63:0] io_counters_11_eventSel,
  input  [1:0]  io_counters_11_inc,
  output [63:0] io_counters_12_eventSel,
  input  [1:0]  io_counters_12_inc,
  output [63:0] io_counters_13_eventSel,
  input  [1:0]  io_counters_13_inc,
  output [63:0] io_counters_14_eventSel,
  input  [1:0]  io_counters_14_inc,
  output [63:0] io_counters_15_eventSel,
  input  [1:0]  io_counters_15_inc,
  output [63:0] io_counters_16_eventSel,
  input  [1:0]  io_counters_16_inc,
  output [63:0] io_counters_17_eventSel,
  input  [1:0]  io_counters_17_inc,
  output [63:0] io_counters_18_eventSel,
  input  [1:0]  io_counters_18_inc,
  output [63:0] io_counters_19_eventSel,
  input  [1:0]  io_counters_19_inc,
  output [63:0] io_counters_20_eventSel,
  input  [1:0]  io_counters_20_inc,
  output [63:0] io_counters_21_eventSel,
  input  [1:0]  io_counters_21_inc,
  output [63:0] io_counters_22_eventSel,
  input  [1:0]  io_counters_22_inc,
  output [63:0] io_counters_23_eventSel,
  input  [1:0]  io_counters_23_inc,
  output [63:0] io_counters_24_eventSel,
  input  [1:0]  io_counters_24_inc,
  output [63:0] io_counters_25_eventSel,
  input  [1:0]  io_counters_25_inc,
  output [63:0] io_counters_26_eventSel,
  input  [1:0]  io_counters_26_inc,
  output [63:0] io_counters_27_eventSel,
  input  [1:0]  io_counters_27_inc,
  output [63:0] io_counters_28_eventSel,
  input  [1:0]  io_counters_28_inc
);
  reg [1:0] reg_mstatus_prv;
  reg [31:0] _RAND_0;
  reg  reg_mstatus_tsr;
  reg [31:0] _RAND_1;
  reg  reg_mstatus_tw;
  reg [31:0] _RAND_2;
  reg  reg_mstatus_tvm;
  reg [31:0] _RAND_3;
  reg  reg_mstatus_mxr;
  reg [31:0] _RAND_4;
  reg  reg_mstatus_sum;
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mprv;
  reg [31:0] _RAND_6;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] _RAND_7;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] _RAND_8;
  reg  reg_mstatus_spp;
  reg [31:0] _RAND_9;
  reg  reg_mstatus_mpie;
  reg [31:0] _RAND_10;
  reg  reg_mstatus_spie;
  reg [31:0] _RAND_11;
  reg  reg_mstatus_mie;
  reg [31:0] _RAND_12;
  reg  reg_mstatus_sie;
  reg [31:0] _RAND_13;
  wire [1:0] new_prv;
  wire  _T_194;
  wire [1:0] _T_196;
  reg  reg_dcsr_ebreakm;
  reg [31:0] _RAND_14;
  reg  reg_dcsr_ebreaks;
  reg [31:0] _RAND_15;
  reg  reg_dcsr_ebreaku;
  reg [31:0] _RAND_16;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] _RAND_17;
  reg  reg_dcsr_step;
  reg [31:0] _RAND_18;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] _RAND_19;
  reg  reg_debug;
  reg [31:0] _RAND_20;
  reg [39:0] reg_dpc;
  reg [63:0] _RAND_21;
  reg [63:0] reg_dscratch;
  reg [63:0] _RAND_22;
  reg  reg_singleStepped;
  reg [31:0] _RAND_23;
  reg  reg_bp_0_control_dmode;
  reg [31:0] _RAND_24;
  reg  reg_bp_0_control_action;
  reg [31:0] _RAND_25;
  reg [1:0] reg_bp_0_control_tmatch;
  reg [31:0] _RAND_26;
  reg  reg_bp_0_control_m;
  reg [31:0] _RAND_27;
  reg  reg_bp_0_control_s;
  reg [31:0] _RAND_28;
  reg  reg_bp_0_control_u;
  reg [31:0] _RAND_29;
  reg  reg_bp_0_control_x;
  reg [31:0] _RAND_30;
  reg  reg_bp_0_control_w;
  reg [31:0] _RAND_31;
  reg  reg_bp_0_control_r;
  reg [31:0] _RAND_32;
  reg [38:0] reg_bp_0_address;
  reg [63:0] _RAND_33;
  reg [63:0] reg_mie;
  reg [63:0] _RAND_34;
  reg [63:0] reg_mideleg;
  reg [63:0] _RAND_35;
  reg [63:0] reg_medeleg;
  reg [63:0] _RAND_36;
  reg  reg_mip_seip;
  reg [31:0] _RAND_37;
  reg  reg_mip_stip;
  reg [31:0] _RAND_38;
  reg  reg_mip_ssip;
  reg [31:0] _RAND_39;
  reg [39:0] reg_mepc;
  reg [63:0] _RAND_40;
  reg [63:0] reg_mcause;
  reg [63:0] _RAND_41;
  reg [39:0] reg_mbadaddr;
  reg [63:0] _RAND_42;
  reg [63:0] reg_mscratch;
  reg [63:0] _RAND_43;
  reg [31:0] reg_mtvec;
  reg [31:0] _RAND_44;
  reg [31:0] reg_mcounteren;
  reg [31:0] _RAND_45;
  reg [31:0] reg_scounteren;
  reg [31:0] _RAND_46;
  reg [39:0] reg_sepc;
  reg [63:0] _RAND_47;
  reg [63:0] reg_scause;
  reg [63:0] _RAND_48;
  reg [39:0] reg_sbadaddr;
  reg [63:0] _RAND_49;
  reg [63:0] reg_sscratch;
  reg [63:0] _RAND_50;
  reg [38:0] reg_stvec;
  reg [63:0] _RAND_51;
  reg [3:0] reg_sptbr_mode;
  reg [31:0] _RAND_52;
  reg [43:0] reg_sptbr_ppn;
  reg [63:0] _RAND_53;
  reg  reg_wfi;
  reg [31:0] _RAND_54;
  reg [4:0] reg_fflags;
  reg [31:0] _RAND_55;
  reg [2:0] reg_frm;
  reg [31:0] _RAND_56;
  reg [5:0] _T_328;
  reg [31:0] _RAND_57;
  wire [5:0] _GEN_0;
  wire [6:0] _T_329;
  reg [57:0] _T_332;
  reg [63:0] _RAND_58;
  wire  _T_333;
  wire [58:0] _T_335;
  wire [57:0] _T_336;
  wire [57:0] _GEN_36;
  wire [63:0] _T_337;
  reg [5:0] _T_341;
  reg [31:0] _RAND_59;
  wire [6:0] _T_342;
  reg [57:0] _T_345;
  reg [63:0] _RAND_60;
  wire  _T_346;
  wire [58:0] _T_348;
  wire [57:0] _T_349;
  wire [57:0] _GEN_37;
  wire [63:0] _T_350;
  reg [63:0] reg_hpmevent_0;
  reg [63:0] _RAND_61;
  reg [63:0] reg_hpmevent_1;
  reg [63:0] _RAND_62;
  reg [63:0] reg_hpmevent_2;
  reg [63:0] _RAND_63;
  reg [63:0] reg_hpmevent_3;
  reg [63:0] _RAND_64;
  reg [63:0] reg_hpmevent_4;
  reg [63:0] _RAND_65;
  reg [63:0] reg_hpmevent_5;
  reg [63:0] _RAND_66;
  reg [63:0] reg_hpmevent_6;
  reg [63:0] _RAND_67;
  reg [63:0] reg_hpmevent_7;
  reg [63:0] _RAND_68;
  reg [63:0] reg_hpmevent_8;
  reg [63:0] _RAND_69;
  reg [63:0] reg_hpmevent_9;
  reg [63:0] _RAND_70;
  reg [63:0] reg_hpmevent_10;
  reg [63:0] _RAND_71;
  reg [63:0] reg_hpmevent_11;
  reg [63:0] _RAND_72;
  reg [63:0] reg_hpmevent_12;
  reg [63:0] _RAND_73;
  reg [63:0] reg_hpmevent_13;
  reg [63:0] _RAND_74;
  reg [63:0] reg_hpmevent_14;
  reg [63:0] _RAND_75;
  reg [63:0] reg_hpmevent_15;
  reg [63:0] _RAND_76;
  reg [63:0] reg_hpmevent_16;
  reg [63:0] _RAND_77;
  reg [63:0] reg_hpmevent_17;
  reg [63:0] _RAND_78;
  reg [63:0] reg_hpmevent_18;
  reg [63:0] _RAND_79;
  reg [63:0] reg_hpmevent_19;
  reg [63:0] _RAND_80;
  reg [63:0] reg_hpmevent_20;
  reg [63:0] _RAND_81;
  reg [63:0] reg_hpmevent_21;
  reg [63:0] _RAND_82;
  reg [63:0] reg_hpmevent_22;
  reg [63:0] _RAND_83;
  reg [63:0] reg_hpmevent_23;
  reg [63:0] _RAND_84;
  reg [63:0] reg_hpmevent_24;
  reg [63:0] _RAND_85;
  reg [63:0] reg_hpmevent_25;
  reg [63:0] _RAND_86;
  reg [63:0] reg_hpmevent_26;
  reg [63:0] _RAND_87;
  reg [63:0] reg_hpmevent_27;
  reg [63:0] _RAND_88;
  reg [63:0] reg_hpmevent_28;
  reg [63:0] _RAND_89;
  reg [5:0] _T_410;
  reg [31:0] _RAND_90;
  wire [5:0] _GEN_1;
  wire [6:0] _T_411;
  reg [33:0] _T_413;
  reg [63:0] _RAND_91;
  wire  _T_414;
  wire [34:0] _T_416;
  wire [33:0] _T_417;
  wire [33:0] _GEN_38;
  wire [39:0] _T_418;
  reg [5:0] _T_420;
  reg [31:0] _RAND_92;
  wire [5:0] _GEN_2;
  wire [6:0] _T_421;
  reg [33:0] _T_423;
  reg [63:0] _RAND_93;
  wire  _T_424;
  wire [34:0] _T_426;
  wire [33:0] _T_427;
  wire [33:0] _GEN_39;
  wire [39:0] _T_428;
  reg [5:0] _T_430;
  reg [31:0] _RAND_94;
  wire [5:0] _GEN_3;
  wire [6:0] _T_431;
  reg [33:0] _T_433;
  reg [63:0] _RAND_95;
  wire  _T_434;
  wire [34:0] _T_436;
  wire [33:0] _T_437;
  wire [33:0] _GEN_40;
  wire [39:0] _T_438;
  reg [5:0] _T_440;
  reg [31:0] _RAND_96;
  wire [5:0] _GEN_4;
  wire [6:0] _T_441;
  reg [33:0] _T_443;
  reg [63:0] _RAND_97;
  wire  _T_444;
  wire [34:0] _T_446;
  wire [33:0] _T_447;
  wire [33:0] _GEN_41;
  wire [39:0] _T_448;
  reg [5:0] _T_450;
  reg [31:0] _RAND_98;
  wire [5:0] _GEN_5;
  wire [6:0] _T_451;
  reg [33:0] _T_453;
  reg [63:0] _RAND_99;
  wire  _T_454;
  wire [34:0] _T_456;
  wire [33:0] _T_457;
  wire [33:0] _GEN_42;
  wire [39:0] _T_458;
  reg [5:0] _T_460;
  reg [31:0] _RAND_100;
  wire [5:0] _GEN_6;
  wire [6:0] _T_461;
  reg [33:0] _T_463;
  reg [63:0] _RAND_101;
  wire  _T_464;
  wire [34:0] _T_466;
  wire [33:0] _T_467;
  wire [33:0] _GEN_43;
  wire [39:0] _T_468;
  reg [5:0] _T_470;
  reg [31:0] _RAND_102;
  wire [5:0] _GEN_7;
  wire [6:0] _T_471;
  reg [33:0] _T_473;
  reg [63:0] _RAND_103;
  wire  _T_474;
  wire [34:0] _T_476;
  wire [33:0] _T_477;
  wire [33:0] _GEN_44;
  wire [39:0] _T_478;
  reg [5:0] _T_480;
  reg [31:0] _RAND_104;
  wire [5:0] _GEN_8;
  wire [6:0] _T_481;
  reg [33:0] _T_483;
  reg [63:0] _RAND_105;
  wire  _T_484;
  wire [34:0] _T_486;
  wire [33:0] _T_487;
  wire [33:0] _GEN_45;
  wire [39:0] _T_488;
  reg [5:0] _T_490;
  reg [31:0] _RAND_106;
  wire [5:0] _GEN_9;
  wire [6:0] _T_491;
  reg [33:0] _T_493;
  reg [63:0] _RAND_107;
  wire  _T_494;
  wire [34:0] _T_496;
  wire [33:0] _T_497;
  wire [33:0] _GEN_46;
  wire [39:0] _T_498;
  reg [5:0] _T_500;
  reg [31:0] _RAND_108;
  wire [5:0] _GEN_10;
  wire [6:0] _T_501;
  reg [33:0] _T_503;
  reg [63:0] _RAND_109;
  wire  _T_504;
  wire [34:0] _T_506;
  wire [33:0] _T_507;
  wire [33:0] _GEN_47;
  wire [39:0] _T_508;
  reg [5:0] _T_510;
  reg [31:0] _RAND_110;
  wire [5:0] _GEN_11;
  wire [6:0] _T_511;
  reg [33:0] _T_513;
  reg [63:0] _RAND_111;
  wire  _T_514;
  wire [34:0] _T_516;
  wire [33:0] _T_517;
  wire [33:0] _GEN_48;
  wire [39:0] _T_518;
  reg [5:0] _T_520;
  reg [31:0] _RAND_112;
  wire [5:0] _GEN_12;
  wire [6:0] _T_521;
  reg [33:0] _T_523;
  reg [63:0] _RAND_113;
  wire  _T_524;
  wire [34:0] _T_526;
  wire [33:0] _T_527;
  wire [33:0] _GEN_49;
  wire [39:0] _T_528;
  reg [5:0] _T_530;
  reg [31:0] _RAND_114;
  wire [5:0] _GEN_13;
  wire [6:0] _T_531;
  reg [33:0] _T_533;
  reg [63:0] _RAND_115;
  wire  _T_534;
  wire [34:0] _T_536;
  wire [33:0] _T_537;
  wire [33:0] _GEN_50;
  wire [39:0] _T_538;
  reg [5:0] _T_540;
  reg [31:0] _RAND_116;
  wire [5:0] _GEN_14;
  wire [6:0] _T_541;
  reg [33:0] _T_543;
  reg [63:0] _RAND_117;
  wire  _T_544;
  wire [34:0] _T_546;
  wire [33:0] _T_547;
  wire [33:0] _GEN_51;
  wire [39:0] _T_548;
  reg [5:0] _T_550;
  reg [31:0] _RAND_118;
  wire [5:0] _GEN_15;
  wire [6:0] _T_551;
  reg [33:0] _T_553;
  reg [63:0] _RAND_119;
  wire  _T_554;
  wire [34:0] _T_556;
  wire [33:0] _T_557;
  wire [33:0] _GEN_52;
  wire [39:0] _T_558;
  reg [5:0] _T_560;
  reg [31:0] _RAND_120;
  wire [5:0] _GEN_16;
  wire [6:0] _T_561;
  reg [33:0] _T_563;
  reg [63:0] _RAND_121;
  wire  _T_564;
  wire [34:0] _T_566;
  wire [33:0] _T_567;
  wire [33:0] _GEN_53;
  wire [39:0] _T_568;
  reg [5:0] _T_570;
  reg [31:0] _RAND_122;
  wire [5:0] _GEN_17;
  wire [6:0] _T_571;
  reg [33:0] _T_573;
  reg [63:0] _RAND_123;
  wire  _T_574;
  wire [34:0] _T_576;
  wire [33:0] _T_577;
  wire [33:0] _GEN_54;
  wire [39:0] _T_578;
  reg [5:0] _T_580;
  reg [31:0] _RAND_124;
  wire [5:0] _GEN_589;
  wire [6:0] _T_581;
  reg [33:0] _T_583;
  reg [63:0] _RAND_125;
  wire  _T_584;
  wire [34:0] _T_586;
  wire [33:0] _T_587;
  wire [33:0] _GEN_55;
  wire [39:0] _T_588;
  reg [5:0] _T_590;
  reg [31:0] _RAND_126;
  wire [5:0] _GEN_590;
  wire [6:0] _T_591;
  reg [33:0] _T_593;
  reg [63:0] _RAND_127;
  wire  _T_594;
  wire [34:0] _T_596;
  wire [33:0] _T_597;
  wire [33:0] _GEN_56;
  wire [39:0] _T_598;
  reg [5:0] _T_600;
  reg [31:0] _RAND_128;
  wire [5:0] _GEN_591;
  wire [6:0] _T_601;
  reg [33:0] _T_603;
  reg [63:0] _RAND_129;
  wire  _T_604;
  wire [34:0] _T_606;
  wire [33:0] _T_607;
  wire [33:0] _GEN_57;
  wire [39:0] _T_608;
  reg [5:0] _T_610;
  reg [31:0] _RAND_130;
  wire [5:0] _GEN_592;
  wire [6:0] _T_611;
  reg [33:0] _T_613;
  reg [63:0] _RAND_131;
  wire  _T_614;
  wire [34:0] _T_616;
  wire [33:0] _T_617;
  wire [33:0] _GEN_58;
  wire [39:0] _T_618;
  reg [5:0] _T_620;
  reg [31:0] _RAND_132;
  wire [5:0] _GEN_593;
  wire [6:0] _T_621;
  reg [33:0] _T_623;
  reg [63:0] _RAND_133;
  wire  _T_624;
  wire [34:0] _T_626;
  wire [33:0] _T_627;
  wire [33:0] _GEN_59;
  wire [39:0] _T_628;
  reg [5:0] _T_630;
  reg [31:0] _RAND_134;
  wire [5:0] _GEN_594;
  wire [6:0] _T_631;
  reg [33:0] _T_633;
  reg [63:0] _RAND_135;
  wire  _T_634;
  wire [34:0] _T_636;
  wire [33:0] _T_637;
  wire [33:0] _GEN_60;
  wire [39:0] _T_638;
  reg [5:0] _T_640;
  reg [31:0] _RAND_136;
  wire [5:0] _GEN_595;
  wire [6:0] _T_641;
  reg [33:0] _T_643;
  reg [63:0] _RAND_137;
  wire  _T_644;
  wire [34:0] _T_646;
  wire [33:0] _T_647;
  wire [33:0] _GEN_61;
  wire [39:0] _T_648;
  reg [5:0] _T_650;
  reg [31:0] _RAND_138;
  wire [5:0] _GEN_596;
  wire [6:0] _T_651;
  reg [33:0] _T_653;
  reg [63:0] _RAND_139;
  wire  _T_654;
  wire [34:0] _T_656;
  wire [33:0] _T_657;
  wire [33:0] _GEN_62;
  wire [39:0] _T_658;
  reg [5:0] _T_660;
  reg [31:0] _RAND_140;
  wire [5:0] _GEN_597;
  wire [6:0] _T_661;
  reg [33:0] _T_663;
  reg [63:0] _RAND_141;
  wire  _T_664;
  wire [34:0] _T_666;
  wire [33:0] _T_667;
  wire [33:0] _GEN_63;
  wire [39:0] _T_668;
  reg [5:0] _T_670;
  reg [31:0] _RAND_142;
  wire [5:0] _GEN_598;
  wire [6:0] _T_671;
  reg [33:0] _T_673;
  reg [63:0] _RAND_143;
  wire  _T_674;
  wire [34:0] _T_676;
  wire [33:0] _T_677;
  wire [33:0] _GEN_64;
  wire [39:0] _T_678;
  reg [5:0] _T_680;
  reg [31:0] _RAND_144;
  wire [5:0] _GEN_599;
  wire [6:0] _T_681;
  reg [33:0] _T_683;
  reg [63:0] _RAND_145;
  wire  _T_684;
  wire [34:0] _T_686;
  wire [33:0] _T_687;
  wire [33:0] _GEN_65;
  wire [39:0] _T_688;
  reg [5:0] _T_690;
  reg [31:0] _RAND_146;
  wire [5:0] _GEN_600;
  wire [6:0] _T_691;
  reg [33:0] _T_693;
  reg [63:0] _RAND_147;
  wire  _T_694;
  wire [34:0] _T_696;
  wire [33:0] _T_697;
  wire [33:0] _GEN_66;
  wire [39:0] _T_698;
  wire  _T_701;
  wire [31:0] _T_704;
  wire [31:0] hpm_mask;
  wire  mip_meip;
  wire  mip_seip;
  wire  mip_mtip;
  wire  mip_stip;
  wire  mip_msip;
  wire  mip_ssip;
  reg  _T_711;
  reg [31:0] _RAND_148;
  wire  _T_712;
  wire [1:0] _T_713;
  wire [1:0] _T_714;
  wire [3:0] _T_715;
  wire [1:0] _T_716;
  wire [1:0] _T_717;
  wire [3:0] _T_718;
  wire [7:0] _T_719;
  wire [1:0] _T_720;
  wire [1:0] _T_721;
  wire [3:0] _T_722;
  wire [7:0] _T_726;
  wire [15:0] _T_727;
  wire [15:0] read_mip;
  wire [63:0] _GEN_601;
  wire [63:0] pending_interrupts;
  wire [14:0] _GEN_602;
  wire [14:0] d_interrupts;
  wire  _T_730;
  wire  _T_731;
  wire [63:0] _T_732;
  wire [63:0] _T_733;
  wire [63:0] _T_734;
  wire [63:0] m_interrupts;
  wire  _T_737;
  wire  _T_740;
  wire  _T_741;
  wire [63:0] _T_742;
  wire [63:0] s_interrupts;
  wire  _T_744;
  wire  _T_745;
  wire  _T_746;
  wire  _T_747;
  wire  _T_748;
  wire  _T_749;
  wire  _T_750;
  wire  _T_751;
  wire  _T_752;
  wire  _T_753;
  wire  _T_754;
  wire  _T_755;
  wire  _T_756;
  wire  _T_757;
  wire  _T_758;
  wire  _T_759;
  wire  _T_760;
  wire  _T_761;
  wire  _T_762;
  wire  _T_763;
  wire  _T_764;
  wire  _T_765;
  wire  _T_766;
  wire  _T_767;
  wire  _T_768;
  wire  _T_769;
  wire  _T_770;
  wire  _T_771;
  wire  _T_772;
  wire  _T_773;
  wire  _T_774;
  wire  _T_775;
  wire  _T_776;
  wire  _T_777;
  wire  _T_778;
  wire  _T_779;
  wire  _T_780;
  wire  _T_781;
  wire  _T_782;
  wire  _T_783;
  wire  _T_784;
  wire  _T_785;
  wire  _T_786;
  wire  _T_787;
  wire  _T_788;
  wire  _T_789;
  wire  _T_790;
  wire  _T_791;
  wire  _T_792;
  wire  _T_793;
  wire  _T_794;
  wire  _T_795;
  wire  _T_796;
  wire  _T_797;
  wire  _T_798;
  wire  _T_799;
  wire  _T_800;
  wire  _T_801;
  wire  _T_802;
  wire  _T_803;
  wire  _T_804;
  wire  _T_805;
  wire  _T_806;
  wire  _T_807;
  wire  _T_808;
  wire  _T_809;
  wire  _T_810;
  wire  _T_811;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_817;
  wire  anyInterrupt;
  wire [2:0] _T_894;
  wire [3:0] _T_895;
  wire [3:0] _T_896;
  wire [3:0] _T_897;
  wire [3:0] _T_898;
  wire [3:0] _T_899;
  wire [3:0] _T_900;
  wire [3:0] _T_901;
  wire [3:0] _T_902;
  wire [3:0] _T_903;
  wire [3:0] _T_904;
  wire [3:0] _T_905;
  wire [3:0] _T_906;
  wire [3:0] _T_907;
  wire [3:0] _T_908;
  wire [3:0] _T_909;
  wire [3:0] _T_910;
  wire [3:0] _T_911;
  wire [3:0] _T_912;
  wire [3:0] _T_913;
  wire [3:0] _T_914;
  wire [3:0] _T_915;
  wire [3:0] _T_916;
  wire [3:0] _T_917;
  wire [3:0] _T_918;
  wire [3:0] _T_919;
  wire [3:0] _T_920;
  wire [3:0] _T_921;
  wire [3:0] _T_922;
  wire [3:0] _T_923;
  wire [3:0] _T_924;
  wire [3:0] _T_925;
  wire [3:0] _T_926;
  wire [3:0] _T_927;
  wire [3:0] _T_928;
  wire [3:0] _T_929;
  wire [3:0] whichInterrupt;
  wire [63:0] _GEN_603;
  wire [64:0] _T_931;
  wire [63:0] interruptCause;
  wire  _T_933;
  wire  _T_934;
  wire  _T_936;
  wire  _T_937;
  wire  _T_938;
  reg [63:0] reg_misa;
  reg [63:0] _RAND_149;
  wire [1:0] _T_941;
  wire [2:0] _T_942;
  wire [1:0] _T_943;
  wire [1:0] _T_944;
  wire [3:0] _T_945;
  wire [6:0] _T_946;
  wire [2:0] _T_947;
  wire [3:0] _T_948;
  wire [3:0] _T_949;
  wire [2:0] _T_950;
  wire [6:0] _T_951;
  wire [10:0] _T_952;
  wire [17:0] _T_953;
  wire [1:0] _T_954;
  wire [2:0] _T_955;
  wire [1:0] _T_956;
  wire [8:0] _T_957;
  wire [10:0] _T_958;
  wire [13:0] _T_959;
  wire [3:0] _T_960;
  wire [27:0] _T_961;
  wire [31:0] _T_962;
  wire [3:0] _T_963;
  wire [32:0] _T_964;
  wire [36:0] _T_965;
  wire [68:0] _T_966;
  wire [82:0] _T_967;
  wire [100:0] _T_968;
  wire [63:0] read_mstatus;
  wire  _GEN_0_control_x;
  wire  _GEN_1_control_w;
  wire [1:0] _T_970;
  wire  _GEN_2_control_r;
  wire [2:0] _T_971;
  wire  _GEN_3_control_s;
  wire  _GEN_4_control_u;
  wire [1:0] _T_972;
  wire  _GEN_5_control_m;
  wire [1:0] _T_973;
  wire [3:0] _T_974;
  wire [6:0] _T_975;
  wire [1:0] _GEN_8_control_tmatch;
  wire [3:0] _T_976;
  wire  _GEN_9_control_action;
  wire [1:0] _T_977;
  wire [5:0] _T_978;
  wire  _GEN_14_control_dmode;
  wire [4:0] _T_980;
  wire [50:0] _T_981;
  wire [56:0] _T_982;
  wire [63:0] _T_983;
  wire [38:0] _GEN_15_address;
  wire  _T_985;
  wire [24:0] _T_989;
  wire [38:0] _GEN_16_address;
  wire [63:0] _T_990;
  wire  _T_994;
  wire [23:0] _T_998;
  wire [63:0] _T_999;
  wire  _T_1000;
  wire [23:0] _T_1004;
  wire [63:0] _T_1005;
  wire [3:0] _T_1006;
  wire [5:0] _T_1007;
  wire [3:0] _T_1008;
  wire [5:0] _T_1010;
  wire [11:0] _T_1011;
  wire [1:0] _T_1012;
  wire [2:0] _T_1013;
  wire [12:0] _T_1014;
  wire [16:0] _T_1016;
  wire [19:0] _T_1017;
  wire [31:0] _T_1018;
  wire [7:0] _T_1019;
  wire [63:0] _T_1022;
  wire [63:0] _T_1023;
  wire  _T_1060_sd;
  wire [1:0] _T_1060_uxl;
  wire  _T_1060_sd_rv32;
  wire  _T_1060_mxr;
  wire  _T_1060_sum;
  wire [1:0] _T_1060_xs;
  wire [1:0] _T_1060_fs;
  wire  _T_1060_spp;
  wire  _T_1060_spie;
  wire  _T_1060_sie;
  wire [1:0] _T_1061;
  wire [2:0] _T_1062;
  wire [1:0] _T_1064;
  wire [3:0] _T_1065;
  wire [6:0] _T_1066;
  wire [2:0] _T_1067;
  wire [3:0] _T_1068;
  wire [3:0] _T_1069;
  wire [2:0] _T_1070;
  wire [6:0] _T_1071;
  wire [10:0] _T_1072;
  wire [17:0] _T_1073;
  wire [1:0] _T_1074;
  wire [2:0] _T_1075;
  wire [8:0] _T_1077;
  wire [10:0] _T_1078;
  wire [13:0] _T_1079;
  wire [3:0] _T_1080;
  wire [27:0] _T_1081;
  wire [31:0] _T_1082;
  wire [68:0] _T_1086;
  wire [82:0] _T_1087;
  wire [100:0] _T_1088;
  wire [63:0] _T_1089;
  wire  _T_1090;
  wire [23:0] _T_1094;
  wire [63:0] _T_1095;
  wire [19:0] _T_1096;
  wire [63:0] _T_1097;
  wire  _T_1098;
  wire [23:0] _T_1102;
  wire [63:0] _T_1103;
  wire  _T_1104;
  wire [24:0] _T_1108;
  wire [63:0] _T_1109;
  wire  _T_1114;
  wire  _T_1116;
  wire  _T_1124;
  wire  _T_1126;
  wire  _T_1128;
  wire  _T_1130;
  wire  _T_1132;
  wire  _T_1134;
  wire  _T_1136;
  wire  _T_1138;
  wire  _T_1140;
  wire  _T_1144;
  wire  _T_1146;
  wire  _T_1148;
  wire  _T_1150;
  wire  _T_1152;
  wire  _T_1154;
  wire  _T_1156;
  wire  _T_1158;
  wire  _T_1160;
  wire  _T_1162;
  wire  _T_1164;
  wire  _T_1166;
  wire  _T_1168;
  wire  _T_1170;
  wire  _T_1172;
  wire  _T_1174;
  wire  _T_1176;
  wire  _T_1178;
  wire  _T_1180;
  wire  _T_1182;
  wire  _T_1184;
  wire  _T_1186;
  wire  _T_1188;
  wire  _T_1190;
  wire  _T_1192;
  wire  _T_1194;
  wire  _T_1196;
  wire  _T_1198;
  wire  _T_1200;
  wire  _T_1202;
  wire  _T_1204;
  wire  _T_1206;
  wire  _T_1208;
  wire  _T_1210;
  wire  _T_1212;
  wire  _T_1214;
  wire  _T_1216;
  wire  _T_1218;
  wire  _T_1220;
  wire  _T_1222;
  wire  _T_1224;
  wire  _T_1226;
  wire  _T_1228;
  wire  _T_1230;
  wire  _T_1232;
  wire  _T_1234;
  wire  _T_1236;
  wire  _T_1238;
  wire  _T_1240;
  wire  _T_1242;
  wire  _T_1244;
  wire  _T_1246;
  wire  _T_1248;
  wire  _T_1250;
  wire  _T_1252;
  wire  _T_1254;
  wire  _T_1256;
  wire  _T_1258;
  wire  _T_1260;
  wire  _T_1262;
  wire  _T_1264;
  wire  _T_1266;
  wire  _T_1268;
  wire  _T_1270;
  wire  _T_1272;
  wire  _T_1274;
  wire  _T_1276;
  wire  _T_1278;
  wire  _T_1280;
  wire  _T_1282;
  wire  _T_1284;
  wire  _T_1286;
  wire  _T_1288;
  wire  _T_1290;
  wire  _T_1292;
  wire  _T_1294;
  wire  _T_1296;
  wire  _T_1298;
  wire  _T_1300;
  wire  _T_1302;
  wire  _T_1304;
  wire  _T_1306;
  wire  _T_1308;
  wire  _T_1310;
  wire  _T_1312;
  wire  _T_1314;
  wire  _T_1316;
  wire  _T_1318;
  wire  _T_1320;
  wire  _T_1322;
  wire  _T_1324;
  wire  _T_1326;
  wire  _T_1328;
  wire  _T_1330;
  wire  _T_1332;
  wire  _T_1334;
  wire  _T_1336;
  wire  _T_1338;
  wire  _T_1340;
  wire  _T_1342;
  wire  _T_1344;
  wire  _T_1346;
  wire  _T_1348;
  wire  _T_1350;
  wire  _T_1352;
  wire  _T_1354;
  wire  _T_1356;
  wire  _T_1358;
  wire  _T_1360;
  wire  _T_1362;
  wire  _T_1365;
  wire  _T_1366;
  wire  _T_1367;
  wire [63:0] _T_1369;
  wire [63:0] _T_1370;
  wire [63:0] _T_1374;
  wire [63:0] _T_1375;
  wire [63:0] wdata;
  wire  system_insn;
  wire [2:0] _T_1378;
  wire [7:0] opcode;
  wire  _T_1379;
  wire  insn_call;
  wire  _T_1380;
  wire  insn_break;
  wire  _T_1381;
  wire  insn_ret;
  wire  _T_1382;
  wire  insn_wfi;
  wire  _T_1385;
  wire  _T_1388;
  wire  _T_1389;
  wire  _T_1395;
  wire  _T_1396;
  wire  _T_1402;
  wire  _T_1403;
  wire  _T_1405;
  wire  _T_1406;
  wire  _T_1408;
  wire  _T_1409;
  wire [1:0] _T_1416;
  wire  _T_1417;
  wire  _T_1419;
  wire  _T_1421;
  wire  _T_1423;
  wire  _T_1425;
  wire  _T_1427;
  wire  _T_1429;
  wire  _T_1431;
  wire  _T_1433;
  wire  _T_1435;
  wire  _T_1437;
  wire  _T_1439;
  wire  _T_1441;
  wire  _T_1443;
  wire  _T_1445;
  wire  _T_1447;
  wire  _T_1449;
  wire  _T_1451;
  wire  _T_1453;
  wire  _T_1455;
  wire  _T_1457;
  wire  _T_1459;
  wire  _T_1461;
  wire  _T_1463;
  wire  _T_1465;
  wire  _T_1467;
  wire  _T_1469;
  wire  _T_1471;
  wire  _T_1473;
  wire  _T_1475;
  wire  _T_1477;
  wire  _T_1479;
  wire  _T_1481;
  wire  _T_1483;
  wire  _T_1485;
  wire  _T_1487;
  wire  _T_1489;
  wire  _T_1491;
  wire  _T_1493;
  wire  _T_1495;
  wire  _T_1497;
  wire  _T_1499;
  wire  _T_1501;
  wire  _T_1503;
  wire  _T_1505;
  wire  _T_1507;
  wire  _T_1509;
  wire  _T_1511;
  wire  _T_1513;
  wire  _T_1515;
  wire  _T_1517;
  wire  _T_1519;
  wire  _T_1521;
  wire  _T_1523;
  wire  _T_1525;
  wire  _T_1527;
  wire  _T_1529;
  wire  _T_1531;
  wire  _T_1533;
  wire  _T_1535;
  wire  _T_1537;
  wire  _T_1539;
  wire  _T_1541;
  wire  _T_1543;
  wire  _T_1545;
  wire  _T_1547;
  wire  _T_1549;
  wire  _T_1551;
  wire  _T_1553;
  wire  _T_1555;
  wire  _T_1557;
  wire  _T_1559;
  wire  _T_1561;
  wire  _T_1563;
  wire  _T_1565;
  wire  _T_1567;
  wire  _T_1569;
  wire  _T_1571;
  wire  _T_1573;
  wire  _T_1575;
  wire  _T_1577;
  wire  _T_1579;
  wire  _T_1581;
  wire  _T_1583;
  wire  _T_1585;
  wire  _T_1587;
  wire  _T_1589;
  wire  _T_1591;
  wire  _T_1593;
  wire  _T_1595;
  wire  _T_1597;
  wire  _T_1599;
  wire  _T_1601;
  wire  _T_1603;
  wire  _T_1605;
  wire  _T_1607;
  wire  _T_1609;
  wire  _T_1611;
  wire  _T_1613;
  wire  _T_1615;
  wire  _T_1617;
  wire  _T_1619;
  wire  _T_1621;
  wire  _T_1623;
  wire  _T_1625;
  wire  _T_1627;
  wire  _T_1629;
  wire  _T_1631;
  wire  _T_1633;
  wire  _T_1635;
  wire  _T_1637;
  wire  _T_1639;
  wire  _T_1641;
  wire  _T_1643;
  wire  _T_1645;
  wire  _T_1647;
  wire  _T_1649;
  wire  _T_1651;
  wire  _T_1653;
  wire  _T_1655;
  wire  _T_1657;
  wire  _T_1659;
  wire  _T_1661;
  wire  _T_1663;
  wire  _T_1665;
  wire  _T_1667;
  wire  _T_1669;
  wire  _T_1670;
  wire  _T_1671;
  wire  _T_1672;
  wire  _T_1673;
  wire  _T_1674;
  wire  _T_1675;
  wire  _T_1676;
  wire  _T_1677;
  wire  _T_1678;
  wire  _T_1679;
  wire  _T_1680;
  wire  _T_1681;
  wire  _T_1682;
  wire  _T_1683;
  wire  _T_1684;
  wire  _T_1685;
  wire  _T_1686;
  wire  _T_1687;
  wire  _T_1688;
  wire  _T_1689;
  wire  _T_1690;
  wire  _T_1691;
  wire  _T_1692;
  wire  _T_1693;
  wire  _T_1694;
  wire  _T_1695;
  wire  _T_1696;
  wire  _T_1697;
  wire  _T_1698;
  wire  _T_1699;
  wire  _T_1700;
  wire  _T_1701;
  wire  _T_1702;
  wire  _T_1703;
  wire  _T_1704;
  wire  _T_1705;
  wire  _T_1706;
  wire  _T_1707;
  wire  _T_1708;
  wire  _T_1709;
  wire  _T_1710;
  wire  _T_1711;
  wire  _T_1712;
  wire  _T_1713;
  wire  _T_1714;
  wire  _T_1715;
  wire  _T_1716;
  wire  _T_1717;
  wire  _T_1718;
  wire  _T_1719;
  wire  _T_1720;
  wire  _T_1721;
  wire  _T_1722;
  wire  _T_1723;
  wire  _T_1724;
  wire  _T_1725;
  wire  _T_1726;
  wire  _T_1727;
  wire  _T_1728;
  wire  _T_1729;
  wire  _T_1730;
  wire  _T_1731;
  wire  _T_1732;
  wire  _T_1733;
  wire  _T_1734;
  wire  _T_1735;
  wire  _T_1736;
  wire  _T_1737;
  wire  _T_1738;
  wire  _T_1739;
  wire  _T_1740;
  wire  _T_1741;
  wire  _T_1742;
  wire  _T_1743;
  wire  _T_1744;
  wire  _T_1745;
  wire  _T_1746;
  wire  _T_1747;
  wire  _T_1748;
  wire  _T_1749;
  wire  _T_1750;
  wire  _T_1751;
  wire  _T_1752;
  wire  _T_1753;
  wire  _T_1754;
  wire  _T_1755;
  wire  _T_1756;
  wire  _T_1757;
  wire  _T_1758;
  wire  _T_1759;
  wire  _T_1760;
  wire  _T_1761;
  wire  _T_1762;
  wire  _T_1763;
  wire  _T_1764;
  wire  _T_1765;
  wire  _T_1766;
  wire  _T_1767;
  wire  _T_1768;
  wire  _T_1769;
  wire  _T_1770;
  wire  _T_1771;
  wire  _T_1772;
  wire  _T_1773;
  wire  _T_1774;
  wire  _T_1775;
  wire  _T_1776;
  wire  _T_1777;
  wire  _T_1778;
  wire  _T_1779;
  wire  _T_1780;
  wire  _T_1781;
  wire  _T_1782;
  wire  _T_1783;
  wire  _T_1784;
  wire  _T_1785;
  wire  _T_1786;
  wire  _T_1787;
  wire  _T_1788;
  wire  _T_1789;
  wire  _T_1790;
  wire  _T_1791;
  wire  _T_1792;
  wire  _T_1793;
  wire  _T_1794;
  wire  _T_1796;
  wire  _T_1797;
  wire  _T_1801;
  wire  _T_1802;
  wire  _T_1803;
  wire  _T_1806;
  wire  _T_1807;
  wire  _T_1808;
  wire  _T_1811;
  wire  _T_1812;
  wire  _T_1813;
  wire  _T_1814;
  wire  _T_1817;
  wire [31:0] _T_1819;
  wire  _T_1820;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1830;
  wire  _T_1831;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1844;
  wire  _T_1845;
  wire  _T_1847;
  wire  _T_1848;
  wire [1:0] _T_1849;
  wire [1:0] _T_1850;
  wire  _T_1852;
  wire  _T_1854;
  wire  _T_1856;
  wire  _T_1857;
  wire  _T_1859;
  wire  _T_1861;
  wire  _T_1862;
  wire  _T_1863;
  wire  _T_1865;
  wire  _T_1868;
  wire  _T_1870;
  wire  _T_1871;
  wire  _T_1872;
  wire  _T_1874;
  wire  _T_1875;
  wire  _T_1876;
  wire  _T_1880;
  wire  _T_1881;
  wire  _T_1883;
  wire  _T_1884;
  wire  _T_1885;
  wire  _T_1889;
  wire  _T_1890;
  wire [1:0] _T_1924;
  wire  _T_1925;
  wire  _T_1927;
  wire  _T_1929;
  wire  _T_1931;
  wire  _T_1933;
  wire  _T_1935;
  wire  _T_1937;
  wire  _T_1939;
  wire  _T_1941;
  wire  _T_1943;
  wire  _T_1945;
  wire  _T_1947;
  wire  _T_1949;
  wire  _T_1951;
  wire  _T_1953;
  wire  _T_1955;
  wire  _T_1957;
  wire  _T_1959;
  wire  _T_1961;
  wire  _T_1963;
  wire  _T_1965;
  wire  _T_1967;
  wire  _T_1969;
  wire  _T_1971;
  wire  _T_1973;
  wire  _T_1975;
  wire  _T_1977;
  wire  _T_1979;
  wire  _T_1981;
  wire  _T_1983;
  wire  _T_1985;
  wire  _T_1987;
  wire  _T_1989;
  wire  _T_1991;
  wire  _T_1993;
  wire  _T_1995;
  wire  _T_1997;
  wire  _T_1999;
  wire  _T_2001;
  wire  _T_2003;
  wire  _T_2005;
  wire  _T_2007;
  wire  _T_2009;
  wire  _T_2011;
  wire  _T_2013;
  wire  _T_2015;
  wire  _T_2017;
  wire  _T_2019;
  wire  _T_2021;
  wire  _T_2023;
  wire  _T_2025;
  wire  _T_2027;
  wire  _T_2029;
  wire  _T_2031;
  wire  _T_2033;
  wire  _T_2035;
  wire  _T_2037;
  wire  _T_2039;
  wire  _T_2041;
  wire  _T_2043;
  wire  _T_2045;
  wire  _T_2047;
  wire  _T_2049;
  wire  _T_2051;
  wire  _T_2053;
  wire  _T_2055;
  wire  _T_2057;
  wire  _T_2059;
  wire  _T_2061;
  wire  _T_2063;
  wire  _T_2065;
  wire  _T_2067;
  wire  _T_2069;
  wire  _T_2071;
  wire  _T_2073;
  wire  _T_2075;
  wire  _T_2077;
  wire  _T_2079;
  wire  _T_2081;
  wire  _T_2083;
  wire  _T_2085;
  wire  _T_2087;
  wire  _T_2089;
  wire  _T_2091;
  wire  _T_2093;
  wire  _T_2095;
  wire  _T_2097;
  wire  _T_2099;
  wire  _T_2101;
  wire  _T_2103;
  wire  _T_2105;
  wire  _T_2107;
  wire  _T_2109;
  wire  _T_2111;
  wire  _T_2113;
  wire  _T_2115;
  wire  _T_2117;
  wire  _T_2119;
  wire  _T_2121;
  wire  _T_2123;
  wire  _T_2125;
  wire  _T_2127;
  wire  _T_2129;
  wire  _T_2131;
  wire  _T_2133;
  wire  _T_2135;
  wire  _T_2137;
  wire  _T_2139;
  wire  _T_2141;
  wire  _T_2143;
  wire  _T_2145;
  wire  _T_2147;
  wire  _T_2149;
  wire  _T_2151;
  wire  _T_2153;
  wire  _T_2155;
  wire  _T_2157;
  wire  _T_2159;
  wire  _T_2161;
  wire  _T_2163;
  wire  _T_2165;
  wire  _T_2167;
  wire  _T_2169;
  wire  _T_2171;
  wire  _T_2173;
  wire  _T_2175;
  wire  _T_2177;
  wire  _T_2178;
  wire  _T_2179;
  wire  _T_2180;
  wire  _T_2181;
  wire  _T_2182;
  wire  _T_2183;
  wire  _T_2184;
  wire  _T_2185;
  wire  _T_2186;
  wire  _T_2187;
  wire  _T_2188;
  wire  _T_2189;
  wire  _T_2190;
  wire  _T_2191;
  wire  _T_2192;
  wire  _T_2193;
  wire  _T_2194;
  wire  _T_2195;
  wire  _T_2196;
  wire  _T_2197;
  wire  _T_2198;
  wire  _T_2199;
  wire  _T_2200;
  wire  _T_2201;
  wire  _T_2202;
  wire  _T_2203;
  wire  _T_2204;
  wire  _T_2205;
  wire  _T_2206;
  wire  _T_2207;
  wire  _T_2208;
  wire  _T_2209;
  wire  _T_2210;
  wire  _T_2211;
  wire  _T_2212;
  wire  _T_2213;
  wire  _T_2214;
  wire  _T_2215;
  wire  _T_2216;
  wire  _T_2217;
  wire  _T_2218;
  wire  _T_2219;
  wire  _T_2220;
  wire  _T_2221;
  wire  _T_2222;
  wire  _T_2223;
  wire  _T_2224;
  wire  _T_2225;
  wire  _T_2226;
  wire  _T_2227;
  wire  _T_2228;
  wire  _T_2229;
  wire  _T_2230;
  wire  _T_2231;
  wire  _T_2232;
  wire  _T_2233;
  wire  _T_2234;
  wire  _T_2235;
  wire  _T_2236;
  wire  _T_2237;
  wire  _T_2238;
  wire  _T_2239;
  wire  _T_2240;
  wire  _T_2241;
  wire  _T_2242;
  wire  _T_2243;
  wire  _T_2244;
  wire  _T_2245;
  wire  _T_2246;
  wire  _T_2247;
  wire  _T_2248;
  wire  _T_2249;
  wire  _T_2250;
  wire  _T_2251;
  wire  _T_2252;
  wire  _T_2253;
  wire  _T_2254;
  wire  _T_2255;
  wire  _T_2256;
  wire  _T_2257;
  wire  _T_2258;
  wire  _T_2259;
  wire  _T_2260;
  wire  _T_2261;
  wire  _T_2262;
  wire  _T_2263;
  wire  _T_2264;
  wire  _T_2265;
  wire  _T_2266;
  wire  _T_2267;
  wire  _T_2268;
  wire  _T_2269;
  wire  _T_2270;
  wire  _T_2271;
  wire  _T_2272;
  wire  _T_2273;
  wire  _T_2274;
  wire  _T_2275;
  wire  _T_2276;
  wire  _T_2277;
  wire  _T_2278;
  wire  _T_2279;
  wire  _T_2280;
  wire  _T_2281;
  wire  _T_2282;
  wire  _T_2283;
  wire  _T_2284;
  wire  _T_2285;
  wire  _T_2286;
  wire  _T_2287;
  wire  _T_2288;
  wire  _T_2289;
  wire  _T_2290;
  wire  _T_2291;
  wire  _T_2292;
  wire  _T_2293;
  wire  _T_2294;
  wire  _T_2295;
  wire  _T_2296;
  wire  _T_2297;
  wire  _T_2298;
  wire  _T_2299;
  wire  _T_2300;
  wire  _T_2301;
  wire  _T_2302;
  wire  _T_2304;
  wire  _T_2305;
  wire  _T_2310;
  wire  _T_2311;
  wire  _T_2314;
  wire  _T_2315;
  wire  _T_2316;
  wire  _T_2319;
  wire  _T_2320;
  wire  _T_2321;
  wire  _T_2322;
  wire  _T_2325;
  wire [31:0] _T_2327;
  wire  _T_2328;
  wire  _T_2329;
  wire  _T_2330;
  wire  _T_2338;
  wire  _T_2339;
  wire  _T_2343;
  wire  _T_2344;
  wire  _T_2352;
  wire  _T_2353;
  wire  _T_2355;
  wire  _T_2356;
  wire [1:0] _T_2357;
  wire [1:0] _T_2358;
  wire  _T_2360;
  wire  _T_2362;
  wire  _T_2364;
  wire  _T_2365;
  wire  _T_2367;
  wire  _T_2369;
  wire  _T_2370;
  wire  _T_2371;
  wire  _T_2373;
  wire  _T_2376;
  wire  _T_2378;
  wire  _T_2379;
  wire  _T_2380;
  wire  _T_2383;
  wire  _T_2384;
  wire  _T_2388;
  wire  _T_2389;
  wire  _T_2392;
  wire  _T_2393;
  wire  _T_2397;
  wire  _T_2398;
  wire [3:0] _GEN_605;
  wire [4:0] _T_2400;
  wire [3:0] _T_2401;
  wire [63:0] _T_2403;
  wire [63:0] cause;
  wire [7:0] cause_lsbs;
  wire  _T_2404;
  wire  _T_2406;
  wire  causeIsDebugInt;
  wire  _T_2409;
  wire  causeIsDebugTrigger;
  wire  _T_2415;
  wire [1:0] _T_2416;
  wire [1:0] _T_2417;
  wire [3:0] _T_2418;
  wire [3:0] _T_2419;
  wire  _T_2420;
  wire  causeIsDebugBreak;
  wire  _T_2422;
  wire  _T_2423;
  wire  _T_2424;
  wire  trapToDebug;
  wire [11:0] _T_2428;
  wire [11:0] debugTVec;
  wire [63:0] _T_2435;
  wire  _T_2436;
  wire [63:0] _T_2437;
  wire  _T_2438;
  wire  _T_2439;
  wire  delegate;
  wire [39:0] _T_2444;
  wire [39:0] _T_2445;
  wire [3:0] _T_2446;
  wire [5:0] _GEN_606;
  wire [5:0] _T_2447;
  wire [33:0] _T_2448;
  wire [39:0] _T_2449;
  wire  _T_2450;
  wire  _T_2452;
  wire [3:0] _T_2453;
  wire  _T_2455;
  wire  _T_2456;
  wire [39:0] notDebugTVec;
  wire [39:0] tvec;
  wire  _T_2457;
  wire  _T_2458;
  wire  _T_2461;
  wire [1:0] _T_2462;
  wire  _T_2464;
  wire [1:0] _T_2465;
  wire  _T_2467;
  wire  _T_2468;
  wire  _T_2473;
  wire [1:0] _T_2474;
  reg [1:0] _T_2476;
  reg [31:0] _RAND_150;
  wire  exception;
  wire [1:0] _T_2478;
  wire [1:0] _T_2479;
  wire [2:0] _T_2480;
  wire  _T_2482;
  wire  _T_2484;
  wire  _T_2486;
  wire  _T_2489;
  wire  _T_2492;
  wire  _GEN_83;
  wire  _T_2495;
  wire  _T_2496;
  wire  _T_2497;
  wire  _GEN_84;
  wire  _T_2500;
  wire  _T_2502;
  wire  _T_2503;
  wire  _T_2505;
  wire  _T_2507;
  wire  _T_2508;
  wire  _T_2509;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _T_2517;
  wire  _T_2518;
  wire  _T_2520;
  wire  _T_2522;
  wire  _T_2524;
  wire  _T_2527;
  wire  _T_2529;
  wire  _T_2531;
  wire [39:0] _T_2532;
  wire [39:0] _T_2534;
  wire [39:0] epc;
  wire  _T_2545;
  wire  _T_2546;
  wire  _T_2547;
  wire  _T_2548;
  wire  _T_2549;
  wire  _T_2550;
  wire  _T_2551;
  wire  _T_2552;
  wire  _T_2553;
  wire  _T_2554;
  wire  _T_2555;
  wire  _T_2556;
  wire  _T_2557;
  wire  _T_2558;
  wire  _T_2559;
  wire  _T_2560;
  wire  _T_2561;
  wire  _T_2562;
  wire  _T_2563;
  wire  write_badaddr;
  wire [39:0] badaddr_value;
  wire [1:0] _T_2572;
  wire [1:0] _T_2573;
  wire [2:0] _T_2574;
  wire  _GEN_87;
  wire [39:0] _GEN_88;
  wire [2:0] _GEN_89;
  wire [1:0] _GEN_90;
  wire [1:0] _GEN_91;
  wire [39:0] _T_2576;
  wire  _T_2577;
  wire  _T_2579;
  wire [1:0] _T_2581;
  wire [39:0] _GEN_607;
  wire [39:0] _T_2582;
  wire [39:0] _T_2583;
  wire [39:0] _GEN_92;
  wire [63:0] _GEN_93;
  wire [39:0] _GEN_94;
  wire  _GEN_95;
  wire [1:0] _GEN_96;
  wire  _GEN_97;
  wire [1:0] _GEN_98;
  wire [39:0] _GEN_99;
  wire [63:0] _GEN_100;
  wire [39:0] _GEN_101;
  wire  _GEN_102;
  wire [1:0] _GEN_103;
  wire  _GEN_104;
  wire  _GEN_105;
  wire [39:0] _GEN_106;
  wire [2:0] _GEN_107;
  wire [1:0] _GEN_108;
  wire [1:0] _GEN_109;
  wire [39:0] _GEN_110;
  wire [63:0] _GEN_111;
  wire [39:0] _GEN_112;
  wire  _GEN_113;
  wire [1:0] _GEN_114;
  wire  _GEN_115;
  wire [39:0] _GEN_116;
  wire [63:0] _GEN_117;
  wire [39:0] _GEN_118;
  wire  _GEN_119;
  wire [1:0] _GEN_120;
  wire  _GEN_121;
  wire  _GEN_122;
  wire [39:0] _GEN_123;
  wire [2:0] _GEN_124;
  wire [1:0] _GEN_125;
  wire [1:0] _GEN_126;
  wire [39:0] _GEN_127;
  wire [63:0] _GEN_128;
  wire [39:0] _GEN_129;
  wire  _GEN_130;
  wire [1:0] _GEN_131;
  wire  _GEN_132;
  wire [39:0] _GEN_133;
  wire [63:0] _GEN_134;
  wire [39:0] _GEN_135;
  wire  _GEN_136;
  wire [1:0] _GEN_137;
  wire  _GEN_138;
  wire  _T_2597;
  wire  _T_2599;
  wire  _T_2604;
  wire [1:0] _GEN_139;
  wire  _GEN_140;
  wire [39:0] _GEN_141;
  wire  _GEN_142;
  wire  _GEN_143;
  wire [1:0] _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire [1:0] _GEN_147;
  wire [1:0] _GEN_148;
  wire [39:0] _GEN_149;
  wire  _GEN_150;
  wire  _GEN_151;
  wire  _GEN_152;
  wire [1:0] _GEN_153;
  wire  _GEN_154;
  wire  _GEN_155;
  wire [1:0] _GEN_156;
  wire [1:0] _GEN_157;
  wire [39:0] _GEN_158;
  wire  _GEN_159;
  wire  _GEN_160;
  wire  _GEN_161;
  wire [1:0] _GEN_162;
  wire [63:0] _T_2617;
  wire [63:0] _T_2619;
  wire [63:0] _T_2627;
  wire [63:0] _T_2629;
  wire [31:0] _T_2631;
  wire [15:0] _T_2633;
  wire [63:0] _T_2635;
  wire [63:0] _T_2637;
  wire [63:0] _T_2639;
  wire [63:0] _T_2641;
  wire [63:0] _T_2643;
  wire [31:0] _T_2647;
  wire [39:0] _T_2649;
  wire [63:0] _T_2651;
  wire [4:0] _T_2653;
  wire [2:0] _T_2655;
  wire [7:0] _T_2657;
  wire [63:0] _T_2659;
  wire [63:0] _T_2661;
  wire [63:0] _T_2663;
  wire [39:0] _T_2665;
  wire [39:0] _T_2667;
  wire [63:0] _T_2669;
  wire [39:0] _T_2671;
  wire [39:0] _T_2673;
  wire [63:0] _T_2675;
  wire [39:0] _T_2677;
  wire [39:0] _T_2679;
  wire [63:0] _T_2681;
  wire [39:0] _T_2683;
  wire [39:0] _T_2685;
  wire [63:0] _T_2687;
  wire [39:0] _T_2689;
  wire [39:0] _T_2691;
  wire [63:0] _T_2693;
  wire [39:0] _T_2695;
  wire [39:0] _T_2697;
  wire [63:0] _T_2699;
  wire [39:0] _T_2701;
  wire [39:0] _T_2703;
  wire [63:0] _T_2705;
  wire [39:0] _T_2707;
  wire [39:0] _T_2709;
  wire [63:0] _T_2711;
  wire [39:0] _T_2713;
  wire [39:0] _T_2715;
  wire [63:0] _T_2717;
  wire [39:0] _T_2719;
  wire [39:0] _T_2721;
  wire [63:0] _T_2723;
  wire [39:0] _T_2725;
  wire [39:0] _T_2727;
  wire [63:0] _T_2729;
  wire [39:0] _T_2731;
  wire [39:0] _T_2733;
  wire [63:0] _T_2735;
  wire [39:0] _T_2737;
  wire [39:0] _T_2739;
  wire [63:0] _T_2741;
  wire [39:0] _T_2743;
  wire [39:0] _T_2745;
  wire [63:0] _T_2747;
  wire [39:0] _T_2749;
  wire [39:0] _T_2751;
  wire [63:0] _T_2753;
  wire [39:0] _T_2755;
  wire [39:0] _T_2757;
  wire [63:0] _T_2759;
  wire [39:0] _T_2761;
  wire [39:0] _T_2763;
  wire [63:0] _T_2765;
  wire [39:0] _T_2767;
  wire [39:0] _T_2769;
  wire [63:0] _T_2771;
  wire [39:0] _T_2773;
  wire [39:0] _T_2775;
  wire [63:0] _T_2777;
  wire [39:0] _T_2779;
  wire [39:0] _T_2781;
  wire [63:0] _T_2783;
  wire [39:0] _T_2785;
  wire [39:0] _T_2787;
  wire [63:0] _T_2789;
  wire [39:0] _T_2791;
  wire [39:0] _T_2793;
  wire [63:0] _T_2795;
  wire [39:0] _T_2797;
  wire [39:0] _T_2799;
  wire [63:0] _T_2801;
  wire [39:0] _T_2803;
  wire [39:0] _T_2805;
  wire [63:0] _T_2807;
  wire [39:0] _T_2809;
  wire [39:0] _T_2811;
  wire [63:0] _T_2813;
  wire [39:0] _T_2815;
  wire [39:0] _T_2817;
  wire [63:0] _T_2819;
  wire [39:0] _T_2821;
  wire [39:0] _T_2823;
  wire [63:0] _T_2825;
  wire [39:0] _T_2827;
  wire [39:0] _T_2829;
  wire [63:0] _T_2831;
  wire [39:0] _T_2833;
  wire [39:0] _T_2835;
  wire [31:0] _T_2837;
  wire [63:0] _T_2839;
  wire [63:0] _T_2841;
  wire [63:0] _T_2843;
  wire [63:0] _T_2845;
  wire [63:0] _T_2847;
  wire [63:0] _T_2849;
  wire [63:0] _T_2851;
  wire [63:0] _T_2853;
  wire [63:0] _T_2855;
  wire [63:0] _T_2857;
  wire [63:0] _T_2859;
  wire [31:0] _T_2861;
  wire [63:0] _T_2863;
  wire [63:0] _T_2865;
  wire [63:0] _T_2867;
  wire [63:0] _T_2871;
  wire [63:0] _T_2872;
  wire [63:0] _GEN_609;
  wire [63:0] _T_2873;
  wire [63:0] _GEN_610;
  wire [63:0] _T_2874;
  wire [63:0] _T_2875;
  wire [63:0] _T_2876;
  wire [63:0] _T_2877;
  wire [63:0] _T_2878;
  wire [63:0] _T_2879;
  wire [63:0] _GEN_611;
  wire [63:0] _T_2881;
  wire [63:0] _GEN_612;
  wire [63:0] _T_2882;
  wire [63:0] _T_2883;
  wire [63:0] _GEN_613;
  wire [63:0] _T_2884;
  wire [63:0] _GEN_614;
  wire [63:0] _T_2885;
  wire [63:0] _GEN_615;
  wire [63:0] _T_2886;
  wire [63:0] _T_2887;
  wire [63:0] _T_2888;
  wire [63:0] _T_2889;
  wire [63:0] _GEN_616;
  wire [63:0] _T_2890;
  wire [63:0] _GEN_617;
  wire [63:0] _T_2891;
  wire [63:0] _T_2892;
  wire [63:0] _GEN_618;
  wire [63:0] _T_2893;
  wire [63:0] _GEN_619;
  wire [63:0] _T_2894;
  wire [63:0] _T_2895;
  wire [63:0] _GEN_620;
  wire [63:0] _T_2896;
  wire [63:0] _GEN_621;
  wire [63:0] _T_2897;
  wire [63:0] _T_2898;
  wire [63:0] _GEN_622;
  wire [63:0] _T_2899;
  wire [63:0] _GEN_623;
  wire [63:0] _T_2900;
  wire [63:0] _T_2901;
  wire [63:0] _GEN_624;
  wire [63:0] _T_2902;
  wire [63:0] _GEN_625;
  wire [63:0] _T_2903;
  wire [63:0] _T_2904;
  wire [63:0] _GEN_626;
  wire [63:0] _T_2905;
  wire [63:0] _GEN_627;
  wire [63:0] _T_2906;
  wire [63:0] _T_2907;
  wire [63:0] _GEN_628;
  wire [63:0] _T_2908;
  wire [63:0] _GEN_629;
  wire [63:0] _T_2909;
  wire [63:0] _T_2910;
  wire [63:0] _GEN_630;
  wire [63:0] _T_2911;
  wire [63:0] _GEN_631;
  wire [63:0] _T_2912;
  wire [63:0] _T_2913;
  wire [63:0] _GEN_632;
  wire [63:0] _T_2914;
  wire [63:0] _GEN_633;
  wire [63:0] _T_2915;
  wire [63:0] _T_2916;
  wire [63:0] _GEN_634;
  wire [63:0] _T_2917;
  wire [63:0] _GEN_635;
  wire [63:0] _T_2918;
  wire [63:0] _T_2919;
  wire [63:0] _GEN_636;
  wire [63:0] _T_2920;
  wire [63:0] _GEN_637;
  wire [63:0] _T_2921;
  wire [63:0] _T_2922;
  wire [63:0] _GEN_638;
  wire [63:0] _T_2923;
  wire [63:0] _GEN_639;
  wire [63:0] _T_2924;
  wire [63:0] _T_2925;
  wire [63:0] _GEN_640;
  wire [63:0] _T_2926;
  wire [63:0] _GEN_641;
  wire [63:0] _T_2927;
  wire [63:0] _T_2928;
  wire [63:0] _GEN_642;
  wire [63:0] _T_2929;
  wire [63:0] _GEN_643;
  wire [63:0] _T_2930;
  wire [63:0] _T_2931;
  wire [63:0] _GEN_644;
  wire [63:0] _T_2932;
  wire [63:0] _GEN_645;
  wire [63:0] _T_2933;
  wire [63:0] _T_2934;
  wire [63:0] _GEN_646;
  wire [63:0] _T_2935;
  wire [63:0] _GEN_647;
  wire [63:0] _T_2936;
  wire [63:0] _T_2937;
  wire [63:0] _GEN_648;
  wire [63:0] _T_2938;
  wire [63:0] _GEN_649;
  wire [63:0] _T_2939;
  wire [63:0] _T_2940;
  wire [63:0] _GEN_650;
  wire [63:0] _T_2941;
  wire [63:0] _GEN_651;
  wire [63:0] _T_2942;
  wire [63:0] _T_2943;
  wire [63:0] _GEN_652;
  wire [63:0] _T_2944;
  wire [63:0] _GEN_653;
  wire [63:0] _T_2945;
  wire [63:0] _T_2946;
  wire [63:0] _GEN_654;
  wire [63:0] _T_2947;
  wire [63:0] _GEN_655;
  wire [63:0] _T_2948;
  wire [63:0] _T_2949;
  wire [63:0] _GEN_656;
  wire [63:0] _T_2950;
  wire [63:0] _GEN_657;
  wire [63:0] _T_2951;
  wire [63:0] _T_2952;
  wire [63:0] _GEN_658;
  wire [63:0] _T_2953;
  wire [63:0] _GEN_659;
  wire [63:0] _T_2954;
  wire [63:0] _T_2955;
  wire [63:0] _GEN_660;
  wire [63:0] _T_2956;
  wire [63:0] _GEN_661;
  wire [63:0] _T_2957;
  wire [63:0] _T_2958;
  wire [63:0] _GEN_662;
  wire [63:0] _T_2959;
  wire [63:0] _GEN_663;
  wire [63:0] _T_2960;
  wire [63:0] _T_2961;
  wire [63:0] _GEN_664;
  wire [63:0] _T_2962;
  wire [63:0] _GEN_665;
  wire [63:0] _T_2963;
  wire [63:0] _T_2964;
  wire [63:0] _GEN_666;
  wire [63:0] _T_2965;
  wire [63:0] _GEN_667;
  wire [63:0] _T_2966;
  wire [63:0] _T_2967;
  wire [63:0] _GEN_668;
  wire [63:0] _T_2968;
  wire [63:0] _GEN_669;
  wire [63:0] _T_2969;
  wire [63:0] _T_2970;
  wire [63:0] _GEN_670;
  wire [63:0] _T_2971;
  wire [63:0] _GEN_671;
  wire [63:0] _T_2972;
  wire [63:0] _T_2973;
  wire [63:0] _GEN_672;
  wire [63:0] _T_2974;
  wire [63:0] _GEN_673;
  wire [63:0] _T_2975;
  wire [63:0] _GEN_674;
  wire [63:0] _T_2976;
  wire [63:0] _T_2977;
  wire [63:0] _T_2978;
  wire [63:0] _T_2979;
  wire [63:0] _T_2980;
  wire [63:0] _T_2981;
  wire [63:0] _T_2982;
  wire [63:0] _T_2983;
  wire [63:0] _T_2984;
  wire [63:0] _T_2985;
  wire [63:0] _T_2986;
  wire [63:0] _T_2987;
  wire [63:0] _GEN_675;
  wire [63:0] _T_2988;
  wire [63:0] _T_2989;
  wire [63:0] _T_2990;
  wire [63:0] _T_2992;
  wire [4:0] _T_2993;
  wire [4:0] _GEN_163;
  wire  _T_2999;
  wire  _T_3001;
  wire  _T_3004_tsr;
  wire  _T_3004_tw;
  wire  _T_3004_tvm;
  wire  _T_3004_mxr;
  wire  _T_3004_sum;
  wire  _T_3004_mprv;
  wire [1:0] _T_3004_fs;
  wire [1:0] _T_3004_mpp;
  wire  _T_3004_spp;
  wire  _T_3004_mpie;
  wire  _T_3004_spie;
  wire  _T_3004_mie;
  wire  _T_3004_sie;
  wire [100:0] _T_3006;
  wire  _T_3008;
  wire  _T_3010;
  wire  _T_3012;
  wire  _T_3014;
  wire  _T_3015;
  wire [1:0] _T_3017;
  wire [1:0] _T_3018;
  wire  _T_3020;
  wire  _T_3021;
  wire  _T_3022;
  wire  _T_3023;
  wire  _T_3024;
  wire  _T_3025;
  wire  _T_3037;
  wire [1:0] _T_3041;
  wire  _GEN_164;
  wire  _GEN_165;
  wire  _GEN_166;
  wire [1:0] _GEN_167;
  wire  _GEN_168;
  wire  _GEN_169;
  wire [1:0] _GEN_170;
  wire  _GEN_171;
  wire  _GEN_172;
  wire  _GEN_173;
  wire  _GEN_174;
  wire  _GEN_175;
  wire [1:0] _GEN_176;
  wire  _T_3043;
  wire [63:0] _T_3044;
  wire  _T_3046;
  wire [3:0] _GEN_676;
  wire [3:0] _T_3047;
  wire [63:0] _GEN_677;
  wire [63:0] _T_3048;
  wire [63:0] _T_3049;
  wire [63:0] _T_3050;
  wire [63:0] _T_3052;
  wire [63:0] _T_3053;
  wire [63:0] _GEN_177;
  wire [1:0] _T_3054;
  wire [3:0] _T_3056;
  wire [1:0] _T_3057;
  wire [3:0] _T_3059;
  wire [7:0] _T_3060;
  wire [1:0] _T_3061;
  wire [3:0] _T_3063;
  wire [7:0] _T_3067;
  wire [15:0] _T_3068;
  wire [15:0] _T_3075;
  wire [63:0] _GEN_678;
  wire [63:0] _T_3076;
  wire [63:0] _T_3082;
  wire  _T_3089_seip;
  wire  _T_3089_stip;
  wire  _T_3089_ssip;
  wire [15:0] _T_3093;
  wire  _T_3095;
  wire  _T_3099;
  wire  _T_3103;
  wire  _GEN_178;
  wire  _GEN_179;
  wire  _GEN_180;
  wire [63:0] _T_3110;
  wire [63:0] _GEN_181;
  wire [63:0] _GEN_679;
  wire [63:0] _T_3117;
  wire [63:0] _T_3118;
  wire [63:0] _GEN_182;
  wire [63:0] _GEN_183;
  wire [63:0] _T_3121;
  wire  _T_3122;
  wire [5:0] _T_3125;
  wire [63:0] _GEN_680;
  wire [63:0] _T_3126;
  wire [63:0] _T_3127;
  wire [63:0] _GEN_184;
  wire [63:0] _T_3129;
  wire [63:0] _GEN_185;
  wire [39:0] _T_3130;
  wire [39:0] _GEN_186;
  wire [33:0] _T_3132;
  wire [39:0] _GEN_187;
  wire [33:0] _GEN_188;
  wire [63:0] _T_3134;
  wire [63:0] _GEN_189;
  wire [39:0] _GEN_190;
  wire [33:0] _GEN_191;
  wire [63:0] _GEN_192;
  wire [39:0] _GEN_193;
  wire [33:0] _GEN_194;
  wire [63:0] _GEN_195;
  wire [39:0] _GEN_196;
  wire [33:0] _GEN_197;
  wire [63:0] _GEN_198;
  wire [39:0] _GEN_199;
  wire [33:0] _GEN_200;
  wire [63:0] _GEN_201;
  wire [39:0] _GEN_202;
  wire [33:0] _GEN_203;
  wire [63:0] _GEN_204;
  wire [39:0] _GEN_205;
  wire [33:0] _GEN_206;
  wire [63:0] _GEN_207;
  wire [39:0] _GEN_208;
  wire [33:0] _GEN_209;
  wire [63:0] _GEN_210;
  wire [39:0] _GEN_211;
  wire [33:0] _GEN_212;
  wire [63:0] _GEN_213;
  wire [39:0] _GEN_214;
  wire [33:0] _GEN_215;
  wire [63:0] _GEN_216;
  wire [39:0] _GEN_217;
  wire [33:0] _GEN_218;
  wire [63:0] _GEN_219;
  wire [39:0] _GEN_220;
  wire [33:0] _GEN_221;
  wire [63:0] _GEN_222;
  wire [39:0] _GEN_223;
  wire [33:0] _GEN_224;
  wire [63:0] _GEN_225;
  wire [39:0] _GEN_226;
  wire [33:0] _GEN_227;
  wire [63:0] _GEN_228;
  wire [39:0] _GEN_229;
  wire [33:0] _GEN_230;
  wire [63:0] _GEN_231;
  wire [39:0] _GEN_232;
  wire [33:0] _GEN_233;
  wire [63:0] _GEN_234;
  wire [39:0] _GEN_235;
  wire [33:0] _GEN_236;
  wire [63:0] _GEN_237;
  wire [39:0] _GEN_238;
  wire [33:0] _GEN_239;
  wire [63:0] _GEN_240;
  wire [39:0] _GEN_241;
  wire [33:0] _GEN_242;
  wire [63:0] _GEN_243;
  wire [39:0] _GEN_244;
  wire [33:0] _GEN_245;
  wire [63:0] _GEN_246;
  wire [39:0] _GEN_247;
  wire [33:0] _GEN_248;
  wire [63:0] _GEN_249;
  wire [39:0] _GEN_250;
  wire [33:0] _GEN_251;
  wire [63:0] _GEN_252;
  wire [39:0] _GEN_253;
  wire [33:0] _GEN_254;
  wire [63:0] _GEN_255;
  wire [39:0] _GEN_256;
  wire [33:0] _GEN_257;
  wire [63:0] _GEN_258;
  wire [39:0] _GEN_259;
  wire [33:0] _GEN_260;
  wire [63:0] _GEN_261;
  wire [39:0] _GEN_262;
  wire [33:0] _GEN_263;
  wire [63:0] _GEN_264;
  wire [39:0] _GEN_265;
  wire [33:0] _GEN_266;
  wire [63:0] _GEN_267;
  wire [39:0] _GEN_268;
  wire [33:0] _GEN_269;
  wire [63:0] _GEN_270;
  wire [39:0] _GEN_271;
  wire [33:0] _GEN_272;
  wire [63:0] _GEN_273;
  wire [57:0] _T_3248;
  wire [63:0] _GEN_274;
  wire [57:0] _GEN_275;
  wire [63:0] _GEN_276;
  wire [57:0] _GEN_277;
  wire [63:0] _GEN_278;
  wire [63:0] _GEN_279;
  wire [58:0] _T_3251;
  wire [63:0] _GEN_280;
  wire [63:0] _GEN_281;
  wire  _T_3254_ebreakm;
  wire  _T_3254_ebreaks;
  wire  _T_3254_ebreaku;
  wire  _T_3254_step;
  wire [1:0] _T_3254_prv;
  wire [31:0] _T_3256;
  wire [1:0] _T_3257;
  wire  _T_3258;
  wire  _T_3264;
  wire  _T_3265;
  wire  _T_3267;
  wire  _GEN_282;
  wire  _GEN_283;
  wire  _GEN_284;
  wire  _GEN_285;
  wire [1:0] _GEN_286;
  wire [63:0] _T_3273;
  wire [63:0] _T_3274;
  wire [63:0] _GEN_287;
  wire [63:0] _GEN_288;
  wire  _T_3277_mxr;
  wire  _T_3277_sum;
  wire [1:0] _T_3277_fs;
  wire  _T_3277_spp;
  wire  _T_3277_spie;
  wire  _T_3277_sie;
  wire [100:0] _T_3279;
  wire  _T_3281;
  wire  _T_3285;
  wire  _T_3288;
  wire [1:0] _T_3291;
  wire  _T_3294;
  wire  _T_3295;
  wire  _T_3310;
  wire [1:0] _T_3314;
  wire  _GEN_289;
  wire  _GEN_290;
  wire [1:0] _GEN_291;
  wire  _GEN_292;
  wire  _GEN_293;
  wire [1:0] _GEN_294;
  wire  _T_3321_ssip;
  wire [15:0] _T_3325;
  wire  _T_3327;
  wire  _GEN_295;
  wire [3:0] _T_3344_mode;
  wire [43:0] _T_3344_ppn;
  wire [63:0] _T_3346;
  wire [43:0] _T_3347;
  wire [3:0] _T_3349;
  wire  _T_3351;
  wire [3:0] _GEN_296;
  wire  _T_3354;
  wire [3:0] _GEN_297;
  wire  _T_3360;
  wire [19:0] _T_3361;
  wire [43:0] _GEN_298;
  wire [3:0] _GEN_299;
  wire [43:0] _GEN_300;
  wire [63:0] _T_3362;
  wire [63:0] _T_3363;
  wire [63:0] _T_3364;
  wire [63:0] _T_3365;
  wire [63:0] _GEN_301;
  wire [63:0] _GEN_302;
  wire [63:0] _GEN_303;
  wire [63:0] _GEN_304;
  wire [63:0] _T_3384;
  wire [63:0] _GEN_305;
  wire [39:0] _GEN_306;
  wire [63:0] _T_3386;
  wire [63:0] _GEN_307;
  wire [63:0] _T_3387;
  wire [63:0] _GEN_308;
  wire [63:0] _T_3389;
  wire [63:0] _GEN_309;
  wire [63:0] _GEN_310;
  wire  _GEN_17_control_dmode;
  wire  _T_3394;
  wire  _T_3395;
  wire  _T_3398_dmode;
  wire  _T_3398_action;
  wire [1:0] _T_3398_tmatch;
  wire  _T_3398_m;
  wire  _T_3398_s;
  wire  _T_3398_u;
  wire  _T_3398_x;
  wire  _T_3398_w;
  wire  _T_3398_r;
  wire [63:0] _T_3400;
  wire  _T_3401;
  wire  _T_3402;
  wire  _T_3403;
  wire  _T_3404;
  wire  _T_3405;
  wire  _T_3407;
  wire [1:0] _T_3408;
  wire  _T_3411;
  wire  _T_3414;
  wire  _T_3416;
  wire [1:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _T_3417;
  wire  _GEN_34;
  wire  _GEN_348;
  wire  _GEN_354;
  wire [1:0] _GEN_360;
  wire  _GEN_362;
  wire  _GEN_366;
  wire  _GEN_368;
  wire  _GEN_370;
  wire  _GEN_372;
  wire  _GEN_374;
  wire [38:0] _GEN_35;
  wire [38:0] _GEN_378;
  wire  _GEN_382;
  wire  _GEN_388;
  wire [1:0] _GEN_394;
  wire  _GEN_396;
  wire  _GEN_400;
  wire  _GEN_402;
  wire  _GEN_404;
  wire  _GEN_406;
  wire  _GEN_408;
  wire [38:0] _GEN_410;
  wire  _GEN_412;
  wire  _GEN_413;
  wire  _GEN_414;
  wire [1:0] _GEN_415;
  wire  _GEN_416;
  wire  _GEN_417;
  wire [1:0] _GEN_418;
  wire  _GEN_419;
  wire  _GEN_420;
  wire  _GEN_421;
  wire  _GEN_422;
  wire  _GEN_423;
  wire [1:0] _GEN_424;
  wire [63:0] _GEN_425;
  wire  _GEN_426;
  wire  _GEN_427;
  wire  _GEN_428;
  wire [63:0] _GEN_429;
  wire [63:0] _GEN_430;
  wire [63:0] _GEN_431;
  wire [63:0] _GEN_432;
  wire [63:0] _GEN_433;
  wire [39:0] _GEN_434;
  wire [39:0] _GEN_435;
  wire [33:0] _GEN_436;
  wire [63:0] _GEN_437;
  wire [39:0] _GEN_438;
  wire [33:0] _GEN_439;
  wire [63:0] _GEN_440;
  wire [39:0] _GEN_441;
  wire [33:0] _GEN_442;
  wire [63:0] _GEN_443;
  wire [39:0] _GEN_444;
  wire [33:0] _GEN_445;
  wire [63:0] _GEN_446;
  wire [39:0] _GEN_447;
  wire [33:0] _GEN_448;
  wire [63:0] _GEN_449;
  wire [39:0] _GEN_450;
  wire [33:0] _GEN_451;
  wire [63:0] _GEN_452;
  wire [39:0] _GEN_453;
  wire [33:0] _GEN_454;
  wire [63:0] _GEN_455;
  wire [39:0] _GEN_456;
  wire [33:0] _GEN_457;
  wire [63:0] _GEN_458;
  wire [39:0] _GEN_459;
  wire [33:0] _GEN_460;
  wire [63:0] _GEN_461;
  wire [39:0] _GEN_462;
  wire [33:0] _GEN_463;
  wire [63:0] _GEN_464;
  wire [39:0] _GEN_465;
  wire [33:0] _GEN_466;
  wire [63:0] _GEN_467;
  wire [39:0] _GEN_468;
  wire [33:0] _GEN_469;
  wire [63:0] _GEN_470;
  wire [39:0] _GEN_471;
  wire [33:0] _GEN_472;
  wire [63:0] _GEN_473;
  wire [39:0] _GEN_474;
  wire [33:0] _GEN_475;
  wire [63:0] _GEN_476;
  wire [39:0] _GEN_477;
  wire [33:0] _GEN_478;
  wire [63:0] _GEN_479;
  wire [39:0] _GEN_480;
  wire [33:0] _GEN_481;
  wire [63:0] _GEN_482;
  wire [39:0] _GEN_483;
  wire [33:0] _GEN_484;
  wire [63:0] _GEN_485;
  wire [39:0] _GEN_486;
  wire [33:0] _GEN_487;
  wire [63:0] _GEN_488;
  wire [39:0] _GEN_489;
  wire [33:0] _GEN_490;
  wire [63:0] _GEN_491;
  wire [39:0] _GEN_492;
  wire [33:0] _GEN_493;
  wire [63:0] _GEN_494;
  wire [39:0] _GEN_495;
  wire [33:0] _GEN_496;
  wire [63:0] _GEN_497;
  wire [39:0] _GEN_498;
  wire [33:0] _GEN_499;
  wire [63:0] _GEN_500;
  wire [39:0] _GEN_501;
  wire [33:0] _GEN_502;
  wire [63:0] _GEN_503;
  wire [39:0] _GEN_504;
  wire [33:0] _GEN_505;
  wire [63:0] _GEN_506;
  wire [39:0] _GEN_507;
  wire [33:0] _GEN_508;
  wire [63:0] _GEN_509;
  wire [39:0] _GEN_510;
  wire [33:0] _GEN_511;
  wire [63:0] _GEN_512;
  wire [39:0] _GEN_513;
  wire [33:0] _GEN_514;
  wire [63:0] _GEN_515;
  wire [39:0] _GEN_516;
  wire [33:0] _GEN_517;
  wire [63:0] _GEN_518;
  wire [39:0] _GEN_519;
  wire [33:0] _GEN_520;
  wire [63:0] _GEN_521;
  wire [63:0] _GEN_522;
  wire [57:0] _GEN_523;
  wire [63:0] _GEN_524;
  wire [57:0] _GEN_525;
  wire [63:0] _GEN_526;
  wire [63:0] _GEN_527;
  wire  _GEN_528;
  wire  _GEN_529;
  wire  _GEN_530;
  wire  _GEN_531;
  wire [1:0] _GEN_532;
  wire [63:0] _GEN_533;
  wire [63:0] _GEN_534;
  wire [3:0] _GEN_535;
  wire [43:0] _GEN_536;
  wire [63:0] _GEN_537;
  wire [63:0] _GEN_538;
  wire [63:0] _GEN_539;
  wire [63:0] _GEN_540;
  wire [39:0] _GEN_541;
  wire [63:0] _GEN_542;
  wire [63:0] _GEN_543;
  wire [63:0] _GEN_544;
  wire [63:0] _GEN_545;
  wire  _GEN_549;
  wire  _GEN_555;
  wire [1:0] _GEN_561;
  wire  _GEN_563;
  wire  _GEN_567;
  wire  _GEN_569;
  wire  _GEN_571;
  wire  _GEN_573;
  wire  _GEN_575;
  wire [38:0] _GEN_577;
  wire  _GEN_579;
  wire  _GEN_580;
  wire  _GEN_581;
  wire  _GEN_582;
  wire  _GEN_583;
  assign _T_194 = new_prv == 2'h2;
  assign _T_196 = _T_194 ? 2'h0 : new_prv;
  assign _GEN_0 = {{4'd0}, io_retire};
  assign _T_329 = _T_328 + _GEN_0;
  assign _T_333 = _T_329[6];
  assign _T_335 = _T_332 + 58'h1;
  assign _T_336 = _T_335[57:0];
  assign _GEN_36 = _T_333 ? _T_336 : _T_332;
  assign _T_337 = {_T_332,_T_328};
  assign _T_342 = _T_341 + 6'h1;
  assign _T_346 = _T_342[6];
  assign _T_348 = _T_345 + 58'h1;
  assign _T_349 = _T_348[57:0];
  assign _GEN_37 = _T_346 ? _T_349 : _T_345;
  assign _T_350 = {_T_345,_T_341};
  assign _GEN_1 = {{4'd0}, io_counters_0_inc};
  assign _T_411 = _T_410 + _GEN_1;
  assign _T_414 = _T_411[6];
  assign _T_416 = _T_413 + 34'h1;
  assign _T_417 = _T_416[33:0];
  assign _GEN_38 = _T_414 ? _T_417 : _T_413;
  assign _T_418 = {_T_413,_T_410};
  assign _GEN_2 = {{4'd0}, io_counters_1_inc};
  assign _T_421 = _T_420 + _GEN_2;
  assign _T_424 = _T_421[6];
  assign _T_426 = _T_423 + 34'h1;
  assign _T_427 = _T_426[33:0];
  assign _GEN_39 = _T_424 ? _T_427 : _T_423;
  assign _T_428 = {_T_423,_T_420};
  assign _GEN_3 = {{4'd0}, io_counters_2_inc};
  assign _T_431 = _T_430 + _GEN_3;
  assign _T_434 = _T_431[6];
  assign _T_436 = _T_433 + 34'h1;
  assign _T_437 = _T_436[33:0];
  assign _GEN_40 = _T_434 ? _T_437 : _T_433;
  assign _T_438 = {_T_433,_T_430};
  assign _GEN_4 = {{4'd0}, io_counters_3_inc};
  assign _T_441 = _T_440 + _GEN_4;
  assign _T_444 = _T_441[6];
  assign _T_446 = _T_443 + 34'h1;
  assign _T_447 = _T_446[33:0];
  assign _GEN_41 = _T_444 ? _T_447 : _T_443;
  assign _T_448 = {_T_443,_T_440};
  assign _GEN_5 = {{4'd0}, io_counters_4_inc};
  assign _T_451 = _T_450 + _GEN_5;
  assign _T_454 = _T_451[6];
  assign _T_456 = _T_453 + 34'h1;
  assign _T_457 = _T_456[33:0];
  assign _GEN_42 = _T_454 ? _T_457 : _T_453;
  assign _T_458 = {_T_453,_T_450};
  assign _GEN_6 = {{4'd0}, io_counters_5_inc};
  assign _T_461 = _T_460 + _GEN_6;
  assign _T_464 = _T_461[6];
  assign _T_466 = _T_463 + 34'h1;
  assign _T_467 = _T_466[33:0];
  assign _GEN_43 = _T_464 ? _T_467 : _T_463;
  assign _T_468 = {_T_463,_T_460};
  assign _GEN_7 = {{4'd0}, io_counters_6_inc};
  assign _T_471 = _T_470 + _GEN_7;
  assign _T_474 = _T_471[6];
  assign _T_476 = _T_473 + 34'h1;
  assign _T_477 = _T_476[33:0];
  assign _GEN_44 = _T_474 ? _T_477 : _T_473;
  assign _T_478 = {_T_473,_T_470};
  assign _GEN_8 = {{4'd0}, io_counters_7_inc};
  assign _T_481 = _T_480 + _GEN_8;
  assign _T_484 = _T_481[6];
  assign _T_486 = _T_483 + 34'h1;
  assign _T_487 = _T_486[33:0];
  assign _GEN_45 = _T_484 ? _T_487 : _T_483;
  assign _T_488 = {_T_483,_T_480};
  assign _GEN_9 = {{4'd0}, io_counters_8_inc};
  assign _T_491 = _T_490 + _GEN_9;
  assign _T_494 = _T_491[6];
  assign _T_496 = _T_493 + 34'h1;
  assign _T_497 = _T_496[33:0];
  assign _GEN_46 = _T_494 ? _T_497 : _T_493;
  assign _T_498 = {_T_493,_T_490};
  assign _GEN_10 = {{4'd0}, io_counters_9_inc};
  assign _T_501 = _T_500 + _GEN_10;
  assign _T_504 = _T_501[6];
  assign _T_506 = _T_503 + 34'h1;
  assign _T_507 = _T_506[33:0];
  assign _GEN_47 = _T_504 ? _T_507 : _T_503;
  assign _T_508 = {_T_503,_T_500};
  assign _GEN_11 = {{4'd0}, io_counters_10_inc};
  assign _T_511 = _T_510 + _GEN_11;
  assign _T_514 = _T_511[6];
  assign _T_516 = _T_513 + 34'h1;
  assign _T_517 = _T_516[33:0];
  assign _GEN_48 = _T_514 ? _T_517 : _T_513;
  assign _T_518 = {_T_513,_T_510};
  assign _GEN_12 = {{4'd0}, io_counters_11_inc};
  assign _T_521 = _T_520 + _GEN_12;
  assign _T_524 = _T_521[6];
  assign _T_526 = _T_523 + 34'h1;
  assign _T_527 = _T_526[33:0];
  assign _GEN_49 = _T_524 ? _T_527 : _T_523;
  assign _T_528 = {_T_523,_T_520};
  assign _GEN_13 = {{4'd0}, io_counters_12_inc};
  assign _T_531 = _T_530 + _GEN_13;
  assign _T_534 = _T_531[6];
  assign _T_536 = _T_533 + 34'h1;
  assign _T_537 = _T_536[33:0];
  assign _GEN_50 = _T_534 ? _T_537 : _T_533;
  assign _T_538 = {_T_533,_T_530};
  assign _GEN_14 = {{4'd0}, io_counters_13_inc};
  assign _T_541 = _T_540 + _GEN_14;
  assign _T_544 = _T_541[6];
  assign _T_546 = _T_543 + 34'h1;
  assign _T_547 = _T_546[33:0];
  assign _GEN_51 = _T_544 ? _T_547 : _T_543;
  assign _T_548 = {_T_543,_T_540};
  assign _GEN_15 = {{4'd0}, io_counters_14_inc};
  assign _T_551 = _T_550 + _GEN_15;
  assign _T_554 = _T_551[6];
  assign _T_556 = _T_553 + 34'h1;
  assign _T_557 = _T_556[33:0];
  assign _GEN_52 = _T_554 ? _T_557 : _T_553;
  assign _T_558 = {_T_553,_T_550};
  assign _GEN_16 = {{4'd0}, io_counters_15_inc};
  assign _T_561 = _T_560 + _GEN_16;
  assign _T_564 = _T_561[6];
  assign _T_566 = _T_563 + 34'h1;
  assign _T_567 = _T_566[33:0];
  assign _GEN_53 = _T_564 ? _T_567 : _T_563;
  assign _T_568 = {_T_563,_T_560};
  assign _GEN_17 = {{4'd0}, io_counters_16_inc};
  assign _T_571 = _T_570 + _GEN_17;
  assign _T_574 = _T_571[6];
  assign _T_576 = _T_573 + 34'h1;
  assign _T_577 = _T_576[33:0];
  assign _GEN_54 = _T_574 ? _T_577 : _T_573;
  assign _T_578 = {_T_573,_T_570};
  assign _GEN_589 = {{4'd0}, io_counters_17_inc};
  assign _T_581 = _T_580 + _GEN_589;
  assign _T_584 = _T_581[6];
  assign _T_586 = _T_583 + 34'h1;
  assign _T_587 = _T_586[33:0];
  assign _GEN_55 = _T_584 ? _T_587 : _T_583;
  assign _T_588 = {_T_583,_T_580};
  assign _GEN_590 = {{4'd0}, io_counters_18_inc};
  assign _T_591 = _T_590 + _GEN_590;
  assign _T_594 = _T_591[6];
  assign _T_596 = _T_593 + 34'h1;
  assign _T_597 = _T_596[33:0];
  assign _GEN_56 = _T_594 ? _T_597 : _T_593;
  assign _T_598 = {_T_593,_T_590};
  assign _GEN_591 = {{4'd0}, io_counters_19_inc};
  assign _T_601 = _T_600 + _GEN_591;
  assign _T_604 = _T_601[6];
  assign _T_606 = _T_603 + 34'h1;
  assign _T_607 = _T_606[33:0];
  assign _GEN_57 = _T_604 ? _T_607 : _T_603;
  assign _T_608 = {_T_603,_T_600};
  assign _GEN_592 = {{4'd0}, io_counters_20_inc};
  assign _T_611 = _T_610 + _GEN_592;
  assign _T_614 = _T_611[6];
  assign _T_616 = _T_613 + 34'h1;
  assign _T_617 = _T_616[33:0];
  assign _GEN_58 = _T_614 ? _T_617 : _T_613;
  assign _T_618 = {_T_613,_T_610};
  assign _GEN_593 = {{4'd0}, io_counters_21_inc};
  assign _T_621 = _T_620 + _GEN_593;
  assign _T_624 = _T_621[6];
  assign _T_626 = _T_623 + 34'h1;
  assign _T_627 = _T_626[33:0];
  assign _GEN_59 = _T_624 ? _T_627 : _T_623;
  assign _T_628 = {_T_623,_T_620};
  assign _GEN_594 = {{4'd0}, io_counters_22_inc};
  assign _T_631 = _T_630 + _GEN_594;
  assign _T_634 = _T_631[6];
  assign _T_636 = _T_633 + 34'h1;
  assign _T_637 = _T_636[33:0];
  assign _GEN_60 = _T_634 ? _T_637 : _T_633;
  assign _T_638 = {_T_633,_T_630};
  assign _GEN_595 = {{4'd0}, io_counters_23_inc};
  assign _T_641 = _T_640 + _GEN_595;
  assign _T_644 = _T_641[6];
  assign _T_646 = _T_643 + 34'h1;
  assign _T_647 = _T_646[33:0];
  assign _GEN_61 = _T_644 ? _T_647 : _T_643;
  assign _T_648 = {_T_643,_T_640};
  assign _GEN_596 = {{4'd0}, io_counters_24_inc};
  assign _T_651 = _T_650 + _GEN_596;
  assign _T_654 = _T_651[6];
  assign _T_656 = _T_653 + 34'h1;
  assign _T_657 = _T_656[33:0];
  assign _GEN_62 = _T_654 ? _T_657 : _T_653;
  assign _T_658 = {_T_653,_T_650};
  assign _GEN_597 = {{4'd0}, io_counters_25_inc};
  assign _T_661 = _T_660 + _GEN_597;
  assign _T_664 = _T_661[6];
  assign _T_666 = _T_663 + 34'h1;
  assign _T_667 = _T_666[33:0];
  assign _GEN_63 = _T_664 ? _T_667 : _T_663;
  assign _T_668 = {_T_663,_T_660};
  assign _GEN_598 = {{4'd0}, io_counters_26_inc};
  assign _T_671 = _T_670 + _GEN_598;
  assign _T_674 = _T_671[6];
  assign _T_676 = _T_673 + 34'h1;
  assign _T_677 = _T_676[33:0];
  assign _GEN_64 = _T_674 ? _T_677 : _T_673;
  assign _T_678 = {_T_673,_T_670};
  assign _GEN_599 = {{4'd0}, io_counters_27_inc};
  assign _T_681 = _T_680 + _GEN_599;
  assign _T_684 = _T_681[6];
  assign _T_686 = _T_683 + 34'h1;
  assign _T_687 = _T_686[33:0];
  assign _GEN_65 = _T_684 ? _T_687 : _T_683;
  assign _T_688 = {_T_683,_T_680};
  assign _GEN_600 = {{4'd0}, io_counters_28_inc};
  assign _T_691 = _T_690 + _GEN_600;
  assign _T_694 = _T_691[6];
  assign _T_696 = _T_693 + 34'h1;
  assign _T_697 = _T_696[33:0];
  assign _GEN_66 = _T_694 ? _T_697 : _T_693;
  assign _T_698 = {_T_693,_T_690};
  assign _T_701 = reg_mstatus_prv == 2'h1;
  assign _T_704 = _T_701 ? 32'hffffffff : reg_scounteren;
  assign hpm_mask = reg_mcounteren & _T_704;
  assign _T_712 = reg_mip_seip | _T_711;
  assign _T_713 = {mip_ssip,1'h0};
  assign _T_714 = {mip_msip,1'h0};
  assign _T_715 = {_T_714,_T_713};
  assign _T_716 = {mip_stip,1'h0};
  assign _T_717 = {mip_mtip,1'h0};
  assign _T_718 = {_T_717,_T_716};
  assign _T_719 = {_T_718,_T_715};
  assign _T_720 = {mip_seip,1'h0};
  assign _T_721 = {mip_meip,1'h0};
  assign _T_722 = {_T_721,_T_720};
  assign _T_726 = {4'h0,_T_722};
  assign _T_727 = {_T_726,_T_719};
  assign read_mip = _T_727 & 16'haaa;
  assign _GEN_601 = {{48'd0}, read_mip};
  assign pending_interrupts = _GEN_601 & reg_mie;
  assign _GEN_602 = {{14'd0}, io_interrupts_debug};
  assign d_interrupts = _GEN_602 << 14;
  assign _T_730 = reg_mstatus_prv <= 2'h1;
  assign _T_731 = _T_730 | reg_mstatus_mie;
  assign _T_732 = ~ pending_interrupts;
  assign _T_733 = _T_732 | reg_mideleg;
  assign _T_734 = ~ _T_733;
  assign m_interrupts = _T_731 ? _T_734 : 64'h0;
  assign _T_737 = reg_mstatus_prv < 2'h1;
  assign _T_740 = _T_701 & reg_mstatus_sie;
  assign _T_741 = _T_737 | _T_740;
  assign _T_742 = pending_interrupts & reg_mideleg;
  assign s_interrupts = _T_741 ? _T_742 : 64'h0;
  assign _T_744 = d_interrupts[14];
  assign _T_745 = d_interrupts[13];
  assign _T_746 = d_interrupts[12];
  assign _T_747 = d_interrupts[11];
  assign _T_748 = d_interrupts[3];
  assign _T_749 = d_interrupts[7];
  assign _T_750 = d_interrupts[9];
  assign _T_751 = d_interrupts[1];
  assign _T_752 = d_interrupts[5];
  assign _T_753 = d_interrupts[8];
  assign _T_754 = d_interrupts[0];
  assign _T_755 = d_interrupts[4];
  assign _T_756 = m_interrupts[15];
  assign _T_757 = m_interrupts[14];
  assign _T_758 = m_interrupts[13];
  assign _T_759 = m_interrupts[12];
  assign _T_760 = m_interrupts[11];
  assign _T_761 = m_interrupts[3];
  assign _T_762 = m_interrupts[7];
  assign _T_763 = m_interrupts[9];
  assign _T_764 = m_interrupts[1];
  assign _T_765 = m_interrupts[5];
  assign _T_766 = m_interrupts[8];
  assign _T_767 = m_interrupts[0];
  assign _T_768 = m_interrupts[4];
  assign _T_769 = s_interrupts[15];
  assign _T_770 = s_interrupts[14];
  assign _T_771 = s_interrupts[13];
  assign _T_772 = s_interrupts[12];
  assign _T_773 = s_interrupts[11];
  assign _T_774 = s_interrupts[3];
  assign _T_775 = s_interrupts[7];
  assign _T_776 = s_interrupts[9];
  assign _T_777 = s_interrupts[1];
  assign _T_778 = s_interrupts[5];
  assign _T_779 = s_interrupts[8];
  assign _T_780 = s_interrupts[0];
  assign _T_781 = s_interrupts[4];
  assign _T_782 = _T_744 | _T_745;
  assign _T_783 = _T_782 | _T_746;
  assign _T_784 = _T_783 | _T_747;
  assign _T_785 = _T_784 | _T_748;
  assign _T_786 = _T_785 | _T_749;
  assign _T_787 = _T_786 | _T_750;
  assign _T_788 = _T_787 | _T_751;
  assign _T_789 = _T_788 | _T_752;
  assign _T_790 = _T_789 | _T_753;
  assign _T_791 = _T_790 | _T_754;
  assign _T_792 = _T_791 | _T_755;
  assign _T_793 = _T_792 | _T_756;
  assign _T_794 = _T_793 | _T_757;
  assign _T_795 = _T_794 | _T_758;
  assign _T_796 = _T_795 | _T_759;
  assign _T_797 = _T_796 | _T_760;
  assign _T_798 = _T_797 | _T_761;
  assign _T_799 = _T_798 | _T_762;
  assign _T_800 = _T_799 | _T_763;
  assign _T_801 = _T_800 | _T_764;
  assign _T_802 = _T_801 | _T_765;
  assign _T_803 = _T_802 | _T_766;
  assign _T_804 = _T_803 | _T_767;
  assign _T_805 = _T_804 | _T_768;
  assign _T_806 = _T_805 | _T_769;
  assign _T_807 = _T_806 | _T_770;
  assign _T_808 = _T_807 | _T_771;
  assign _T_809 = _T_808 | _T_772;
  assign _T_810 = _T_809 | _T_773;
  assign _T_811 = _T_810 | _T_774;
  assign _T_812 = _T_811 | _T_775;
  assign _T_813 = _T_812 | _T_776;
  assign _T_814 = _T_813 | _T_777;
  assign _T_815 = _T_814 | _T_778;
  assign _T_816 = _T_815 | _T_779;
  assign _T_817 = _T_816 | _T_780;
  assign anyInterrupt = _T_817 | _T_781;
  assign _T_894 = _T_780 ? 3'h0 : 3'h4;
  assign _T_895 = _T_779 ? 4'h8 : {{1'd0}, _T_894};
  assign _T_896 = _T_778 ? 4'h5 : _T_895;
  assign _T_897 = _T_777 ? 4'h1 : _T_896;
  assign _T_898 = _T_776 ? 4'h9 : _T_897;
  assign _T_899 = _T_775 ? 4'h7 : _T_898;
  assign _T_900 = _T_774 ? 4'h3 : _T_899;
  assign _T_901 = _T_773 ? 4'hb : _T_900;
  assign _T_902 = _T_772 ? 4'hc : _T_901;
  assign _T_903 = _T_771 ? 4'hd : _T_902;
  assign _T_904 = _T_770 ? 4'he : _T_903;
  assign _T_905 = _T_769 ? 4'hf : _T_904;
  assign _T_906 = _T_768 ? 4'h4 : _T_905;
  assign _T_907 = _T_767 ? 4'h0 : _T_906;
  assign _T_908 = _T_766 ? 4'h8 : _T_907;
  assign _T_909 = _T_765 ? 4'h5 : _T_908;
  assign _T_910 = _T_764 ? 4'h1 : _T_909;
  assign _T_911 = _T_763 ? 4'h9 : _T_910;
  assign _T_912 = _T_762 ? 4'h7 : _T_911;
  assign _T_913 = _T_761 ? 4'h3 : _T_912;
  assign _T_914 = _T_760 ? 4'hb : _T_913;
  assign _T_915 = _T_759 ? 4'hc : _T_914;
  assign _T_916 = _T_758 ? 4'hd : _T_915;
  assign _T_917 = _T_757 ? 4'he : _T_916;
  assign _T_918 = _T_756 ? 4'hf : _T_917;
  assign _T_919 = _T_755 ? 4'h4 : _T_918;
  assign _T_920 = _T_754 ? 4'h0 : _T_919;
  assign _T_921 = _T_753 ? 4'h8 : _T_920;
  assign _T_922 = _T_752 ? 4'h5 : _T_921;
  assign _T_923 = _T_751 ? 4'h1 : _T_922;
  assign _T_924 = _T_750 ? 4'h9 : _T_923;
  assign _T_925 = _T_749 ? 4'h7 : _T_924;
  assign _T_926 = _T_748 ? 4'h3 : _T_925;
  assign _T_927 = _T_747 ? 4'hb : _T_926;
  assign _T_928 = _T_746 ? 4'hc : _T_927;
  assign _T_929 = _T_745 ? 4'hd : _T_928;
  assign whichInterrupt = _T_744 ? 4'he : _T_929;
  assign _GEN_603 = {{60'd0}, whichInterrupt};
  assign _T_931 = 64'h8000000000000000 + _GEN_603;
  assign interruptCause = _T_931[63:0];
  assign _T_933 = reg_debug == 1'h0;
  assign _T_934 = anyInterrupt & _T_933;
  assign _T_936 = io_singleStep == 1'h0;
  assign _T_937 = _T_934 & _T_936;
  assign _T_938 = _T_937 | reg_singleStepped;
  assign _T_941 = {io_status_hie,io_status_sie};
  assign _T_942 = {_T_941,io_status_uie};
  assign _T_943 = {io_status_upie,io_status_mie};
  assign _T_944 = {io_status_hpie,io_status_spie};
  assign _T_945 = {_T_944,_T_943};
  assign _T_946 = {_T_945,_T_942};
  assign _T_947 = {io_status_hpp,io_status_spp};
  assign _T_948 = {_T_947,io_status_mpie};
  assign _T_949 = {io_status_fs,io_status_mpp};
  assign _T_950 = {io_status_mprv,io_status_xs};
  assign _T_951 = {_T_950,_T_949};
  assign _T_952 = {_T_951,_T_948};
  assign _T_953 = {_T_952,_T_946};
  assign _T_954 = {io_status_tvm,io_status_mxr};
  assign _T_955 = {_T_954,io_status_sum};
  assign _T_956 = {io_status_tsr,io_status_tw};
  assign _T_957 = {io_status_sd_rv32,io_status_zero1};
  assign _T_958 = {_T_957,_T_956};
  assign _T_959 = {_T_958,_T_955};
  assign _T_960 = {io_status_sxl,io_status_uxl};
  assign _T_961 = {io_status_sd,io_status_zero2};
  assign _T_962 = {_T_961,_T_960};
  assign _T_963 = {io_status_dprv,io_status_prv};
  assign _T_964 = {io_status_debug,io_status_isa};
  assign _T_965 = {_T_964,_T_963};
  assign _T_966 = {_T_965,_T_962};
  assign _T_967 = {_T_966,_T_959};
  assign _T_968 = {_T_967,_T_953};
  assign read_mstatus = _T_968[63:0];
  assign _T_970 = {_GEN_0_control_x,_GEN_1_control_w};
  assign _T_971 = {_T_970,_GEN_2_control_r};
  assign _T_972 = {_GEN_3_control_s,_GEN_4_control_u};
  assign _T_973 = {_GEN_5_control_m,1'h0};
  assign _T_974 = {_T_973,_T_972};
  assign _T_975 = {_T_974,_T_971};
  assign _T_976 = {2'h0,_GEN_8_control_tmatch};
  assign _T_977 = {_GEN_9_control_action,1'h0};
  assign _T_978 = {_T_977,_T_976};
  assign _T_980 = {4'h2,_GEN_14_control_dmode};
  assign _T_981 = {_T_980,46'h40000000000};
  assign _T_982 = {_T_981,_T_978};
  assign _T_983 = {_T_982,_T_975};
  assign _T_985 = _GEN_15_address[38];
  assign _T_989 = _T_985 ? 25'h1ffffff : 25'h0;
  assign _T_990 = {_T_989,_GEN_16_address};
  assign _T_994 = reg_mepc[39];
  assign _T_998 = _T_994 ? 24'hffffff : 24'h0;
  assign _T_999 = {_T_998,reg_mepc};
  assign _T_1000 = reg_mbadaddr[39];
  assign _T_1004 = _T_1000 ? 24'hffffff : 24'h0;
  assign _T_1005 = {_T_1004,reg_mbadaddr};
  assign _T_1006 = {3'h0,reg_dcsr_step};
  assign _T_1007 = {_T_1006,reg_dcsr_prv};
  assign _T_1008 = {1'h0,reg_dcsr_cause};
  assign _T_1010 = {2'h0,_T_1008};
  assign _T_1011 = {_T_1010,_T_1007};
  assign _T_1012 = {1'h0,reg_dcsr_ebreaks};
  assign _T_1013 = {_T_1012,reg_dcsr_ebreaku};
  assign _T_1014 = {12'h0,reg_dcsr_ebreakm};
  assign _T_1016 = {4'h4,_T_1014};
  assign _T_1017 = {_T_1016,_T_1013};
  assign _T_1018 = {_T_1017,_T_1011};
  assign _T_1019 = {reg_frm,reg_fflags};
  assign _T_1022 = reg_mie & reg_mideleg;
  assign _T_1023 = _GEN_601 & reg_mideleg;
  assign _T_1061 = {1'h0,_T_1060_sie};
  assign _T_1062 = {_T_1061,1'h0};
  assign _T_1064 = {1'h0,_T_1060_spie};
  assign _T_1065 = {_T_1064,2'h0};
  assign _T_1066 = {_T_1065,_T_1062};
  assign _T_1067 = {2'h0,_T_1060_spp};
  assign _T_1068 = {_T_1067,1'h0};
  assign _T_1069 = {_T_1060_fs,2'h0};
  assign _T_1070 = {1'h0,_T_1060_xs};
  assign _T_1071 = {_T_1070,_T_1069};
  assign _T_1072 = {_T_1071,_T_1068};
  assign _T_1073 = {_T_1072,_T_1066};
  assign _T_1074 = {1'h0,_T_1060_mxr};
  assign _T_1075 = {_T_1074,_T_1060_sum};
  assign _T_1077 = {_T_1060_sd_rv32,8'h0};
  assign _T_1078 = {_T_1077,2'h0};
  assign _T_1079 = {_T_1078,_T_1075};
  assign _T_1080 = {2'h0,_T_1060_uxl};
  assign _T_1081 = {_T_1060_sd,27'h0};
  assign _T_1082 = {_T_1081,_T_1080};
  assign _T_1086 = {37'h0,_T_1082};
  assign _T_1087 = {_T_1086,_T_1079};
  assign _T_1088 = {_T_1087,_T_1073};
  assign _T_1089 = _T_1088[63:0];
  assign _T_1090 = reg_sbadaddr[39];
  assign _T_1094 = _T_1090 ? 24'hffffff : 24'h0;
  assign _T_1095 = {_T_1094,reg_sbadaddr};
  assign _T_1096 = {reg_sptbr_mode,16'h0};
  assign _T_1097 = {_T_1096,reg_sptbr_ppn};
  assign _T_1098 = reg_sepc[39];
  assign _T_1102 = _T_1098 ? 24'hffffff : 24'h0;
  assign _T_1103 = {_T_1102,reg_sepc};
  assign _T_1104 = reg_stvec[38];
  assign _T_1108 = _T_1104 ? 25'h1ffffff : 25'h0;
  assign _T_1109 = {_T_1108,reg_stvec};
  assign _T_1114 = io_rw_addr == 12'h7a1;
  assign _T_1116 = io_rw_addr == 12'h7a2;
  assign _T_1124 = io_rw_addr == 12'h301;
  assign _T_1126 = io_rw_addr == 12'h300;
  assign _T_1128 = io_rw_addr == 12'h305;
  assign _T_1130 = io_rw_addr == 12'h344;
  assign _T_1132 = io_rw_addr == 12'h304;
  assign _T_1134 = io_rw_addr == 12'h340;
  assign _T_1136 = io_rw_addr == 12'h341;
  assign _T_1138 = io_rw_addr == 12'h343;
  assign _T_1140 = io_rw_addr == 12'h342;
  assign _T_1144 = io_rw_addr == 12'h7b0;
  assign _T_1146 = io_rw_addr == 12'h7b1;
  assign _T_1148 = io_rw_addr == 12'h7b2;
  assign _T_1150 = io_rw_addr == 12'h1;
  assign _T_1152 = io_rw_addr == 12'h2;
  assign _T_1154 = io_rw_addr == 12'h3;
  assign _T_1156 = io_rw_addr == 12'hb00;
  assign _T_1158 = io_rw_addr == 12'hb02;
  assign _T_1160 = io_rw_addr == 12'h323;
  assign _T_1162 = io_rw_addr == 12'hb03;
  assign _T_1164 = io_rw_addr == 12'hc03;
  assign _T_1166 = io_rw_addr == 12'h324;
  assign _T_1168 = io_rw_addr == 12'hb04;
  assign _T_1170 = io_rw_addr == 12'hc04;
  assign _T_1172 = io_rw_addr == 12'h325;
  assign _T_1174 = io_rw_addr == 12'hb05;
  assign _T_1176 = io_rw_addr == 12'hc05;
  assign _T_1178 = io_rw_addr == 12'h326;
  assign _T_1180 = io_rw_addr == 12'hb06;
  assign _T_1182 = io_rw_addr == 12'hc06;
  assign _T_1184 = io_rw_addr == 12'h327;
  assign _T_1186 = io_rw_addr == 12'hb07;
  assign _T_1188 = io_rw_addr == 12'hc07;
  assign _T_1190 = io_rw_addr == 12'h328;
  assign _T_1192 = io_rw_addr == 12'hb08;
  assign _T_1194 = io_rw_addr == 12'hc08;
  assign _T_1196 = io_rw_addr == 12'h329;
  assign _T_1198 = io_rw_addr == 12'hb09;
  assign _T_1200 = io_rw_addr == 12'hc09;
  assign _T_1202 = io_rw_addr == 12'h32a;
  assign _T_1204 = io_rw_addr == 12'hb0a;
  assign _T_1206 = io_rw_addr == 12'hc0a;
  assign _T_1208 = io_rw_addr == 12'h32b;
  assign _T_1210 = io_rw_addr == 12'hb0b;
  assign _T_1212 = io_rw_addr == 12'hc0b;
  assign _T_1214 = io_rw_addr == 12'h32c;
  assign _T_1216 = io_rw_addr == 12'hb0c;
  assign _T_1218 = io_rw_addr == 12'hc0c;
  assign _T_1220 = io_rw_addr == 12'h32d;
  assign _T_1222 = io_rw_addr == 12'hb0d;
  assign _T_1224 = io_rw_addr == 12'hc0d;
  assign _T_1226 = io_rw_addr == 12'h32e;
  assign _T_1228 = io_rw_addr == 12'hb0e;
  assign _T_1230 = io_rw_addr == 12'hc0e;
  assign _T_1232 = io_rw_addr == 12'h32f;
  assign _T_1234 = io_rw_addr == 12'hb0f;
  assign _T_1236 = io_rw_addr == 12'hc0f;
  assign _T_1238 = io_rw_addr == 12'h330;
  assign _T_1240 = io_rw_addr == 12'hb10;
  assign _T_1242 = io_rw_addr == 12'hc10;
  assign _T_1244 = io_rw_addr == 12'h331;
  assign _T_1246 = io_rw_addr == 12'hb11;
  assign _T_1248 = io_rw_addr == 12'hc11;
  assign _T_1250 = io_rw_addr == 12'h332;
  assign _T_1252 = io_rw_addr == 12'hb12;
  assign _T_1254 = io_rw_addr == 12'hc12;
  assign _T_1256 = io_rw_addr == 12'h333;
  assign _T_1258 = io_rw_addr == 12'hb13;
  assign _T_1260 = io_rw_addr == 12'hc13;
  assign _T_1262 = io_rw_addr == 12'h334;
  assign _T_1264 = io_rw_addr == 12'hb14;
  assign _T_1266 = io_rw_addr == 12'hc14;
  assign _T_1268 = io_rw_addr == 12'h335;
  assign _T_1270 = io_rw_addr == 12'hb15;
  assign _T_1272 = io_rw_addr == 12'hc15;
  assign _T_1274 = io_rw_addr == 12'h336;
  assign _T_1276 = io_rw_addr == 12'hb16;
  assign _T_1278 = io_rw_addr == 12'hc16;
  assign _T_1280 = io_rw_addr == 12'h337;
  assign _T_1282 = io_rw_addr == 12'hb17;
  assign _T_1284 = io_rw_addr == 12'hc17;
  assign _T_1286 = io_rw_addr == 12'h338;
  assign _T_1288 = io_rw_addr == 12'hb18;
  assign _T_1290 = io_rw_addr == 12'hc18;
  assign _T_1292 = io_rw_addr == 12'h339;
  assign _T_1294 = io_rw_addr == 12'hb19;
  assign _T_1296 = io_rw_addr == 12'hc19;
  assign _T_1298 = io_rw_addr == 12'h33a;
  assign _T_1300 = io_rw_addr == 12'hb1a;
  assign _T_1302 = io_rw_addr == 12'hc1a;
  assign _T_1304 = io_rw_addr == 12'h33b;
  assign _T_1306 = io_rw_addr == 12'hb1b;
  assign _T_1308 = io_rw_addr == 12'hc1b;
  assign _T_1310 = io_rw_addr == 12'h33c;
  assign _T_1312 = io_rw_addr == 12'hb1c;
  assign _T_1314 = io_rw_addr == 12'hc1c;
  assign _T_1316 = io_rw_addr == 12'h33d;
  assign _T_1318 = io_rw_addr == 12'hb1d;
  assign _T_1320 = io_rw_addr == 12'hc1d;
  assign _T_1322 = io_rw_addr == 12'h33e;
  assign _T_1324 = io_rw_addr == 12'hb1e;
  assign _T_1326 = io_rw_addr == 12'hc1e;
  assign _T_1328 = io_rw_addr == 12'h33f;
  assign _T_1330 = io_rw_addr == 12'hb1f;
  assign _T_1332 = io_rw_addr == 12'hc1f;
  assign _T_1334 = io_rw_addr == 12'h306;
  assign _T_1336 = io_rw_addr == 12'hc00;
  assign _T_1338 = io_rw_addr == 12'hc02;
  assign _T_1340 = io_rw_addr == 12'h100;
  assign _T_1342 = io_rw_addr == 12'h144;
  assign _T_1344 = io_rw_addr == 12'h104;
  assign _T_1346 = io_rw_addr == 12'h140;
  assign _T_1348 = io_rw_addr == 12'h142;
  assign _T_1350 = io_rw_addr == 12'h143;
  assign _T_1352 = io_rw_addr == 12'h180;
  assign _T_1354 = io_rw_addr == 12'h141;
  assign _T_1356 = io_rw_addr == 12'h105;
  assign _T_1358 = io_rw_addr == 12'h106;
  assign _T_1360 = io_rw_addr == 12'h303;
  assign _T_1362 = io_rw_addr == 12'h302;
  assign _T_1365 = io_rw_cmd == 3'h2;
  assign _T_1366 = io_rw_cmd == 3'h3;
  assign _T_1367 = _T_1365 | _T_1366;
  assign _T_1369 = _T_1367 ? io_rw_rdata : 64'h0;
  assign _T_1370 = _T_1369 | io_rw_wdata;
  assign _T_1374 = _T_1366 ? io_rw_wdata : 64'h0;
  assign _T_1375 = ~ _T_1374;
  assign wdata = _T_1370 & _T_1375;
  assign system_insn = io_rw_cmd == 3'h4;
  assign _T_1378 = io_rw_addr[2:0];
  assign opcode = 8'h1 << _T_1378;
  assign _T_1379 = opcode[0];
  assign insn_call = system_insn & _T_1379;
  assign _T_1380 = opcode[1];
  assign insn_break = system_insn & _T_1380;
  assign _T_1381 = opcode[2];
  assign insn_ret = system_insn & _T_1381;
  assign _T_1382 = opcode[5];
  assign insn_wfi = system_insn & _T_1382;
  assign _T_1385 = reg_mstatus_prv > 2'h1;
  assign _T_1388 = reg_mstatus_tw == 1'h0;
  assign _T_1389 = _T_1385 | _T_1388;
  assign _T_1395 = reg_mstatus_tvm == 1'h0;
  assign _T_1396 = _T_1385 | _T_1395;
  assign _T_1402 = reg_mstatus_tsr == 1'h0;
  assign _T_1403 = _T_1385 | _T_1402;
  assign _T_1405 = io_status_fs == 2'h0;
  assign _T_1406 = reg_misa[5];
  assign _T_1408 = _T_1406 == 1'h0;
  assign _T_1409 = _T_1405 | _T_1408;
  assign _T_1416 = io_decode_0_csr[9:8];
  assign _T_1417 = reg_mstatus_prv < _T_1416;
  assign _T_1419 = io_decode_0_csr == 12'h7a0;
  assign _T_1421 = io_decode_0_csr == 12'h7a1;
  assign _T_1423 = io_decode_0_csr == 12'h7a2;
  assign _T_1425 = io_decode_0_csr == 12'hf13;
  assign _T_1427 = io_decode_0_csr == 12'hf12;
  assign _T_1429 = io_decode_0_csr == 12'hf11;
  assign _T_1431 = io_decode_0_csr == 12'h301;
  assign _T_1433 = io_decode_0_csr == 12'h300;
  assign _T_1435 = io_decode_0_csr == 12'h305;
  assign _T_1437 = io_decode_0_csr == 12'h344;
  assign _T_1439 = io_decode_0_csr == 12'h304;
  assign _T_1441 = io_decode_0_csr == 12'h340;
  assign _T_1443 = io_decode_0_csr == 12'h341;
  assign _T_1445 = io_decode_0_csr == 12'h343;
  assign _T_1447 = io_decode_0_csr == 12'h342;
  assign _T_1449 = io_decode_0_csr == 12'hf14;
  assign _T_1451 = io_decode_0_csr == 12'h7b0;
  assign _T_1453 = io_decode_0_csr == 12'h7b1;
  assign _T_1455 = io_decode_0_csr == 12'h7b2;
  assign _T_1457 = io_decode_0_csr == 12'h1;
  assign _T_1459 = io_decode_0_csr == 12'h2;
  assign _T_1461 = io_decode_0_csr == 12'h3;
  assign _T_1463 = io_decode_0_csr == 12'hb00;
  assign _T_1465 = io_decode_0_csr == 12'hb02;
  assign _T_1467 = io_decode_0_csr == 12'h323;
  assign _T_1469 = io_decode_0_csr == 12'hb03;
  assign _T_1471 = io_decode_0_csr == 12'hc03;
  assign _T_1473 = io_decode_0_csr == 12'h324;
  assign _T_1475 = io_decode_0_csr == 12'hb04;
  assign _T_1477 = io_decode_0_csr == 12'hc04;
  assign _T_1479 = io_decode_0_csr == 12'h325;
  assign _T_1481 = io_decode_0_csr == 12'hb05;
  assign _T_1483 = io_decode_0_csr == 12'hc05;
  assign _T_1485 = io_decode_0_csr == 12'h326;
  assign _T_1487 = io_decode_0_csr == 12'hb06;
  assign _T_1489 = io_decode_0_csr == 12'hc06;
  assign _T_1491 = io_decode_0_csr == 12'h327;
  assign _T_1493 = io_decode_0_csr == 12'hb07;
  assign _T_1495 = io_decode_0_csr == 12'hc07;
  assign _T_1497 = io_decode_0_csr == 12'h328;
  assign _T_1499 = io_decode_0_csr == 12'hb08;
  assign _T_1501 = io_decode_0_csr == 12'hc08;
  assign _T_1503 = io_decode_0_csr == 12'h329;
  assign _T_1505 = io_decode_0_csr == 12'hb09;
  assign _T_1507 = io_decode_0_csr == 12'hc09;
  assign _T_1509 = io_decode_0_csr == 12'h32a;
  assign _T_1511 = io_decode_0_csr == 12'hb0a;
  assign _T_1513 = io_decode_0_csr == 12'hc0a;
  assign _T_1515 = io_decode_0_csr == 12'h32b;
  assign _T_1517 = io_decode_0_csr == 12'hb0b;
  assign _T_1519 = io_decode_0_csr == 12'hc0b;
  assign _T_1521 = io_decode_0_csr == 12'h32c;
  assign _T_1523 = io_decode_0_csr == 12'hb0c;
  assign _T_1525 = io_decode_0_csr == 12'hc0c;
  assign _T_1527 = io_decode_0_csr == 12'h32d;
  assign _T_1529 = io_decode_0_csr == 12'hb0d;
  assign _T_1531 = io_decode_0_csr == 12'hc0d;
  assign _T_1533 = io_decode_0_csr == 12'h32e;
  assign _T_1535 = io_decode_0_csr == 12'hb0e;
  assign _T_1537 = io_decode_0_csr == 12'hc0e;
  assign _T_1539 = io_decode_0_csr == 12'h32f;
  assign _T_1541 = io_decode_0_csr == 12'hb0f;
  assign _T_1543 = io_decode_0_csr == 12'hc0f;
  assign _T_1545 = io_decode_0_csr == 12'h330;
  assign _T_1547 = io_decode_0_csr == 12'hb10;
  assign _T_1549 = io_decode_0_csr == 12'hc10;
  assign _T_1551 = io_decode_0_csr == 12'h331;
  assign _T_1553 = io_decode_0_csr == 12'hb11;
  assign _T_1555 = io_decode_0_csr == 12'hc11;
  assign _T_1557 = io_decode_0_csr == 12'h332;
  assign _T_1559 = io_decode_0_csr == 12'hb12;
  assign _T_1561 = io_decode_0_csr == 12'hc12;
  assign _T_1563 = io_decode_0_csr == 12'h333;
  assign _T_1565 = io_decode_0_csr == 12'hb13;
  assign _T_1567 = io_decode_0_csr == 12'hc13;
  assign _T_1569 = io_decode_0_csr == 12'h334;
  assign _T_1571 = io_decode_0_csr == 12'hb14;
  assign _T_1573 = io_decode_0_csr == 12'hc14;
  assign _T_1575 = io_decode_0_csr == 12'h335;
  assign _T_1577 = io_decode_0_csr == 12'hb15;
  assign _T_1579 = io_decode_0_csr == 12'hc15;
  assign _T_1581 = io_decode_0_csr == 12'h336;
  assign _T_1583 = io_decode_0_csr == 12'hb16;
  assign _T_1585 = io_decode_0_csr == 12'hc16;
  assign _T_1587 = io_decode_0_csr == 12'h337;
  assign _T_1589 = io_decode_0_csr == 12'hb17;
  assign _T_1591 = io_decode_0_csr == 12'hc17;
  assign _T_1593 = io_decode_0_csr == 12'h338;
  assign _T_1595 = io_decode_0_csr == 12'hb18;
  assign _T_1597 = io_decode_0_csr == 12'hc18;
  assign _T_1599 = io_decode_0_csr == 12'h339;
  assign _T_1601 = io_decode_0_csr == 12'hb19;
  assign _T_1603 = io_decode_0_csr == 12'hc19;
  assign _T_1605 = io_decode_0_csr == 12'h33a;
  assign _T_1607 = io_decode_0_csr == 12'hb1a;
  assign _T_1609 = io_decode_0_csr == 12'hc1a;
  assign _T_1611 = io_decode_0_csr == 12'h33b;
  assign _T_1613 = io_decode_0_csr == 12'hb1b;
  assign _T_1615 = io_decode_0_csr == 12'hc1b;
  assign _T_1617 = io_decode_0_csr == 12'h33c;
  assign _T_1619 = io_decode_0_csr == 12'hb1c;
  assign _T_1621 = io_decode_0_csr == 12'hc1c;
  assign _T_1623 = io_decode_0_csr == 12'h33d;
  assign _T_1625 = io_decode_0_csr == 12'hb1d;
  assign _T_1627 = io_decode_0_csr == 12'hc1d;
  assign _T_1629 = io_decode_0_csr == 12'h33e;
  assign _T_1631 = io_decode_0_csr == 12'hb1e;
  assign _T_1633 = io_decode_0_csr == 12'hc1e;
  assign _T_1635 = io_decode_0_csr == 12'h33f;
  assign _T_1637 = io_decode_0_csr == 12'hb1f;
  assign _T_1639 = io_decode_0_csr == 12'hc1f;
  assign _T_1641 = io_decode_0_csr == 12'h306;
  assign _T_1643 = io_decode_0_csr == 12'hc00;
  assign _T_1645 = io_decode_0_csr == 12'hc02;
  assign _T_1647 = io_decode_0_csr == 12'h100;
  assign _T_1649 = io_decode_0_csr == 12'h144;
  assign _T_1651 = io_decode_0_csr == 12'h104;
  assign _T_1653 = io_decode_0_csr == 12'h140;
  assign _T_1655 = io_decode_0_csr == 12'h142;
  assign _T_1657 = io_decode_0_csr == 12'h143;
  assign _T_1659 = io_decode_0_csr == 12'h180;
  assign _T_1661 = io_decode_0_csr == 12'h141;
  assign _T_1663 = io_decode_0_csr == 12'h105;
  assign _T_1665 = io_decode_0_csr == 12'h106;
  assign _T_1667 = io_decode_0_csr == 12'h303;
  assign _T_1669 = io_decode_0_csr == 12'h302;
  assign _T_1670 = _T_1419 | _T_1421;
  assign _T_1671 = _T_1670 | _T_1423;
  assign _T_1672 = _T_1671 | _T_1425;
  assign _T_1673 = _T_1672 | _T_1427;
  assign _T_1674 = _T_1673 | _T_1429;
  assign _T_1675 = _T_1674 | _T_1431;
  assign _T_1676 = _T_1675 | _T_1433;
  assign _T_1677 = _T_1676 | _T_1435;
  assign _T_1678 = _T_1677 | _T_1437;
  assign _T_1679 = _T_1678 | _T_1439;
  assign _T_1680 = _T_1679 | _T_1441;
  assign _T_1681 = _T_1680 | _T_1443;
  assign _T_1682 = _T_1681 | _T_1445;
  assign _T_1683 = _T_1682 | _T_1447;
  assign _T_1684 = _T_1683 | _T_1449;
  assign _T_1685 = _T_1684 | _T_1451;
  assign _T_1686 = _T_1685 | _T_1453;
  assign _T_1687 = _T_1686 | _T_1455;
  assign _T_1688 = _T_1687 | _T_1457;
  assign _T_1689 = _T_1688 | _T_1459;
  assign _T_1690 = _T_1689 | _T_1461;
  assign _T_1691 = _T_1690 | _T_1463;
  assign _T_1692 = _T_1691 | _T_1465;
  assign _T_1693 = _T_1692 | _T_1467;
  assign _T_1694 = _T_1693 | _T_1469;
  assign _T_1695 = _T_1694 | _T_1471;
  assign _T_1696 = _T_1695 | _T_1473;
  assign _T_1697 = _T_1696 | _T_1475;
  assign _T_1698 = _T_1697 | _T_1477;
  assign _T_1699 = _T_1698 | _T_1479;
  assign _T_1700 = _T_1699 | _T_1481;
  assign _T_1701 = _T_1700 | _T_1483;
  assign _T_1702 = _T_1701 | _T_1485;
  assign _T_1703 = _T_1702 | _T_1487;
  assign _T_1704 = _T_1703 | _T_1489;
  assign _T_1705 = _T_1704 | _T_1491;
  assign _T_1706 = _T_1705 | _T_1493;
  assign _T_1707 = _T_1706 | _T_1495;
  assign _T_1708 = _T_1707 | _T_1497;
  assign _T_1709 = _T_1708 | _T_1499;
  assign _T_1710 = _T_1709 | _T_1501;
  assign _T_1711 = _T_1710 | _T_1503;
  assign _T_1712 = _T_1711 | _T_1505;
  assign _T_1713 = _T_1712 | _T_1507;
  assign _T_1714 = _T_1713 | _T_1509;
  assign _T_1715 = _T_1714 | _T_1511;
  assign _T_1716 = _T_1715 | _T_1513;
  assign _T_1717 = _T_1716 | _T_1515;
  assign _T_1718 = _T_1717 | _T_1517;
  assign _T_1719 = _T_1718 | _T_1519;
  assign _T_1720 = _T_1719 | _T_1521;
  assign _T_1721 = _T_1720 | _T_1523;
  assign _T_1722 = _T_1721 | _T_1525;
  assign _T_1723 = _T_1722 | _T_1527;
  assign _T_1724 = _T_1723 | _T_1529;
  assign _T_1725 = _T_1724 | _T_1531;
  assign _T_1726 = _T_1725 | _T_1533;
  assign _T_1727 = _T_1726 | _T_1535;
  assign _T_1728 = _T_1727 | _T_1537;
  assign _T_1729 = _T_1728 | _T_1539;
  assign _T_1730 = _T_1729 | _T_1541;
  assign _T_1731 = _T_1730 | _T_1543;
  assign _T_1732 = _T_1731 | _T_1545;
  assign _T_1733 = _T_1732 | _T_1547;
  assign _T_1734 = _T_1733 | _T_1549;
  assign _T_1735 = _T_1734 | _T_1551;
  assign _T_1736 = _T_1735 | _T_1553;
  assign _T_1737 = _T_1736 | _T_1555;
  assign _T_1738 = _T_1737 | _T_1557;
  assign _T_1739 = _T_1738 | _T_1559;
  assign _T_1740 = _T_1739 | _T_1561;
  assign _T_1741 = _T_1740 | _T_1563;
  assign _T_1742 = _T_1741 | _T_1565;
  assign _T_1743 = _T_1742 | _T_1567;
  assign _T_1744 = _T_1743 | _T_1569;
  assign _T_1745 = _T_1744 | _T_1571;
  assign _T_1746 = _T_1745 | _T_1573;
  assign _T_1747 = _T_1746 | _T_1575;
  assign _T_1748 = _T_1747 | _T_1577;
  assign _T_1749 = _T_1748 | _T_1579;
  assign _T_1750 = _T_1749 | _T_1581;
  assign _T_1751 = _T_1750 | _T_1583;
  assign _T_1752 = _T_1751 | _T_1585;
  assign _T_1753 = _T_1752 | _T_1587;
  assign _T_1754 = _T_1753 | _T_1589;
  assign _T_1755 = _T_1754 | _T_1591;
  assign _T_1756 = _T_1755 | _T_1593;
  assign _T_1757 = _T_1756 | _T_1595;
  assign _T_1758 = _T_1757 | _T_1597;
  assign _T_1759 = _T_1758 | _T_1599;
  assign _T_1760 = _T_1759 | _T_1601;
  assign _T_1761 = _T_1760 | _T_1603;
  assign _T_1762 = _T_1761 | _T_1605;
  assign _T_1763 = _T_1762 | _T_1607;
  assign _T_1764 = _T_1763 | _T_1609;
  assign _T_1765 = _T_1764 | _T_1611;
  assign _T_1766 = _T_1765 | _T_1613;
  assign _T_1767 = _T_1766 | _T_1615;
  assign _T_1768 = _T_1767 | _T_1617;
  assign _T_1769 = _T_1768 | _T_1619;
  assign _T_1770 = _T_1769 | _T_1621;
  assign _T_1771 = _T_1770 | _T_1623;
  assign _T_1772 = _T_1771 | _T_1625;
  assign _T_1773 = _T_1772 | _T_1627;
  assign _T_1774 = _T_1773 | _T_1629;
  assign _T_1775 = _T_1774 | _T_1631;
  assign _T_1776 = _T_1775 | _T_1633;
  assign _T_1777 = _T_1776 | _T_1635;
  assign _T_1778 = _T_1777 | _T_1637;
  assign _T_1779 = _T_1778 | _T_1639;
  assign _T_1780 = _T_1779 | _T_1641;
  assign _T_1781 = _T_1780 | _T_1643;
  assign _T_1782 = _T_1781 | _T_1645;
  assign _T_1783 = _T_1782 | _T_1647;
  assign _T_1784 = _T_1783 | _T_1649;
  assign _T_1785 = _T_1784 | _T_1651;
  assign _T_1786 = _T_1785 | _T_1653;
  assign _T_1787 = _T_1786 | _T_1655;
  assign _T_1788 = _T_1787 | _T_1657;
  assign _T_1789 = _T_1788 | _T_1659;
  assign _T_1790 = _T_1789 | _T_1661;
  assign _T_1791 = _T_1790 | _T_1663;
  assign _T_1792 = _T_1791 | _T_1665;
  assign _T_1793 = _T_1792 | _T_1667;
  assign _T_1794 = _T_1793 | _T_1669;
  assign _T_1796 = _T_1794 == 1'h0;
  assign _T_1797 = _T_1417 | _T_1796;
  assign _T_1801 = _T_1396 == 1'h0;
  assign _T_1802 = _T_1659 & _T_1801;
  assign _T_1803 = _T_1797 | _T_1802;
  assign _T_1806 = io_decode_0_csr >= 12'hc00;
  assign _T_1807 = io_decode_0_csr < 12'hc20;
  assign _T_1808 = _T_1806 & _T_1807;
  assign _T_1811 = io_decode_0_csr >= 12'hc80;
  assign _T_1812 = io_decode_0_csr < 12'hca0;
  assign _T_1813 = _T_1811 & _T_1812;
  assign _T_1814 = _T_1808 | _T_1813;
  assign _T_1817 = _T_1814 & _T_730;
  assign _T_1819 = hpm_mask >> io_decode_0_csr;
  assign _T_1820 = _T_1819[0];
  assign _T_1821 = _T_1817 & _T_1820;
  assign _T_1822 = _T_1803 | _T_1821;
  assign _T_1830 = _T_1451 | _T_1453;
  assign _T_1831 = _T_1830 | _T_1455;
  assign _T_1835 = _T_1831 & _T_933;
  assign _T_1836 = _T_1822 | _T_1835;
  assign _T_1844 = _T_1457 | _T_1459;
  assign _T_1845 = _T_1844 | _T_1461;
  assign _T_1847 = _T_1845 & io_decode_0_fp_illegal;
  assign _T_1848 = _T_1836 | _T_1847;
  assign _T_1849 = io_decode_0_csr[11:10];
  assign _T_1850 = ~ _T_1849;
  assign _T_1852 = _T_1850 == 2'h0;
  assign _T_1854 = io_decode_0_csr >= 12'h340;
  assign _T_1856 = io_decode_0_csr <= 12'h343;
  assign _T_1857 = _T_1854 & _T_1856;
  assign _T_1859 = io_decode_0_csr >= 12'h140;
  assign _T_1861 = io_decode_0_csr <= 12'h143;
  assign _T_1862 = _T_1859 & _T_1861;
  assign _T_1863 = _T_1857 | _T_1862;
  assign _T_1865 = _T_1863 == 1'h0;
  assign _T_1868 = io_decode_0_csr[5];
  assign _T_1870 = _T_1868 == 1'h0;
  assign _T_1871 = io_decode_0_csr[2];
  assign _T_1872 = _T_1870 & _T_1871;
  assign _T_1874 = _T_1389 == 1'h0;
  assign _T_1875 = _T_1872 & _T_1874;
  assign _T_1876 = _T_1417 | _T_1875;
  assign _T_1880 = io_decode_0_csr[1];
  assign _T_1881 = _T_1870 & _T_1880;
  assign _T_1883 = _T_1403 == 1'h0;
  assign _T_1884 = _T_1881 & _T_1883;
  assign _T_1885 = _T_1876 | _T_1884;
  assign _T_1889 = _T_1868 & _T_1801;
  assign _T_1890 = _T_1885 | _T_1889;
  assign _T_1924 = io_decode_1_csr[9:8];
  assign _T_1925 = reg_mstatus_prv < _T_1924;
  assign _T_1927 = io_decode_1_csr == 12'h7a0;
  assign _T_1929 = io_decode_1_csr == 12'h7a1;
  assign _T_1931 = io_decode_1_csr == 12'h7a2;
  assign _T_1933 = io_decode_1_csr == 12'hf13;
  assign _T_1935 = io_decode_1_csr == 12'hf12;
  assign _T_1937 = io_decode_1_csr == 12'hf11;
  assign _T_1939 = io_decode_1_csr == 12'h301;
  assign _T_1941 = io_decode_1_csr == 12'h300;
  assign _T_1943 = io_decode_1_csr == 12'h305;
  assign _T_1945 = io_decode_1_csr == 12'h344;
  assign _T_1947 = io_decode_1_csr == 12'h304;
  assign _T_1949 = io_decode_1_csr == 12'h340;
  assign _T_1951 = io_decode_1_csr == 12'h341;
  assign _T_1953 = io_decode_1_csr == 12'h343;
  assign _T_1955 = io_decode_1_csr == 12'h342;
  assign _T_1957 = io_decode_1_csr == 12'hf14;
  assign _T_1959 = io_decode_1_csr == 12'h7b0;
  assign _T_1961 = io_decode_1_csr == 12'h7b1;
  assign _T_1963 = io_decode_1_csr == 12'h7b2;
  assign _T_1965 = io_decode_1_csr == 12'h1;
  assign _T_1967 = io_decode_1_csr == 12'h2;
  assign _T_1969 = io_decode_1_csr == 12'h3;
  assign _T_1971 = io_decode_1_csr == 12'hb00;
  assign _T_1973 = io_decode_1_csr == 12'hb02;
  assign _T_1975 = io_decode_1_csr == 12'h323;
  assign _T_1977 = io_decode_1_csr == 12'hb03;
  assign _T_1979 = io_decode_1_csr == 12'hc03;
  assign _T_1981 = io_decode_1_csr == 12'h324;
  assign _T_1983 = io_decode_1_csr == 12'hb04;
  assign _T_1985 = io_decode_1_csr == 12'hc04;
  assign _T_1987 = io_decode_1_csr == 12'h325;
  assign _T_1989 = io_decode_1_csr == 12'hb05;
  assign _T_1991 = io_decode_1_csr == 12'hc05;
  assign _T_1993 = io_decode_1_csr == 12'h326;
  assign _T_1995 = io_decode_1_csr == 12'hb06;
  assign _T_1997 = io_decode_1_csr == 12'hc06;
  assign _T_1999 = io_decode_1_csr == 12'h327;
  assign _T_2001 = io_decode_1_csr == 12'hb07;
  assign _T_2003 = io_decode_1_csr == 12'hc07;
  assign _T_2005 = io_decode_1_csr == 12'h328;
  assign _T_2007 = io_decode_1_csr == 12'hb08;
  assign _T_2009 = io_decode_1_csr == 12'hc08;
  assign _T_2011 = io_decode_1_csr == 12'h329;
  assign _T_2013 = io_decode_1_csr == 12'hb09;
  assign _T_2015 = io_decode_1_csr == 12'hc09;
  assign _T_2017 = io_decode_1_csr == 12'h32a;
  assign _T_2019 = io_decode_1_csr == 12'hb0a;
  assign _T_2021 = io_decode_1_csr == 12'hc0a;
  assign _T_2023 = io_decode_1_csr == 12'h32b;
  assign _T_2025 = io_decode_1_csr == 12'hb0b;
  assign _T_2027 = io_decode_1_csr == 12'hc0b;
  assign _T_2029 = io_decode_1_csr == 12'h32c;
  assign _T_2031 = io_decode_1_csr == 12'hb0c;
  assign _T_2033 = io_decode_1_csr == 12'hc0c;
  assign _T_2035 = io_decode_1_csr == 12'h32d;
  assign _T_2037 = io_decode_1_csr == 12'hb0d;
  assign _T_2039 = io_decode_1_csr == 12'hc0d;
  assign _T_2041 = io_decode_1_csr == 12'h32e;
  assign _T_2043 = io_decode_1_csr == 12'hb0e;
  assign _T_2045 = io_decode_1_csr == 12'hc0e;
  assign _T_2047 = io_decode_1_csr == 12'h32f;
  assign _T_2049 = io_decode_1_csr == 12'hb0f;
  assign _T_2051 = io_decode_1_csr == 12'hc0f;
  assign _T_2053 = io_decode_1_csr == 12'h330;
  assign _T_2055 = io_decode_1_csr == 12'hb10;
  assign _T_2057 = io_decode_1_csr == 12'hc10;
  assign _T_2059 = io_decode_1_csr == 12'h331;
  assign _T_2061 = io_decode_1_csr == 12'hb11;
  assign _T_2063 = io_decode_1_csr == 12'hc11;
  assign _T_2065 = io_decode_1_csr == 12'h332;
  assign _T_2067 = io_decode_1_csr == 12'hb12;
  assign _T_2069 = io_decode_1_csr == 12'hc12;
  assign _T_2071 = io_decode_1_csr == 12'h333;
  assign _T_2073 = io_decode_1_csr == 12'hb13;
  assign _T_2075 = io_decode_1_csr == 12'hc13;
  assign _T_2077 = io_decode_1_csr == 12'h334;
  assign _T_2079 = io_decode_1_csr == 12'hb14;
  assign _T_2081 = io_decode_1_csr == 12'hc14;
  assign _T_2083 = io_decode_1_csr == 12'h335;
  assign _T_2085 = io_decode_1_csr == 12'hb15;
  assign _T_2087 = io_decode_1_csr == 12'hc15;
  assign _T_2089 = io_decode_1_csr == 12'h336;
  assign _T_2091 = io_decode_1_csr == 12'hb16;
  assign _T_2093 = io_decode_1_csr == 12'hc16;
  assign _T_2095 = io_decode_1_csr == 12'h337;
  assign _T_2097 = io_decode_1_csr == 12'hb17;
  assign _T_2099 = io_decode_1_csr == 12'hc17;
  assign _T_2101 = io_decode_1_csr == 12'h338;
  assign _T_2103 = io_decode_1_csr == 12'hb18;
  assign _T_2105 = io_decode_1_csr == 12'hc18;
  assign _T_2107 = io_decode_1_csr == 12'h339;
  assign _T_2109 = io_decode_1_csr == 12'hb19;
  assign _T_2111 = io_decode_1_csr == 12'hc19;
  assign _T_2113 = io_decode_1_csr == 12'h33a;
  assign _T_2115 = io_decode_1_csr == 12'hb1a;
  assign _T_2117 = io_decode_1_csr == 12'hc1a;
  assign _T_2119 = io_decode_1_csr == 12'h33b;
  assign _T_2121 = io_decode_1_csr == 12'hb1b;
  assign _T_2123 = io_decode_1_csr == 12'hc1b;
  assign _T_2125 = io_decode_1_csr == 12'h33c;
  assign _T_2127 = io_decode_1_csr == 12'hb1c;
  assign _T_2129 = io_decode_1_csr == 12'hc1c;
  assign _T_2131 = io_decode_1_csr == 12'h33d;
  assign _T_2133 = io_decode_1_csr == 12'hb1d;
  assign _T_2135 = io_decode_1_csr == 12'hc1d;
  assign _T_2137 = io_decode_1_csr == 12'h33e;
  assign _T_2139 = io_decode_1_csr == 12'hb1e;
  assign _T_2141 = io_decode_1_csr == 12'hc1e;
  assign _T_2143 = io_decode_1_csr == 12'h33f;
  assign _T_2145 = io_decode_1_csr == 12'hb1f;
  assign _T_2147 = io_decode_1_csr == 12'hc1f;
  assign _T_2149 = io_decode_1_csr == 12'h306;
  assign _T_2151 = io_decode_1_csr == 12'hc00;
  assign _T_2153 = io_decode_1_csr == 12'hc02;
  assign _T_2155 = io_decode_1_csr == 12'h100;
  assign _T_2157 = io_decode_1_csr == 12'h144;
  assign _T_2159 = io_decode_1_csr == 12'h104;
  assign _T_2161 = io_decode_1_csr == 12'h140;
  assign _T_2163 = io_decode_1_csr == 12'h142;
  assign _T_2165 = io_decode_1_csr == 12'h143;
  assign _T_2167 = io_decode_1_csr == 12'h180;
  assign _T_2169 = io_decode_1_csr == 12'h141;
  assign _T_2171 = io_decode_1_csr == 12'h105;
  assign _T_2173 = io_decode_1_csr == 12'h106;
  assign _T_2175 = io_decode_1_csr == 12'h303;
  assign _T_2177 = io_decode_1_csr == 12'h302;
  assign _T_2178 = _T_1927 | _T_1929;
  assign _T_2179 = _T_2178 | _T_1931;
  assign _T_2180 = _T_2179 | _T_1933;
  assign _T_2181 = _T_2180 | _T_1935;
  assign _T_2182 = _T_2181 | _T_1937;
  assign _T_2183 = _T_2182 | _T_1939;
  assign _T_2184 = _T_2183 | _T_1941;
  assign _T_2185 = _T_2184 | _T_1943;
  assign _T_2186 = _T_2185 | _T_1945;
  assign _T_2187 = _T_2186 | _T_1947;
  assign _T_2188 = _T_2187 | _T_1949;
  assign _T_2189 = _T_2188 | _T_1951;
  assign _T_2190 = _T_2189 | _T_1953;
  assign _T_2191 = _T_2190 | _T_1955;
  assign _T_2192 = _T_2191 | _T_1957;
  assign _T_2193 = _T_2192 | _T_1959;
  assign _T_2194 = _T_2193 | _T_1961;
  assign _T_2195 = _T_2194 | _T_1963;
  assign _T_2196 = _T_2195 | _T_1965;
  assign _T_2197 = _T_2196 | _T_1967;
  assign _T_2198 = _T_2197 | _T_1969;
  assign _T_2199 = _T_2198 | _T_1971;
  assign _T_2200 = _T_2199 | _T_1973;
  assign _T_2201 = _T_2200 | _T_1975;
  assign _T_2202 = _T_2201 | _T_1977;
  assign _T_2203 = _T_2202 | _T_1979;
  assign _T_2204 = _T_2203 | _T_1981;
  assign _T_2205 = _T_2204 | _T_1983;
  assign _T_2206 = _T_2205 | _T_1985;
  assign _T_2207 = _T_2206 | _T_1987;
  assign _T_2208 = _T_2207 | _T_1989;
  assign _T_2209 = _T_2208 | _T_1991;
  assign _T_2210 = _T_2209 | _T_1993;
  assign _T_2211 = _T_2210 | _T_1995;
  assign _T_2212 = _T_2211 | _T_1997;
  assign _T_2213 = _T_2212 | _T_1999;
  assign _T_2214 = _T_2213 | _T_2001;
  assign _T_2215 = _T_2214 | _T_2003;
  assign _T_2216 = _T_2215 | _T_2005;
  assign _T_2217 = _T_2216 | _T_2007;
  assign _T_2218 = _T_2217 | _T_2009;
  assign _T_2219 = _T_2218 | _T_2011;
  assign _T_2220 = _T_2219 | _T_2013;
  assign _T_2221 = _T_2220 | _T_2015;
  assign _T_2222 = _T_2221 | _T_2017;
  assign _T_2223 = _T_2222 | _T_2019;
  assign _T_2224 = _T_2223 | _T_2021;
  assign _T_2225 = _T_2224 | _T_2023;
  assign _T_2226 = _T_2225 | _T_2025;
  assign _T_2227 = _T_2226 | _T_2027;
  assign _T_2228 = _T_2227 | _T_2029;
  assign _T_2229 = _T_2228 | _T_2031;
  assign _T_2230 = _T_2229 | _T_2033;
  assign _T_2231 = _T_2230 | _T_2035;
  assign _T_2232 = _T_2231 | _T_2037;
  assign _T_2233 = _T_2232 | _T_2039;
  assign _T_2234 = _T_2233 | _T_2041;
  assign _T_2235 = _T_2234 | _T_2043;
  assign _T_2236 = _T_2235 | _T_2045;
  assign _T_2237 = _T_2236 | _T_2047;
  assign _T_2238 = _T_2237 | _T_2049;
  assign _T_2239 = _T_2238 | _T_2051;
  assign _T_2240 = _T_2239 | _T_2053;
  assign _T_2241 = _T_2240 | _T_2055;
  assign _T_2242 = _T_2241 | _T_2057;
  assign _T_2243 = _T_2242 | _T_2059;
  assign _T_2244 = _T_2243 | _T_2061;
  assign _T_2245 = _T_2244 | _T_2063;
  assign _T_2246 = _T_2245 | _T_2065;
  assign _T_2247 = _T_2246 | _T_2067;
  assign _T_2248 = _T_2247 | _T_2069;
  assign _T_2249 = _T_2248 | _T_2071;
  assign _T_2250 = _T_2249 | _T_2073;
  assign _T_2251 = _T_2250 | _T_2075;
  assign _T_2252 = _T_2251 | _T_2077;
  assign _T_2253 = _T_2252 | _T_2079;
  assign _T_2254 = _T_2253 | _T_2081;
  assign _T_2255 = _T_2254 | _T_2083;
  assign _T_2256 = _T_2255 | _T_2085;
  assign _T_2257 = _T_2256 | _T_2087;
  assign _T_2258 = _T_2257 | _T_2089;
  assign _T_2259 = _T_2258 | _T_2091;
  assign _T_2260 = _T_2259 | _T_2093;
  assign _T_2261 = _T_2260 | _T_2095;
  assign _T_2262 = _T_2261 | _T_2097;
  assign _T_2263 = _T_2262 | _T_2099;
  assign _T_2264 = _T_2263 | _T_2101;
  assign _T_2265 = _T_2264 | _T_2103;
  assign _T_2266 = _T_2265 | _T_2105;
  assign _T_2267 = _T_2266 | _T_2107;
  assign _T_2268 = _T_2267 | _T_2109;
  assign _T_2269 = _T_2268 | _T_2111;
  assign _T_2270 = _T_2269 | _T_2113;
  assign _T_2271 = _T_2270 | _T_2115;
  assign _T_2272 = _T_2271 | _T_2117;
  assign _T_2273 = _T_2272 | _T_2119;
  assign _T_2274 = _T_2273 | _T_2121;
  assign _T_2275 = _T_2274 | _T_2123;
  assign _T_2276 = _T_2275 | _T_2125;
  assign _T_2277 = _T_2276 | _T_2127;
  assign _T_2278 = _T_2277 | _T_2129;
  assign _T_2279 = _T_2278 | _T_2131;
  assign _T_2280 = _T_2279 | _T_2133;
  assign _T_2281 = _T_2280 | _T_2135;
  assign _T_2282 = _T_2281 | _T_2137;
  assign _T_2283 = _T_2282 | _T_2139;
  assign _T_2284 = _T_2283 | _T_2141;
  assign _T_2285 = _T_2284 | _T_2143;
  assign _T_2286 = _T_2285 | _T_2145;
  assign _T_2287 = _T_2286 | _T_2147;
  assign _T_2288 = _T_2287 | _T_2149;
  assign _T_2289 = _T_2288 | _T_2151;
  assign _T_2290 = _T_2289 | _T_2153;
  assign _T_2291 = _T_2290 | _T_2155;
  assign _T_2292 = _T_2291 | _T_2157;
  assign _T_2293 = _T_2292 | _T_2159;
  assign _T_2294 = _T_2293 | _T_2161;
  assign _T_2295 = _T_2294 | _T_2163;
  assign _T_2296 = _T_2295 | _T_2165;
  assign _T_2297 = _T_2296 | _T_2167;
  assign _T_2298 = _T_2297 | _T_2169;
  assign _T_2299 = _T_2298 | _T_2171;
  assign _T_2300 = _T_2299 | _T_2173;
  assign _T_2301 = _T_2300 | _T_2175;
  assign _T_2302 = _T_2301 | _T_2177;
  assign _T_2304 = _T_2302 == 1'h0;
  assign _T_2305 = _T_1925 | _T_2304;
  assign _T_2310 = _T_2167 & _T_1801;
  assign _T_2311 = _T_2305 | _T_2310;
  assign _T_2314 = io_decode_1_csr >= 12'hc00;
  assign _T_2315 = io_decode_1_csr < 12'hc20;
  assign _T_2316 = _T_2314 & _T_2315;
  assign _T_2319 = io_decode_1_csr >= 12'hc80;
  assign _T_2320 = io_decode_1_csr < 12'hca0;
  assign _T_2321 = _T_2319 & _T_2320;
  assign _T_2322 = _T_2316 | _T_2321;
  assign _T_2325 = _T_2322 & _T_730;
  assign _T_2327 = hpm_mask >> io_decode_1_csr;
  assign _T_2328 = _T_2327[0];
  assign _T_2329 = _T_2325 & _T_2328;
  assign _T_2330 = _T_2311 | _T_2329;
  assign _T_2338 = _T_1959 | _T_1961;
  assign _T_2339 = _T_2338 | _T_1963;
  assign _T_2343 = _T_2339 & _T_933;
  assign _T_2344 = _T_2330 | _T_2343;
  assign _T_2352 = _T_1965 | _T_1967;
  assign _T_2353 = _T_2352 | _T_1969;
  assign _T_2355 = _T_2353 & io_decode_1_fp_illegal;
  assign _T_2356 = _T_2344 | _T_2355;
  assign _T_2357 = io_decode_1_csr[11:10];
  assign _T_2358 = ~ _T_2357;
  assign _T_2360 = _T_2358 == 2'h0;
  assign _T_2362 = io_decode_1_csr >= 12'h340;
  assign _T_2364 = io_decode_1_csr <= 12'h343;
  assign _T_2365 = _T_2362 & _T_2364;
  assign _T_2367 = io_decode_1_csr >= 12'h140;
  assign _T_2369 = io_decode_1_csr <= 12'h143;
  assign _T_2370 = _T_2367 & _T_2369;
  assign _T_2371 = _T_2365 | _T_2370;
  assign _T_2373 = _T_2371 == 1'h0;
  assign _T_2376 = io_decode_1_csr[5];
  assign _T_2378 = _T_2376 == 1'h0;
  assign _T_2379 = io_decode_1_csr[2];
  assign _T_2380 = _T_2378 & _T_2379;
  assign _T_2383 = _T_2380 & _T_1874;
  assign _T_2384 = _T_1925 | _T_2383;
  assign _T_2388 = io_decode_1_csr[1];
  assign _T_2389 = _T_2378 & _T_2388;
  assign _T_2392 = _T_2389 & _T_1883;
  assign _T_2393 = _T_2384 | _T_2392;
  assign _T_2397 = _T_2376 & _T_1801;
  assign _T_2398 = _T_2393 | _T_2397;
  assign _GEN_605 = {{2'd0}, reg_mstatus_prv};
  assign _T_2400 = _GEN_605 + 4'h8;
  assign _T_2401 = _T_2400[3:0];
  assign _T_2403 = insn_break ? 64'h3 : io_cause;
  assign cause = insn_call ? {{60'd0}, _T_2401} : _T_2403;
  assign cause_lsbs = cause[7:0];
  assign _T_2404 = cause[63];
  assign _T_2406 = cause_lsbs == 8'he;
  assign causeIsDebugInt = _T_2404 & _T_2406;
  assign _T_2409 = _T_2404 == 1'h0;
  assign causeIsDebugTrigger = _T_2409 & _T_2406;
  assign _T_2415 = _T_2409 & insn_break;
  assign _T_2416 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign _T_2417 = {reg_dcsr_ebreakm,1'h0};
  assign _T_2418 = {_T_2417,_T_2416};
  assign _T_2419 = _T_2418 >> reg_mstatus_prv;
  assign _T_2420 = _T_2419[0];
  assign causeIsDebugBreak = _T_2415 & _T_2420;
  assign _T_2422 = reg_singleStepped | causeIsDebugInt;
  assign _T_2423 = _T_2422 | causeIsDebugTrigger;
  assign _T_2424 = _T_2423 | causeIsDebugBreak;
  assign trapToDebug = _T_2424 | reg_debug;
  assign _T_2428 = insn_break ? 12'h800 : 12'h808;
  assign debugTVec = reg_debug ? _T_2428 : 12'h800;
  assign _T_2435 = reg_mideleg >> cause_lsbs;
  assign _T_2436 = _T_2435[0];
  assign _T_2437 = reg_medeleg >> cause_lsbs;
  assign _T_2438 = _T_2437[0];
  assign _T_2439 = _T_2404 ? _T_2436 : _T_2438;
  assign delegate = _T_730 & _T_2439;
  assign _T_2444 = {_T_1104,reg_stvec};
  assign _T_2445 = delegate ? _T_2444 : {{8'd0}, reg_mtvec};
  assign _T_2446 = cause[3:0];
  assign _GEN_606 = {{2'd0}, _T_2446};
  assign _T_2447 = _GEN_606 << 2;
  assign _T_2448 = _T_2445[39:6];
  assign _T_2449 = {_T_2448,_T_2447};
  assign _T_2450 = _T_2445[0];
  assign _T_2452 = _T_2450 & _T_2404;
  assign _T_2453 = cause_lsbs[7:4];
  assign _T_2455 = _T_2453 == 4'h0;
  assign _T_2456 = _T_2452 & _T_2455;
  assign notDebugTVec = _T_2456 ? _T_2449 : _T_2445;
  assign tvec = trapToDebug ? {{28'd0}, debugTVec} : notDebugTVec;
  assign _T_2457 = insn_call | insn_break;
  assign _T_2458 = _T_2457 | insn_ret;
  assign _T_2461 = reg_dcsr_step & _T_933;
  assign _T_2462 = ~ io_status_fs;
  assign _T_2464 = _T_2462 == 2'h0;
  assign _T_2465 = ~ io_status_xs;
  assign _T_2467 = _T_2465 == 2'h0;
  assign _T_2468 = _T_2464 | _T_2467;
  assign _T_2473 = reg_mstatus_mprv & _T_933;
  assign _T_2474 = _T_2473 ? reg_mstatus_mpp : reg_mstatus_prv;
  assign exception = _T_2457 | io_exception;
  assign _T_2478 = insn_ret + insn_call;
  assign _T_2479 = insn_break + io_exception;
  assign _T_2480 = _T_2478 + _T_2479;
  assign _T_2482 = _T_2480 <= 3'h1;
  assign _T_2484 = _T_2482 | reset;
  assign _T_2486 = _T_2484 == 1'h0;
  assign _T_2489 = insn_wfi & _T_936;
  assign _T_2492 = _T_2489 & _T_933;
  assign _GEN_83 = _T_2492 ? 1'h1 : reg_wfi;
  assign _T_2495 = pending_interrupts != 64'h0;
  assign _T_2496 = _T_2495 | exception;
  assign _T_2497 = _T_2496 | io_interrupts_debug;
  assign _GEN_84 = _T_2497 ? 1'h0 : _GEN_83;
  assign _T_2500 = reg_wfi == 1'h0;
  assign _T_2502 = io_retire == 2'h0;
  assign _T_2503 = _T_2500 | _T_2502;
  assign _T_2505 = _T_2503 | reset;
  assign _T_2507 = _T_2505 == 1'h0;
  assign _T_2508 = io_retire[0];
  assign _T_2509 = _T_2508 | exception;
  assign _GEN_85 = _T_2509 ? 1'h1 : reg_singleStepped;
  assign _GEN_86 = _T_936 ? 1'h0 : _GEN_85;
  assign _T_2517 = io_retire <= 2'h1;
  assign _T_2518 = _T_936 | _T_2517;
  assign _T_2520 = _T_2518 | reset;
  assign _T_2522 = _T_2520 == 1'h0;
  assign _T_2524 = reg_singleStepped == 1'h0;
  assign _T_2527 = _T_2524 | _T_2502;
  assign _T_2529 = _T_2527 | reset;
  assign _T_2531 = _T_2529 == 1'h0;
  assign _T_2532 = ~ io_pc;
  assign _T_2534 = _T_2532 | 40'h3;
  assign epc = ~ _T_2534;
  assign _T_2545 = cause == 64'h2;
  assign _T_2546 = cause == 64'h3;
  assign _T_2547 = cause == 64'h4;
  assign _T_2548 = cause == 64'h6;
  assign _T_2549 = cause == 64'h5;
  assign _T_2550 = cause == 64'h7;
  assign _T_2551 = cause == 64'h1;
  assign _T_2552 = cause == 64'hd;
  assign _T_2553 = cause == 64'hf;
  assign _T_2554 = cause == 64'hc;
  assign _T_2555 = _T_2545 | _T_2546;
  assign _T_2556 = _T_2555 | _T_2547;
  assign _T_2557 = _T_2556 | _T_2548;
  assign _T_2558 = _T_2557 | _T_2549;
  assign _T_2559 = _T_2558 | _T_2550;
  assign _T_2560 = _T_2559 | _T_2551;
  assign _T_2561 = _T_2560 | _T_2552;
  assign _T_2562 = _T_2561 | _T_2553;
  assign _T_2563 = _T_2562 | _T_2554;
  assign write_badaddr = exception & _T_2563;
  assign badaddr_value = write_badaddr ? io_badaddr : 40'h0;
  assign _T_2572 = causeIsDebugTrigger ? 2'h2 : 2'h1;
  assign _T_2573 = causeIsDebugInt ? 2'h3 : _T_2572;
  assign _T_2574 = reg_singleStepped ? 3'h4 : {{1'd0}, _T_2573};
  assign _GEN_87 = _T_933 ? 1'h1 : reg_debug;
  assign _GEN_88 = _T_933 ? epc : reg_dpc;
  assign _GEN_89 = _T_933 ? _T_2574 : reg_dcsr_cause;
  assign _GEN_90 = _T_933 ? reg_mstatus_prv : reg_dcsr_prv;
  assign _GEN_91 = _T_933 ? 2'h3 : reg_mstatus_prv;
  assign _T_2576 = ~ epc;
  assign _T_2577 = reg_misa[2];
  assign _T_2579 = _T_2577 == 1'h0;
  assign _T_2581 = {_T_2579,1'h1};
  assign _GEN_607 = {{38'd0}, _T_2581};
  assign _T_2582 = _T_2576 | _GEN_607;
  assign _T_2583 = ~ _T_2582;
  assign _GEN_92 = delegate ? _T_2583 : reg_sepc;
  assign _GEN_93 = delegate ? cause : reg_scause;
  assign _GEN_94 = delegate ? badaddr_value : reg_sbadaddr;
  assign _GEN_95 = delegate ? reg_mstatus_sie : reg_mstatus_spie;
  assign _GEN_96 = delegate ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp};
  assign _GEN_97 = delegate ? 1'h0 : reg_mstatus_sie;
  assign _GEN_98 = delegate ? 2'h1 : 2'h3;
  assign _GEN_99 = delegate ? reg_mepc : _T_2583;
  assign _GEN_100 = delegate ? reg_mcause : cause;
  assign _GEN_101 = delegate ? reg_mbadaddr : badaddr_value;
  assign _GEN_102 = delegate ? reg_mstatus_mpie : reg_mstatus_mie;
  assign _GEN_103 = delegate ? reg_mstatus_mpp : reg_mstatus_prv;
  assign _GEN_104 = delegate ? reg_mstatus_mie : 1'h0;
  assign _GEN_105 = trapToDebug ? _GEN_87 : reg_debug;
  assign _GEN_106 = trapToDebug ? _GEN_88 : reg_dpc;
  assign _GEN_107 = trapToDebug ? _GEN_89 : reg_dcsr_cause;
  assign _GEN_108 = trapToDebug ? _GEN_90 : reg_dcsr_prv;
  assign _GEN_109 = trapToDebug ? _GEN_91 : _GEN_98;
  assign _GEN_110 = trapToDebug ? reg_sepc : _GEN_92;
  assign _GEN_111 = trapToDebug ? reg_scause : _GEN_93;
  assign _GEN_112 = trapToDebug ? reg_sbadaddr : _GEN_94;
  assign _GEN_113 = trapToDebug ? reg_mstatus_spie : _GEN_95;
  assign _GEN_114 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_96;
  assign _GEN_115 = trapToDebug ? reg_mstatus_sie : _GEN_97;
  assign _GEN_116 = trapToDebug ? reg_mepc : _GEN_99;
  assign _GEN_117 = trapToDebug ? reg_mcause : _GEN_100;
  assign _GEN_118 = trapToDebug ? reg_mbadaddr : _GEN_101;
  assign _GEN_119 = trapToDebug ? reg_mstatus_mpie : _GEN_102;
  assign _GEN_120 = trapToDebug ? reg_mstatus_mpp : _GEN_103;
  assign _GEN_121 = trapToDebug ? reg_mstatus_mie : _GEN_104;
  assign _GEN_122 = exception ? _GEN_105 : reg_debug;
  assign _GEN_123 = exception ? _GEN_106 : reg_dpc;
  assign _GEN_124 = exception ? _GEN_107 : reg_dcsr_cause;
  assign _GEN_125 = exception ? _GEN_108 : reg_dcsr_prv;
  assign _GEN_126 = exception ? _GEN_109 : reg_mstatus_prv;
  assign _GEN_127 = exception ? _GEN_110 : reg_sepc;
  assign _GEN_128 = exception ? _GEN_111 : reg_scause;
  assign _GEN_129 = exception ? _GEN_112 : reg_sbadaddr;
  assign _GEN_130 = exception ? _GEN_113 : reg_mstatus_spie;
  assign _GEN_131 = exception ? _GEN_114 : {{1'd0}, reg_mstatus_spp};
  assign _GEN_132 = exception ? _GEN_115 : reg_mstatus_sie;
  assign _GEN_133 = exception ? _GEN_116 : reg_mepc;
  assign _GEN_134 = exception ? _GEN_117 : reg_mcause;
  assign _GEN_135 = exception ? _GEN_118 : reg_mbadaddr;
  assign _GEN_136 = exception ? _GEN_119 : reg_mstatus_mpie;
  assign _GEN_137 = exception ? _GEN_120 : reg_mstatus_mpp;
  assign _GEN_138 = exception ? _GEN_121 : reg_mstatus_mie;
  assign _T_2597 = io_rw_addr[9];
  assign _T_2599 = _T_2597 == 1'h0;
  assign _T_2604 = io_rw_addr[10];
  assign _GEN_139 = _T_2604 ? reg_dcsr_prv : reg_mstatus_mpp;
  assign _GEN_140 = _T_2604 ? 1'h0 : _GEN_122;
  assign _GEN_141 = _T_2604 ? reg_dpc : reg_mepc;
  assign _GEN_142 = _T_2604 ? _GEN_138 : reg_mstatus_mpie;
  assign _GEN_143 = _T_2604 ? _GEN_136 : 1'h1;
  assign _GEN_144 = _T_2604 ? _GEN_137 : 2'h0;
  assign _GEN_145 = _T_2599 ? reg_mstatus_spie : _GEN_132;
  assign _GEN_146 = _T_2599 ? 1'h1 : _GEN_130;
  assign _GEN_147 = _T_2599 ? 2'h0 : _GEN_131;
  assign _GEN_148 = _T_2599 ? {{1'd0}, reg_mstatus_spp} : _GEN_139;
  assign _GEN_149 = _T_2599 ? reg_sepc : _GEN_141;
  assign _GEN_150 = _T_2599 ? _GEN_122 : _GEN_140;
  assign _GEN_151 = _T_2599 ? _GEN_138 : _GEN_142;
  assign _GEN_152 = _T_2599 ? _GEN_136 : _GEN_143;
  assign _GEN_153 = _T_2599 ? _GEN_137 : _GEN_144;
  assign _GEN_154 = insn_ret ? _GEN_145 : _GEN_132;
  assign _GEN_155 = insn_ret ? _GEN_146 : _GEN_130;
  assign _GEN_156 = insn_ret ? _GEN_147 : _GEN_131;
  assign _GEN_157 = insn_ret ? _GEN_148 : _GEN_126;
  assign _GEN_158 = insn_ret ? _GEN_149 : tvec;
  assign _GEN_159 = insn_ret ? _GEN_150 : _GEN_122;
  assign _GEN_160 = insn_ret ? _GEN_151 : _GEN_138;
  assign _GEN_161 = insn_ret ? _GEN_152 : _GEN_136;
  assign _GEN_162 = insn_ret ? _GEN_153 : _GEN_137;
  assign _T_2617 = _T_1114 ? _T_983 : 64'h0;
  assign _T_2619 = _T_1116 ? _T_990 : 64'h0;
  assign _T_2627 = _T_1124 ? reg_misa : 64'h0;
  assign _T_2629 = _T_1126 ? read_mstatus : 64'h0;
  assign _T_2631 = _T_1128 ? reg_mtvec : 32'h0;
  assign _T_2633 = _T_1130 ? read_mip : 16'h0;
  assign _T_2635 = _T_1132 ? reg_mie : 64'h0;
  assign _T_2637 = _T_1134 ? reg_mscratch : 64'h0;
  assign _T_2639 = _T_1136 ? _T_999 : 64'h0;
  assign _T_2641 = _T_1138 ? _T_1005 : 64'h0;
  assign _T_2643 = _T_1140 ? reg_mcause : 64'h0;
  assign _T_2647 = _T_1144 ? _T_1018 : 32'h0;
  assign _T_2649 = _T_1146 ? reg_dpc : 40'h0;
  assign _T_2651 = _T_1148 ? reg_dscratch : 64'h0;
  assign _T_2653 = _T_1150 ? reg_fflags : 5'h0;
  assign _T_2655 = _T_1152 ? reg_frm : 3'h0;
  assign _T_2657 = _T_1154 ? _T_1019 : 8'h0;
  assign _T_2659 = _T_1156 ? _T_350 : 64'h0;
  assign _T_2661 = _T_1158 ? _T_337 : 64'h0;
  assign _T_2663 = _T_1160 ? reg_hpmevent_0 : 64'h0;
  assign _T_2665 = _T_1162 ? _T_418 : 40'h0;
  assign _T_2667 = _T_1164 ? _T_418 : 40'h0;
  assign _T_2669 = _T_1166 ? reg_hpmevent_1 : 64'h0;
  assign _T_2671 = _T_1168 ? _T_428 : 40'h0;
  assign _T_2673 = _T_1170 ? _T_428 : 40'h0;
  assign _T_2675 = _T_1172 ? reg_hpmevent_2 : 64'h0;
  assign _T_2677 = _T_1174 ? _T_438 : 40'h0;
  assign _T_2679 = _T_1176 ? _T_438 : 40'h0;
  assign _T_2681 = _T_1178 ? reg_hpmevent_3 : 64'h0;
  assign _T_2683 = _T_1180 ? _T_448 : 40'h0;
  assign _T_2685 = _T_1182 ? _T_448 : 40'h0;
  assign _T_2687 = _T_1184 ? reg_hpmevent_4 : 64'h0;
  assign _T_2689 = _T_1186 ? _T_458 : 40'h0;
  assign _T_2691 = _T_1188 ? _T_458 : 40'h0;
  assign _T_2693 = _T_1190 ? reg_hpmevent_5 : 64'h0;
  assign _T_2695 = _T_1192 ? _T_468 : 40'h0;
  assign _T_2697 = _T_1194 ? _T_468 : 40'h0;
  assign _T_2699 = _T_1196 ? reg_hpmevent_6 : 64'h0;
  assign _T_2701 = _T_1198 ? _T_478 : 40'h0;
  assign _T_2703 = _T_1200 ? _T_478 : 40'h0;
  assign _T_2705 = _T_1202 ? reg_hpmevent_7 : 64'h0;
  assign _T_2707 = _T_1204 ? _T_488 : 40'h0;
  assign _T_2709 = _T_1206 ? _T_488 : 40'h0;
  assign _T_2711 = _T_1208 ? reg_hpmevent_8 : 64'h0;
  assign _T_2713 = _T_1210 ? _T_498 : 40'h0;
  assign _T_2715 = _T_1212 ? _T_498 : 40'h0;
  assign _T_2717 = _T_1214 ? reg_hpmevent_9 : 64'h0;
  assign _T_2719 = _T_1216 ? _T_508 : 40'h0;
  assign _T_2721 = _T_1218 ? _T_508 : 40'h0;
  assign _T_2723 = _T_1220 ? reg_hpmevent_10 : 64'h0;
  assign _T_2725 = _T_1222 ? _T_518 : 40'h0;
  assign _T_2727 = _T_1224 ? _T_518 : 40'h0;
  assign _T_2729 = _T_1226 ? reg_hpmevent_11 : 64'h0;
  assign _T_2731 = _T_1228 ? _T_528 : 40'h0;
  assign _T_2733 = _T_1230 ? _T_528 : 40'h0;
  assign _T_2735 = _T_1232 ? reg_hpmevent_12 : 64'h0;
  assign _T_2737 = _T_1234 ? _T_538 : 40'h0;
  assign _T_2739 = _T_1236 ? _T_538 : 40'h0;
  assign _T_2741 = _T_1238 ? reg_hpmevent_13 : 64'h0;
  assign _T_2743 = _T_1240 ? _T_548 : 40'h0;
  assign _T_2745 = _T_1242 ? _T_548 : 40'h0;
  assign _T_2747 = _T_1244 ? reg_hpmevent_14 : 64'h0;
  assign _T_2749 = _T_1246 ? _T_558 : 40'h0;
  assign _T_2751 = _T_1248 ? _T_558 : 40'h0;
  assign _T_2753 = _T_1250 ? reg_hpmevent_15 : 64'h0;
  assign _T_2755 = _T_1252 ? _T_568 : 40'h0;
  assign _T_2757 = _T_1254 ? _T_568 : 40'h0;
  assign _T_2759 = _T_1256 ? reg_hpmevent_16 : 64'h0;
  assign _T_2761 = _T_1258 ? _T_578 : 40'h0;
  assign _T_2763 = _T_1260 ? _T_578 : 40'h0;
  assign _T_2765 = _T_1262 ? reg_hpmevent_17 : 64'h0;
  assign _T_2767 = _T_1264 ? _T_588 : 40'h0;
  assign _T_2769 = _T_1266 ? _T_588 : 40'h0;
  assign _T_2771 = _T_1268 ? reg_hpmevent_18 : 64'h0;
  assign _T_2773 = _T_1270 ? _T_598 : 40'h0;
  assign _T_2775 = _T_1272 ? _T_598 : 40'h0;
  assign _T_2777 = _T_1274 ? reg_hpmevent_19 : 64'h0;
  assign _T_2779 = _T_1276 ? _T_608 : 40'h0;
  assign _T_2781 = _T_1278 ? _T_608 : 40'h0;
  assign _T_2783 = _T_1280 ? reg_hpmevent_20 : 64'h0;
  assign _T_2785 = _T_1282 ? _T_618 : 40'h0;
  assign _T_2787 = _T_1284 ? _T_618 : 40'h0;
  assign _T_2789 = _T_1286 ? reg_hpmevent_21 : 64'h0;
  assign _T_2791 = _T_1288 ? _T_628 : 40'h0;
  assign _T_2793 = _T_1290 ? _T_628 : 40'h0;
  assign _T_2795 = _T_1292 ? reg_hpmevent_22 : 64'h0;
  assign _T_2797 = _T_1294 ? _T_638 : 40'h0;
  assign _T_2799 = _T_1296 ? _T_638 : 40'h0;
  assign _T_2801 = _T_1298 ? reg_hpmevent_23 : 64'h0;
  assign _T_2803 = _T_1300 ? _T_648 : 40'h0;
  assign _T_2805 = _T_1302 ? _T_648 : 40'h0;
  assign _T_2807 = _T_1304 ? reg_hpmevent_24 : 64'h0;
  assign _T_2809 = _T_1306 ? _T_658 : 40'h0;
  assign _T_2811 = _T_1308 ? _T_658 : 40'h0;
  assign _T_2813 = _T_1310 ? reg_hpmevent_25 : 64'h0;
  assign _T_2815 = _T_1312 ? _T_668 : 40'h0;
  assign _T_2817 = _T_1314 ? _T_668 : 40'h0;
  assign _T_2819 = _T_1316 ? reg_hpmevent_26 : 64'h0;
  assign _T_2821 = _T_1318 ? _T_678 : 40'h0;
  assign _T_2823 = _T_1320 ? _T_678 : 40'h0;
  assign _T_2825 = _T_1322 ? reg_hpmevent_27 : 64'h0;
  assign _T_2827 = _T_1324 ? _T_688 : 40'h0;
  assign _T_2829 = _T_1326 ? _T_688 : 40'h0;
  assign _T_2831 = _T_1328 ? reg_hpmevent_28 : 64'h0;
  assign _T_2833 = _T_1330 ? _T_698 : 40'h0;
  assign _T_2835 = _T_1332 ? _T_698 : 40'h0;
  assign _T_2837 = _T_1334 ? reg_mcounteren : 32'h0;
  assign _T_2839 = _T_1336 ? _T_350 : 64'h0;
  assign _T_2841 = _T_1338 ? _T_337 : 64'h0;
  assign _T_2843 = _T_1340 ? _T_1089 : 64'h0;
  assign _T_2845 = _T_1342 ? _T_1023 : 64'h0;
  assign _T_2847 = _T_1344 ? _T_1022 : 64'h0;
  assign _T_2849 = _T_1346 ? reg_sscratch : 64'h0;
  assign _T_2851 = _T_1348 ? reg_scause : 64'h0;
  assign _T_2853 = _T_1350 ? _T_1095 : 64'h0;
  assign _T_2855 = _T_1352 ? _T_1097 : 64'h0;
  assign _T_2857 = _T_1354 ? _T_1103 : 64'h0;
  assign _T_2859 = _T_1356 ? _T_1109 : 64'h0;
  assign _T_2861 = _T_1358 ? reg_scounteren : 32'h0;
  assign _T_2863 = _T_1360 ? reg_mideleg : 64'h0;
  assign _T_2865 = _T_1362 ? reg_medeleg : 64'h0;
  assign _T_2867 = _T_2617 | _T_2619;
  assign _T_2871 = _T_2867 | _T_2627;
  assign _T_2872 = _T_2871 | _T_2629;
  assign _GEN_609 = {{32'd0}, _T_2631};
  assign _T_2873 = _T_2872 | _GEN_609;
  assign _GEN_610 = {{48'd0}, _T_2633};
  assign _T_2874 = _T_2873 | _GEN_610;
  assign _T_2875 = _T_2874 | _T_2635;
  assign _T_2876 = _T_2875 | _T_2637;
  assign _T_2877 = _T_2876 | _T_2639;
  assign _T_2878 = _T_2877 | _T_2641;
  assign _T_2879 = _T_2878 | _T_2643;
  assign _GEN_611 = {{32'd0}, _T_2647};
  assign _T_2881 = _T_2879 | _GEN_611;
  assign _GEN_612 = {{24'd0}, _T_2649};
  assign _T_2882 = _T_2881 | _GEN_612;
  assign _T_2883 = _T_2882 | _T_2651;
  assign _GEN_613 = {{59'd0}, _T_2653};
  assign _T_2884 = _T_2883 | _GEN_613;
  assign _GEN_614 = {{61'd0}, _T_2655};
  assign _T_2885 = _T_2884 | _GEN_614;
  assign _GEN_615 = {{56'd0}, _T_2657};
  assign _T_2886 = _T_2885 | _GEN_615;
  assign _T_2887 = _T_2886 | _T_2659;
  assign _T_2888 = _T_2887 | _T_2661;
  assign _T_2889 = _T_2888 | _T_2663;
  assign _GEN_616 = {{24'd0}, _T_2665};
  assign _T_2890 = _T_2889 | _GEN_616;
  assign _GEN_617 = {{24'd0}, _T_2667};
  assign _T_2891 = _T_2890 | _GEN_617;
  assign _T_2892 = _T_2891 | _T_2669;
  assign _GEN_618 = {{24'd0}, _T_2671};
  assign _T_2893 = _T_2892 | _GEN_618;
  assign _GEN_619 = {{24'd0}, _T_2673};
  assign _T_2894 = _T_2893 | _GEN_619;
  assign _T_2895 = _T_2894 | _T_2675;
  assign _GEN_620 = {{24'd0}, _T_2677};
  assign _T_2896 = _T_2895 | _GEN_620;
  assign _GEN_621 = {{24'd0}, _T_2679};
  assign _T_2897 = _T_2896 | _GEN_621;
  assign _T_2898 = _T_2897 | _T_2681;
  assign _GEN_622 = {{24'd0}, _T_2683};
  assign _T_2899 = _T_2898 | _GEN_622;
  assign _GEN_623 = {{24'd0}, _T_2685};
  assign _T_2900 = _T_2899 | _GEN_623;
  assign _T_2901 = _T_2900 | _T_2687;
  assign _GEN_624 = {{24'd0}, _T_2689};
  assign _T_2902 = _T_2901 | _GEN_624;
  assign _GEN_625 = {{24'd0}, _T_2691};
  assign _T_2903 = _T_2902 | _GEN_625;
  assign _T_2904 = _T_2903 | _T_2693;
  assign _GEN_626 = {{24'd0}, _T_2695};
  assign _T_2905 = _T_2904 | _GEN_626;
  assign _GEN_627 = {{24'd0}, _T_2697};
  assign _T_2906 = _T_2905 | _GEN_627;
  assign _T_2907 = _T_2906 | _T_2699;
  assign _GEN_628 = {{24'd0}, _T_2701};
  assign _T_2908 = _T_2907 | _GEN_628;
  assign _GEN_629 = {{24'd0}, _T_2703};
  assign _T_2909 = _T_2908 | _GEN_629;
  assign _T_2910 = _T_2909 | _T_2705;
  assign _GEN_630 = {{24'd0}, _T_2707};
  assign _T_2911 = _T_2910 | _GEN_630;
  assign _GEN_631 = {{24'd0}, _T_2709};
  assign _T_2912 = _T_2911 | _GEN_631;
  assign _T_2913 = _T_2912 | _T_2711;
  assign _GEN_632 = {{24'd0}, _T_2713};
  assign _T_2914 = _T_2913 | _GEN_632;
  assign _GEN_633 = {{24'd0}, _T_2715};
  assign _T_2915 = _T_2914 | _GEN_633;
  assign _T_2916 = _T_2915 | _T_2717;
  assign _GEN_634 = {{24'd0}, _T_2719};
  assign _T_2917 = _T_2916 | _GEN_634;
  assign _GEN_635 = {{24'd0}, _T_2721};
  assign _T_2918 = _T_2917 | _GEN_635;
  assign _T_2919 = _T_2918 | _T_2723;
  assign _GEN_636 = {{24'd0}, _T_2725};
  assign _T_2920 = _T_2919 | _GEN_636;
  assign _GEN_637 = {{24'd0}, _T_2727};
  assign _T_2921 = _T_2920 | _GEN_637;
  assign _T_2922 = _T_2921 | _T_2729;
  assign _GEN_638 = {{24'd0}, _T_2731};
  assign _T_2923 = _T_2922 | _GEN_638;
  assign _GEN_639 = {{24'd0}, _T_2733};
  assign _T_2924 = _T_2923 | _GEN_639;
  assign _T_2925 = _T_2924 | _T_2735;
  assign _GEN_640 = {{24'd0}, _T_2737};
  assign _T_2926 = _T_2925 | _GEN_640;
  assign _GEN_641 = {{24'd0}, _T_2739};
  assign _T_2927 = _T_2926 | _GEN_641;
  assign _T_2928 = _T_2927 | _T_2741;
  assign _GEN_642 = {{24'd0}, _T_2743};
  assign _T_2929 = _T_2928 | _GEN_642;
  assign _GEN_643 = {{24'd0}, _T_2745};
  assign _T_2930 = _T_2929 | _GEN_643;
  assign _T_2931 = _T_2930 | _T_2747;
  assign _GEN_644 = {{24'd0}, _T_2749};
  assign _T_2932 = _T_2931 | _GEN_644;
  assign _GEN_645 = {{24'd0}, _T_2751};
  assign _T_2933 = _T_2932 | _GEN_645;
  assign _T_2934 = _T_2933 | _T_2753;
  assign _GEN_646 = {{24'd0}, _T_2755};
  assign _T_2935 = _T_2934 | _GEN_646;
  assign _GEN_647 = {{24'd0}, _T_2757};
  assign _T_2936 = _T_2935 | _GEN_647;
  assign _T_2937 = _T_2936 | _T_2759;
  assign _GEN_648 = {{24'd0}, _T_2761};
  assign _T_2938 = _T_2937 | _GEN_648;
  assign _GEN_649 = {{24'd0}, _T_2763};
  assign _T_2939 = _T_2938 | _GEN_649;
  assign _T_2940 = _T_2939 | _T_2765;
  assign _GEN_650 = {{24'd0}, _T_2767};
  assign _T_2941 = _T_2940 | _GEN_650;
  assign _GEN_651 = {{24'd0}, _T_2769};
  assign _T_2942 = _T_2941 | _GEN_651;
  assign _T_2943 = _T_2942 | _T_2771;
  assign _GEN_652 = {{24'd0}, _T_2773};
  assign _T_2944 = _T_2943 | _GEN_652;
  assign _GEN_653 = {{24'd0}, _T_2775};
  assign _T_2945 = _T_2944 | _GEN_653;
  assign _T_2946 = _T_2945 | _T_2777;
  assign _GEN_654 = {{24'd0}, _T_2779};
  assign _T_2947 = _T_2946 | _GEN_654;
  assign _GEN_655 = {{24'd0}, _T_2781};
  assign _T_2948 = _T_2947 | _GEN_655;
  assign _T_2949 = _T_2948 | _T_2783;
  assign _GEN_656 = {{24'd0}, _T_2785};
  assign _T_2950 = _T_2949 | _GEN_656;
  assign _GEN_657 = {{24'd0}, _T_2787};
  assign _T_2951 = _T_2950 | _GEN_657;
  assign _T_2952 = _T_2951 | _T_2789;
  assign _GEN_658 = {{24'd0}, _T_2791};
  assign _T_2953 = _T_2952 | _GEN_658;
  assign _GEN_659 = {{24'd0}, _T_2793};
  assign _T_2954 = _T_2953 | _GEN_659;
  assign _T_2955 = _T_2954 | _T_2795;
  assign _GEN_660 = {{24'd0}, _T_2797};
  assign _T_2956 = _T_2955 | _GEN_660;
  assign _GEN_661 = {{24'd0}, _T_2799};
  assign _T_2957 = _T_2956 | _GEN_661;
  assign _T_2958 = _T_2957 | _T_2801;
  assign _GEN_662 = {{24'd0}, _T_2803};
  assign _T_2959 = _T_2958 | _GEN_662;
  assign _GEN_663 = {{24'd0}, _T_2805};
  assign _T_2960 = _T_2959 | _GEN_663;
  assign _T_2961 = _T_2960 | _T_2807;
  assign _GEN_664 = {{24'd0}, _T_2809};
  assign _T_2962 = _T_2961 | _GEN_664;
  assign _GEN_665 = {{24'd0}, _T_2811};
  assign _T_2963 = _T_2962 | _GEN_665;
  assign _T_2964 = _T_2963 | _T_2813;
  assign _GEN_666 = {{24'd0}, _T_2815};
  assign _T_2965 = _T_2964 | _GEN_666;
  assign _GEN_667 = {{24'd0}, _T_2817};
  assign _T_2966 = _T_2965 | _GEN_667;
  assign _T_2967 = _T_2966 | _T_2819;
  assign _GEN_668 = {{24'd0}, _T_2821};
  assign _T_2968 = _T_2967 | _GEN_668;
  assign _GEN_669 = {{24'd0}, _T_2823};
  assign _T_2969 = _T_2968 | _GEN_669;
  assign _T_2970 = _T_2969 | _T_2825;
  assign _GEN_670 = {{24'd0}, _T_2827};
  assign _T_2971 = _T_2970 | _GEN_670;
  assign _GEN_671 = {{24'd0}, _T_2829};
  assign _T_2972 = _T_2971 | _GEN_671;
  assign _T_2973 = _T_2972 | _T_2831;
  assign _GEN_672 = {{24'd0}, _T_2833};
  assign _T_2974 = _T_2973 | _GEN_672;
  assign _GEN_673 = {{24'd0}, _T_2835};
  assign _T_2975 = _T_2974 | _GEN_673;
  assign _GEN_674 = {{32'd0}, _T_2837};
  assign _T_2976 = _T_2975 | _GEN_674;
  assign _T_2977 = _T_2976 | _T_2839;
  assign _T_2978 = _T_2977 | _T_2841;
  assign _T_2979 = _T_2978 | _T_2843;
  assign _T_2980 = _T_2979 | _T_2845;
  assign _T_2981 = _T_2980 | _T_2847;
  assign _T_2982 = _T_2981 | _T_2849;
  assign _T_2983 = _T_2982 | _T_2851;
  assign _T_2984 = _T_2983 | _T_2853;
  assign _T_2985 = _T_2984 | _T_2855;
  assign _T_2986 = _T_2985 | _T_2857;
  assign _T_2987 = _T_2986 | _T_2859;
  assign _GEN_675 = {{32'd0}, _T_2861};
  assign _T_2988 = _T_2987 | _GEN_675;
  assign _T_2989 = _T_2988 | _T_2863;
  assign _T_2990 = _T_2989 | _T_2865;
  assign _T_2993 = reg_fflags | io_fcsr_flags_bits;
  assign _GEN_163 = io_fcsr_flags_valid ? _T_2993 : reg_fflags;
  assign _T_2999 = io_rw_cmd == 3'h1;
  assign _T_3001 = _T_1367 | _T_2999;
  assign _T_3008 = _T_3006[1];
  assign _T_3010 = _T_3006[3];
  assign _T_3012 = _T_3006[5];
  assign _T_3014 = _T_3006[7];
  assign _T_3015 = _T_3006[8];
  assign _T_3017 = _T_3006[12:11];
  assign _T_3018 = _T_3006[14:13];
  assign _T_3020 = _T_3006[17];
  assign _T_3021 = _T_3006[18];
  assign _T_3022 = _T_3006[19];
  assign _T_3023 = _T_3006[20];
  assign _T_3024 = _T_3006[21];
  assign _T_3025 = _T_3006[22];
  assign _T_3037 = _T_3004_fs != 2'h0;
  assign _T_3041 = _T_3037 ? 2'h3 : 2'h0;
  assign _GEN_164 = _T_1126 ? _T_3004_mie : _GEN_160;
  assign _GEN_165 = _T_1126 ? _T_3004_mpie : _GEN_161;
  assign _GEN_166 = _T_1126 ? _T_3004_mprv : reg_mstatus_mprv;
  assign _GEN_167 = _T_1126 ? _T_3004_mpp : _GEN_162;
  assign _GEN_168 = _T_1126 ? _T_3004_mxr : reg_mstatus_mxr;
  assign _GEN_169 = _T_1126 ? _T_3004_sum : reg_mstatus_sum;
  assign _GEN_170 = _T_1126 ? {{1'd0}, _T_3004_spp} : _GEN_156;
  assign _GEN_171 = _T_1126 ? _T_3004_spie : _GEN_155;
  assign _GEN_172 = _T_1126 ? _T_3004_sie : _GEN_154;
  assign _GEN_173 = _T_1126 ? _T_3004_tw : reg_mstatus_tw;
  assign _GEN_174 = _T_1126 ? _T_3004_tvm : reg_mstatus_tvm;
  assign _GEN_175 = _T_1126 ? _T_3004_tsr : reg_mstatus_tsr;
  assign _GEN_176 = _T_1126 ? _T_3041 : reg_mstatus_fs;
  assign _T_3043 = wdata[5];
  assign _T_3044 = ~ wdata;
  assign _T_3046 = _T_3043 == 1'h0;
  assign _GEN_676 = {{3'd0}, _T_3046};
  assign _T_3047 = _GEN_676 << 3;
  assign _GEN_677 = {{60'd0}, _T_3047};
  assign _T_3048 = _T_3044 | _GEN_677;
  assign _T_3049 = ~ _T_3048;
  assign _T_3050 = _T_3049 & 64'h1029;
  assign _T_3052 = reg_misa & 64'hffffffffffffefd6;
  assign _T_3053 = _T_3050 | _T_3052;
  assign _GEN_177 = _T_1124 ? _T_3053 : reg_misa;
  assign _T_3054 = {reg_mip_ssip,1'h0};
  assign _T_3056 = {2'h0,_T_3054};
  assign _T_3057 = {reg_mip_stip,1'h0};
  assign _T_3059 = {2'h0,_T_3057};
  assign _T_3060 = {_T_3059,_T_3056};
  assign _T_3061 = {reg_mip_seip,1'h0};
  assign _T_3063 = {2'h0,_T_3061};
  assign _T_3067 = {4'h0,_T_3063};
  assign _T_3068 = {_T_3067,_T_3060};
  assign _T_3075 = _T_1367 ? _T_3068 : 16'h0;
  assign _GEN_678 = {{48'd0}, _T_3075};
  assign _T_3076 = _GEN_678 | io_rw_wdata;
  assign _T_3082 = _T_3076 & _T_1375;
  assign _T_3095 = _T_3093[1];
  assign _T_3099 = _T_3093[5];
  assign _T_3103 = _T_3093[9];
  assign _GEN_178 = _T_1130 ? _T_3089_ssip : reg_mip_ssip;
  assign _GEN_179 = _T_1130 ? _T_3089_stip : reg_mip_stip;
  assign _GEN_180 = _T_1130 ? _T_3089_seip : reg_mip_seip;
  assign _T_3110 = wdata & 64'haaa;
  assign _GEN_181 = _T_1132 ? _T_3110 : reg_mie;
  assign _GEN_679 = {{62'd0}, _T_2581};
  assign _T_3117 = _T_3044 | _GEN_679;
  assign _T_3118 = ~ _T_3117;
  assign _GEN_182 = _T_1136 ? _T_3118 : {{24'd0}, _GEN_133};
  assign _GEN_183 = _T_1134 ? wdata : reg_mscratch;
  assign _T_3121 = _T_3044 | 64'h2;
  assign _T_3122 = wdata[0];
  assign _T_3125 = _T_3122 ? 6'h3c : 6'h0;
  assign _GEN_680 = {{58'd0}, _T_3125};
  assign _T_3126 = _T_3121 | _GEN_680;
  assign _T_3127 = ~ _T_3126;
  assign _GEN_184 = _T_1128 ? _T_3127 : {{32'd0}, reg_mtvec};
  assign _T_3129 = wdata & 64'h800000000000000f;
  assign _GEN_185 = _T_1140 ? _T_3129 : _GEN_134;
  assign _T_3130 = wdata[39:0];
  assign _GEN_186 = _T_1138 ? _T_3130 : _GEN_135;
  assign _T_3132 = _T_3130[39:6];
  assign _GEN_187 = _T_1162 ? _T_3130 : {{33'd0}, _T_411};
  assign _GEN_188 = _T_1162 ? _T_3132 : _GEN_38;
  assign _T_3134 = wdata & 64'h3f03;
  assign _GEN_189 = _T_1160 ? _T_3134 : reg_hpmevent_0;
  assign _GEN_190 = _T_1168 ? _T_3130 : {{33'd0}, _T_421};
  assign _GEN_191 = _T_1168 ? _T_3132 : _GEN_39;
  assign _GEN_192 = _T_1166 ? _T_3134 : reg_hpmevent_1;
  assign _GEN_193 = _T_1174 ? _T_3130 : {{33'd0}, _T_431};
  assign _GEN_194 = _T_1174 ? _T_3132 : _GEN_40;
  assign _GEN_195 = _T_1172 ? _T_3134 : reg_hpmevent_2;
  assign _GEN_196 = _T_1180 ? _T_3130 : {{33'd0}, _T_441};
  assign _GEN_197 = _T_1180 ? _T_3132 : _GEN_41;
  assign _GEN_198 = _T_1178 ? _T_3134 : reg_hpmevent_3;
  assign _GEN_199 = _T_1186 ? _T_3130 : {{33'd0}, _T_451};
  assign _GEN_200 = _T_1186 ? _T_3132 : _GEN_42;
  assign _GEN_201 = _T_1184 ? _T_3134 : reg_hpmevent_4;
  assign _GEN_202 = _T_1192 ? _T_3130 : {{33'd0}, _T_461};
  assign _GEN_203 = _T_1192 ? _T_3132 : _GEN_43;
  assign _GEN_204 = _T_1190 ? _T_3134 : reg_hpmevent_5;
  assign _GEN_205 = _T_1198 ? _T_3130 : {{33'd0}, _T_471};
  assign _GEN_206 = _T_1198 ? _T_3132 : _GEN_44;
  assign _GEN_207 = _T_1196 ? _T_3134 : reg_hpmevent_6;
  assign _GEN_208 = _T_1204 ? _T_3130 : {{33'd0}, _T_481};
  assign _GEN_209 = _T_1204 ? _T_3132 : _GEN_45;
  assign _GEN_210 = _T_1202 ? _T_3134 : reg_hpmevent_7;
  assign _GEN_211 = _T_1210 ? _T_3130 : {{33'd0}, _T_491};
  assign _GEN_212 = _T_1210 ? _T_3132 : _GEN_46;
  assign _GEN_213 = _T_1208 ? _T_3134 : reg_hpmevent_8;
  assign _GEN_214 = _T_1216 ? _T_3130 : {{33'd0}, _T_501};
  assign _GEN_215 = _T_1216 ? _T_3132 : _GEN_47;
  assign _GEN_216 = _T_1214 ? _T_3134 : reg_hpmevent_9;
  assign _GEN_217 = _T_1222 ? _T_3130 : {{33'd0}, _T_511};
  assign _GEN_218 = _T_1222 ? _T_3132 : _GEN_48;
  assign _GEN_219 = _T_1220 ? _T_3134 : reg_hpmevent_10;
  assign _GEN_220 = _T_1228 ? _T_3130 : {{33'd0}, _T_521};
  assign _GEN_221 = _T_1228 ? _T_3132 : _GEN_49;
  assign _GEN_222 = _T_1226 ? _T_3134 : reg_hpmevent_11;
  assign _GEN_223 = _T_1234 ? _T_3130 : {{33'd0}, _T_531};
  assign _GEN_224 = _T_1234 ? _T_3132 : _GEN_50;
  assign _GEN_225 = _T_1232 ? _T_3134 : reg_hpmevent_12;
  assign _GEN_226 = _T_1240 ? _T_3130 : {{33'd0}, _T_541};
  assign _GEN_227 = _T_1240 ? _T_3132 : _GEN_51;
  assign _GEN_228 = _T_1238 ? _T_3134 : reg_hpmevent_13;
  assign _GEN_229 = _T_1246 ? _T_3130 : {{33'd0}, _T_551};
  assign _GEN_230 = _T_1246 ? _T_3132 : _GEN_52;
  assign _GEN_231 = _T_1244 ? _T_3134 : reg_hpmevent_14;
  assign _GEN_232 = _T_1252 ? _T_3130 : {{33'd0}, _T_561};
  assign _GEN_233 = _T_1252 ? _T_3132 : _GEN_53;
  assign _GEN_234 = _T_1250 ? _T_3134 : reg_hpmevent_15;
  assign _GEN_235 = _T_1258 ? _T_3130 : {{33'd0}, _T_571};
  assign _GEN_236 = _T_1258 ? _T_3132 : _GEN_54;
  assign _GEN_237 = _T_1256 ? _T_3134 : reg_hpmevent_16;
  assign _GEN_238 = _T_1264 ? _T_3130 : {{33'd0}, _T_581};
  assign _GEN_239 = _T_1264 ? _T_3132 : _GEN_55;
  assign _GEN_240 = _T_1262 ? _T_3134 : reg_hpmevent_17;
  assign _GEN_241 = _T_1270 ? _T_3130 : {{33'd0}, _T_591};
  assign _GEN_242 = _T_1270 ? _T_3132 : _GEN_56;
  assign _GEN_243 = _T_1268 ? _T_3134 : reg_hpmevent_18;
  assign _GEN_244 = _T_1276 ? _T_3130 : {{33'd0}, _T_601};
  assign _GEN_245 = _T_1276 ? _T_3132 : _GEN_57;
  assign _GEN_246 = _T_1274 ? _T_3134 : reg_hpmevent_19;
  assign _GEN_247 = _T_1282 ? _T_3130 : {{33'd0}, _T_611};
  assign _GEN_248 = _T_1282 ? _T_3132 : _GEN_58;
  assign _GEN_249 = _T_1280 ? _T_3134 : reg_hpmevent_20;
  assign _GEN_250 = _T_1288 ? _T_3130 : {{33'd0}, _T_621};
  assign _GEN_251 = _T_1288 ? _T_3132 : _GEN_59;
  assign _GEN_252 = _T_1286 ? _T_3134 : reg_hpmevent_21;
  assign _GEN_253 = _T_1294 ? _T_3130 : {{33'd0}, _T_631};
  assign _GEN_254 = _T_1294 ? _T_3132 : _GEN_60;
  assign _GEN_255 = _T_1292 ? _T_3134 : reg_hpmevent_22;
  assign _GEN_256 = _T_1300 ? _T_3130 : {{33'd0}, _T_641};
  assign _GEN_257 = _T_1300 ? _T_3132 : _GEN_61;
  assign _GEN_258 = _T_1298 ? _T_3134 : reg_hpmevent_23;
  assign _GEN_259 = _T_1306 ? _T_3130 : {{33'd0}, _T_651};
  assign _GEN_260 = _T_1306 ? _T_3132 : _GEN_62;
  assign _GEN_261 = _T_1304 ? _T_3134 : reg_hpmevent_24;
  assign _GEN_262 = _T_1312 ? _T_3130 : {{33'd0}, _T_661};
  assign _GEN_263 = _T_1312 ? _T_3132 : _GEN_63;
  assign _GEN_264 = _T_1310 ? _T_3134 : reg_hpmevent_25;
  assign _GEN_265 = _T_1318 ? _T_3130 : {{33'd0}, _T_671};
  assign _GEN_266 = _T_1318 ? _T_3132 : _GEN_64;
  assign _GEN_267 = _T_1316 ? _T_3134 : reg_hpmevent_26;
  assign _GEN_268 = _T_1324 ? _T_3130 : {{33'd0}, _T_681};
  assign _GEN_269 = _T_1324 ? _T_3132 : _GEN_65;
  assign _GEN_270 = _T_1322 ? _T_3134 : reg_hpmevent_27;
  assign _GEN_271 = _T_1330 ? _T_3130 : {{33'd0}, _T_691};
  assign _GEN_272 = _T_1330 ? _T_3132 : _GEN_66;
  assign _GEN_273 = _T_1328 ? _T_3134 : reg_hpmevent_28;
  assign _T_3248 = wdata[63:6];
  assign _GEN_274 = _T_1156 ? wdata : {{57'd0}, _T_342};
  assign _GEN_275 = _T_1156 ? _T_3248 : _GEN_37;
  assign _GEN_276 = _T_1158 ? wdata : {{57'd0}, _T_329};
  assign _GEN_277 = _T_1158 ? _T_3248 : _GEN_36;
  assign _GEN_278 = _T_1150 ? wdata : {{59'd0}, _GEN_163};
  assign _GEN_279 = _T_1152 ? wdata : {{61'd0}, reg_frm};
  assign _T_3251 = wdata[63:5];
  assign _GEN_280 = _T_1154 ? wdata : _GEN_278;
  assign _GEN_281 = _T_1154 ? {{5'd0}, _T_3251} : _GEN_279;
  assign _T_3257 = _T_3256[1:0];
  assign _T_3258 = _T_3256[2];
  assign _T_3264 = _T_3256[12];
  assign _T_3265 = _T_3256[13];
  assign _T_3267 = _T_3256[15];
  assign _GEN_282 = _T_1144 ? _T_3254_step : reg_dcsr_step;
  assign _GEN_283 = _T_1144 ? _T_3254_ebreakm : reg_dcsr_ebreakm;
  assign _GEN_284 = _T_1144 ? _T_3254_ebreaks : reg_dcsr_ebreaks;
  assign _GEN_285 = _T_1144 ? _T_3254_ebreaku : reg_dcsr_ebreaku;
  assign _GEN_286 = _T_1144 ? _T_3254_prv : _GEN_125;
  assign _T_3273 = _T_3044 | 64'h3;
  assign _T_3274 = ~ _T_3273;
  assign _GEN_287 = _T_1146 ? _T_3274 : {{24'd0}, _GEN_123};
  assign _GEN_288 = _T_1148 ? wdata : reg_dscratch;
  assign _T_3281 = _T_3279[1];
  assign _T_3285 = _T_3279[5];
  assign _T_3288 = _T_3279[8];
  assign _T_3291 = _T_3279[14:13];
  assign _T_3294 = _T_3279[18];
  assign _T_3295 = _T_3279[19];
  assign _T_3310 = _T_3277_fs != 2'h0;
  assign _T_3314 = _T_3310 ? 2'h3 : 2'h0;
  assign _GEN_289 = _T_1340 ? _T_3277_sie : _GEN_172;
  assign _GEN_290 = _T_1340 ? _T_3277_spie : _GEN_171;
  assign _GEN_291 = _T_1340 ? {{1'd0}, _T_3277_spp} : _GEN_170;
  assign _GEN_292 = _T_1340 ? _T_3277_mxr : _GEN_168;
  assign _GEN_293 = _T_1340 ? _T_3277_sum : _GEN_169;
  assign _GEN_294 = _T_1340 ? _T_3314 : _GEN_176;
  assign _T_3327 = _T_3325[1];
  assign _GEN_295 = _T_1342 ? _T_3321_ssip : _GEN_178;
  assign _T_3347 = _T_3346[43:0];
  assign _T_3349 = _T_3346[63:60];
  assign _T_3351 = _T_3344_mode == 4'h0;
  assign _GEN_296 = _T_3351 ? 4'h0 : reg_sptbr_mode;
  assign _T_3354 = _T_3344_mode == 4'h8;
  assign _GEN_297 = _T_3354 ? 4'h8 : _GEN_296;
  assign _T_3360 = _T_3351 | _T_3354;
  assign _T_3361 = _T_3344_ppn[19:0];
  assign _GEN_298 = _T_3360 ? {{24'd0}, _T_3361} : reg_sptbr_ppn;
  assign _GEN_299 = _T_1352 ? _GEN_297 : reg_sptbr_mode;
  assign _GEN_300 = _T_1352 ? _GEN_298 : reg_sptbr_ppn;
  assign _T_3362 = ~ reg_mideleg;
  assign _T_3363 = reg_mie & _T_3362;
  assign _T_3364 = wdata & reg_mideleg;
  assign _T_3365 = _T_3363 | _T_3364;
  assign _GEN_301 = _T_1344 ? _T_3365 : _GEN_181;
  assign _GEN_302 = _T_1346 ? wdata : reg_sscratch;
  assign _GEN_303 = _T_1354 ? _T_3118 : {{24'd0}, _GEN_127};
  assign _GEN_304 = _T_1356 ? _T_3127 : {{25'd0}, reg_stvec};
  assign _T_3384 = wdata & 64'h800000000000001f;
  assign _GEN_305 = _T_1348 ? _T_3384 : _GEN_128;
  assign _GEN_306 = _T_1350 ? _T_3130 : _GEN_129;
  assign _T_3386 = wdata & 64'h222;
  assign _GEN_307 = _T_1360 ? _T_3386 : reg_mideleg;
  assign _T_3387 = wdata & 64'hb109;
  assign _GEN_308 = _T_1362 ? _T_3387 : reg_medeleg;
  assign _T_3389 = wdata & 64'hffffffff;
  assign _GEN_309 = _T_1358 ? _T_3389 : {{32'd0}, reg_scounteren};
  assign _GEN_310 = _T_1334 ? _T_3389 : {{32'd0}, reg_mcounteren};
  assign _T_3394 = _GEN_17_control_dmode == 1'h0;
  assign _T_3395 = _T_3394 | reg_debug;
  assign _T_3401 = _T_3400[0];
  assign _T_3402 = _T_3400[1];
  assign _T_3403 = _T_3400[2];
  assign _T_3404 = _T_3400[3];
  assign _T_3405 = _T_3400[4];
  assign _T_3407 = _T_3400[6];
  assign _T_3408 = _T_3400[8:7];
  assign _T_3411 = _T_3400[12];
  assign _T_3414 = _T_3400[59];
  assign _T_3416 = _T_3398_dmode & reg_debug;
  assign _T_3417 = _T_3416 & _T_3398_action;
  assign _GEN_348 = _T_1114 ? _GEN_33 : reg_bp_0_control_dmode;
  assign _GEN_354 = _T_1114 ? _GEN_34 : reg_bp_0_control_action;
  assign _GEN_360 = _T_1114 ? _GEN_25 : reg_bp_0_control_tmatch;
  assign _GEN_362 = _T_1114 ? _GEN_26 : reg_bp_0_control_m;
  assign _GEN_366 = _T_1114 ? _GEN_28 : reg_bp_0_control_s;
  assign _GEN_368 = _T_1114 ? _GEN_29 : reg_bp_0_control_u;
  assign _GEN_370 = _T_1114 ? _GEN_30 : reg_bp_0_control_x;
  assign _GEN_372 = _T_1114 ? _GEN_31 : reg_bp_0_control_w;
  assign _GEN_374 = _T_1114 ? _GEN_32 : reg_bp_0_control_r;
  assign _GEN_378 = _T_1116 ? _GEN_35 : reg_bp_0_address;
  assign _GEN_382 = _T_3395 ? _GEN_348 : reg_bp_0_control_dmode;
  assign _GEN_388 = _T_3395 ? _GEN_354 : reg_bp_0_control_action;
  assign _GEN_394 = _T_3395 ? _GEN_360 : reg_bp_0_control_tmatch;
  assign _GEN_396 = _T_3395 ? _GEN_362 : reg_bp_0_control_m;
  assign _GEN_400 = _T_3395 ? _GEN_366 : reg_bp_0_control_s;
  assign _GEN_402 = _T_3395 ? _GEN_368 : reg_bp_0_control_u;
  assign _GEN_404 = _T_3395 ? _GEN_370 : reg_bp_0_control_x;
  assign _GEN_406 = _T_3395 ? _GEN_372 : reg_bp_0_control_w;
  assign _GEN_408 = _T_3395 ? _GEN_374 : reg_bp_0_control_r;
  assign _GEN_410 = _T_3395 ? _GEN_378 : reg_bp_0_address;
  assign _GEN_412 = _T_3001 ? _GEN_164 : _GEN_160;
  assign _GEN_413 = _T_3001 ? _GEN_165 : _GEN_161;
  assign _GEN_414 = _T_3001 ? _GEN_166 : reg_mstatus_mprv;
  assign _GEN_415 = _T_3001 ? _GEN_167 : _GEN_162;
  assign _GEN_416 = _T_3001 ? _GEN_292 : reg_mstatus_mxr;
  assign _GEN_417 = _T_3001 ? _GEN_293 : reg_mstatus_sum;
  assign _GEN_418 = _T_3001 ? _GEN_291 : _GEN_156;
  assign _GEN_419 = _T_3001 ? _GEN_290 : _GEN_155;
  assign _GEN_420 = _T_3001 ? _GEN_289 : _GEN_154;
  assign _GEN_421 = _T_3001 ? _GEN_173 : reg_mstatus_tw;
  assign _GEN_422 = _T_3001 ? _GEN_174 : reg_mstatus_tvm;
  assign _GEN_423 = _T_3001 ? _GEN_175 : reg_mstatus_tsr;
  assign _GEN_424 = _T_3001 ? _GEN_294 : reg_mstatus_fs;
  assign _GEN_425 = _T_3001 ? _GEN_177 : reg_misa;
  assign _GEN_426 = _T_3001 ? _GEN_295 : reg_mip_ssip;
  assign _GEN_427 = _T_3001 ? _GEN_179 : reg_mip_stip;
  assign _GEN_428 = _T_3001 ? _GEN_180 : reg_mip_seip;
  assign _GEN_429 = _T_3001 ? _GEN_301 : reg_mie;
  assign _GEN_430 = _T_3001 ? _GEN_182 : {{24'd0}, _GEN_133};
  assign _GEN_431 = _T_3001 ? _GEN_183 : reg_mscratch;
  assign _GEN_432 = _T_3001 ? _GEN_184 : {{32'd0}, reg_mtvec};
  assign _GEN_433 = _T_3001 ? _GEN_185 : _GEN_134;
  assign _GEN_434 = _T_3001 ? _GEN_186 : _GEN_135;
  assign _GEN_435 = _T_3001 ? _GEN_187 : {{33'd0}, _T_411};
  assign _GEN_436 = _T_3001 ? _GEN_188 : _GEN_38;
  assign _GEN_437 = _T_3001 ? _GEN_189 : reg_hpmevent_0;
  assign _GEN_438 = _T_3001 ? _GEN_190 : {{33'd0}, _T_421};
  assign _GEN_439 = _T_3001 ? _GEN_191 : _GEN_39;
  assign _GEN_440 = _T_3001 ? _GEN_192 : reg_hpmevent_1;
  assign _GEN_441 = _T_3001 ? _GEN_193 : {{33'd0}, _T_431};
  assign _GEN_442 = _T_3001 ? _GEN_194 : _GEN_40;
  assign _GEN_443 = _T_3001 ? _GEN_195 : reg_hpmevent_2;
  assign _GEN_444 = _T_3001 ? _GEN_196 : {{33'd0}, _T_441};
  assign _GEN_445 = _T_3001 ? _GEN_197 : _GEN_41;
  assign _GEN_446 = _T_3001 ? _GEN_198 : reg_hpmevent_3;
  assign _GEN_447 = _T_3001 ? _GEN_199 : {{33'd0}, _T_451};
  assign _GEN_448 = _T_3001 ? _GEN_200 : _GEN_42;
  assign _GEN_449 = _T_3001 ? _GEN_201 : reg_hpmevent_4;
  assign _GEN_450 = _T_3001 ? _GEN_202 : {{33'd0}, _T_461};
  assign _GEN_451 = _T_3001 ? _GEN_203 : _GEN_43;
  assign _GEN_452 = _T_3001 ? _GEN_204 : reg_hpmevent_5;
  assign _GEN_453 = _T_3001 ? _GEN_205 : {{33'd0}, _T_471};
  assign _GEN_454 = _T_3001 ? _GEN_206 : _GEN_44;
  assign _GEN_455 = _T_3001 ? _GEN_207 : reg_hpmevent_6;
  assign _GEN_456 = _T_3001 ? _GEN_208 : {{33'd0}, _T_481};
  assign _GEN_457 = _T_3001 ? _GEN_209 : _GEN_45;
  assign _GEN_458 = _T_3001 ? _GEN_210 : reg_hpmevent_7;
  assign _GEN_459 = _T_3001 ? _GEN_211 : {{33'd0}, _T_491};
  assign _GEN_460 = _T_3001 ? _GEN_212 : _GEN_46;
  assign _GEN_461 = _T_3001 ? _GEN_213 : reg_hpmevent_8;
  assign _GEN_462 = _T_3001 ? _GEN_214 : {{33'd0}, _T_501};
  assign _GEN_463 = _T_3001 ? _GEN_215 : _GEN_47;
  assign _GEN_464 = _T_3001 ? _GEN_216 : reg_hpmevent_9;
  assign _GEN_465 = _T_3001 ? _GEN_217 : {{33'd0}, _T_511};
  assign _GEN_466 = _T_3001 ? _GEN_218 : _GEN_48;
  assign _GEN_467 = _T_3001 ? _GEN_219 : reg_hpmevent_10;
  assign _GEN_468 = _T_3001 ? _GEN_220 : {{33'd0}, _T_521};
  assign _GEN_469 = _T_3001 ? _GEN_221 : _GEN_49;
  assign _GEN_470 = _T_3001 ? _GEN_222 : reg_hpmevent_11;
  assign _GEN_471 = _T_3001 ? _GEN_223 : {{33'd0}, _T_531};
  assign _GEN_472 = _T_3001 ? _GEN_224 : _GEN_50;
  assign _GEN_473 = _T_3001 ? _GEN_225 : reg_hpmevent_12;
  assign _GEN_474 = _T_3001 ? _GEN_226 : {{33'd0}, _T_541};
  assign _GEN_475 = _T_3001 ? _GEN_227 : _GEN_51;
  assign _GEN_476 = _T_3001 ? _GEN_228 : reg_hpmevent_13;
  assign _GEN_477 = _T_3001 ? _GEN_229 : {{33'd0}, _T_551};
  assign _GEN_478 = _T_3001 ? _GEN_230 : _GEN_52;
  assign _GEN_479 = _T_3001 ? _GEN_231 : reg_hpmevent_14;
  assign _GEN_480 = _T_3001 ? _GEN_232 : {{33'd0}, _T_561};
  assign _GEN_481 = _T_3001 ? _GEN_233 : _GEN_53;
  assign _GEN_482 = _T_3001 ? _GEN_234 : reg_hpmevent_15;
  assign _GEN_483 = _T_3001 ? _GEN_235 : {{33'd0}, _T_571};
  assign _GEN_484 = _T_3001 ? _GEN_236 : _GEN_54;
  assign _GEN_485 = _T_3001 ? _GEN_237 : reg_hpmevent_16;
  assign _GEN_486 = _T_3001 ? _GEN_238 : {{33'd0}, _T_581};
  assign _GEN_487 = _T_3001 ? _GEN_239 : _GEN_55;
  assign _GEN_488 = _T_3001 ? _GEN_240 : reg_hpmevent_17;
  assign _GEN_489 = _T_3001 ? _GEN_241 : {{33'd0}, _T_591};
  assign _GEN_490 = _T_3001 ? _GEN_242 : _GEN_56;
  assign _GEN_491 = _T_3001 ? _GEN_243 : reg_hpmevent_18;
  assign _GEN_492 = _T_3001 ? _GEN_244 : {{33'd0}, _T_601};
  assign _GEN_493 = _T_3001 ? _GEN_245 : _GEN_57;
  assign _GEN_494 = _T_3001 ? _GEN_246 : reg_hpmevent_19;
  assign _GEN_495 = _T_3001 ? _GEN_247 : {{33'd0}, _T_611};
  assign _GEN_496 = _T_3001 ? _GEN_248 : _GEN_58;
  assign _GEN_497 = _T_3001 ? _GEN_249 : reg_hpmevent_20;
  assign _GEN_498 = _T_3001 ? _GEN_250 : {{33'd0}, _T_621};
  assign _GEN_499 = _T_3001 ? _GEN_251 : _GEN_59;
  assign _GEN_500 = _T_3001 ? _GEN_252 : reg_hpmevent_21;
  assign _GEN_501 = _T_3001 ? _GEN_253 : {{33'd0}, _T_631};
  assign _GEN_502 = _T_3001 ? _GEN_254 : _GEN_60;
  assign _GEN_503 = _T_3001 ? _GEN_255 : reg_hpmevent_22;
  assign _GEN_504 = _T_3001 ? _GEN_256 : {{33'd0}, _T_641};
  assign _GEN_505 = _T_3001 ? _GEN_257 : _GEN_61;
  assign _GEN_506 = _T_3001 ? _GEN_258 : reg_hpmevent_23;
  assign _GEN_507 = _T_3001 ? _GEN_259 : {{33'd0}, _T_651};
  assign _GEN_508 = _T_3001 ? _GEN_260 : _GEN_62;
  assign _GEN_509 = _T_3001 ? _GEN_261 : reg_hpmevent_24;
  assign _GEN_510 = _T_3001 ? _GEN_262 : {{33'd0}, _T_661};
  assign _GEN_511 = _T_3001 ? _GEN_263 : _GEN_63;
  assign _GEN_512 = _T_3001 ? _GEN_264 : reg_hpmevent_25;
  assign _GEN_513 = _T_3001 ? _GEN_265 : {{33'd0}, _T_671};
  assign _GEN_514 = _T_3001 ? _GEN_266 : _GEN_64;
  assign _GEN_515 = _T_3001 ? _GEN_267 : reg_hpmevent_26;
  assign _GEN_516 = _T_3001 ? _GEN_268 : {{33'd0}, _T_681};
  assign _GEN_517 = _T_3001 ? _GEN_269 : _GEN_65;
  assign _GEN_518 = _T_3001 ? _GEN_270 : reg_hpmevent_27;
  assign _GEN_519 = _T_3001 ? _GEN_271 : {{33'd0}, _T_691};
  assign _GEN_520 = _T_3001 ? _GEN_272 : _GEN_66;
  assign _GEN_521 = _T_3001 ? _GEN_273 : reg_hpmevent_28;
  assign _GEN_522 = _T_3001 ? _GEN_274 : {{57'd0}, _T_342};
  assign _GEN_523 = _T_3001 ? _GEN_275 : _GEN_37;
  assign _GEN_524 = _T_3001 ? _GEN_276 : {{57'd0}, _T_329};
  assign _GEN_525 = _T_3001 ? _GEN_277 : _GEN_36;
  assign _GEN_526 = _T_3001 ? _GEN_280 : {{59'd0}, _GEN_163};
  assign _GEN_527 = _T_3001 ? _GEN_281 : {{61'd0}, reg_frm};
  assign _GEN_528 = _T_3001 ? _GEN_282 : reg_dcsr_step;
  assign _GEN_529 = _T_3001 ? _GEN_283 : reg_dcsr_ebreakm;
  assign _GEN_530 = _T_3001 ? _GEN_284 : reg_dcsr_ebreaks;
  assign _GEN_531 = _T_3001 ? _GEN_285 : reg_dcsr_ebreaku;
  assign _GEN_532 = _T_3001 ? _GEN_286 : _GEN_125;
  assign _GEN_533 = _T_3001 ? _GEN_287 : {{24'd0}, _GEN_123};
  assign _GEN_534 = _T_3001 ? _GEN_288 : reg_dscratch;
  assign _GEN_535 = _T_3001 ? _GEN_299 : reg_sptbr_mode;
  assign _GEN_536 = _T_3001 ? _GEN_300 : reg_sptbr_ppn;
  assign _GEN_537 = _T_3001 ? _GEN_302 : reg_sscratch;
  assign _GEN_538 = _T_3001 ? _GEN_303 : {{24'd0}, _GEN_127};
  assign _GEN_539 = _T_3001 ? _GEN_304 : {{25'd0}, reg_stvec};
  assign _GEN_540 = _T_3001 ? _GEN_305 : _GEN_128;
  assign _GEN_541 = _T_3001 ? _GEN_306 : _GEN_129;
  assign _GEN_542 = _T_3001 ? _GEN_307 : reg_mideleg;
  assign _GEN_543 = _T_3001 ? _GEN_308 : reg_medeleg;
  assign _GEN_544 = _T_3001 ? _GEN_309 : {{32'd0}, reg_scounteren};
  assign _GEN_545 = _T_3001 ? _GEN_310 : {{32'd0}, reg_mcounteren};
  assign _GEN_549 = _T_3001 ? _GEN_382 : reg_bp_0_control_dmode;
  assign _GEN_555 = _T_3001 ? _GEN_388 : reg_bp_0_control_action;
  assign _GEN_561 = _T_3001 ? _GEN_394 : reg_bp_0_control_tmatch;
  assign _GEN_563 = _T_3001 ? _GEN_396 : reg_bp_0_control_m;
  assign _GEN_567 = _T_3001 ? _GEN_400 : reg_bp_0_control_s;
  assign _GEN_569 = _T_3001 ? _GEN_402 : reg_bp_0_control_u;
  assign _GEN_571 = _T_3001 ? _GEN_404 : reg_bp_0_control_x;
  assign _GEN_573 = _T_3001 ? _GEN_406 : reg_bp_0_control_w;
  assign _GEN_575 = _T_3001 ? _GEN_408 : reg_bp_0_control_r;
  assign _GEN_577 = _T_3001 ? _GEN_410 : reg_bp_0_address;
  assign _GEN_579 = reset ? 1'h0 : _GEN_555;
  assign _GEN_580 = reset ? 1'h0 : _GEN_549;
  assign _GEN_581 = reset ? 1'h0 : _GEN_575;
  assign _GEN_582 = reset ? 1'h0 : _GEN_573;
  assign _GEN_583 = reset ? 1'h0 : _GEN_571;
  assign io_rw_rdata = _T_2992;
  assign io_decode_0_fp_illegal = _T_1409;
  assign io_decode_0_read_illegal = _T_1848;
  assign io_decode_0_write_illegal = _T_1852;
  assign io_decode_0_write_flush = _T_1865;
  assign io_decode_0_system_illegal = _T_1890;
  assign io_decode_1_fp_illegal = _T_1409;
  assign io_decode_1_read_illegal = _T_2356;
  assign io_decode_1_write_illegal = _T_2360;
  assign io_decode_1_write_flush = _T_2373;
  assign io_decode_1_system_illegal = _T_2398;
  assign io_csr_stall = reg_wfi;
  assign io_eret = _T_2458;
  assign io_singleStep = _T_2461;
  assign io_status_debug = reg_debug;
  assign io_status_isa = reg_misa[31:0];
  assign io_status_dprv = _T_2476;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = _T_2468;
  assign io_status_zero2 = 27'h0;
  assign io_status_sxl = 2'h2;
  assign io_status_uxl = 2'h2;
  assign io_status_sd_rv32 = 1'h0;
  assign io_status_zero1 = 8'h0;
  assign io_status_tsr = reg_mstatus_tsr;
  assign io_status_tw = reg_mstatus_tw;
  assign io_status_tvm = reg_mstatus_tvm;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_sum = reg_mstatus_sum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = 2'h0;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = 2'h0;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = 1'h0;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = 1'h0;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = 1'h0;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = 1'h0;
  assign io_ptbr_mode = reg_sptbr_mode;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = _GEN_158;
  assign io_fcsr_rm = reg_frm;
  assign io_interrupt = _T_938;
  assign io_interrupt_cause = interruptCause;
  assign io_counters_0_eventSel = reg_hpmevent_0;
  assign io_counters_1_eventSel = reg_hpmevent_1;
  assign io_counters_2_eventSel = reg_hpmevent_2;
  assign io_counters_3_eventSel = reg_hpmevent_3;
  assign io_counters_4_eventSel = reg_hpmevent_4;
  assign io_counters_5_eventSel = reg_hpmevent_5;
  assign io_counters_6_eventSel = reg_hpmevent_6;
  assign io_counters_7_eventSel = reg_hpmevent_7;
  assign io_counters_8_eventSel = reg_hpmevent_8;
  assign io_counters_9_eventSel = reg_hpmevent_9;
  assign io_counters_10_eventSel = reg_hpmevent_10;
  assign io_counters_11_eventSel = reg_hpmevent_11;
  assign io_counters_12_eventSel = reg_hpmevent_12;
  assign io_counters_13_eventSel = reg_hpmevent_13;
  assign io_counters_14_eventSel = reg_hpmevent_14;
  assign io_counters_15_eventSel = reg_hpmevent_15;
  assign io_counters_16_eventSel = reg_hpmevent_16;
  assign io_counters_17_eventSel = reg_hpmevent_17;
  assign io_counters_18_eventSel = reg_hpmevent_18;
  assign io_counters_19_eventSel = reg_hpmevent_19;
  assign io_counters_20_eventSel = reg_hpmevent_20;
  assign io_counters_21_eventSel = reg_hpmevent_21;
  assign io_counters_22_eventSel = reg_hpmevent_22;
  assign io_counters_23_eventSel = reg_hpmevent_23;
  assign io_counters_24_eventSel = reg_hpmevent_24;
  assign io_counters_25_eventSel = reg_hpmevent_25;
  assign io_counters_26_eventSel = reg_hpmevent_26;
  assign io_counters_27_eventSel = reg_hpmevent_27;
  assign io_counters_28_eventSel = reg_hpmevent_28;
  assign new_prv = _GEN_157;
  assign mip_meip = io_interrupts_meip;
  assign mip_seip = _T_712;
  assign mip_mtip = io_interrupts_mtip;
  assign mip_stip = reg_mip_stip;
  assign mip_msip = io_interrupts_msip;
  assign mip_ssip = reg_mip_ssip;
  assign _GEN_0_control_x = reg_bp_0_control_x;
  assign _GEN_1_control_w = reg_bp_0_control_w;
  assign _GEN_2_control_r = reg_bp_0_control_r;
  assign _GEN_3_control_s = reg_bp_0_control_s;
  assign _GEN_4_control_u = reg_bp_0_control_u;
  assign _GEN_5_control_m = reg_bp_0_control_m;
  assign _GEN_8_control_tmatch = reg_bp_0_control_tmatch;
  assign _GEN_9_control_action = reg_bp_0_control_action;
  assign _GEN_14_control_dmode = reg_bp_0_control_dmode;
  assign _GEN_15_address = reg_bp_0_address;
  assign _GEN_16_address = reg_bp_0_address;
  assign _T_1060_sd = io_status_sd;
  assign _T_1060_uxl = io_status_uxl;
  assign _T_1060_sd_rv32 = io_status_sd_rv32;
  assign _T_1060_mxr = io_status_mxr;
  assign _T_1060_sum = io_status_sum;
  assign _T_1060_xs = io_status_xs;
  assign _T_1060_fs = io_status_fs;
  assign _T_1060_spp = io_status_spp;
  assign _T_1060_spie = io_status_spie;
  assign _T_1060_sie = io_status_sie;
  assign _T_2992 = _T_2990;
  assign _T_3004_tsr = _T_3025;
  assign _T_3004_tw = _T_3024;
  assign _T_3004_tvm = _T_3023;
  assign _T_3004_mxr = _T_3022;
  assign _T_3004_sum = _T_3021;
  assign _T_3004_mprv = _T_3020;
  assign _T_3004_fs = _T_3018;
  assign _T_3004_mpp = _T_3017;
  assign _T_3004_spp = _T_3015;
  assign _T_3004_mpie = _T_3014;
  assign _T_3004_spie = _T_3012;
  assign _T_3004_mie = _T_3010;
  assign _T_3004_sie = _T_3008;
  assign _T_3006 = {{37'd0}, wdata};
  assign _T_3089_seip = _T_3103;
  assign _T_3089_stip = _T_3099;
  assign _T_3089_ssip = _T_3095;
  assign _T_3093 = _T_3082[15:0];
  assign _T_3254_ebreakm = _T_3267;
  assign _T_3254_ebreaks = _T_3265;
  assign _T_3254_ebreaku = _T_3264;
  assign _T_3254_step = _T_3258;
  assign _T_3254_prv = _T_3257;
  assign _T_3256 = wdata[31:0];
  assign _T_3277_mxr = _T_3295;
  assign _T_3277_sum = _T_3294;
  assign _T_3277_fs = _T_3291;
  assign _T_3277_spp = _T_3288;
  assign _T_3277_spie = _T_3285;
  assign _T_3277_sie = _T_3281;
  assign _T_3279 = {{37'd0}, wdata};
  assign _T_3321_ssip = _T_3327;
  assign _T_3325 = wdata[15:0];
  assign _T_3344_mode = _T_3349;
  assign _T_3344_ppn = _T_3347;
  assign _T_3346 = wdata;
  assign _GEN_17_control_dmode = reg_bp_0_control_dmode;
  assign _T_3398_dmode = _T_3414;
  assign _T_3398_action = _T_3411;
  assign _T_3398_tmatch = _T_3408;
  assign _T_3398_m = _T_3407;
  assign _T_3398_s = _T_3405;
  assign _T_3398_u = _T_3404;
  assign _T_3398_x = _T_3403;
  assign _T_3398_w = _T_3402;
  assign _T_3398_r = _T_3401;
  assign _T_3400 = wdata;
  assign _GEN_25 = _T_3398_tmatch;
  assign _GEN_26 = _T_3398_m;
  assign _GEN_28 = _T_3398_s;
  assign _GEN_29 = _T_3398_u;
  assign _GEN_30 = _T_3398_x;
  assign _GEN_31 = _T_3398_w;
  assign _GEN_32 = _T_3398_r;
  assign _GEN_33 = _T_3416;
  assign _GEN_34 = _T_3417;
  assign _GEN_35 = wdata[38:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_mstatus_tsr = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_mstatus_tw = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_mstatus_tvm = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_mstatus_mxr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_mstatus_sum = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_mstatus_mprv = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_mstatus_fs = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_mstatus_mpp = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_mstatus_spp = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_mstatus_mpie = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  reg_mstatus_spie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  reg_mstatus_mie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  reg_mstatus_sie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  reg_dcsr_ebreakm = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  reg_dcsr_ebreaks = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  reg_dcsr_ebreaku = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  reg_dcsr_cause = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  reg_dcsr_step = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  reg_dcsr_prv = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  reg_debug = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{$random}};
  reg_dpc = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{$random}};
  reg_dscratch = _RAND_22[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  reg_singleStepped = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  reg_bp_0_control_dmode = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  reg_bp_0_control_action = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  reg_bp_0_control_tmatch = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  reg_bp_0_control_m = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  reg_bp_0_control_s = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  reg_bp_0_control_u = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  reg_bp_0_control_x = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  reg_bp_0_control_w = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  reg_bp_0_control_r = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{$random}};
  reg_bp_0_address = _RAND_33[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{$random}};
  reg_mie = _RAND_34[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{$random}};
  reg_mideleg = _RAND_35[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{$random}};
  reg_medeleg = _RAND_36[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  reg_mip_seip = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  reg_mip_stip = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  reg_mip_ssip = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{$random}};
  reg_mepc = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{$random}};
  reg_mcause = _RAND_41[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{$random}};
  reg_mbadaddr = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{$random}};
  reg_mscratch = _RAND_43[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  reg_mtvec = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  reg_mcounteren = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  reg_scounteren = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{$random}};
  reg_sepc = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{$random}};
  reg_scause = _RAND_48[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{$random}};
  reg_sbadaddr = _RAND_49[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{$random}};
  reg_sscratch = _RAND_50[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{$random}};
  reg_stvec = _RAND_51[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  reg_sptbr_mode = _RAND_52[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{$random}};
  reg_sptbr_ppn = _RAND_53[43:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  reg_wfi = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  reg_fflags = _RAND_55[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  reg_frm = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_328 = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{$random}};
  _T_332 = _RAND_58[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_341 = _RAND_59[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{$random}};
  _T_345 = _RAND_60[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{$random}};
  reg_hpmevent_0 = _RAND_61[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{$random}};
  reg_hpmevent_1 = _RAND_62[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{$random}};
  reg_hpmevent_2 = _RAND_63[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{$random}};
  reg_hpmevent_3 = _RAND_64[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{$random}};
  reg_hpmevent_4 = _RAND_65[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{$random}};
  reg_hpmevent_5 = _RAND_66[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{$random}};
  reg_hpmevent_6 = _RAND_67[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {2{$random}};
  reg_hpmevent_7 = _RAND_68[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{$random}};
  reg_hpmevent_8 = _RAND_69[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{$random}};
  reg_hpmevent_9 = _RAND_70[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {2{$random}};
  reg_hpmevent_10 = _RAND_71[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {2{$random}};
  reg_hpmevent_11 = _RAND_72[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{$random}};
  reg_hpmevent_12 = _RAND_73[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{$random}};
  reg_hpmevent_13 = _RAND_74[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {2{$random}};
  reg_hpmevent_14 = _RAND_75[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{$random}};
  reg_hpmevent_15 = _RAND_76[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{$random}};
  reg_hpmevent_16 = _RAND_77[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{$random}};
  reg_hpmevent_17 = _RAND_78[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{$random}};
  reg_hpmevent_18 = _RAND_79[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {2{$random}};
  reg_hpmevent_19 = _RAND_80[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {2{$random}};
  reg_hpmevent_20 = _RAND_81[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{$random}};
  reg_hpmevent_21 = _RAND_82[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {2{$random}};
  reg_hpmevent_22 = _RAND_83[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{$random}};
  reg_hpmevent_23 = _RAND_84[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {2{$random}};
  reg_hpmevent_24 = _RAND_85[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{$random}};
  reg_hpmevent_25 = _RAND_86[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{$random}};
  reg_hpmevent_26 = _RAND_87[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{$random}};
  reg_hpmevent_27 = _RAND_88[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{$random}};
  reg_hpmevent_28 = _RAND_89[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_410 = _RAND_90[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{$random}};
  _T_413 = _RAND_91[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_420 = _RAND_92[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {2{$random}};
  _T_423 = _RAND_93[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_430 = _RAND_94[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {2{$random}};
  _T_433 = _RAND_95[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_440 = _RAND_96[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{$random}};
  _T_443 = _RAND_97[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_450 = _RAND_98[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{$random}};
  _T_453 = _RAND_99[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_460 = _RAND_100[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {2{$random}};
  _T_463 = _RAND_101[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_470 = _RAND_102[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {2{$random}};
  _T_473 = _RAND_103[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_480 = _RAND_104[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {2{$random}};
  _T_483 = _RAND_105[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_490 = _RAND_106[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {2{$random}};
  _T_493 = _RAND_107[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_500 = _RAND_108[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {2{$random}};
  _T_503 = _RAND_109[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_510 = _RAND_110[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {2{$random}};
  _T_513 = _RAND_111[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_520 = _RAND_112[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {2{$random}};
  _T_523 = _RAND_113[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_530 = _RAND_114[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {2{$random}};
  _T_533 = _RAND_115[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_540 = _RAND_116[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {2{$random}};
  _T_543 = _RAND_117[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_550 = _RAND_118[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {2{$random}};
  _T_553 = _RAND_119[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_560 = _RAND_120[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {2{$random}};
  _T_563 = _RAND_121[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_570 = _RAND_122[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {2{$random}};
  _T_573 = _RAND_123[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_580 = _RAND_124[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {2{$random}};
  _T_583 = _RAND_125[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_590 = _RAND_126[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {2{$random}};
  _T_593 = _RAND_127[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_600 = _RAND_128[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {2{$random}};
  _T_603 = _RAND_129[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_610 = _RAND_130[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {2{$random}};
  _T_613 = _RAND_131[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_620 = _RAND_132[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {2{$random}};
  _T_623 = _RAND_133[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_630 = _RAND_134[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {2{$random}};
  _T_633 = _RAND_135[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_640 = _RAND_136[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {2{$random}};
  _T_643 = _RAND_137[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_650 = _RAND_138[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {2{$random}};
  _T_653 = _RAND_139[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_660 = _RAND_140[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {2{$random}};
  _T_663 = _RAND_141[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_670 = _RAND_142[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {2{$random}};
  _T_673 = _RAND_143[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_680 = _RAND_144[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {2{$random}};
  _T_683 = _RAND_145[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_690 = _RAND_146[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {2{$random}};
  _T_693 = _RAND_147[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_711 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {2{$random}};
  reg_misa = _RAND_149[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_2476 = _RAND_150[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_194) begin
        reg_mstatus_prv <= 2'h0;
      end else begin
        reg_mstatus_prv <= new_prv;
      end
    end
    if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_tsr <= _T_3004_tsr;
        end
      end
    end
    if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_tw <= _T_3004_tw;
        end
      end
    end
    if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_tvm <= _T_3004_tvm;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1340) begin
          reg_mstatus_mxr <= _T_3277_mxr;
        end else begin
          if (_T_1126) begin
            reg_mstatus_mxr <= _T_3004_mxr;
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1340) begin
          reg_mstatus_sum <= _T_3277_sum;
        end else begin
          if (_T_1126) begin
            reg_mstatus_sum <= _T_3004_sum;
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_mprv <= _T_3004_mprv;
        end
      end
    end
    if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1340) begin
          if (_T_3310) begin
            reg_mstatus_fs <= 2'h3;
          end else begin
            reg_mstatus_fs <= 2'h0;
          end
        end else begin
          if (_T_1126) begin
            if (_T_3037) begin
              reg_mstatus_fs <= 2'h3;
            end else begin
              reg_mstatus_fs <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_mpp <= _T_3004_mpp;
        end else begin
          if (insn_ret) begin
            if (_T_2599) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (!(delegate)) begin
                    reg_mstatus_mpp <= reg_mstatus_prv;
                  end
                end
              end
            end else begin
              if (_T_2604) begin
                if (exception) begin
                  if (!(trapToDebug)) begin
                    if (!(delegate)) begin
                      reg_mstatus_mpp <= reg_mstatus_prv;
                    end
                  end
                end
              end else begin
                reg_mstatus_mpp <= 2'h0;
              end
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mpp <= reg_mstatus_prv;
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2599) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mpp <= reg_mstatus_prv;
                end
              end
            end
          end else begin
            if (_T_2604) begin
              reg_mstatus_mpp <= _GEN_137;
            end else begin
              reg_mstatus_mpp <= 2'h0;
            end
          end
        end else begin
          reg_mstatus_mpp <= _GEN_137;
        end
      end
    end
    if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_418[0];
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_mpie <= _T_3004_mpie;
        end else begin
          if (insn_ret) begin
            if (_T_2599) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (!(delegate)) begin
                    reg_mstatus_mpie <= reg_mstatus_mie;
                  end
                end
              end
            end else begin
              if (_T_2604) begin
                if (exception) begin
                  if (!(trapToDebug)) begin
                    if (!(delegate)) begin
                      reg_mstatus_mpie <= reg_mstatus_mie;
                    end
                  end
                end
              end else begin
                reg_mstatus_mpie <= 1'h1;
              end
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mpie <= reg_mstatus_mie;
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2599) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mpie <= reg_mstatus_mie;
                end
              end
            end
          end else begin
            if (_T_2604) begin
              reg_mstatus_mpie <= _GEN_136;
            end else begin
              reg_mstatus_mpie <= 1'h1;
            end
          end
        end else begin
          reg_mstatus_mpie <= _GEN_136;
        end
      end
    end
    if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1340) begin
          reg_mstatus_spie <= _T_3277_spie;
        end else begin
          if (_T_1126) begin
            reg_mstatus_spie <= _T_3004_spie;
          end else begin
            if (insn_ret) begin
              if (_T_2599) begin
                reg_mstatus_spie <= 1'h1;
              end else begin
                if (exception) begin
                  if (!(trapToDebug)) begin
                    if (delegate) begin
                      reg_mstatus_spie <= reg_mstatus_sie;
                    end
                  end
                end
              end
            end else begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (delegate) begin
                    reg_mstatus_spie <= reg_mstatus_sie;
                  end
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2599) begin
            reg_mstatus_spie <= 1'h1;
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (delegate) begin
                  reg_mstatus_spie <= reg_mstatus_sie;
                end
              end
            end
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (delegate) begin
                reg_mstatus_spie <= reg_mstatus_sie;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1126) begin
          reg_mstatus_mie <= _T_3004_mie;
        end else begin
          if (insn_ret) begin
            if (_T_2599) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (!(delegate)) begin
                    reg_mstatus_mie <= 1'h0;
                  end
                end
              end
            end else begin
              if (_T_2604) begin
                if (exception) begin
                  if (!(trapToDebug)) begin
                    if (!(delegate)) begin
                      reg_mstatus_mie <= 1'h0;
                    end
                  end
                end
              end else begin
                reg_mstatus_mie <= reg_mstatus_mpie;
              end
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2599) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (!(delegate)) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if (_T_2604) begin
              reg_mstatus_mie <= _GEN_138;
            end else begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end
          end
        end else begin
          reg_mstatus_mie <= _GEN_138;
        end
      end
    end
    if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1340) begin
          reg_mstatus_sie <= _T_3277_sie;
        end else begin
          if (_T_1126) begin
            reg_mstatus_sie <= _T_3004_sie;
          end else begin
            if (insn_ret) begin
              if (_T_2599) begin
                reg_mstatus_sie <= reg_mstatus_spie;
              end else begin
                if (exception) begin
                  if (!(trapToDebug)) begin
                    if (delegate) begin
                      reg_mstatus_sie <= 1'h0;
                    end
                  end
                end
              end
            end else begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  if (delegate) begin
                    reg_mstatus_sie <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2599) begin
            reg_mstatus_sie <= reg_mstatus_spie;
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                if (delegate) begin
                  reg_mstatus_sie <= 1'h0;
                end
              end
            end
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (delegate) begin
                reg_mstatus_sie <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1144) begin
          reg_dcsr_ebreakm <= _T_3254_ebreakm;
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1144) begin
          reg_dcsr_ebreaks <= _T_3254_ebreaks;
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1144) begin
          reg_dcsr_ebreaku <= _T_3254_ebreaku;
        end
      end
    end
    if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else begin
      if (exception) begin
        if (trapToDebug) begin
          if (_T_933) begin
            if (reg_singleStepped) begin
              reg_dcsr_cause <= 3'h4;
            end else begin
              reg_dcsr_cause <= {{1'd0}, _T_2573};
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1144) begin
          reg_dcsr_step <= _T_3254_step;
        end
      end
    end
    if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else begin
      if (_T_3001) begin
        if (_T_1144) begin
          reg_dcsr_prv <= _T_3254_prv;
        end else begin
          if (exception) begin
            if (trapToDebug) begin
              if (_T_933) begin
                reg_dcsr_prv <= reg_mstatus_prv;
              end
            end
          end
        end
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_933) begin
              reg_dcsr_prv <= reg_mstatus_prv;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_debug <= 1'h0;
    end else begin
      if (insn_ret) begin
        if (_T_2599) begin
          if (exception) begin
            if (trapToDebug) begin
              if (_T_933) begin
                reg_debug <= 1'h1;
              end
            end
          end
        end else begin
          if (_T_2604) begin
            reg_debug <= 1'h0;
          end else begin
            if (exception) begin
              if (trapToDebug) begin
                if (_T_933) begin
                  reg_debug <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_933) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end
    end
    reg_dpc <= _GEN_533[39:0];
    if (_T_3001) begin
      if (_T_1148) begin
        reg_dscratch <= wdata;
      end
    end
    if (_T_936) begin
      reg_singleStepped <= 1'h0;
    end else begin
      if (_T_2509) begin
        reg_singleStepped <= 1'h1;
      end
    end
    if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_3395) begin
          if (_T_1114) begin
            reg_bp_0_control_dmode <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_3395) begin
          if (_T_1114) begin
            reg_bp_0_control_action <= _GEN_34;
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_3395) begin
        if (_T_1114) begin
          reg_bp_0_control_tmatch <= _GEN_25;
        end
      end
    end
    if (_T_3001) begin
      if (_T_3395) begin
        if (_T_1114) begin
          reg_bp_0_control_m <= _GEN_26;
        end
      end
    end
    if (_T_3001) begin
      if (_T_3395) begin
        if (_T_1114) begin
          reg_bp_0_control_s <= _GEN_28;
        end
      end
    end
    if (_T_3001) begin
      if (_T_3395) begin
        if (_T_1114) begin
          reg_bp_0_control_u <= _GEN_29;
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_3395) begin
          if (_T_1114) begin
            reg_bp_0_control_x <= _GEN_30;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_3395) begin
          if (_T_1114) begin
            reg_bp_0_control_w <= _GEN_31;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else begin
      if (_T_3001) begin
        if (_T_3395) begin
          if (_T_1114) begin
            reg_bp_0_control_r <= _GEN_32;
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_3395) begin
        if (_T_1116) begin
          reg_bp_0_address <= _GEN_35;
        end
      end
    end
    if (_T_3001) begin
      if (_T_1344) begin
        reg_mie <= _T_3365;
      end else begin
        if (_T_1132) begin
          reg_mie <= _T_3110;
        end
      end
    end
    if (_T_3001) begin
      if (_T_1360) begin
        reg_mideleg <= _T_3386;
      end
    end
    if (_T_3001) begin
      if (_T_1362) begin
        reg_medeleg <= _T_3387;
      end
    end
    if (_T_3001) begin
      if (_T_1130) begin
        reg_mip_seip <= _T_3089_seip;
      end
    end
    if (_T_3001) begin
      if (_T_1130) begin
        reg_mip_stip <= _T_3089_stip;
      end
    end
    if (_T_3001) begin
      if (_T_1342) begin
        reg_mip_ssip <= _T_3321_ssip;
      end else begin
        if (_T_1130) begin
          reg_mip_ssip <= _T_3089_ssip;
        end
      end
    end
    reg_mepc <= _GEN_430[39:0];
    if (_T_3001) begin
      if (_T_1140) begin
        reg_mcause <= _T_3129;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              if (insn_call) begin
                reg_mcause <= {{60'd0}, _T_2401};
              end else begin
                if (insn_break) begin
                  reg_mcause <= 64'h3;
                end else begin
                  reg_mcause <= io_cause;
                end
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            if (insn_call) begin
              reg_mcause <= {{60'd0}, _T_2401};
            end else begin
              if (insn_break) begin
                reg_mcause <= 64'h3;
              end else begin
                reg_mcause <= io_cause;
              end
            end
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_1138) begin
        reg_mbadaddr <= _T_3130;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(delegate)) begin
              if (write_badaddr) begin
                reg_mbadaddr <= io_badaddr;
              end else begin
                reg_mbadaddr <= 40'h0;
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (!(delegate)) begin
            if (write_badaddr) begin
              reg_mbadaddr <= io_badaddr;
            end else begin
              reg_mbadaddr <= 40'h0;
            end
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_1134) begin
        reg_mscratch <= wdata;
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      reg_mtvec <= _GEN_432[31:0];
    end
    reg_mcounteren <= _GEN_545[31:0];
    reg_scounteren <= _GEN_544[31:0];
    reg_sepc <= _GEN_538[39:0];
    if (_T_3001) begin
      if (_T_1348) begin
        reg_scause <= _T_3384;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (delegate) begin
              if (insn_call) begin
                reg_scause <= {{60'd0}, _T_2401};
              end else begin
                if (insn_break) begin
                  reg_scause <= 64'h3;
                end else begin
                  reg_scause <= io_cause;
                end
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            if (insn_call) begin
              reg_scause <= {{60'd0}, _T_2401};
            end else begin
              if (insn_break) begin
                reg_scause <= 64'h3;
              end else begin
                reg_scause <= io_cause;
              end
            end
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_1350) begin
        reg_sbadaddr <= _T_3130;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (delegate) begin
              if (write_badaddr) begin
                reg_sbadaddr <= io_badaddr;
              end else begin
                reg_sbadaddr <= 40'h0;
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (delegate) begin
            if (write_badaddr) begin
              reg_sbadaddr <= io_badaddr;
            end else begin
              reg_sbadaddr <= 40'h0;
            end
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_1346) begin
        reg_sscratch <= wdata;
      end
    end
    reg_stvec <= _GEN_539[38:0];
    if (_T_3001) begin
      if (_T_1352) begin
        if (_T_3354) begin
          reg_sptbr_mode <= 4'h8;
        end else begin
          if (_T_3351) begin
            reg_sptbr_mode <= 4'h0;
          end
        end
      end
    end
    if (_T_3001) begin
      if (_T_1352) begin
        if (_T_3360) begin
          reg_sptbr_ppn <= {{24'd0}, _T_3361};
        end
      end
    end
    if (reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if (_T_2497) begin
        reg_wfi <= 1'h0;
      end else begin
        if (_T_2492) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    reg_fflags <= _GEN_526[4:0];
    reg_frm <= _GEN_527[2:0];
    if (reset) begin
      _T_328 <= 6'h0;
    end else begin
      _T_328 <= _GEN_524[5:0];
    end
    if (reset) begin
      _T_332 <= 58'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1158) begin
          _T_332 <= _T_3248;
        end else begin
          if (_T_333) begin
            _T_332 <= _T_336;
          end
        end
      end else begin
        if (_T_333) begin
          _T_332 <= _T_336;
        end
      end
    end
    if (reset) begin
      _T_341 <= 6'h0;
    end else begin
      _T_341 <= _GEN_522[5:0];
    end
    if (reset) begin
      _T_345 <= 58'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1156) begin
          _T_345 <= _T_3248;
        end else begin
          if (_T_346) begin
            _T_345 <= _T_349;
          end
        end
      end else begin
        if (_T_346) begin
          _T_345 <= _T_349;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_0 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1160) begin
          reg_hpmevent_0 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_1 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1166) begin
          reg_hpmevent_1 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_2 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1172) begin
          reg_hpmevent_2 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_3 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1178) begin
          reg_hpmevent_3 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_4 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1184) begin
          reg_hpmevent_4 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_5 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1190) begin
          reg_hpmevent_5 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_6 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1196) begin
          reg_hpmevent_6 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_7 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1202) begin
          reg_hpmevent_7 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_8 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1208) begin
          reg_hpmevent_8 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_9 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1214) begin
          reg_hpmevent_9 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_10 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1220) begin
          reg_hpmevent_10 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_11 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1226) begin
          reg_hpmevent_11 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_12 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1232) begin
          reg_hpmevent_12 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_13 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1238) begin
          reg_hpmevent_13 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_14 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1244) begin
          reg_hpmevent_14 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_15 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1250) begin
          reg_hpmevent_15 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_16 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1256) begin
          reg_hpmevent_16 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_17 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1262) begin
          reg_hpmevent_17 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_18 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1268) begin
          reg_hpmevent_18 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_19 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1274) begin
          reg_hpmevent_19 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_20 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1280) begin
          reg_hpmevent_20 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_21 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1286) begin
          reg_hpmevent_21 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_22 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1292) begin
          reg_hpmevent_22 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_23 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1298) begin
          reg_hpmevent_23 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_24 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1304) begin
          reg_hpmevent_24 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_25 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1310) begin
          reg_hpmevent_25 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_26 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1316) begin
          reg_hpmevent_26 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_27 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1322) begin
          reg_hpmevent_27 <= _T_3134;
        end
      end
    end
    if (reset) begin
      reg_hpmevent_28 <= 64'h0;
    end else begin
      if (_T_3001) begin
        if (_T_1328) begin
          reg_hpmevent_28 <= _T_3134;
        end
      end
    end
    _T_410 <= _GEN_435[5:0];
    if (_T_3001) begin
      if (_T_1162) begin
        _T_413 <= _T_3132;
      end else begin
        if (_T_414) begin
          _T_413 <= _T_417;
        end
      end
    end else begin
      if (_T_414) begin
        _T_413 <= _T_417;
      end
    end
    _T_420 <= _GEN_438[5:0];
    if (_T_3001) begin
      if (_T_1168) begin
        _T_423 <= _T_3132;
      end else begin
        if (_T_424) begin
          _T_423 <= _T_427;
        end
      end
    end else begin
      if (_T_424) begin
        _T_423 <= _T_427;
      end
    end
    _T_430 <= _GEN_441[5:0];
    if (_T_3001) begin
      if (_T_1174) begin
        _T_433 <= _T_3132;
      end else begin
        if (_T_434) begin
          _T_433 <= _T_437;
        end
      end
    end else begin
      if (_T_434) begin
        _T_433 <= _T_437;
      end
    end
    _T_440 <= _GEN_444[5:0];
    if (_T_3001) begin
      if (_T_1180) begin
        _T_443 <= _T_3132;
      end else begin
        if (_T_444) begin
          _T_443 <= _T_447;
        end
      end
    end else begin
      if (_T_444) begin
        _T_443 <= _T_447;
      end
    end
    _T_450 <= _GEN_447[5:0];
    if (_T_3001) begin
      if (_T_1186) begin
        _T_453 <= _T_3132;
      end else begin
        if (_T_454) begin
          _T_453 <= _T_457;
        end
      end
    end else begin
      if (_T_454) begin
        _T_453 <= _T_457;
      end
    end
    _T_460 <= _GEN_450[5:0];
    if (_T_3001) begin
      if (_T_1192) begin
        _T_463 <= _T_3132;
      end else begin
        if (_T_464) begin
          _T_463 <= _T_467;
        end
      end
    end else begin
      if (_T_464) begin
        _T_463 <= _T_467;
      end
    end
    _T_470 <= _GEN_453[5:0];
    if (_T_3001) begin
      if (_T_1198) begin
        _T_473 <= _T_3132;
      end else begin
        if (_T_474) begin
          _T_473 <= _T_477;
        end
      end
    end else begin
      if (_T_474) begin
        _T_473 <= _T_477;
      end
    end
    _T_480 <= _GEN_456[5:0];
    if (_T_3001) begin
      if (_T_1204) begin
        _T_483 <= _T_3132;
      end else begin
        if (_T_484) begin
          _T_483 <= _T_487;
        end
      end
    end else begin
      if (_T_484) begin
        _T_483 <= _T_487;
      end
    end
    _T_490 <= _GEN_459[5:0];
    if (_T_3001) begin
      if (_T_1210) begin
        _T_493 <= _T_3132;
      end else begin
        if (_T_494) begin
          _T_493 <= _T_497;
        end
      end
    end else begin
      if (_T_494) begin
        _T_493 <= _T_497;
      end
    end
    _T_500 <= _GEN_462[5:0];
    if (_T_3001) begin
      if (_T_1216) begin
        _T_503 <= _T_3132;
      end else begin
        if (_T_504) begin
          _T_503 <= _T_507;
        end
      end
    end else begin
      if (_T_504) begin
        _T_503 <= _T_507;
      end
    end
    _T_510 <= _GEN_465[5:0];
    if (_T_3001) begin
      if (_T_1222) begin
        _T_513 <= _T_3132;
      end else begin
        if (_T_514) begin
          _T_513 <= _T_517;
        end
      end
    end else begin
      if (_T_514) begin
        _T_513 <= _T_517;
      end
    end
    _T_520 <= _GEN_468[5:0];
    if (_T_3001) begin
      if (_T_1228) begin
        _T_523 <= _T_3132;
      end else begin
        if (_T_524) begin
          _T_523 <= _T_527;
        end
      end
    end else begin
      if (_T_524) begin
        _T_523 <= _T_527;
      end
    end
    _T_530 <= _GEN_471[5:0];
    if (_T_3001) begin
      if (_T_1234) begin
        _T_533 <= _T_3132;
      end else begin
        if (_T_534) begin
          _T_533 <= _T_537;
        end
      end
    end else begin
      if (_T_534) begin
        _T_533 <= _T_537;
      end
    end
    _T_540 <= _GEN_474[5:0];
    if (_T_3001) begin
      if (_T_1240) begin
        _T_543 <= _T_3132;
      end else begin
        if (_T_544) begin
          _T_543 <= _T_547;
        end
      end
    end else begin
      if (_T_544) begin
        _T_543 <= _T_547;
      end
    end
    _T_550 <= _GEN_477[5:0];
    if (_T_3001) begin
      if (_T_1246) begin
        _T_553 <= _T_3132;
      end else begin
        if (_T_554) begin
          _T_553 <= _T_557;
        end
      end
    end else begin
      if (_T_554) begin
        _T_553 <= _T_557;
      end
    end
    _T_560 <= _GEN_480[5:0];
    if (_T_3001) begin
      if (_T_1252) begin
        _T_563 <= _T_3132;
      end else begin
        if (_T_564) begin
          _T_563 <= _T_567;
        end
      end
    end else begin
      if (_T_564) begin
        _T_563 <= _T_567;
      end
    end
    _T_570 <= _GEN_483[5:0];
    if (_T_3001) begin
      if (_T_1258) begin
        _T_573 <= _T_3132;
      end else begin
        if (_T_574) begin
          _T_573 <= _T_577;
        end
      end
    end else begin
      if (_T_574) begin
        _T_573 <= _T_577;
      end
    end
    _T_580 <= _GEN_486[5:0];
    if (_T_3001) begin
      if (_T_1264) begin
        _T_583 <= _T_3132;
      end else begin
        if (_T_584) begin
          _T_583 <= _T_587;
        end
      end
    end else begin
      if (_T_584) begin
        _T_583 <= _T_587;
      end
    end
    _T_590 <= _GEN_489[5:0];
    if (_T_3001) begin
      if (_T_1270) begin
        _T_593 <= _T_3132;
      end else begin
        if (_T_594) begin
          _T_593 <= _T_597;
        end
      end
    end else begin
      if (_T_594) begin
        _T_593 <= _T_597;
      end
    end
    _T_600 <= _GEN_492[5:0];
    if (_T_3001) begin
      if (_T_1276) begin
        _T_603 <= _T_3132;
      end else begin
        if (_T_604) begin
          _T_603 <= _T_607;
        end
      end
    end else begin
      if (_T_604) begin
        _T_603 <= _T_607;
      end
    end
    _T_610 <= _GEN_495[5:0];
    if (_T_3001) begin
      if (_T_1282) begin
        _T_613 <= _T_3132;
      end else begin
        if (_T_614) begin
          _T_613 <= _T_617;
        end
      end
    end else begin
      if (_T_614) begin
        _T_613 <= _T_617;
      end
    end
    _T_620 <= _GEN_498[5:0];
    if (_T_3001) begin
      if (_T_1288) begin
        _T_623 <= _T_3132;
      end else begin
        if (_T_624) begin
          _T_623 <= _T_627;
        end
      end
    end else begin
      if (_T_624) begin
        _T_623 <= _T_627;
      end
    end
    _T_630 <= _GEN_501[5:0];
    if (_T_3001) begin
      if (_T_1294) begin
        _T_633 <= _T_3132;
      end else begin
        if (_T_634) begin
          _T_633 <= _T_637;
        end
      end
    end else begin
      if (_T_634) begin
        _T_633 <= _T_637;
      end
    end
    _T_640 <= _GEN_504[5:0];
    if (_T_3001) begin
      if (_T_1300) begin
        _T_643 <= _T_3132;
      end else begin
        if (_T_644) begin
          _T_643 <= _T_647;
        end
      end
    end else begin
      if (_T_644) begin
        _T_643 <= _T_647;
      end
    end
    _T_650 <= _GEN_507[5:0];
    if (_T_3001) begin
      if (_T_1306) begin
        _T_653 <= _T_3132;
      end else begin
        if (_T_654) begin
          _T_653 <= _T_657;
        end
      end
    end else begin
      if (_T_654) begin
        _T_653 <= _T_657;
      end
    end
    _T_660 <= _GEN_510[5:0];
    if (_T_3001) begin
      if (_T_1312) begin
        _T_663 <= _T_3132;
      end else begin
        if (_T_664) begin
          _T_663 <= _T_667;
        end
      end
    end else begin
      if (_T_664) begin
        _T_663 <= _T_667;
      end
    end
    _T_670 <= _GEN_513[5:0];
    if (_T_3001) begin
      if (_T_1318) begin
        _T_673 <= _T_3132;
      end else begin
        if (_T_674) begin
          _T_673 <= _T_677;
        end
      end
    end else begin
      if (_T_674) begin
        _T_673 <= _T_677;
      end
    end
    _T_680 <= _GEN_516[5:0];
    if (_T_3001) begin
      if (_T_1324) begin
        _T_683 <= _T_3132;
      end else begin
        if (_T_684) begin
          _T_683 <= _T_687;
        end
      end
    end else begin
      if (_T_684) begin
        _T_683 <= _T_687;
      end
    end
    _T_690 <= _GEN_519[5:0];
    if (_T_3001) begin
      if (_T_1330) begin
        _T_693 <= _T_3132;
      end else begin
        if (_T_694) begin
          _T_693 <= _T_697;
        end
      end
    end else begin
      if (_T_694) begin
        _T_693 <= _T_697;
      end
    end
    _T_711 <= io_interrupts_seip;
    if (reset) begin
      reg_misa <= 64'h8000000000141129;
    end else begin
      if (_T_3001) begin
        if (_T_1124) begin
          reg_misa <= _T_3053;
        end
      end
    end
    if (_T_2473) begin
      _T_2476 <= reg_mstatus_mpp;
    end else begin
      _T_2476 <= reg_mstatus_prv;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2486) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:517 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2486) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2507) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:521 assert(!reg_wfi || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2507) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2522) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:525 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2531) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:526 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2531) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BoomCore(
  input         clock,
  input         reset,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  output        io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_sfence_bits_rs2,
  output [38:0] io_imem_sfence_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [39:0] io_imem_resp_bits_pc,
  input  [63:0] io_imem_resp_bits_data,
  input  [1:0]  io_imem_resp_bits_mask,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_flush_icache,
  input         io_imem_perf_acquire,
  input         io_imem_perf_tlbMiss,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [2:0]  io_dmem_req_bits_typ,
  output        io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [63:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_has_data,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  output        io_dmem_invalidate_lr,
  input         io_dmem_ordered,
  input         io_dmem_perf_acquire,
  input         io_dmem_perf_release,
  input         io_dmem_perf_tlbMiss,
  output [3:0]  io_ptw_ptbr_mode,
  output [43:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output [1:0]  io_ptw_status_dprv,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  input         io_ptw_tlb_req_ready,
  output        io_ptw_tlb_req_valid,
  output [26:0] io_ptw_tlb_req_bits_addr,
  input         io_ptw_tlb_resp_valid,
  input         io_ptw_tlb_resp_bits_ae,
  input  [53:0] io_ptw_tlb_resp_bits_pte_ppn,
  input         io_ptw_tlb_resp_bits_pte_d,
  input         io_ptw_tlb_resp_bits_pte_a,
  input         io_ptw_tlb_resp_bits_pte_g,
  input         io_ptw_tlb_resp_bits_pte_u,
  input         io_ptw_tlb_resp_bits_pte_x,
  input         io_ptw_tlb_resp_bits_pte_w,
  input         io_ptw_tlb_resp_bits_pte_r,
  input         io_ptw_tlb_resp_bits_pte_v,
  input  [1:0]  io_ptw_tlb_resp_bits_level,
  input         io_ptw_tlb_resp_bits_homogeneous,
  input  [3:0]  io_ptw_tlb_ptbr_mode,
  input  [1:0]  io_ptw_tlb_status_dprv,
  input         io_ptw_tlb_status_mxr,
  input         io_ptw_tlb_status_sum
);
  wire  mem_unit_clock;
  wire  mem_unit_reset;
  wire  mem_unit_io_req_valid;
  wire [8:0] mem_unit_io_req_bits_uop_uopc;
  wire  mem_unit_io_req_bits_uop_ctrl_is_load;
  wire  mem_unit_io_req_bits_uop_ctrl_is_sta;
  wire  mem_unit_io_req_bits_uop_ctrl_is_std;
  wire [7:0] mem_unit_io_req_bits_uop_br_mask;
  wire [19:0] mem_unit_io_req_bits_uop_imm_packed;
  wire [6:0] mem_unit_io_req_bits_uop_rob_idx;
  wire [3:0] mem_unit_io_req_bits_uop_ldq_idx;
  wire [3:0] mem_unit_io_req_bits_uop_stq_idx;
  wire [6:0] mem_unit_io_req_bits_uop_pdst;
  wire [4:0] mem_unit_io_req_bits_uop_mem_cmd;
  wire [2:0] mem_unit_io_req_bits_uop_mem_typ;
  wire  mem_unit_io_req_bits_uop_is_fence;
  wire  mem_unit_io_req_bits_uop_is_store;
  wire  mem_unit_io_req_bits_uop_is_amo;
  wire  mem_unit_io_req_bits_uop_is_load;
  wire [1:0] mem_unit_io_req_bits_uop_dst_rtype;
  wire  mem_unit_io_req_bits_uop_fp_val;
  wire [64:0] mem_unit_io_req_bits_rs1_data;
  wire [64:0] mem_unit_io_req_bits_rs2_data;
  wire  mem_unit_io_resp_0_valid;
  wire [8:0] mem_unit_io_resp_0_bits_uop_uopc;
  wire  mem_unit_io_resp_0_bits_uop_ctrl_rf_wen;
  wire [6:0] mem_unit_io_resp_0_bits_uop_rob_idx;
  wire [6:0] mem_unit_io_resp_0_bits_uop_pdst;
  wire [2:0] mem_unit_io_resp_0_bits_uop_mem_typ;
  wire  mem_unit_io_resp_0_bits_uop_is_store;
  wire  mem_unit_io_resp_0_bits_uop_is_amo;
  wire [1:0] mem_unit_io_resp_0_bits_uop_dst_rtype;
  wire  mem_unit_io_resp_0_bits_uop_fp_val;
  wire [64:0] mem_unit_io_resp_0_bits_data;
  wire  mem_unit_io_brinfo_valid;
  wire  mem_unit_io_brinfo_mispredict;
  wire [7:0] mem_unit_io_brinfo_mask;
  wire  mem_unit_io_lsu_io_exe_resp_valid;
  wire [8:0] mem_unit_io_lsu_io_exe_resp_bits_uop_uopc;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_load;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_sta;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_std;
  wire [7:0] mem_unit_io_lsu_io_exe_resp_bits_uop_br_mask;
  wire [6:0] mem_unit_io_lsu_io_exe_resp_bits_uop_rob_idx;
  wire [3:0] mem_unit_io_lsu_io_exe_resp_bits_uop_ldq_idx;
  wire [3:0] mem_unit_io_lsu_io_exe_resp_bits_uop_stq_idx;
  wire [6:0] mem_unit_io_lsu_io_exe_resp_bits_uop_pdst;
  wire [4:0] mem_unit_io_lsu_io_exe_resp_bits_uop_mem_cmd;
  wire [2:0] mem_unit_io_lsu_io_exe_resp_bits_uop_mem_typ;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_is_fence;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_is_store;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_is_amo;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_is_load;
  wire [1:0] mem_unit_io_lsu_io_exe_resp_bits_uop_dst_rtype;
  wire  mem_unit_io_lsu_io_exe_resp_bits_uop_fp_val;
  wire [63:0] mem_unit_io_lsu_io_exe_resp_bits_data;
  wire [39:0] mem_unit_io_lsu_io_exe_resp_bits_addr;
  wire  mem_unit_io_lsu_io_exe_resp_bits_mxcpt_valid;
  wire [16:0] mem_unit_io_lsu_io_exe_resp_bits_mxcpt_bits;
  wire  mem_unit_io_lsu_io_exe_resp_bits_sfence_valid;
  wire  mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs1;
  wire  mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs2;
  wire [38:0] mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_addr;
  wire  mem_unit_io_lsu_io_memreq_val;
  wire [31:0] mem_unit_io_lsu_io_memreq_addr;
  wire [63:0] mem_unit_io_lsu_io_memreq_wdata;
  wire [8:0] mem_unit_io_lsu_io_memreq_uop_uopc;
  wire [7:0] mem_unit_io_lsu_io_memreq_uop_br_mask;
  wire [6:0] mem_unit_io_lsu_io_memreq_uop_rob_idx;
  wire [3:0] mem_unit_io_lsu_io_memreq_uop_ldq_idx;
  wire [3:0] mem_unit_io_lsu_io_memreq_uop_stq_idx;
  wire [6:0] mem_unit_io_lsu_io_memreq_uop_pdst;
  wire [4:0] mem_unit_io_lsu_io_memreq_uop_mem_cmd;
  wire [2:0] mem_unit_io_lsu_io_memreq_uop_mem_typ;
  wire  mem_unit_io_lsu_io_memreq_uop_is_store;
  wire  mem_unit_io_lsu_io_memreq_uop_is_amo;
  wire  mem_unit_io_lsu_io_memreq_uop_is_load;
  wire [1:0] mem_unit_io_lsu_io_memreq_uop_dst_rtype;
  wire  mem_unit_io_lsu_io_memreq_uop_fp_val;
  wire  mem_unit_io_lsu_io_memreq_kill;
  wire  mem_unit_io_lsu_io_forward_val;
  wire [63:0] mem_unit_io_lsu_io_forward_data;
  wire [8:0] mem_unit_io_lsu_io_forward_uop_uopc;
  wire [6:0] mem_unit_io_lsu_io_forward_uop_rob_idx;
  wire [3:0] mem_unit_io_lsu_io_forward_uop_ldq_idx;
  wire [3:0] mem_unit_io_lsu_io_forward_uop_stq_idx;
  wire [6:0] mem_unit_io_lsu_io_forward_uop_pdst;
  wire [2:0] mem_unit_io_lsu_io_forward_uop_mem_typ;
  wire  mem_unit_io_lsu_io_forward_uop_is_store;
  wire  mem_unit_io_lsu_io_forward_uop_is_amo;
  wire  mem_unit_io_lsu_io_forward_uop_is_load;
  wire [1:0] mem_unit_io_lsu_io_forward_uop_dst_rtype;
  wire  mem_unit_io_lsu_io_forward_uop_fp_val;
  wire  mem_unit_io_lsu_io_memresp_valid;
  wire [3:0] mem_unit_io_lsu_io_memresp_bits_ldq_idx;
  wire [3:0] mem_unit_io_lsu_io_memresp_bits_stq_idx;
  wire  mem_unit_io_lsu_io_memresp_bits_is_load;
  wire  mem_unit_io_dmem_req_valid;
  wire [39:0] mem_unit_io_dmem_req_bits_addr;
  wire [8:0] mem_unit_io_dmem_req_bits_uop_uopc;
  wire [7:0] mem_unit_io_dmem_req_bits_uop_br_mask;
  wire [6:0] mem_unit_io_dmem_req_bits_uop_rob_idx;
  wire [3:0] mem_unit_io_dmem_req_bits_uop_ldq_idx;
  wire [3:0] mem_unit_io_dmem_req_bits_uop_stq_idx;
  wire [6:0] mem_unit_io_dmem_req_bits_uop_pdst;
  wire [4:0] mem_unit_io_dmem_req_bits_uop_mem_cmd;
  wire [2:0] mem_unit_io_dmem_req_bits_uop_mem_typ;
  wire  mem_unit_io_dmem_req_bits_uop_is_store;
  wire  mem_unit_io_dmem_req_bits_uop_is_amo;
  wire  mem_unit_io_dmem_req_bits_uop_is_load;
  wire [1:0] mem_unit_io_dmem_req_bits_uop_dst_rtype;
  wire  mem_unit_io_dmem_req_bits_uop_fp_val;
  wire [63:0] mem_unit_io_dmem_req_bits_data;
  wire  mem_unit_io_dmem_req_bits_kill;
  wire  mem_unit_io_dmem_resp_valid;
  wire [63:0] mem_unit_io_dmem_resp_bits_data_subword;
  wire [8:0] mem_unit_io_dmem_resp_bits_uop_uopc;
  wire [6:0] mem_unit_io_dmem_resp_bits_uop_rob_idx;
  wire [3:0] mem_unit_io_dmem_resp_bits_uop_ldq_idx;
  wire [3:0] mem_unit_io_dmem_resp_bits_uop_stq_idx;
  wire [6:0] mem_unit_io_dmem_resp_bits_uop_pdst;
  wire [4:0] mem_unit_io_dmem_resp_bits_uop_mem_cmd;
  wire [2:0] mem_unit_io_dmem_resp_bits_uop_mem_typ;
  wire  mem_unit_io_dmem_resp_bits_uop_is_store;
  wire  mem_unit_io_dmem_resp_bits_uop_is_amo;
  wire  mem_unit_io_dmem_resp_bits_uop_is_load;
  wire [1:0] mem_unit_io_dmem_resp_bits_uop_dst_rtype;
  wire  mem_unit_io_dmem_resp_bits_uop_fp_val;
  wire  mem_unit_io_com_exception;
  wire  csr_exe_unit_clock;
  wire  csr_exe_unit_reset;
  wire [9:0] csr_exe_unit_io_fu_types;
  wire  csr_exe_unit_io_req_valid;
  wire  csr_exe_unit_io_req_bits_uop_valid;
  wire [1:0] csr_exe_unit_io_req_bits_uop_iw_state;
  wire [8:0] csr_exe_unit_io_req_bits_uop_uopc;
  wire [31:0] csr_exe_unit_io_req_bits_uop_inst;
  wire [39:0] csr_exe_unit_io_req_bits_uop_pc;
  wire [1:0] csr_exe_unit_io_req_bits_uop_iqtype;
  wire [9:0] csr_exe_unit_io_req_bits_uop_fu_code;
  wire [3:0] csr_exe_unit_io_req_bits_uop_ctrl_br_type;
  wire [1:0] csr_exe_unit_io_req_bits_uop_ctrl_op1_sel;
  wire [2:0] csr_exe_unit_io_req_bits_uop_ctrl_op2_sel;
  wire [2:0] csr_exe_unit_io_req_bits_uop_ctrl_imm_sel;
  wire [3:0] csr_exe_unit_io_req_bits_uop_ctrl_op_fcn;
  wire  csr_exe_unit_io_req_bits_uop_ctrl_fcn_dw;
  wire  csr_exe_unit_io_req_bits_uop_ctrl_rf_wen;
  wire [2:0] csr_exe_unit_io_req_bits_uop_ctrl_csr_cmd;
  wire  csr_exe_unit_io_req_bits_uop_ctrl_is_load;
  wire  csr_exe_unit_io_req_bits_uop_ctrl_is_sta;
  wire  csr_exe_unit_io_req_bits_uop_ctrl_is_std;
  wire  csr_exe_unit_io_req_bits_uop_allocate_brtag;
  wire  csr_exe_unit_io_req_bits_uop_is_br_or_jmp;
  wire  csr_exe_unit_io_req_bits_uop_is_jump;
  wire  csr_exe_unit_io_req_bits_uop_is_jal;
  wire  csr_exe_unit_io_req_bits_uop_is_ret;
  wire  csr_exe_unit_io_req_bits_uop_is_call;
  wire [7:0] csr_exe_unit_io_req_bits_uop_br_mask;
  wire [2:0] csr_exe_unit_io_req_bits_uop_br_tag;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_btb_blame;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_btb_hit;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_btb_taken;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_bpd_blame;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_bpd_hit;
  wire  csr_exe_unit_io_req_bits_uop_br_prediction_bpd_taken;
  wire [1:0] csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_value;
  wire [5:0] csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_takens;
  wire [14:0] csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history;
  wire [14:0] csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_info;
  wire  csr_exe_unit_io_req_bits_uop_stat_brjmp_mispredicted;
  wire  csr_exe_unit_io_req_bits_uop_stat_btb_made_pred;
  wire  csr_exe_unit_io_req_bits_uop_stat_btb_mispredicted;
  wire  csr_exe_unit_io_req_bits_uop_stat_bpd_made_pred;
  wire  csr_exe_unit_io_req_bits_uop_stat_bpd_mispredicted;
  wire [2:0] csr_exe_unit_io_req_bits_uop_fetch_pc_lob;
  wire [19:0] csr_exe_unit_io_req_bits_uop_imm_packed;
  wire [11:0] csr_exe_unit_io_req_bits_uop_csr_addr;
  wire [6:0] csr_exe_unit_io_req_bits_uop_rob_idx;
  wire [3:0] csr_exe_unit_io_req_bits_uop_ldq_idx;
  wire [3:0] csr_exe_unit_io_req_bits_uop_stq_idx;
  wire [5:0] csr_exe_unit_io_req_bits_uop_brob_idx;
  wire [6:0] csr_exe_unit_io_req_bits_uop_pdst;
  wire [6:0] csr_exe_unit_io_req_bits_uop_pop1;
  wire [6:0] csr_exe_unit_io_req_bits_uop_pop2;
  wire [6:0] csr_exe_unit_io_req_bits_uop_pop3;
  wire  csr_exe_unit_io_req_bits_uop_prs1_busy;
  wire  csr_exe_unit_io_req_bits_uop_prs2_busy;
  wire  csr_exe_unit_io_req_bits_uop_prs3_busy;
  wire [6:0] csr_exe_unit_io_req_bits_uop_stale_pdst;
  wire  csr_exe_unit_io_req_bits_uop_exception;
  wire [63:0] csr_exe_unit_io_req_bits_uop_exc_cause;
  wire  csr_exe_unit_io_req_bits_uop_bypassable;
  wire [4:0] csr_exe_unit_io_req_bits_uop_mem_cmd;
  wire [2:0] csr_exe_unit_io_req_bits_uop_mem_typ;
  wire  csr_exe_unit_io_req_bits_uop_is_fence;
  wire  csr_exe_unit_io_req_bits_uop_is_fencei;
  wire  csr_exe_unit_io_req_bits_uop_is_store;
  wire  csr_exe_unit_io_req_bits_uop_is_amo;
  wire  csr_exe_unit_io_req_bits_uop_is_load;
  wire  csr_exe_unit_io_req_bits_uop_is_sys_pc2epc;
  wire  csr_exe_unit_io_req_bits_uop_is_unique;
  wire  csr_exe_unit_io_req_bits_uop_flush_on_commit;
  wire [5:0] csr_exe_unit_io_req_bits_uop_ldst;
  wire [5:0] csr_exe_unit_io_req_bits_uop_lrs1;
  wire [5:0] csr_exe_unit_io_req_bits_uop_lrs2;
  wire [5:0] csr_exe_unit_io_req_bits_uop_lrs3;
  wire  csr_exe_unit_io_req_bits_uop_ldst_val;
  wire [1:0] csr_exe_unit_io_req_bits_uop_dst_rtype;
  wire [1:0] csr_exe_unit_io_req_bits_uop_lrs1_rtype;
  wire [1:0] csr_exe_unit_io_req_bits_uop_lrs2_rtype;
  wire  csr_exe_unit_io_req_bits_uop_frs3_en;
  wire  csr_exe_unit_io_req_bits_uop_fp_val;
  wire  csr_exe_unit_io_req_bits_uop_fp_single;
  wire  csr_exe_unit_io_req_bits_uop_xcpt_pf_if;
  wire  csr_exe_unit_io_req_bits_uop_xcpt_ae_if;
  wire  csr_exe_unit_io_req_bits_uop_replay_if;
  wire  csr_exe_unit_io_req_bits_uop_xcpt_ma_if;
  wire [63:0] csr_exe_unit_io_req_bits_uop_debug_wdata;
  wire [31:0] csr_exe_unit_io_req_bits_uop_debug_events_fetch_seq;
  wire [63:0] csr_exe_unit_io_req_bits_rs1_data;
  wire [63:0] csr_exe_unit_io_req_bits_rs2_data;
  wire  csr_exe_unit_io_req_bits_kill;
  wire  csr_exe_unit_io_resp_0_valid;
  wire  csr_exe_unit_io_resp_0_bits_uop_ctrl_rf_wen;
  wire [2:0] csr_exe_unit_io_resp_0_bits_uop_ctrl_csr_cmd;
  wire [11:0] csr_exe_unit_io_resp_0_bits_uop_csr_addr;
  wire [6:0] csr_exe_unit_io_resp_0_bits_uop_rob_idx;
  wire [6:0] csr_exe_unit_io_resp_0_bits_uop_pdst;
  wire  csr_exe_unit_io_resp_0_bits_uop_bypassable;
  wire  csr_exe_unit_io_resp_0_bits_uop_is_store;
  wire  csr_exe_unit_io_resp_0_bits_uop_is_amo;
  wire [1:0] csr_exe_unit_io_resp_0_bits_uop_dst_rtype;
  wire [63:0] csr_exe_unit_io_resp_0_bits_data;
  wire  csr_exe_unit_io_bypass_valid_0;
  wire  csr_exe_unit_io_bypass_valid_1;
  wire  csr_exe_unit_io_bypass_valid_2;
  wire  csr_exe_unit_io_bypass_uop_0_ctrl_rf_wen;
  wire [6:0] csr_exe_unit_io_bypass_uop_0_pdst;
  wire [1:0] csr_exe_unit_io_bypass_uop_0_dst_rtype;
  wire  csr_exe_unit_io_bypass_uop_1_ctrl_rf_wen;
  wire [6:0] csr_exe_unit_io_bypass_uop_1_pdst;
  wire [1:0] csr_exe_unit_io_bypass_uop_1_dst_rtype;
  wire  csr_exe_unit_io_bypass_uop_2_ctrl_rf_wen;
  wire [6:0] csr_exe_unit_io_bypass_uop_2_pdst;
  wire [1:0] csr_exe_unit_io_bypass_uop_2_dst_rtype;
  wire [63:0] csr_exe_unit_io_bypass_data_0;
  wire [63:0] csr_exe_unit_io_bypass_data_1;
  wire [63:0] csr_exe_unit_io_bypass_data_2;
  wire  csr_exe_unit_io_brinfo_valid;
  wire  csr_exe_unit_io_brinfo_mispredict;
  wire [7:0] csr_exe_unit_io_brinfo_mask;
  wire  csr_exe_unit_io_br_unit_take_pc;
  wire [39:0] csr_exe_unit_io_br_unit_target;
  wire  csr_exe_unit_io_br_unit_brinfo_valid;
  wire  csr_exe_unit_io_br_unit_brinfo_mispredict;
  wire [7:0] csr_exe_unit_io_br_unit_brinfo_mask;
  wire [2:0] csr_exe_unit_io_br_unit_brinfo_tag;
  wire [7:0] csr_exe_unit_io_br_unit_brinfo_exe_mask;
  wire [6:0] csr_exe_unit_io_br_unit_brinfo_rob_idx;
  wire [3:0] csr_exe_unit_io_br_unit_brinfo_ldq_idx;
  wire [3:0] csr_exe_unit_io_br_unit_brinfo_stq_idx;
  wire  csr_exe_unit_io_br_unit_brinfo_is_jr;
  wire  csr_exe_unit_io_br_unit_btb_update_valid;
  wire [38:0] csr_exe_unit_io_br_unit_btb_update_bits_pc;
  wire [38:0] csr_exe_unit_io_br_unit_btb_update_bits_target;
  wire [38:0] csr_exe_unit_io_br_unit_btb_update_bits_cfi_pc;
  wire [2:0] csr_exe_unit_io_br_unit_btb_update_bits_bpd_type;
  wire [2:0] csr_exe_unit_io_br_unit_btb_update_bits_cfi_type;
  wire  csr_exe_unit_io_br_unit_bim_update_valid;
  wire  csr_exe_unit_io_br_unit_bim_update_bits_taken;
  wire [1:0] csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_value;
  wire [5:0] csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_entry_idx;
  wire [1:0] csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_way_idx;
  wire  csr_exe_unit_io_br_unit_bpd_update_valid;
  wire [2:0] csr_exe_unit_io_br_unit_bpd_update_bits_br_pc;
  wire [5:0] csr_exe_unit_io_br_unit_bpd_update_bits_brob_idx;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_mispredict;
  wire [14:0] csr_exe_unit_io_br_unit_bpd_update_bits_history;
  wire [7:0] csr_exe_unit_io_br_unit_bpd_update_bits_history_ptr;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_bpd_predict_val;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_bpd_mispredict;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_taken;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_is_br;
  wire  csr_exe_unit_io_br_unit_bpd_update_bits_new_pc_same_packet;
  wire  csr_exe_unit_io_br_unit_xcpt_valid;
  wire [7:0] csr_exe_unit_io_br_unit_xcpt_bits_uop_br_mask;
  wire [6:0] csr_exe_unit_io_br_unit_xcpt_bits_uop_rob_idx;
  wire [39:0] csr_exe_unit_io_br_unit_xcpt_bits_badvaddr;
  wire [39:0] csr_exe_unit_io_get_rob_pc_curr_pc;
  wire [5:0] csr_exe_unit_io_get_rob_pc_curr_brob_idx;
  wire  csr_exe_unit_io_get_rob_pc_next_val;
  wire [39:0] csr_exe_unit_io_get_rob_pc_next_pc;
  wire [1:0] csr_exe_unit_io_get_pred_info_bim_resp_value;
  wire [5:0] csr_exe_unit_io_get_pred_info_bim_resp_entry_idx;
  wire [1:0] csr_exe_unit_io_get_pred_info_bim_resp_way_idx;
  wire [14:0] csr_exe_unit_io_get_pred_info_bpd_resp_history;
  wire [7:0] csr_exe_unit_io_get_pred_info_bpd_resp_history_ptr;
  wire  csr_exe_unit_io_status_debug;
  wire  ALUExeUnit_clock;
  wire  ALUExeUnit_reset;
  wire  ALUExeUnit_io_req_valid;
  wire  ALUExeUnit_io_req_bits_uop_valid;
  wire [1:0] ALUExeUnit_io_req_bits_uop_iw_state;
  wire [8:0] ALUExeUnit_io_req_bits_uop_uopc;
  wire [31:0] ALUExeUnit_io_req_bits_uop_inst;
  wire [39:0] ALUExeUnit_io_req_bits_uop_pc;
  wire [1:0] ALUExeUnit_io_req_bits_uop_iqtype;
  wire [9:0] ALUExeUnit_io_req_bits_uop_fu_code;
  wire [1:0] ALUExeUnit_io_req_bits_uop_ctrl_op1_sel;
  wire [2:0] ALUExeUnit_io_req_bits_uop_ctrl_op2_sel;
  wire [2:0] ALUExeUnit_io_req_bits_uop_ctrl_imm_sel;
  wire [3:0] ALUExeUnit_io_req_bits_uop_ctrl_op_fcn;
  wire  ALUExeUnit_io_req_bits_uop_ctrl_fcn_dw;
  wire  ALUExeUnit_io_req_bits_uop_ctrl_rf_wen;
  wire  ALUExeUnit_io_req_bits_uop_ctrl_is_load;
  wire  ALUExeUnit_io_req_bits_uop_ctrl_is_sta;
  wire  ALUExeUnit_io_req_bits_uop_ctrl_is_std;
  wire  ALUExeUnit_io_req_bits_uop_allocate_brtag;
  wire  ALUExeUnit_io_req_bits_uop_is_br_or_jmp;
  wire  ALUExeUnit_io_req_bits_uop_is_jump;
  wire  ALUExeUnit_io_req_bits_uop_is_jal;
  wire  ALUExeUnit_io_req_bits_uop_is_ret;
  wire  ALUExeUnit_io_req_bits_uop_is_call;
  wire [7:0] ALUExeUnit_io_req_bits_uop_br_mask;
  wire [2:0] ALUExeUnit_io_req_bits_uop_br_tag;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_btb_blame;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_btb_hit;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_btb_taken;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_bpd_blame;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_bpd_hit;
  wire  ALUExeUnit_io_req_bits_uop_br_prediction_bpd_taken;
  wire [1:0] ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_value;
  wire [5:0] ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_takens;
  wire [14:0] ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history;
  wire [14:0] ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_info;
  wire  ALUExeUnit_io_req_bits_uop_stat_brjmp_mispredicted;
  wire  ALUExeUnit_io_req_bits_uop_stat_btb_made_pred;
  wire  ALUExeUnit_io_req_bits_uop_stat_btb_mispredicted;
  wire  ALUExeUnit_io_req_bits_uop_stat_bpd_made_pred;
  wire  ALUExeUnit_io_req_bits_uop_stat_bpd_mispredicted;
  wire [2:0] ALUExeUnit_io_req_bits_uop_fetch_pc_lob;
  wire [19:0] ALUExeUnit_io_req_bits_uop_imm_packed;
  wire [11:0] ALUExeUnit_io_req_bits_uop_csr_addr;
  wire [6:0] ALUExeUnit_io_req_bits_uop_rob_idx;
  wire [3:0] ALUExeUnit_io_req_bits_uop_ldq_idx;
  wire [3:0] ALUExeUnit_io_req_bits_uop_stq_idx;
  wire [5:0] ALUExeUnit_io_req_bits_uop_brob_idx;
  wire [6:0] ALUExeUnit_io_req_bits_uop_pdst;
  wire [6:0] ALUExeUnit_io_req_bits_uop_pop1;
  wire [6:0] ALUExeUnit_io_req_bits_uop_pop2;
  wire [6:0] ALUExeUnit_io_req_bits_uop_pop3;
  wire  ALUExeUnit_io_req_bits_uop_prs1_busy;
  wire  ALUExeUnit_io_req_bits_uop_prs2_busy;
  wire  ALUExeUnit_io_req_bits_uop_prs3_busy;
  wire [6:0] ALUExeUnit_io_req_bits_uop_stale_pdst;
  wire  ALUExeUnit_io_req_bits_uop_exception;
  wire [63:0] ALUExeUnit_io_req_bits_uop_exc_cause;
  wire  ALUExeUnit_io_req_bits_uop_bypassable;
  wire [4:0] ALUExeUnit_io_req_bits_uop_mem_cmd;
  wire [2:0] ALUExeUnit_io_req_bits_uop_mem_typ;
  wire  ALUExeUnit_io_req_bits_uop_is_fence;
  wire  ALUExeUnit_io_req_bits_uop_is_fencei;
  wire  ALUExeUnit_io_req_bits_uop_is_store;
  wire  ALUExeUnit_io_req_bits_uop_is_amo;
  wire  ALUExeUnit_io_req_bits_uop_is_load;
  wire  ALUExeUnit_io_req_bits_uop_is_sys_pc2epc;
  wire  ALUExeUnit_io_req_bits_uop_is_unique;
  wire  ALUExeUnit_io_req_bits_uop_flush_on_commit;
  wire [5:0] ALUExeUnit_io_req_bits_uop_ldst;
  wire [5:0] ALUExeUnit_io_req_bits_uop_lrs1;
  wire [5:0] ALUExeUnit_io_req_bits_uop_lrs2;
  wire [5:0] ALUExeUnit_io_req_bits_uop_lrs3;
  wire  ALUExeUnit_io_req_bits_uop_ldst_val;
  wire [1:0] ALUExeUnit_io_req_bits_uop_dst_rtype;
  wire [1:0] ALUExeUnit_io_req_bits_uop_lrs1_rtype;
  wire [1:0] ALUExeUnit_io_req_bits_uop_lrs2_rtype;
  wire  ALUExeUnit_io_req_bits_uop_frs3_en;
  wire  ALUExeUnit_io_req_bits_uop_fp_val;
  wire  ALUExeUnit_io_req_bits_uop_fp_single;
  wire  ALUExeUnit_io_req_bits_uop_xcpt_pf_if;
  wire  ALUExeUnit_io_req_bits_uop_xcpt_ae_if;
  wire  ALUExeUnit_io_req_bits_uop_replay_if;
  wire  ALUExeUnit_io_req_bits_uop_xcpt_ma_if;
  wire [63:0] ALUExeUnit_io_req_bits_uop_debug_wdata;
  wire [31:0] ALUExeUnit_io_req_bits_uop_debug_events_fetch_seq;
  wire [63:0] ALUExeUnit_io_req_bits_rs1_data;
  wire [63:0] ALUExeUnit_io_req_bits_rs2_data;
  wire  ALUExeUnit_io_req_bits_kill;
  wire  ALUExeUnit_io_resp_0_valid;
  wire  ALUExeUnit_io_resp_0_bits_uop_ctrl_rf_wen;
  wire [6:0] ALUExeUnit_io_resp_0_bits_uop_rob_idx;
  wire [6:0] ALUExeUnit_io_resp_0_bits_uop_pdst;
  wire  ALUExeUnit_io_resp_0_bits_uop_bypassable;
  wire  ALUExeUnit_io_resp_0_bits_uop_is_store;
  wire  ALUExeUnit_io_resp_0_bits_uop_is_amo;
  wire [1:0] ALUExeUnit_io_resp_0_bits_uop_dst_rtype;
  wire [63:0] ALUExeUnit_io_resp_0_bits_data;
  wire  ALUExeUnit_io_bypass_valid_0;
  wire  ALUExeUnit_io_bypass_uop_0_ctrl_rf_wen;
  wire [6:0] ALUExeUnit_io_bypass_uop_0_pdst;
  wire [1:0] ALUExeUnit_io_bypass_uop_0_dst_rtype;
  wire [63:0] ALUExeUnit_io_bypass_data_0;
  wire  ALUExeUnit_io_brinfo_valid;
  wire  ALUExeUnit_io_brinfo_mispredict;
  wire [7:0] ALUExeUnit_io_brinfo_mask;
  wire  fp_pipeline_clock;
  wire  fp_pipeline_reset;
  wire  fp_pipeline_io_brinfo_valid;
  wire  fp_pipeline_io_brinfo_mispredict;
  wire [7:0] fp_pipeline_io_brinfo_mask;
  wire  fp_pipeline_io_flush_pipeline;
  wire [2:0] fp_pipeline_io_fcsr_rm;
  wire  fp_pipeline_io_dis_valids_0;
  wire  fp_pipeline_io_dis_valids_1;
  wire  fp_pipeline_io_dis_uops_0_valid;
  wire [8:0] fp_pipeline_io_dis_uops_0_uopc;
  wire [31:0] fp_pipeline_io_dis_uops_0_inst;
  wire [39:0] fp_pipeline_io_dis_uops_0_pc;
  wire [1:0] fp_pipeline_io_dis_uops_0_iqtype;
  wire [9:0] fp_pipeline_io_dis_uops_0_fu_code;
  wire  fp_pipeline_io_dis_uops_0_allocate_brtag;
  wire  fp_pipeline_io_dis_uops_0_is_br_or_jmp;
  wire  fp_pipeline_io_dis_uops_0_is_jump;
  wire  fp_pipeline_io_dis_uops_0_is_jal;
  wire  fp_pipeline_io_dis_uops_0_is_ret;
  wire  fp_pipeline_io_dis_uops_0_is_call;
  wire [7:0] fp_pipeline_io_dis_uops_0_br_mask;
  wire [2:0] fp_pipeline_io_dis_uops_0_br_tag;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_btb_blame;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_btb_hit;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_btb_taken;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_bpd_blame;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_bpd_hit;
  wire  fp_pipeline_io_dis_uops_0_br_prediction_bpd_taken;
  wire [1:0] fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_value;
  wire [5:0] fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_info;
  wire  fp_pipeline_io_dis_uops_0_stat_brjmp_mispredicted;
  wire  fp_pipeline_io_dis_uops_0_stat_btb_made_pred;
  wire  fp_pipeline_io_dis_uops_0_stat_btb_mispredicted;
  wire  fp_pipeline_io_dis_uops_0_stat_bpd_made_pred;
  wire  fp_pipeline_io_dis_uops_0_stat_bpd_mispredicted;
  wire [2:0] fp_pipeline_io_dis_uops_0_fetch_pc_lob;
  wire [19:0] fp_pipeline_io_dis_uops_0_imm_packed;
  wire [11:0] fp_pipeline_io_dis_uops_0_csr_addr;
  wire [6:0] fp_pipeline_io_dis_uops_0_rob_idx;
  wire [3:0] fp_pipeline_io_dis_uops_0_ldq_idx;
  wire [3:0] fp_pipeline_io_dis_uops_0_stq_idx;
  wire [5:0] fp_pipeline_io_dis_uops_0_brob_idx;
  wire [6:0] fp_pipeline_io_dis_uops_0_pdst;
  wire [6:0] fp_pipeline_io_dis_uops_0_pop1;
  wire [6:0] fp_pipeline_io_dis_uops_0_pop2;
  wire [6:0] fp_pipeline_io_dis_uops_0_pop3;
  wire  fp_pipeline_io_dis_uops_0_prs1_busy;
  wire  fp_pipeline_io_dis_uops_0_prs2_busy;
  wire  fp_pipeline_io_dis_uops_0_prs3_busy;
  wire [6:0] fp_pipeline_io_dis_uops_0_stale_pdst;
  wire  fp_pipeline_io_dis_uops_0_exception;
  wire [63:0] fp_pipeline_io_dis_uops_0_exc_cause;
  wire  fp_pipeline_io_dis_uops_0_bypassable;
  wire [4:0] fp_pipeline_io_dis_uops_0_mem_cmd;
  wire [2:0] fp_pipeline_io_dis_uops_0_mem_typ;
  wire  fp_pipeline_io_dis_uops_0_is_fence;
  wire  fp_pipeline_io_dis_uops_0_is_fencei;
  wire  fp_pipeline_io_dis_uops_0_is_store;
  wire  fp_pipeline_io_dis_uops_0_is_amo;
  wire  fp_pipeline_io_dis_uops_0_is_load;
  wire  fp_pipeline_io_dis_uops_0_is_sys_pc2epc;
  wire  fp_pipeline_io_dis_uops_0_is_unique;
  wire  fp_pipeline_io_dis_uops_0_flush_on_commit;
  wire [5:0] fp_pipeline_io_dis_uops_0_ldst;
  wire [5:0] fp_pipeline_io_dis_uops_0_lrs1;
  wire [5:0] fp_pipeline_io_dis_uops_0_lrs2;
  wire [5:0] fp_pipeline_io_dis_uops_0_lrs3;
  wire  fp_pipeline_io_dis_uops_0_ldst_val;
  wire [1:0] fp_pipeline_io_dis_uops_0_dst_rtype;
  wire [1:0] fp_pipeline_io_dis_uops_0_lrs1_rtype;
  wire [1:0] fp_pipeline_io_dis_uops_0_lrs2_rtype;
  wire  fp_pipeline_io_dis_uops_0_frs3_en;
  wire  fp_pipeline_io_dis_uops_0_fp_val;
  wire  fp_pipeline_io_dis_uops_0_fp_single;
  wire  fp_pipeline_io_dis_uops_0_xcpt_pf_if;
  wire  fp_pipeline_io_dis_uops_0_xcpt_ae_if;
  wire  fp_pipeline_io_dis_uops_0_replay_if;
  wire  fp_pipeline_io_dis_uops_0_xcpt_ma_if;
  wire [63:0] fp_pipeline_io_dis_uops_0_debug_wdata;
  wire [31:0] fp_pipeline_io_dis_uops_0_debug_events_fetch_seq;
  wire  fp_pipeline_io_dis_uops_1_valid;
  wire [8:0] fp_pipeline_io_dis_uops_1_uopc;
  wire [31:0] fp_pipeline_io_dis_uops_1_inst;
  wire [39:0] fp_pipeline_io_dis_uops_1_pc;
  wire [1:0] fp_pipeline_io_dis_uops_1_iqtype;
  wire [9:0] fp_pipeline_io_dis_uops_1_fu_code;
  wire  fp_pipeline_io_dis_uops_1_allocate_brtag;
  wire  fp_pipeline_io_dis_uops_1_is_br_or_jmp;
  wire  fp_pipeline_io_dis_uops_1_is_jump;
  wire  fp_pipeline_io_dis_uops_1_is_jal;
  wire  fp_pipeline_io_dis_uops_1_is_ret;
  wire  fp_pipeline_io_dis_uops_1_is_call;
  wire [7:0] fp_pipeline_io_dis_uops_1_br_mask;
  wire [2:0] fp_pipeline_io_dis_uops_1_br_tag;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_btb_blame;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_btb_hit;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_btb_taken;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_bpd_blame;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_bpd_hit;
  wire  fp_pipeline_io_dis_uops_1_br_prediction_bpd_taken;
  wire [1:0] fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_value;
  wire [5:0] fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_info;
  wire  fp_pipeline_io_dis_uops_1_stat_brjmp_mispredicted;
  wire  fp_pipeline_io_dis_uops_1_stat_btb_made_pred;
  wire  fp_pipeline_io_dis_uops_1_stat_btb_mispredicted;
  wire  fp_pipeline_io_dis_uops_1_stat_bpd_made_pred;
  wire  fp_pipeline_io_dis_uops_1_stat_bpd_mispredicted;
  wire [2:0] fp_pipeline_io_dis_uops_1_fetch_pc_lob;
  wire [19:0] fp_pipeline_io_dis_uops_1_imm_packed;
  wire [11:0] fp_pipeline_io_dis_uops_1_csr_addr;
  wire [6:0] fp_pipeline_io_dis_uops_1_rob_idx;
  wire [3:0] fp_pipeline_io_dis_uops_1_ldq_idx;
  wire [3:0] fp_pipeline_io_dis_uops_1_stq_idx;
  wire [5:0] fp_pipeline_io_dis_uops_1_brob_idx;
  wire [6:0] fp_pipeline_io_dis_uops_1_pdst;
  wire [6:0] fp_pipeline_io_dis_uops_1_pop1;
  wire [6:0] fp_pipeline_io_dis_uops_1_pop2;
  wire [6:0] fp_pipeline_io_dis_uops_1_pop3;
  wire  fp_pipeline_io_dis_uops_1_prs1_busy;
  wire  fp_pipeline_io_dis_uops_1_prs2_busy;
  wire  fp_pipeline_io_dis_uops_1_prs3_busy;
  wire [6:0] fp_pipeline_io_dis_uops_1_stale_pdst;
  wire  fp_pipeline_io_dis_uops_1_exception;
  wire [63:0] fp_pipeline_io_dis_uops_1_exc_cause;
  wire  fp_pipeline_io_dis_uops_1_bypassable;
  wire [4:0] fp_pipeline_io_dis_uops_1_mem_cmd;
  wire [2:0] fp_pipeline_io_dis_uops_1_mem_typ;
  wire  fp_pipeline_io_dis_uops_1_is_fence;
  wire  fp_pipeline_io_dis_uops_1_is_fencei;
  wire  fp_pipeline_io_dis_uops_1_is_store;
  wire  fp_pipeline_io_dis_uops_1_is_amo;
  wire  fp_pipeline_io_dis_uops_1_is_load;
  wire  fp_pipeline_io_dis_uops_1_is_sys_pc2epc;
  wire  fp_pipeline_io_dis_uops_1_is_unique;
  wire  fp_pipeline_io_dis_uops_1_flush_on_commit;
  wire [5:0] fp_pipeline_io_dis_uops_1_ldst;
  wire [5:0] fp_pipeline_io_dis_uops_1_lrs1;
  wire [5:0] fp_pipeline_io_dis_uops_1_lrs2;
  wire [5:0] fp_pipeline_io_dis_uops_1_lrs3;
  wire  fp_pipeline_io_dis_uops_1_ldst_val;
  wire [1:0] fp_pipeline_io_dis_uops_1_dst_rtype;
  wire [1:0] fp_pipeline_io_dis_uops_1_lrs1_rtype;
  wire [1:0] fp_pipeline_io_dis_uops_1_lrs2_rtype;
  wire  fp_pipeline_io_dis_uops_1_frs3_en;
  wire  fp_pipeline_io_dis_uops_1_fp_val;
  wire  fp_pipeline_io_dis_uops_1_fp_single;
  wire  fp_pipeline_io_dis_uops_1_xcpt_pf_if;
  wire  fp_pipeline_io_dis_uops_1_xcpt_ae_if;
  wire  fp_pipeline_io_dis_uops_1_replay_if;
  wire  fp_pipeline_io_dis_uops_1_xcpt_ma_if;
  wire [63:0] fp_pipeline_io_dis_uops_1_debug_wdata;
  wire [31:0] fp_pipeline_io_dis_uops_1_debug_events_fetch_seq;
  wire  fp_pipeline_io_dis_readys_0;
  wire  fp_pipeline_io_dis_readys_1;
  wire  fp_pipeline_io_ll_wport_valid;
  wire [6:0] fp_pipeline_io_ll_wport_bits_uop_rob_idx;
  wire [6:0] fp_pipeline_io_ll_wport_bits_uop_pdst;
  wire [2:0] fp_pipeline_io_ll_wport_bits_uop_mem_typ;
  wire [1:0] fp_pipeline_io_ll_wport_bits_uop_dst_rtype;
  wire  fp_pipeline_io_ll_wport_bits_uop_fp_val;
  wire [64:0] fp_pipeline_io_ll_wport_bits_data;
  wire  fp_pipeline_io_fromint_valid;
  wire [8:0] fp_pipeline_io_fromint_bits_uop_uopc;
  wire  fp_pipeline_io_fromint_bits_uop_ctrl_rf_wen;
  wire [7:0] fp_pipeline_io_fromint_bits_uop_br_mask;
  wire [19:0] fp_pipeline_io_fromint_bits_uop_imm_packed;
  wire [6:0] fp_pipeline_io_fromint_bits_uop_rob_idx;
  wire [6:0] fp_pipeline_io_fromint_bits_uop_pdst;
  wire [1:0] fp_pipeline_io_fromint_bits_uop_dst_rtype;
  wire  fp_pipeline_io_fromint_bits_uop_fp_val;
  wire [64:0] fp_pipeline_io_fromint_bits_rs1_data;
  wire  fp_pipeline_io_tosdq_valid;
  wire [7:0] fp_pipeline_io_tosdq_bits_uop_br_mask;
  wire [6:0] fp_pipeline_io_tosdq_bits_uop_rob_idx;
  wire [3:0] fp_pipeline_io_tosdq_bits_uop_stq_idx;
  wire  fp_pipeline_io_tosdq_bits_uop_is_amo;
  wire [63:0] fp_pipeline_io_tosdq_bits_data;
  wire  fp_pipeline_io_toint_ready;
  wire  fp_pipeline_io_toint_valid;
  wire [6:0] fp_pipeline_io_toint_bits_uop_rob_idx;
  wire [6:0] fp_pipeline_io_toint_bits_uop_pdst;
  wire  fp_pipeline_io_toint_bits_uop_is_store;
  wire  fp_pipeline_io_toint_bits_uop_is_amo;
  wire [1:0] fp_pipeline_io_toint_bits_uop_dst_rtype;
  wire [63:0] fp_pipeline_io_toint_bits_data;
  wire  fp_pipeline_io_wakeups_0_valid;
  wire [6:0] fp_pipeline_io_wakeups_0_bits_uop_rob_idx;
  wire [6:0] fp_pipeline_io_wakeups_0_bits_uop_pdst;
  wire [1:0] fp_pipeline_io_wakeups_0_bits_uop_dst_rtype;
  wire  fp_pipeline_io_wakeups_0_bits_uop_fp_val;
  wire  fp_pipeline_io_wakeups_0_bits_fflags_valid;
  wire [6:0] fp_pipeline_io_wakeups_0_bits_fflags_bits_uop_rob_idx;
  wire [4:0] fp_pipeline_io_wakeups_0_bits_fflags_bits_flags;
  wire  fp_pipeline_io_wakeups_1_valid;
  wire [6:0] fp_pipeline_io_wakeups_1_bits_uop_rob_idx;
  wire [6:0] fp_pipeline_io_wakeups_1_bits_uop_pdst;
  wire [1:0] fp_pipeline_io_wakeups_1_bits_uop_dst_rtype;
  wire  fp_pipeline_io_wakeups_1_bits_uop_fp_val;
  wire  fp_pipeline_io_wakeups_1_bits_fflags_valid;
  wire [6:0] fp_pipeline_io_wakeups_1_bits_fflags_bits_uop_rob_idx;
  wire [4:0] fp_pipeline_io_wakeups_1_bits_fflags_bits_flags;
  wire  fetch_unit_clock;
  wire  fetch_unit_reset;
  wire  fetch_unit_io_imem_req_valid;
  wire [39:0] fetch_unit_io_imem_req_bits_pc;
  wire  fetch_unit_io_imem_req_bits_speculative;
  wire  fetch_unit_io_imem_resp_ready;
  wire  fetch_unit_io_imem_resp_valid;
  wire [39:0] fetch_unit_io_imem_resp_bits_pc;
  wire [63:0] fetch_unit_io_imem_resp_bits_data;
  wire [1:0] fetch_unit_io_imem_resp_bits_mask;
  wire  fetch_unit_io_imem_resp_bits_xcpt_pf_inst;
  wire  fetch_unit_io_imem_resp_bits_xcpt_ae_inst;
  wire  fetch_unit_io_imem_resp_bits_replay;
  wire [1:0] fetch_unit_io_f2_btb_resp_bits_bim_resp_value;
  wire [5:0] fetch_unit_io_f2_btb_resp_bits_bim_resp_entry_idx;
  wire [1:0] fetch_unit_io_f2_btb_resp_bits_bim_resp_way_idx;
  wire [1:0] fetch_unit_io_f2_bpd_resp_bits_takens;
  wire [14:0] fetch_unit_io_f2_bpd_resp_bits_info;
  wire [14:0] fetch_unit_io_f3_bpd_resp_bits_history;
  wire [7:0] fetch_unit_io_f3_bpd_resp_bits_history_ptr;
  wire  fetch_unit_io_f3_btb_update_valid;
  wire [38:0] fetch_unit_io_f3_btb_update_bits_pc;
  wire [38:0] fetch_unit_io_f3_btb_update_bits_target;
  wire [38:0] fetch_unit_io_f3_btb_update_bits_cfi_pc;
  wire [2:0] fetch_unit_io_f3_btb_update_bits_bpd_type;
  wire [2:0] fetch_unit_io_f3_btb_update_bits_cfi_type;
  wire  fetch_unit_io_f3_hist_update_valid;
  wire  fetch_unit_io_f3_hist_update_bits_taken;
  wire  fetch_unit_io_f3_bim_update_valid;
  wire  fetch_unit_io_f3_bim_update_bits_taken;
  wire [1:0] fetch_unit_io_f3_bim_update_bits_bim_resp_value;
  wire [5:0] fetch_unit_io_f3_bim_update_bits_bim_resp_entry_idx;
  wire [1:0] fetch_unit_io_f3_bim_update_bits_bim_resp_way_idx;
  wire  fetch_unit_io_br_unit_take_pc;
  wire [39:0] fetch_unit_io_br_unit_target;
  wire  fetch_unit_io_clear_fetchbuffer;
  wire  fetch_unit_io_flush_take_pc;
  wire [39:0] fetch_unit_io_flush_pc;
  wire  fetch_unit_io_sfence_take_pc;
  wire [39:0] fetch_unit_io_sfence_addr;
  wire  fetch_unit_io_resp_ready;
  wire  fetch_unit_io_resp_valid;
  wire [39:0] fetch_unit_io_resp_bits_pc;
  wire [31:0] fetch_unit_io_resp_bits_insts_0;
  wire [31:0] fetch_unit_io_resp_bits_insts_1;
  wire [1:0] fetch_unit_io_resp_bits_mask;
  wire  fetch_unit_io_resp_bits_xcpt_pf_if;
  wire  fetch_unit_io_resp_bits_xcpt_ae_if;
  wire  fetch_unit_io_resp_bits_replay_if;
  wire [1:0] fetch_unit_io_resp_bits_xcpt_ma_if_oh;
  wire  fetch_unit_io_resp_bits_bpu_info_0_btb_blame;
  wire  fetch_unit_io_resp_bits_bpu_info_0_btb_hit;
  wire  fetch_unit_io_resp_bits_bpu_info_0_btb_taken;
  wire  fetch_unit_io_resp_bits_bpu_info_0_bpd_blame;
  wire  fetch_unit_io_resp_bits_bpu_info_0_bpd_hit;
  wire  fetch_unit_io_resp_bits_bpu_info_0_bpd_taken;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_0_bim_resp_value;
  wire [5:0] fetch_unit_io_resp_bits_bpu_info_0_bim_resp_entry_idx;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_0_bim_resp_way_idx;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_takens;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_u;
  wire [7:0] fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_ptr;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_info;
  wire  fetch_unit_io_resp_bits_bpu_info_1_btb_blame;
  wire  fetch_unit_io_resp_bits_bpu_info_1_btb_hit;
  wire  fetch_unit_io_resp_bits_bpu_info_1_btb_taken;
  wire  fetch_unit_io_resp_bits_bpu_info_1_bpd_blame;
  wire  fetch_unit_io_resp_bits_bpu_info_1_bpd_hit;
  wire  fetch_unit_io_resp_bits_bpu_info_1_bpd_taken;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_1_bim_resp_value;
  wire [5:0] fetch_unit_io_resp_bits_bpu_info_1_bim_resp_entry_idx;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_1_bim_resp_way_idx;
  wire [1:0] fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_takens;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_u;
  wire [7:0] fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_ptr;
  wire [14:0] fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_info;
  wire [31:0] fetch_unit_io_resp_bits_debug_events_0_fetch_seq;
  wire [31:0] fetch_unit_io_resp_bits_debug_events_1_fetch_seq;
  wire  fetch_unit_io_stalled;
  wire  bpd_stage_clock;
  wire  bpd_stage_reset;
  wire  bpd_stage_io_fetch_stalled;
  wire [1:0] bpd_stage_io_f2_btb_resp_bits_bim_resp_value;
  wire [5:0] bpd_stage_io_f2_btb_resp_bits_bim_resp_entry_idx;
  wire [1:0] bpd_stage_io_f2_btb_resp_bits_bim_resp_way_idx;
  wire [1:0] bpd_stage_io_f2_bpd_resp_bits_takens;
  wire [14:0] bpd_stage_io_f2_bpd_resp_bits_info;
  wire [14:0] bpd_stage_io_f3_bpd_resp_bits_history;
  wire [7:0] bpd_stage_io_f3_bpd_resp_bits_history_ptr;
  wire  bpd_stage_io_f3_btb_update_valid;
  wire [38:0] bpd_stage_io_f3_btb_update_bits_pc;
  wire [38:0] bpd_stage_io_f3_btb_update_bits_target;
  wire [38:0] bpd_stage_io_f3_btb_update_bits_cfi_pc;
  wire [2:0] bpd_stage_io_f3_btb_update_bits_bpd_type;
  wire [2:0] bpd_stage_io_f3_btb_update_bits_cfi_type;
  wire  bpd_stage_io_f3_hist_update_valid;
  wire  bpd_stage_io_f3_hist_update_bits_taken;
  wire  bpd_stage_io_f3_bim_update_valid;
  wire  bpd_stage_io_f3_bim_update_bits_taken;
  wire [1:0] bpd_stage_io_f3_bim_update_bits_bim_resp_value;
  wire [5:0] bpd_stage_io_f3_bim_update_bits_bim_resp_entry_idx;
  wire [1:0] bpd_stage_io_f3_bim_update_bits_bim_resp_way_idx;
  wire  bpd_stage_io_br_unit_btb_update_valid;
  wire [38:0] bpd_stage_io_br_unit_btb_update_bits_pc;
  wire [38:0] bpd_stage_io_br_unit_btb_update_bits_target;
  wire [38:0] bpd_stage_io_br_unit_btb_update_bits_cfi_pc;
  wire [2:0] bpd_stage_io_br_unit_btb_update_bits_bpd_type;
  wire [2:0] bpd_stage_io_br_unit_btb_update_bits_cfi_type;
  wire  bpd_stage_io_br_unit_bim_update_valid;
  wire  bpd_stage_io_br_unit_bim_update_bits_taken;
  wire [1:0] bpd_stage_io_br_unit_bim_update_bits_bim_resp_value;
  wire [5:0] bpd_stage_io_br_unit_bim_update_bits_bim_resp_entry_idx;
  wire [1:0] bpd_stage_io_br_unit_bim_update_bits_bim_resp_way_idx;
  wire  bpd_stage_io_br_unit_bpd_update_valid;
  wire  bpd_stage_io_br_unit_bpd_update_bits_mispredict;
  wire [14:0] bpd_stage_io_br_unit_bpd_update_bits_history;
  wire [7:0] bpd_stage_io_br_unit_bpd_update_bits_history_ptr;
  wire  bpd_stage_io_br_unit_bpd_update_bits_bpd_mispredict;
  wire  bpd_stage_io_br_unit_bpd_update_bits_taken;
  wire  bpd_stage_io_br_unit_bpd_update_bits_new_pc_same_packet;
  wire  bpd_stage_io_brob_allocate_ready;
  wire  bpd_stage_io_brob_allocate_valid;
  wire [5:0] bpd_stage_io_brob_allocate_bits_ctrl_brob_idx;
  wire [14:0] bpd_stage_io_brob_allocate_bits_info_info;
  wire [5:0] bpd_stage_io_brob_allocate_brob_tail;
  wire  bpd_stage_io_brob_deallocate_valid;
  wire [5:0] bpd_stage_io_brob_deallocate_bits_brob_idx;
  wire  bpd_stage_io_brob_bpd_update_valid;
  wire [2:0] bpd_stage_io_brob_bpd_update_bits_br_pc;
  wire [5:0] bpd_stage_io_brob_bpd_update_bits_brob_idx;
  wire  bpd_stage_io_brob_bpd_update_bits_mispredict;
  wire  bpd_stage_io_brob_bpd_update_bits_bpd_predict_val;
  wire  bpd_stage_io_brob_bpd_update_bits_bpd_mispredict;
  wire  bpd_stage_io_brob_bpd_update_bits_taken;
  wire  bpd_stage_io_brob_bpd_update_bits_is_br;
  wire  bpd_stage_io_brob_flush;
  wire  bpd_stage_io_flush;
  wire  bpd_stage_io_redirect;
  wire  bpd_stage_io_status_debug;
  wire  dec_serializer_io_enq_ready;
  wire  dec_serializer_io_enq_valid;
  wire [39:0] dec_serializer_io_enq_bits_pc;
  wire [31:0] dec_serializer_io_enq_bits_insts_0;
  wire [31:0] dec_serializer_io_enq_bits_insts_1;
  wire [1:0] dec_serializer_io_enq_bits_mask;
  wire  dec_serializer_io_enq_bits_xcpt_pf_if;
  wire  dec_serializer_io_enq_bits_xcpt_ae_if;
  wire  dec_serializer_io_enq_bits_replay_if;
  wire [1:0] dec_serializer_io_enq_bits_xcpt_ma_if_oh;
  wire  dec_serializer_io_enq_bits_bpu_info_0_btb_blame;
  wire  dec_serializer_io_enq_bits_bpu_info_0_btb_hit;
  wire  dec_serializer_io_enq_bits_bpu_info_0_btb_taken;
  wire  dec_serializer_io_enq_bits_bpu_info_0_bpd_blame;
  wire  dec_serializer_io_enq_bits_bpu_info_0_bpd_hit;
  wire  dec_serializer_io_enq_bits_bpu_info_0_bpd_taken;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_0_bim_resp_value;
  wire [5:0] dec_serializer_io_enq_bits_bpu_info_0_bim_resp_entry_idx;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_0_bim_resp_way_idx;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_takens;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_u;
  wire [7:0] dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_ptr;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_info;
  wire  dec_serializer_io_enq_bits_bpu_info_1_btb_blame;
  wire  dec_serializer_io_enq_bits_bpu_info_1_btb_hit;
  wire  dec_serializer_io_enq_bits_bpu_info_1_btb_taken;
  wire  dec_serializer_io_enq_bits_bpu_info_1_bpd_blame;
  wire  dec_serializer_io_enq_bits_bpu_info_1_bpd_hit;
  wire  dec_serializer_io_enq_bits_bpu_info_1_bpd_taken;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_1_bim_resp_value;
  wire [5:0] dec_serializer_io_enq_bits_bpu_info_1_bim_resp_entry_idx;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_1_bim_resp_way_idx;
  wire [1:0] dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_takens;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_u;
  wire [7:0] dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_ptr;
  wire [14:0] dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_info;
  wire [31:0] dec_serializer_io_enq_bits_debug_events_0_fetch_seq;
  wire [31:0] dec_serializer_io_enq_bits_debug_events_1_fetch_seq;
  wire  dec_serializer_io_deq_ready;
  wire  dec_serializer_io_deq_valid;
  wire  dec_serializer_io_deq_bits_uops_0_valid;
  wire [31:0] dec_serializer_io_deq_bits_uops_0_inst;
  wire [39:0] dec_serializer_io_deq_bits_uops_0_pc;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_btb_blame;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_btb_hit;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_btb_taken;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_blame;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_hit;
  wire  dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_taken;
  wire [1:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_value;
  wire [5:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_info;
  wire [2:0] dec_serializer_io_deq_bits_uops_0_fetch_pc_lob;
  wire  dec_serializer_io_deq_bits_uops_0_xcpt_pf_if;
  wire  dec_serializer_io_deq_bits_uops_0_xcpt_ae_if;
  wire  dec_serializer_io_deq_bits_uops_0_replay_if;
  wire  dec_serializer_io_deq_bits_uops_0_xcpt_ma_if;
  wire [31:0] dec_serializer_io_deq_bits_uops_0_debug_events_fetch_seq;
  wire  dec_serializer_io_deq_bits_uops_1_valid;
  wire [31:0] dec_serializer_io_deq_bits_uops_1_inst;
  wire [39:0] dec_serializer_io_deq_bits_uops_1_pc;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_btb_blame;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_btb_hit;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_btb_taken;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_blame;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_hit;
  wire  dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_taken;
  wire [1:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_value;
  wire [5:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_info;
  wire [2:0] dec_serializer_io_deq_bits_uops_1_fetch_pc_lob;
  wire  dec_serializer_io_deq_bits_uops_1_xcpt_pf_if;
  wire  dec_serializer_io_deq_bits_uops_1_xcpt_ae_if;
  wire  dec_serializer_io_deq_bits_uops_1_replay_if;
  wire  dec_serializer_io_deq_bits_uops_1_xcpt_ma_if;
  wire [31:0] dec_serializer_io_deq_bits_uops_1_debug_events_fetch_seq;
  wire [14:0] dec_serializer_io_deq_bits_bpd_resp_info;
  wire  decode_units_0_io_enq_uop_valid;
  wire [31:0] decode_units_0_io_enq_uop_inst;
  wire [39:0] decode_units_0_io_enq_uop_pc;
  wire  decode_units_0_io_enq_uop_br_prediction_btb_blame;
  wire  decode_units_0_io_enq_uop_br_prediction_btb_hit;
  wire  decode_units_0_io_enq_uop_br_prediction_btb_taken;
  wire  decode_units_0_io_enq_uop_br_prediction_bpd_blame;
  wire  decode_units_0_io_enq_uop_br_prediction_bpd_hit;
  wire  decode_units_0_io_enq_uop_br_prediction_bpd_taken;
  wire [1:0] decode_units_0_io_enq_uop_br_prediction_bim_resp_value;
  wire [5:0] decode_units_0_io_enq_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] decode_units_0_io_enq_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] decode_units_0_io_enq_uop_br_prediction_bpd_resp_takens;
  wire [14:0] decode_units_0_io_enq_uop_br_prediction_bpd_resp_history;
  wire [14:0] decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] decode_units_0_io_enq_uop_br_prediction_bpd_resp_info;
  wire [2:0] decode_units_0_io_enq_uop_fetch_pc_lob;
  wire  decode_units_0_io_enq_uop_xcpt_pf_if;
  wire  decode_units_0_io_enq_uop_xcpt_ae_if;
  wire  decode_units_0_io_enq_uop_replay_if;
  wire  decode_units_0_io_enq_uop_xcpt_ma_if;
  wire [31:0] decode_units_0_io_enq_uop_debug_events_fetch_seq;
  wire  decode_units_0_io_deq_uop_valid;
  wire [8:0] decode_units_0_io_deq_uop_uopc;
  wire [31:0] decode_units_0_io_deq_uop_inst;
  wire [39:0] decode_units_0_io_deq_uop_pc;
  wire [1:0] decode_units_0_io_deq_uop_iqtype;
  wire [9:0] decode_units_0_io_deq_uop_fu_code;
  wire  decode_units_0_io_deq_uop_allocate_brtag;
  wire  decode_units_0_io_deq_uop_is_br_or_jmp;
  wire  decode_units_0_io_deq_uop_is_jump;
  wire  decode_units_0_io_deq_uop_is_jal;
  wire  decode_units_0_io_deq_uop_is_ret;
  wire  decode_units_0_io_deq_uop_is_call;
  wire  decode_units_0_io_deq_uop_br_prediction_btb_blame;
  wire  decode_units_0_io_deq_uop_br_prediction_btb_hit;
  wire  decode_units_0_io_deq_uop_br_prediction_btb_taken;
  wire  decode_units_0_io_deq_uop_br_prediction_bpd_blame;
  wire  decode_units_0_io_deq_uop_br_prediction_bpd_hit;
  wire  decode_units_0_io_deq_uop_br_prediction_bpd_taken;
  wire [1:0] decode_units_0_io_deq_uop_br_prediction_bim_resp_value;
  wire [5:0] decode_units_0_io_deq_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] decode_units_0_io_deq_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] decode_units_0_io_deq_uop_br_prediction_bpd_resp_takens;
  wire [14:0] decode_units_0_io_deq_uop_br_prediction_bpd_resp_history;
  wire [14:0] decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] decode_units_0_io_deq_uop_br_prediction_bpd_resp_info;
  wire [2:0] decode_units_0_io_deq_uop_fetch_pc_lob;
  wire [19:0] decode_units_0_io_deq_uop_imm_packed;
  wire  decode_units_0_io_deq_uop_exception;
  wire [63:0] decode_units_0_io_deq_uop_exc_cause;
  wire  decode_units_0_io_deq_uop_bypassable;
  wire [4:0] decode_units_0_io_deq_uop_mem_cmd;
  wire [2:0] decode_units_0_io_deq_uop_mem_typ;
  wire  decode_units_0_io_deq_uop_is_fence;
  wire  decode_units_0_io_deq_uop_is_fencei;
  wire  decode_units_0_io_deq_uop_is_store;
  wire  decode_units_0_io_deq_uop_is_amo;
  wire  decode_units_0_io_deq_uop_is_load;
  wire  decode_units_0_io_deq_uop_is_sys_pc2epc;
  wire  decode_units_0_io_deq_uop_is_unique;
  wire  decode_units_0_io_deq_uop_flush_on_commit;
  wire [5:0] decode_units_0_io_deq_uop_ldst;
  wire [5:0] decode_units_0_io_deq_uop_lrs1;
  wire [5:0] decode_units_0_io_deq_uop_lrs2;
  wire [5:0] decode_units_0_io_deq_uop_lrs3;
  wire  decode_units_0_io_deq_uop_ldst_val;
  wire [1:0] decode_units_0_io_deq_uop_dst_rtype;
  wire [1:0] decode_units_0_io_deq_uop_lrs1_rtype;
  wire [1:0] decode_units_0_io_deq_uop_lrs2_rtype;
  wire  decode_units_0_io_deq_uop_frs3_en;
  wire  decode_units_0_io_deq_uop_fp_val;
  wire  decode_units_0_io_deq_uop_fp_single;
  wire  decode_units_0_io_deq_uop_xcpt_pf_if;
  wire  decode_units_0_io_deq_uop_xcpt_ae_if;
  wire  decode_units_0_io_deq_uop_replay_if;
  wire  decode_units_0_io_deq_uop_xcpt_ma_if;
  wire [31:0] decode_units_0_io_deq_uop_debug_events_fetch_seq;
  wire [31:0] decode_units_0_io_status_isa;
  wire [11:0] decode_units_0_io_csr_decode_csr;
  wire  decode_units_0_io_csr_decode_fp_illegal;
  wire  decode_units_0_io_csr_decode_read_illegal;
  wire  decode_units_0_io_csr_decode_write_illegal;
  wire  decode_units_0_io_csr_decode_write_flush;
  wire  decode_units_0_io_csr_decode_system_illegal;
  wire  decode_units_0_io_interrupt;
  wire [63:0] decode_units_0_io_interrupt_cause;
  wire  decode_units_1_io_enq_uop_valid;
  wire [31:0] decode_units_1_io_enq_uop_inst;
  wire [39:0] decode_units_1_io_enq_uop_pc;
  wire  decode_units_1_io_enq_uop_br_prediction_btb_blame;
  wire  decode_units_1_io_enq_uop_br_prediction_btb_hit;
  wire  decode_units_1_io_enq_uop_br_prediction_btb_taken;
  wire  decode_units_1_io_enq_uop_br_prediction_bpd_blame;
  wire  decode_units_1_io_enq_uop_br_prediction_bpd_hit;
  wire  decode_units_1_io_enq_uop_br_prediction_bpd_taken;
  wire [1:0] decode_units_1_io_enq_uop_br_prediction_bim_resp_value;
  wire [5:0] decode_units_1_io_enq_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] decode_units_1_io_enq_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] decode_units_1_io_enq_uop_br_prediction_bpd_resp_takens;
  wire [14:0] decode_units_1_io_enq_uop_br_prediction_bpd_resp_history;
  wire [14:0] decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] decode_units_1_io_enq_uop_br_prediction_bpd_resp_info;
  wire [2:0] decode_units_1_io_enq_uop_fetch_pc_lob;
  wire  decode_units_1_io_enq_uop_xcpt_pf_if;
  wire  decode_units_1_io_enq_uop_xcpt_ae_if;
  wire  decode_units_1_io_enq_uop_replay_if;
  wire  decode_units_1_io_enq_uop_xcpt_ma_if;
  wire [31:0] decode_units_1_io_enq_uop_debug_events_fetch_seq;
  wire  decode_units_1_io_deq_uop_valid;
  wire [8:0] decode_units_1_io_deq_uop_uopc;
  wire [31:0] decode_units_1_io_deq_uop_inst;
  wire [39:0] decode_units_1_io_deq_uop_pc;
  wire [1:0] decode_units_1_io_deq_uop_iqtype;
  wire [9:0] decode_units_1_io_deq_uop_fu_code;
  wire  decode_units_1_io_deq_uop_allocate_brtag;
  wire  decode_units_1_io_deq_uop_is_br_or_jmp;
  wire  decode_units_1_io_deq_uop_is_jump;
  wire  decode_units_1_io_deq_uop_is_jal;
  wire  decode_units_1_io_deq_uop_is_ret;
  wire  decode_units_1_io_deq_uop_is_call;
  wire  decode_units_1_io_deq_uop_br_prediction_btb_blame;
  wire  decode_units_1_io_deq_uop_br_prediction_btb_hit;
  wire  decode_units_1_io_deq_uop_br_prediction_btb_taken;
  wire  decode_units_1_io_deq_uop_br_prediction_bpd_blame;
  wire  decode_units_1_io_deq_uop_br_prediction_bpd_hit;
  wire  decode_units_1_io_deq_uop_br_prediction_bpd_taken;
  wire [1:0] decode_units_1_io_deq_uop_br_prediction_bim_resp_value;
  wire [5:0] decode_units_1_io_deq_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] decode_units_1_io_deq_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] decode_units_1_io_deq_uop_br_prediction_bpd_resp_takens;
  wire [14:0] decode_units_1_io_deq_uop_br_prediction_bpd_resp_history;
  wire [14:0] decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] decode_units_1_io_deq_uop_br_prediction_bpd_resp_info;
  wire [2:0] decode_units_1_io_deq_uop_fetch_pc_lob;
  wire [19:0] decode_units_1_io_deq_uop_imm_packed;
  wire  decode_units_1_io_deq_uop_exception;
  wire [63:0] decode_units_1_io_deq_uop_exc_cause;
  wire  decode_units_1_io_deq_uop_bypassable;
  wire [4:0] decode_units_1_io_deq_uop_mem_cmd;
  wire [2:0] decode_units_1_io_deq_uop_mem_typ;
  wire  decode_units_1_io_deq_uop_is_fence;
  wire  decode_units_1_io_deq_uop_is_fencei;
  wire  decode_units_1_io_deq_uop_is_store;
  wire  decode_units_1_io_deq_uop_is_amo;
  wire  decode_units_1_io_deq_uop_is_load;
  wire  decode_units_1_io_deq_uop_is_sys_pc2epc;
  wire  decode_units_1_io_deq_uop_is_unique;
  wire  decode_units_1_io_deq_uop_flush_on_commit;
  wire [5:0] decode_units_1_io_deq_uop_ldst;
  wire [5:0] decode_units_1_io_deq_uop_lrs1;
  wire [5:0] decode_units_1_io_deq_uop_lrs2;
  wire [5:0] decode_units_1_io_deq_uop_lrs3;
  wire  decode_units_1_io_deq_uop_ldst_val;
  wire [1:0] decode_units_1_io_deq_uop_dst_rtype;
  wire [1:0] decode_units_1_io_deq_uop_lrs1_rtype;
  wire [1:0] decode_units_1_io_deq_uop_lrs2_rtype;
  wire  decode_units_1_io_deq_uop_frs3_en;
  wire  decode_units_1_io_deq_uop_fp_val;
  wire  decode_units_1_io_deq_uop_fp_single;
  wire  decode_units_1_io_deq_uop_xcpt_pf_if;
  wire  decode_units_1_io_deq_uop_xcpt_ae_if;
  wire  decode_units_1_io_deq_uop_replay_if;
  wire  decode_units_1_io_deq_uop_xcpt_ma_if;
  wire [31:0] decode_units_1_io_deq_uop_debug_events_fetch_seq;
  wire [31:0] decode_units_1_io_status_isa;
  wire [11:0] decode_units_1_io_csr_decode_csr;
  wire  decode_units_1_io_csr_decode_fp_illegal;
  wire  decode_units_1_io_csr_decode_read_illegal;
  wire  decode_units_1_io_csr_decode_write_illegal;
  wire  decode_units_1_io_csr_decode_write_flush;
  wire  decode_units_1_io_csr_decode_system_illegal;
  wire  decode_units_1_io_interrupt;
  wire [63:0] decode_units_1_io_interrupt_cause;
  wire  dec_brmask_logic_clock;
  wire  dec_brmask_logic_reset;
  wire  dec_brmask_logic_io_is_branch_0;
  wire  dec_brmask_logic_io_is_branch_1;
  wire  dec_brmask_logic_io_will_fire_0;
  wire  dec_brmask_logic_io_will_fire_1;
  wire [2:0] dec_brmask_logic_io_br_tag_0;
  wire [2:0] dec_brmask_logic_io_br_tag_1;
  wire [7:0] dec_brmask_logic_io_br_mask_0;
  wire [7:0] dec_brmask_logic_io_br_mask_1;
  wire  dec_brmask_logic_io_is_full_0;
  wire  dec_brmask_logic_io_is_full_1;
  wire  dec_brmask_logic_io_brinfo_valid;
  wire  dec_brmask_logic_io_brinfo_mispredict;
  wire [7:0] dec_brmask_logic_io_brinfo_mask;
  wire [7:0] dec_brmask_logic_io_brinfo_exe_mask;
  wire  dec_brmask_logic_io_flush_pipeline;
  wire  rename_stage_clock;
  wire  rename_stage_reset;
  wire  rename_stage_io_inst_can_proceed_0;
  wire  rename_stage_io_inst_can_proceed_1;
  wire  rename_stage_io_kill;
  wire  rename_stage_io_dec_will_fire_0;
  wire  rename_stage_io_dec_will_fire_1;
  wire  rename_stage_io_dec_uops_0_valid;
  wire [8:0] rename_stage_io_dec_uops_0_uopc;
  wire [31:0] rename_stage_io_dec_uops_0_inst;
  wire [39:0] rename_stage_io_dec_uops_0_pc;
  wire [1:0] rename_stage_io_dec_uops_0_iqtype;
  wire [9:0] rename_stage_io_dec_uops_0_fu_code;
  wire  rename_stage_io_dec_uops_0_allocate_brtag;
  wire  rename_stage_io_dec_uops_0_is_br_or_jmp;
  wire  rename_stage_io_dec_uops_0_is_jump;
  wire  rename_stage_io_dec_uops_0_is_jal;
  wire  rename_stage_io_dec_uops_0_is_ret;
  wire  rename_stage_io_dec_uops_0_is_call;
  wire [7:0] rename_stage_io_dec_uops_0_br_mask;
  wire [2:0] rename_stage_io_dec_uops_0_br_tag;
  wire  rename_stage_io_dec_uops_0_br_prediction_btb_blame;
  wire  rename_stage_io_dec_uops_0_br_prediction_btb_hit;
  wire  rename_stage_io_dec_uops_0_br_prediction_btb_taken;
  wire  rename_stage_io_dec_uops_0_br_prediction_bpd_blame;
  wire  rename_stage_io_dec_uops_0_br_prediction_bpd_hit;
  wire  rename_stage_io_dec_uops_0_br_prediction_bpd_taken;
  wire [1:0] rename_stage_io_dec_uops_0_br_prediction_bim_resp_value;
  wire [5:0] rename_stage_io_dec_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_dec_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] rename_stage_io_dec_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] rename_stage_io_dec_uops_0_br_prediction_bpd_resp_info;
  wire [2:0] rename_stage_io_dec_uops_0_fetch_pc_lob;
  wire [19:0] rename_stage_io_dec_uops_0_imm_packed;
  wire [6:0] rename_stage_io_dec_uops_0_rob_idx;
  wire [3:0] rename_stage_io_dec_uops_0_ldq_idx;
  wire [3:0] rename_stage_io_dec_uops_0_stq_idx;
  wire [5:0] rename_stage_io_dec_uops_0_brob_idx;
  wire  rename_stage_io_dec_uops_0_exception;
  wire [63:0] rename_stage_io_dec_uops_0_exc_cause;
  wire  rename_stage_io_dec_uops_0_bypassable;
  wire [4:0] rename_stage_io_dec_uops_0_mem_cmd;
  wire [2:0] rename_stage_io_dec_uops_0_mem_typ;
  wire  rename_stage_io_dec_uops_0_is_fence;
  wire  rename_stage_io_dec_uops_0_is_fencei;
  wire  rename_stage_io_dec_uops_0_is_store;
  wire  rename_stage_io_dec_uops_0_is_amo;
  wire  rename_stage_io_dec_uops_0_is_load;
  wire  rename_stage_io_dec_uops_0_is_sys_pc2epc;
  wire  rename_stage_io_dec_uops_0_is_unique;
  wire  rename_stage_io_dec_uops_0_flush_on_commit;
  wire [5:0] rename_stage_io_dec_uops_0_ldst;
  wire [5:0] rename_stage_io_dec_uops_0_lrs1;
  wire [5:0] rename_stage_io_dec_uops_0_lrs2;
  wire [5:0] rename_stage_io_dec_uops_0_lrs3;
  wire  rename_stage_io_dec_uops_0_ldst_val;
  wire [1:0] rename_stage_io_dec_uops_0_dst_rtype;
  wire [1:0] rename_stage_io_dec_uops_0_lrs1_rtype;
  wire [1:0] rename_stage_io_dec_uops_0_lrs2_rtype;
  wire  rename_stage_io_dec_uops_0_frs3_en;
  wire  rename_stage_io_dec_uops_0_fp_val;
  wire  rename_stage_io_dec_uops_0_fp_single;
  wire  rename_stage_io_dec_uops_0_xcpt_pf_if;
  wire  rename_stage_io_dec_uops_0_xcpt_ae_if;
  wire  rename_stage_io_dec_uops_0_replay_if;
  wire  rename_stage_io_dec_uops_0_xcpt_ma_if;
  wire [31:0] rename_stage_io_dec_uops_0_debug_events_fetch_seq;
  wire  rename_stage_io_dec_uops_1_valid;
  wire [8:0] rename_stage_io_dec_uops_1_uopc;
  wire [31:0] rename_stage_io_dec_uops_1_inst;
  wire [39:0] rename_stage_io_dec_uops_1_pc;
  wire [1:0] rename_stage_io_dec_uops_1_iqtype;
  wire [9:0] rename_stage_io_dec_uops_1_fu_code;
  wire  rename_stage_io_dec_uops_1_allocate_brtag;
  wire  rename_stage_io_dec_uops_1_is_br_or_jmp;
  wire  rename_stage_io_dec_uops_1_is_jump;
  wire  rename_stage_io_dec_uops_1_is_jal;
  wire  rename_stage_io_dec_uops_1_is_ret;
  wire  rename_stage_io_dec_uops_1_is_call;
  wire [7:0] rename_stage_io_dec_uops_1_br_mask;
  wire [2:0] rename_stage_io_dec_uops_1_br_tag;
  wire  rename_stage_io_dec_uops_1_br_prediction_btb_blame;
  wire  rename_stage_io_dec_uops_1_br_prediction_btb_hit;
  wire  rename_stage_io_dec_uops_1_br_prediction_btb_taken;
  wire  rename_stage_io_dec_uops_1_br_prediction_bpd_blame;
  wire  rename_stage_io_dec_uops_1_br_prediction_bpd_hit;
  wire  rename_stage_io_dec_uops_1_br_prediction_bpd_taken;
  wire [1:0] rename_stage_io_dec_uops_1_br_prediction_bim_resp_value;
  wire [5:0] rename_stage_io_dec_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_dec_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] rename_stage_io_dec_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] rename_stage_io_dec_uops_1_br_prediction_bpd_resp_info;
  wire [2:0] rename_stage_io_dec_uops_1_fetch_pc_lob;
  wire [19:0] rename_stage_io_dec_uops_1_imm_packed;
  wire [6:0] rename_stage_io_dec_uops_1_rob_idx;
  wire [3:0] rename_stage_io_dec_uops_1_ldq_idx;
  wire [3:0] rename_stage_io_dec_uops_1_stq_idx;
  wire [5:0] rename_stage_io_dec_uops_1_brob_idx;
  wire  rename_stage_io_dec_uops_1_exception;
  wire [63:0] rename_stage_io_dec_uops_1_exc_cause;
  wire  rename_stage_io_dec_uops_1_bypassable;
  wire [4:0] rename_stage_io_dec_uops_1_mem_cmd;
  wire [2:0] rename_stage_io_dec_uops_1_mem_typ;
  wire  rename_stage_io_dec_uops_1_is_fence;
  wire  rename_stage_io_dec_uops_1_is_fencei;
  wire  rename_stage_io_dec_uops_1_is_store;
  wire  rename_stage_io_dec_uops_1_is_amo;
  wire  rename_stage_io_dec_uops_1_is_load;
  wire  rename_stage_io_dec_uops_1_is_sys_pc2epc;
  wire  rename_stage_io_dec_uops_1_is_unique;
  wire  rename_stage_io_dec_uops_1_flush_on_commit;
  wire [5:0] rename_stage_io_dec_uops_1_ldst;
  wire [5:0] rename_stage_io_dec_uops_1_lrs1;
  wire [5:0] rename_stage_io_dec_uops_1_lrs2;
  wire [5:0] rename_stage_io_dec_uops_1_lrs3;
  wire  rename_stage_io_dec_uops_1_ldst_val;
  wire [1:0] rename_stage_io_dec_uops_1_dst_rtype;
  wire [1:0] rename_stage_io_dec_uops_1_lrs1_rtype;
  wire [1:0] rename_stage_io_dec_uops_1_lrs2_rtype;
  wire  rename_stage_io_dec_uops_1_frs3_en;
  wire  rename_stage_io_dec_uops_1_fp_val;
  wire  rename_stage_io_dec_uops_1_fp_single;
  wire  rename_stage_io_dec_uops_1_xcpt_pf_if;
  wire  rename_stage_io_dec_uops_1_xcpt_ae_if;
  wire  rename_stage_io_dec_uops_1_replay_if;
  wire  rename_stage_io_dec_uops_1_xcpt_ma_if;
  wire [31:0] rename_stage_io_dec_uops_1_debug_events_fetch_seq;
  wire  rename_stage_io_ren1_mask_0;
  wire  rename_stage_io_ren1_mask_1;
  wire [39:0] rename_stage_io_ren1_uops_0_pc;
  wire [7:0] rename_stage_io_ren1_uops_0_br_mask;
  wire [6:0] rename_stage_io_ren1_uops_0_rob_idx;
  wire [5:0] rename_stage_io_ren1_uops_0_brob_idx;
  wire [6:0] rename_stage_io_ren1_uops_0_pdst;
  wire [6:0] rename_stage_io_ren1_uops_0_stale_pdst;
  wire  rename_stage_io_ren1_uops_0_exception;
  wire [63:0] rename_stage_io_ren1_uops_0_exc_cause;
  wire  rename_stage_io_ren1_uops_0_is_fence;
  wire  rename_stage_io_ren1_uops_0_is_fencei;
  wire  rename_stage_io_ren1_uops_0_is_store;
  wire  rename_stage_io_ren1_uops_0_is_load;
  wire  rename_stage_io_ren1_uops_0_is_sys_pc2epc;
  wire  rename_stage_io_ren1_uops_0_is_unique;
  wire  rename_stage_io_ren1_uops_0_flush_on_commit;
  wire [5:0] rename_stage_io_ren1_uops_0_ldst;
  wire  rename_stage_io_ren1_uops_0_ldst_val;
  wire [1:0] rename_stage_io_ren1_uops_0_dst_rtype;
  wire  rename_stage_io_ren1_uops_0_fp_val;
  wire [7:0] rename_stage_io_ren1_uops_1_br_mask;
  wire [6:0] rename_stage_io_ren1_uops_1_rob_idx;
  wire [6:0] rename_stage_io_ren1_uops_1_pdst;
  wire [6:0] rename_stage_io_ren1_uops_1_stale_pdst;
  wire  rename_stage_io_ren1_uops_1_exception;
  wire [63:0] rename_stage_io_ren1_uops_1_exc_cause;
  wire  rename_stage_io_ren1_uops_1_is_fence;
  wire  rename_stage_io_ren1_uops_1_is_fencei;
  wire  rename_stage_io_ren1_uops_1_is_store;
  wire  rename_stage_io_ren1_uops_1_is_load;
  wire  rename_stage_io_ren1_uops_1_is_sys_pc2epc;
  wire  rename_stage_io_ren1_uops_1_is_unique;
  wire  rename_stage_io_ren1_uops_1_flush_on_commit;
  wire [5:0] rename_stage_io_ren1_uops_1_ldst;
  wire  rename_stage_io_ren1_uops_1_ldst_val;
  wire [1:0] rename_stage_io_ren1_uops_1_dst_rtype;
  wire  rename_stage_io_ren1_uops_1_fp_val;
  wire  rename_stage_io_ren2_mask_0;
  wire  rename_stage_io_ren2_mask_1;
  wire  rename_stage_io_ren2_uops_0_valid;
  wire [8:0] rename_stage_io_ren2_uops_0_uopc;
  wire [31:0] rename_stage_io_ren2_uops_0_inst;
  wire [39:0] rename_stage_io_ren2_uops_0_pc;
  wire [1:0] rename_stage_io_ren2_uops_0_iqtype;
  wire [9:0] rename_stage_io_ren2_uops_0_fu_code;
  wire  rename_stage_io_ren2_uops_0_allocate_brtag;
  wire  rename_stage_io_ren2_uops_0_is_br_or_jmp;
  wire  rename_stage_io_ren2_uops_0_is_jump;
  wire  rename_stage_io_ren2_uops_0_is_jal;
  wire  rename_stage_io_ren2_uops_0_is_ret;
  wire  rename_stage_io_ren2_uops_0_is_call;
  wire [7:0] rename_stage_io_ren2_uops_0_br_mask;
  wire [2:0] rename_stage_io_ren2_uops_0_br_tag;
  wire  rename_stage_io_ren2_uops_0_br_prediction_btb_blame;
  wire  rename_stage_io_ren2_uops_0_br_prediction_btb_hit;
  wire  rename_stage_io_ren2_uops_0_br_prediction_btb_taken;
  wire  rename_stage_io_ren2_uops_0_br_prediction_bpd_blame;
  wire  rename_stage_io_ren2_uops_0_br_prediction_bpd_hit;
  wire  rename_stage_io_ren2_uops_0_br_prediction_bpd_taken;
  wire [1:0] rename_stage_io_ren2_uops_0_br_prediction_bim_resp_value;
  wire [5:0] rename_stage_io_ren2_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_ren2_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_info;
  wire  rename_stage_io_ren2_uops_0_stat_brjmp_mispredicted;
  wire  rename_stage_io_ren2_uops_0_stat_btb_made_pred;
  wire  rename_stage_io_ren2_uops_0_stat_btb_mispredicted;
  wire  rename_stage_io_ren2_uops_0_stat_bpd_made_pred;
  wire  rename_stage_io_ren2_uops_0_stat_bpd_mispredicted;
  wire [2:0] rename_stage_io_ren2_uops_0_fetch_pc_lob;
  wire [19:0] rename_stage_io_ren2_uops_0_imm_packed;
  wire [11:0] rename_stage_io_ren2_uops_0_csr_addr;
  wire [6:0] rename_stage_io_ren2_uops_0_rob_idx;
  wire [3:0] rename_stage_io_ren2_uops_0_ldq_idx;
  wire [3:0] rename_stage_io_ren2_uops_0_stq_idx;
  wire [5:0] rename_stage_io_ren2_uops_0_brob_idx;
  wire [6:0] rename_stage_io_ren2_uops_0_pdst;
  wire [6:0] rename_stage_io_ren2_uops_0_pop1;
  wire [6:0] rename_stage_io_ren2_uops_0_pop2;
  wire [6:0] rename_stage_io_ren2_uops_0_pop3;
  wire  rename_stage_io_ren2_uops_0_prs1_busy;
  wire  rename_stage_io_ren2_uops_0_prs2_busy;
  wire  rename_stage_io_ren2_uops_0_prs3_busy;
  wire [6:0] rename_stage_io_ren2_uops_0_stale_pdst;
  wire  rename_stage_io_ren2_uops_0_exception;
  wire [63:0] rename_stage_io_ren2_uops_0_exc_cause;
  wire  rename_stage_io_ren2_uops_0_bypassable;
  wire [4:0] rename_stage_io_ren2_uops_0_mem_cmd;
  wire [2:0] rename_stage_io_ren2_uops_0_mem_typ;
  wire  rename_stage_io_ren2_uops_0_is_fence;
  wire  rename_stage_io_ren2_uops_0_is_fencei;
  wire  rename_stage_io_ren2_uops_0_is_store;
  wire  rename_stage_io_ren2_uops_0_is_amo;
  wire  rename_stage_io_ren2_uops_0_is_load;
  wire  rename_stage_io_ren2_uops_0_is_sys_pc2epc;
  wire  rename_stage_io_ren2_uops_0_is_unique;
  wire  rename_stage_io_ren2_uops_0_flush_on_commit;
  wire [5:0] rename_stage_io_ren2_uops_0_ldst;
  wire [5:0] rename_stage_io_ren2_uops_0_lrs1;
  wire [5:0] rename_stage_io_ren2_uops_0_lrs2;
  wire [5:0] rename_stage_io_ren2_uops_0_lrs3;
  wire  rename_stage_io_ren2_uops_0_ldst_val;
  wire [1:0] rename_stage_io_ren2_uops_0_dst_rtype;
  wire [1:0] rename_stage_io_ren2_uops_0_lrs1_rtype;
  wire [1:0] rename_stage_io_ren2_uops_0_lrs2_rtype;
  wire  rename_stage_io_ren2_uops_0_frs3_en;
  wire  rename_stage_io_ren2_uops_0_fp_val;
  wire  rename_stage_io_ren2_uops_0_fp_single;
  wire  rename_stage_io_ren2_uops_0_xcpt_pf_if;
  wire  rename_stage_io_ren2_uops_0_xcpt_ae_if;
  wire  rename_stage_io_ren2_uops_0_replay_if;
  wire  rename_stage_io_ren2_uops_0_xcpt_ma_if;
  wire [63:0] rename_stage_io_ren2_uops_0_debug_wdata;
  wire [31:0] rename_stage_io_ren2_uops_0_debug_events_fetch_seq;
  wire  rename_stage_io_ren2_uops_1_valid;
  wire [8:0] rename_stage_io_ren2_uops_1_uopc;
  wire [31:0] rename_stage_io_ren2_uops_1_inst;
  wire [39:0] rename_stage_io_ren2_uops_1_pc;
  wire [1:0] rename_stage_io_ren2_uops_1_iqtype;
  wire [9:0] rename_stage_io_ren2_uops_1_fu_code;
  wire  rename_stage_io_ren2_uops_1_allocate_brtag;
  wire  rename_stage_io_ren2_uops_1_is_br_or_jmp;
  wire  rename_stage_io_ren2_uops_1_is_jump;
  wire  rename_stage_io_ren2_uops_1_is_jal;
  wire  rename_stage_io_ren2_uops_1_is_ret;
  wire  rename_stage_io_ren2_uops_1_is_call;
  wire [7:0] rename_stage_io_ren2_uops_1_br_mask;
  wire [2:0] rename_stage_io_ren2_uops_1_br_tag;
  wire  rename_stage_io_ren2_uops_1_br_prediction_btb_blame;
  wire  rename_stage_io_ren2_uops_1_br_prediction_btb_hit;
  wire  rename_stage_io_ren2_uops_1_br_prediction_btb_taken;
  wire  rename_stage_io_ren2_uops_1_br_prediction_bpd_blame;
  wire  rename_stage_io_ren2_uops_1_br_prediction_bpd_hit;
  wire  rename_stage_io_ren2_uops_1_br_prediction_bpd_taken;
  wire [1:0] rename_stage_io_ren2_uops_1_br_prediction_bim_resp_value;
  wire [5:0] rename_stage_io_ren2_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_ren2_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_info;
  wire  rename_stage_io_ren2_uops_1_stat_brjmp_mispredicted;
  wire  rename_stage_io_ren2_uops_1_stat_btb_made_pred;
  wire  rename_stage_io_ren2_uops_1_stat_btb_mispredicted;
  wire  rename_stage_io_ren2_uops_1_stat_bpd_made_pred;
  wire  rename_stage_io_ren2_uops_1_stat_bpd_mispredicted;
  wire [2:0] rename_stage_io_ren2_uops_1_fetch_pc_lob;
  wire [19:0] rename_stage_io_ren2_uops_1_imm_packed;
  wire [11:0] rename_stage_io_ren2_uops_1_csr_addr;
  wire [6:0] rename_stage_io_ren2_uops_1_rob_idx;
  wire [3:0] rename_stage_io_ren2_uops_1_ldq_idx;
  wire [3:0] rename_stage_io_ren2_uops_1_stq_idx;
  wire [5:0] rename_stage_io_ren2_uops_1_brob_idx;
  wire [6:0] rename_stage_io_ren2_uops_1_pdst;
  wire [6:0] rename_stage_io_ren2_uops_1_pop1;
  wire [6:0] rename_stage_io_ren2_uops_1_pop2;
  wire [6:0] rename_stage_io_ren2_uops_1_pop3;
  wire  rename_stage_io_ren2_uops_1_prs1_busy;
  wire  rename_stage_io_ren2_uops_1_prs2_busy;
  wire  rename_stage_io_ren2_uops_1_prs3_busy;
  wire [6:0] rename_stage_io_ren2_uops_1_stale_pdst;
  wire  rename_stage_io_ren2_uops_1_exception;
  wire [63:0] rename_stage_io_ren2_uops_1_exc_cause;
  wire  rename_stage_io_ren2_uops_1_bypassable;
  wire [4:0] rename_stage_io_ren2_uops_1_mem_cmd;
  wire [2:0] rename_stage_io_ren2_uops_1_mem_typ;
  wire  rename_stage_io_ren2_uops_1_is_fence;
  wire  rename_stage_io_ren2_uops_1_is_fencei;
  wire  rename_stage_io_ren2_uops_1_is_store;
  wire  rename_stage_io_ren2_uops_1_is_amo;
  wire  rename_stage_io_ren2_uops_1_is_load;
  wire  rename_stage_io_ren2_uops_1_is_sys_pc2epc;
  wire  rename_stage_io_ren2_uops_1_is_unique;
  wire  rename_stage_io_ren2_uops_1_flush_on_commit;
  wire [5:0] rename_stage_io_ren2_uops_1_ldst;
  wire [5:0] rename_stage_io_ren2_uops_1_lrs1;
  wire [5:0] rename_stage_io_ren2_uops_1_lrs2;
  wire [5:0] rename_stage_io_ren2_uops_1_lrs3;
  wire  rename_stage_io_ren2_uops_1_ldst_val;
  wire [1:0] rename_stage_io_ren2_uops_1_dst_rtype;
  wire [1:0] rename_stage_io_ren2_uops_1_lrs1_rtype;
  wire [1:0] rename_stage_io_ren2_uops_1_lrs2_rtype;
  wire  rename_stage_io_ren2_uops_1_frs3_en;
  wire  rename_stage_io_ren2_uops_1_fp_val;
  wire  rename_stage_io_ren2_uops_1_fp_single;
  wire  rename_stage_io_ren2_uops_1_xcpt_pf_if;
  wire  rename_stage_io_ren2_uops_1_xcpt_ae_if;
  wire  rename_stage_io_ren2_uops_1_replay_if;
  wire  rename_stage_io_ren2_uops_1_xcpt_ma_if;
  wire [63:0] rename_stage_io_ren2_uops_1_debug_wdata;
  wire [31:0] rename_stage_io_ren2_uops_1_debug_events_fetch_seq;
  wire [1:0] rename_stage_io_ren_pred_info_0_bim_resp_value;
  wire [5:0] rename_stage_io_ren_pred_info_0_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_ren_pred_info_0_bim_resp_way_idx;
  wire [14:0] rename_stage_io_ren_pred_info_0_bpd_resp_history;
  wire [7:0] rename_stage_io_ren_pred_info_0_bpd_resp_history_ptr;
  wire [1:0] rename_stage_io_ren_pred_info_1_bim_resp_value;
  wire [5:0] rename_stage_io_ren_pred_info_1_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_ren_pred_info_1_bim_resp_way_idx;
  wire [14:0] rename_stage_io_ren_pred_info_1_bpd_resp_history;
  wire [7:0] rename_stage_io_ren_pred_info_1_bpd_resp_history_ptr;
  wire  rename_stage_io_brinfo_valid;
  wire  rename_stage_io_brinfo_mispredict;
  wire [7:0] rename_stage_io_brinfo_mask;
  wire [2:0] rename_stage_io_brinfo_tag;
  wire [2:0] rename_stage_io_get_pred_br_tag;
  wire [1:0] rename_stage_io_get_pred_info_bim_resp_value;
  wire [5:0] rename_stage_io_get_pred_info_bim_resp_entry_idx;
  wire [1:0] rename_stage_io_get_pred_info_bim_resp_way_idx;
  wire [14:0] rename_stage_io_get_pred_info_bpd_resp_history;
  wire [7:0] rename_stage_io_get_pred_info_bpd_resp_history_ptr;
  wire  rename_stage_io_dis_inst_can_proceed_0;
  wire  rename_stage_io_dis_inst_can_proceed_1;
  wire  rename_stage_io_int_wakeups_0_valid;
  wire [6:0] rename_stage_io_int_wakeups_0_bits_uop_pdst;
  wire [1:0] rename_stage_io_int_wakeups_0_bits_uop_dst_rtype;
  wire  rename_stage_io_int_wakeups_1_valid;
  wire [6:0] rename_stage_io_int_wakeups_1_bits_uop_pdst;
  wire [1:0] rename_stage_io_int_wakeups_1_bits_uop_dst_rtype;
  wire  rename_stage_io_int_wakeups_2_valid;
  wire [6:0] rename_stage_io_int_wakeups_2_bits_uop_pdst;
  wire [1:0] rename_stage_io_int_wakeups_2_bits_uop_dst_rtype;
  wire  rename_stage_io_int_wakeups_3_valid;
  wire [6:0] rename_stage_io_int_wakeups_3_bits_uop_pdst;
  wire [1:0] rename_stage_io_int_wakeups_3_bits_uop_dst_rtype;
  wire  rename_stage_io_int_wakeups_4_valid;
  wire [6:0] rename_stage_io_int_wakeups_4_bits_uop_pdst;
  wire [1:0] rename_stage_io_int_wakeups_4_bits_uop_dst_rtype;
  wire  rename_stage_io_fp_wakeups_0_valid;
  wire [6:0] rename_stage_io_fp_wakeups_0_bits_uop_pdst;
  wire [1:0] rename_stage_io_fp_wakeups_0_bits_uop_dst_rtype;
  wire  rename_stage_io_fp_wakeups_1_valid;
  wire [6:0] rename_stage_io_fp_wakeups_1_bits_uop_pdst;
  wire [1:0] rename_stage_io_fp_wakeups_1_bits_uop_dst_rtype;
  wire  rename_stage_io_com_valids_0;
  wire  rename_stage_io_com_valids_1;
  wire [6:0] rename_stage_io_com_uops_0_pdst;
  wire [6:0] rename_stage_io_com_uops_0_stale_pdst;
  wire [5:0] rename_stage_io_com_uops_0_ldst;
  wire [1:0] rename_stage_io_com_uops_0_dst_rtype;
  wire [6:0] rename_stage_io_com_uops_1_pdst;
  wire [6:0] rename_stage_io_com_uops_1_stale_pdst;
  wire [5:0] rename_stage_io_com_uops_1_ldst;
  wire [1:0] rename_stage_io_com_uops_1_dst_rtype;
  wire  rename_stage_io_com_rbk_valids_0;
  wire  rename_stage_io_com_rbk_valids_1;
  wire  rename_stage_io_debug_rob_empty;
  wire  issue_units_0_clock;
  wire  issue_units_0_reset;
  wire  issue_units_0_io_dis_valids_0;
  wire  issue_units_0_io_dis_valids_1;
  wire  issue_units_0_io_dis_uops_0_valid;
  wire [8:0] issue_units_0_io_dis_uops_0_uopc;
  wire [31:0] issue_units_0_io_dis_uops_0_inst;
  wire [39:0] issue_units_0_io_dis_uops_0_pc;
  wire [1:0] issue_units_0_io_dis_uops_0_iqtype;
  wire [9:0] issue_units_0_io_dis_uops_0_fu_code;
  wire  issue_units_0_io_dis_uops_0_allocate_brtag;
  wire  issue_units_0_io_dis_uops_0_is_br_or_jmp;
  wire  issue_units_0_io_dis_uops_0_is_jump;
  wire  issue_units_0_io_dis_uops_0_is_jal;
  wire  issue_units_0_io_dis_uops_0_is_ret;
  wire  issue_units_0_io_dis_uops_0_is_call;
  wire [7:0] issue_units_0_io_dis_uops_0_br_mask;
  wire [2:0] issue_units_0_io_dis_uops_0_br_tag;
  wire  issue_units_0_io_dis_uops_0_br_prediction_btb_blame;
  wire  issue_units_0_io_dis_uops_0_br_prediction_btb_hit;
  wire  issue_units_0_io_dis_uops_0_br_prediction_btb_taken;
  wire  issue_units_0_io_dis_uops_0_br_prediction_bpd_blame;
  wire  issue_units_0_io_dis_uops_0_br_prediction_bpd_hit;
  wire  issue_units_0_io_dis_uops_0_br_prediction_bpd_taken;
  wire [1:0] issue_units_0_io_dis_uops_0_br_prediction_bim_resp_value;
  wire [5:0] issue_units_0_io_dis_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_0_io_dis_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_info;
  wire  issue_units_0_io_dis_uops_0_stat_brjmp_mispredicted;
  wire  issue_units_0_io_dis_uops_0_stat_btb_made_pred;
  wire  issue_units_0_io_dis_uops_0_stat_btb_mispredicted;
  wire  issue_units_0_io_dis_uops_0_stat_bpd_made_pred;
  wire  issue_units_0_io_dis_uops_0_stat_bpd_mispredicted;
  wire [2:0] issue_units_0_io_dis_uops_0_fetch_pc_lob;
  wire [19:0] issue_units_0_io_dis_uops_0_imm_packed;
  wire [11:0] issue_units_0_io_dis_uops_0_csr_addr;
  wire [6:0] issue_units_0_io_dis_uops_0_rob_idx;
  wire [3:0] issue_units_0_io_dis_uops_0_ldq_idx;
  wire [3:0] issue_units_0_io_dis_uops_0_stq_idx;
  wire [5:0] issue_units_0_io_dis_uops_0_brob_idx;
  wire [6:0] issue_units_0_io_dis_uops_0_pdst;
  wire [6:0] issue_units_0_io_dis_uops_0_pop1;
  wire [6:0] issue_units_0_io_dis_uops_0_pop2;
  wire [6:0] issue_units_0_io_dis_uops_0_pop3;
  wire  issue_units_0_io_dis_uops_0_prs1_busy;
  wire  issue_units_0_io_dis_uops_0_prs2_busy;
  wire  issue_units_0_io_dis_uops_0_prs3_busy;
  wire [6:0] issue_units_0_io_dis_uops_0_stale_pdst;
  wire  issue_units_0_io_dis_uops_0_exception;
  wire [63:0] issue_units_0_io_dis_uops_0_exc_cause;
  wire  issue_units_0_io_dis_uops_0_bypassable;
  wire [4:0] issue_units_0_io_dis_uops_0_mem_cmd;
  wire [2:0] issue_units_0_io_dis_uops_0_mem_typ;
  wire  issue_units_0_io_dis_uops_0_is_fence;
  wire  issue_units_0_io_dis_uops_0_is_fencei;
  wire  issue_units_0_io_dis_uops_0_is_store;
  wire  issue_units_0_io_dis_uops_0_is_amo;
  wire  issue_units_0_io_dis_uops_0_is_load;
  wire  issue_units_0_io_dis_uops_0_is_sys_pc2epc;
  wire  issue_units_0_io_dis_uops_0_is_unique;
  wire  issue_units_0_io_dis_uops_0_flush_on_commit;
  wire [5:0] issue_units_0_io_dis_uops_0_ldst;
  wire [5:0] issue_units_0_io_dis_uops_0_lrs1;
  wire [5:0] issue_units_0_io_dis_uops_0_lrs2;
  wire [5:0] issue_units_0_io_dis_uops_0_lrs3;
  wire  issue_units_0_io_dis_uops_0_ldst_val;
  wire [1:0] issue_units_0_io_dis_uops_0_dst_rtype;
  wire [1:0] issue_units_0_io_dis_uops_0_lrs1_rtype;
  wire [1:0] issue_units_0_io_dis_uops_0_lrs2_rtype;
  wire  issue_units_0_io_dis_uops_0_frs3_en;
  wire  issue_units_0_io_dis_uops_0_fp_val;
  wire  issue_units_0_io_dis_uops_0_fp_single;
  wire  issue_units_0_io_dis_uops_0_xcpt_pf_if;
  wire  issue_units_0_io_dis_uops_0_xcpt_ae_if;
  wire  issue_units_0_io_dis_uops_0_replay_if;
  wire  issue_units_0_io_dis_uops_0_xcpt_ma_if;
  wire [63:0] issue_units_0_io_dis_uops_0_debug_wdata;
  wire [31:0] issue_units_0_io_dis_uops_0_debug_events_fetch_seq;
  wire  issue_units_0_io_dis_uops_1_valid;
  wire [8:0] issue_units_0_io_dis_uops_1_uopc;
  wire [31:0] issue_units_0_io_dis_uops_1_inst;
  wire [39:0] issue_units_0_io_dis_uops_1_pc;
  wire [1:0] issue_units_0_io_dis_uops_1_iqtype;
  wire [9:0] issue_units_0_io_dis_uops_1_fu_code;
  wire  issue_units_0_io_dis_uops_1_allocate_brtag;
  wire  issue_units_0_io_dis_uops_1_is_br_or_jmp;
  wire  issue_units_0_io_dis_uops_1_is_jump;
  wire  issue_units_0_io_dis_uops_1_is_jal;
  wire  issue_units_0_io_dis_uops_1_is_ret;
  wire  issue_units_0_io_dis_uops_1_is_call;
  wire [7:0] issue_units_0_io_dis_uops_1_br_mask;
  wire [2:0] issue_units_0_io_dis_uops_1_br_tag;
  wire  issue_units_0_io_dis_uops_1_br_prediction_btb_blame;
  wire  issue_units_0_io_dis_uops_1_br_prediction_btb_hit;
  wire  issue_units_0_io_dis_uops_1_br_prediction_btb_taken;
  wire  issue_units_0_io_dis_uops_1_br_prediction_bpd_blame;
  wire  issue_units_0_io_dis_uops_1_br_prediction_bpd_hit;
  wire  issue_units_0_io_dis_uops_1_br_prediction_bpd_taken;
  wire [1:0] issue_units_0_io_dis_uops_1_br_prediction_bim_resp_value;
  wire [5:0] issue_units_0_io_dis_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_0_io_dis_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_info;
  wire  issue_units_0_io_dis_uops_1_stat_brjmp_mispredicted;
  wire  issue_units_0_io_dis_uops_1_stat_btb_made_pred;
  wire  issue_units_0_io_dis_uops_1_stat_btb_mispredicted;
  wire  issue_units_0_io_dis_uops_1_stat_bpd_made_pred;
  wire  issue_units_0_io_dis_uops_1_stat_bpd_mispredicted;
  wire [2:0] issue_units_0_io_dis_uops_1_fetch_pc_lob;
  wire [19:0] issue_units_0_io_dis_uops_1_imm_packed;
  wire [11:0] issue_units_0_io_dis_uops_1_csr_addr;
  wire [6:0] issue_units_0_io_dis_uops_1_rob_idx;
  wire [3:0] issue_units_0_io_dis_uops_1_ldq_idx;
  wire [3:0] issue_units_0_io_dis_uops_1_stq_idx;
  wire [5:0] issue_units_0_io_dis_uops_1_brob_idx;
  wire [6:0] issue_units_0_io_dis_uops_1_pdst;
  wire [6:0] issue_units_0_io_dis_uops_1_pop1;
  wire [6:0] issue_units_0_io_dis_uops_1_pop2;
  wire [6:0] issue_units_0_io_dis_uops_1_pop3;
  wire  issue_units_0_io_dis_uops_1_prs1_busy;
  wire  issue_units_0_io_dis_uops_1_prs2_busy;
  wire  issue_units_0_io_dis_uops_1_prs3_busy;
  wire [6:0] issue_units_0_io_dis_uops_1_stale_pdst;
  wire  issue_units_0_io_dis_uops_1_exception;
  wire [63:0] issue_units_0_io_dis_uops_1_exc_cause;
  wire  issue_units_0_io_dis_uops_1_bypassable;
  wire [4:0] issue_units_0_io_dis_uops_1_mem_cmd;
  wire [2:0] issue_units_0_io_dis_uops_1_mem_typ;
  wire  issue_units_0_io_dis_uops_1_is_fence;
  wire  issue_units_0_io_dis_uops_1_is_fencei;
  wire  issue_units_0_io_dis_uops_1_is_store;
  wire  issue_units_0_io_dis_uops_1_is_amo;
  wire  issue_units_0_io_dis_uops_1_is_load;
  wire  issue_units_0_io_dis_uops_1_is_sys_pc2epc;
  wire  issue_units_0_io_dis_uops_1_is_unique;
  wire  issue_units_0_io_dis_uops_1_flush_on_commit;
  wire [5:0] issue_units_0_io_dis_uops_1_ldst;
  wire [5:0] issue_units_0_io_dis_uops_1_lrs1;
  wire [5:0] issue_units_0_io_dis_uops_1_lrs2;
  wire [5:0] issue_units_0_io_dis_uops_1_lrs3;
  wire  issue_units_0_io_dis_uops_1_ldst_val;
  wire [1:0] issue_units_0_io_dis_uops_1_dst_rtype;
  wire [1:0] issue_units_0_io_dis_uops_1_lrs1_rtype;
  wire [1:0] issue_units_0_io_dis_uops_1_lrs2_rtype;
  wire  issue_units_0_io_dis_uops_1_frs3_en;
  wire  issue_units_0_io_dis_uops_1_fp_val;
  wire  issue_units_0_io_dis_uops_1_fp_single;
  wire  issue_units_0_io_dis_uops_1_xcpt_pf_if;
  wire  issue_units_0_io_dis_uops_1_xcpt_ae_if;
  wire  issue_units_0_io_dis_uops_1_replay_if;
  wire  issue_units_0_io_dis_uops_1_xcpt_ma_if;
  wire [63:0] issue_units_0_io_dis_uops_1_debug_wdata;
  wire [31:0] issue_units_0_io_dis_uops_1_debug_events_fetch_seq;
  wire  issue_units_0_io_dis_readys_0;
  wire  issue_units_0_io_dis_readys_1;
  wire  issue_units_0_io_iss_valids_0;
  wire [8:0] issue_units_0_io_iss_uops_0_uopc;
  wire [7:0] issue_units_0_io_iss_uops_0_br_mask;
  wire [19:0] issue_units_0_io_iss_uops_0_imm_packed;
  wire [6:0] issue_units_0_io_iss_uops_0_rob_idx;
  wire [3:0] issue_units_0_io_iss_uops_0_ldq_idx;
  wire [3:0] issue_units_0_io_iss_uops_0_stq_idx;
  wire [6:0] issue_units_0_io_iss_uops_0_pdst;
  wire [6:0] issue_units_0_io_iss_uops_0_pop1;
  wire [6:0] issue_units_0_io_iss_uops_0_pop2;
  wire [4:0] issue_units_0_io_iss_uops_0_mem_cmd;
  wire [2:0] issue_units_0_io_iss_uops_0_mem_typ;
  wire  issue_units_0_io_iss_uops_0_is_fence;
  wire  issue_units_0_io_iss_uops_0_is_store;
  wire  issue_units_0_io_iss_uops_0_is_amo;
  wire  issue_units_0_io_iss_uops_0_is_load;
  wire [1:0] issue_units_0_io_iss_uops_0_dst_rtype;
  wire [1:0] issue_units_0_io_iss_uops_0_lrs1_rtype;
  wire [1:0] issue_units_0_io_iss_uops_0_lrs2_rtype;
  wire  issue_units_0_io_iss_uops_0_fp_val;
  wire  issue_units_0_io_wakeup_pdsts_0_valid;
  wire [6:0] issue_units_0_io_wakeup_pdsts_0_bits;
  wire  issue_units_0_io_wakeup_pdsts_1_valid;
  wire [6:0] issue_units_0_io_wakeup_pdsts_1_bits;
  wire  issue_units_0_io_wakeup_pdsts_2_valid;
  wire [6:0] issue_units_0_io_wakeup_pdsts_2_bits;
  wire  issue_units_0_io_wakeup_pdsts_3_valid;
  wire [6:0] issue_units_0_io_wakeup_pdsts_3_bits;
  wire  issue_units_0_io_wakeup_pdsts_4_valid;
  wire [6:0] issue_units_0_io_wakeup_pdsts_4_bits;
  wire  issue_units_0_io_brinfo_valid;
  wire  issue_units_0_io_brinfo_mispredict;
  wire [7:0] issue_units_0_io_brinfo_mask;
  wire  issue_units_0_io_flush_pipeline;
  wire  issue_units_1_clock;
  wire  issue_units_1_reset;
  wire  issue_units_1_io_dis_valids_0;
  wire  issue_units_1_io_dis_valids_1;
  wire  issue_units_1_io_dis_uops_0_valid;
  wire [8:0] issue_units_1_io_dis_uops_0_uopc;
  wire [31:0] issue_units_1_io_dis_uops_0_inst;
  wire [39:0] issue_units_1_io_dis_uops_0_pc;
  wire [1:0] issue_units_1_io_dis_uops_0_iqtype;
  wire [9:0] issue_units_1_io_dis_uops_0_fu_code;
  wire  issue_units_1_io_dis_uops_0_allocate_brtag;
  wire  issue_units_1_io_dis_uops_0_is_br_or_jmp;
  wire  issue_units_1_io_dis_uops_0_is_jump;
  wire  issue_units_1_io_dis_uops_0_is_jal;
  wire  issue_units_1_io_dis_uops_0_is_ret;
  wire  issue_units_1_io_dis_uops_0_is_call;
  wire [7:0] issue_units_1_io_dis_uops_0_br_mask;
  wire [2:0] issue_units_1_io_dis_uops_0_br_tag;
  wire  issue_units_1_io_dis_uops_0_br_prediction_btb_blame;
  wire  issue_units_1_io_dis_uops_0_br_prediction_btb_hit;
  wire  issue_units_1_io_dis_uops_0_br_prediction_btb_taken;
  wire  issue_units_1_io_dis_uops_0_br_prediction_bpd_blame;
  wire  issue_units_1_io_dis_uops_0_br_prediction_bpd_hit;
  wire  issue_units_1_io_dis_uops_0_br_prediction_bpd_taken;
  wire [1:0] issue_units_1_io_dis_uops_0_br_prediction_bim_resp_value;
  wire [5:0] issue_units_1_io_dis_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_1_io_dis_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_info;
  wire  issue_units_1_io_dis_uops_0_stat_brjmp_mispredicted;
  wire  issue_units_1_io_dis_uops_0_stat_btb_made_pred;
  wire  issue_units_1_io_dis_uops_0_stat_btb_mispredicted;
  wire  issue_units_1_io_dis_uops_0_stat_bpd_made_pred;
  wire  issue_units_1_io_dis_uops_0_stat_bpd_mispredicted;
  wire [2:0] issue_units_1_io_dis_uops_0_fetch_pc_lob;
  wire [19:0] issue_units_1_io_dis_uops_0_imm_packed;
  wire [11:0] issue_units_1_io_dis_uops_0_csr_addr;
  wire [6:0] issue_units_1_io_dis_uops_0_rob_idx;
  wire [3:0] issue_units_1_io_dis_uops_0_ldq_idx;
  wire [3:0] issue_units_1_io_dis_uops_0_stq_idx;
  wire [5:0] issue_units_1_io_dis_uops_0_brob_idx;
  wire [6:0] issue_units_1_io_dis_uops_0_pdst;
  wire [6:0] issue_units_1_io_dis_uops_0_pop1;
  wire [6:0] issue_units_1_io_dis_uops_0_pop2;
  wire [6:0] issue_units_1_io_dis_uops_0_pop3;
  wire  issue_units_1_io_dis_uops_0_prs1_busy;
  wire  issue_units_1_io_dis_uops_0_prs2_busy;
  wire  issue_units_1_io_dis_uops_0_prs3_busy;
  wire [6:0] issue_units_1_io_dis_uops_0_stale_pdst;
  wire  issue_units_1_io_dis_uops_0_exception;
  wire [63:0] issue_units_1_io_dis_uops_0_exc_cause;
  wire  issue_units_1_io_dis_uops_0_bypassable;
  wire [4:0] issue_units_1_io_dis_uops_0_mem_cmd;
  wire [2:0] issue_units_1_io_dis_uops_0_mem_typ;
  wire  issue_units_1_io_dis_uops_0_is_fence;
  wire  issue_units_1_io_dis_uops_0_is_fencei;
  wire  issue_units_1_io_dis_uops_0_is_store;
  wire  issue_units_1_io_dis_uops_0_is_amo;
  wire  issue_units_1_io_dis_uops_0_is_load;
  wire  issue_units_1_io_dis_uops_0_is_sys_pc2epc;
  wire  issue_units_1_io_dis_uops_0_is_unique;
  wire  issue_units_1_io_dis_uops_0_flush_on_commit;
  wire [5:0] issue_units_1_io_dis_uops_0_ldst;
  wire [5:0] issue_units_1_io_dis_uops_0_lrs1;
  wire [5:0] issue_units_1_io_dis_uops_0_lrs2;
  wire [5:0] issue_units_1_io_dis_uops_0_lrs3;
  wire  issue_units_1_io_dis_uops_0_ldst_val;
  wire [1:0] issue_units_1_io_dis_uops_0_dst_rtype;
  wire [1:0] issue_units_1_io_dis_uops_0_lrs1_rtype;
  wire [1:0] issue_units_1_io_dis_uops_0_lrs2_rtype;
  wire  issue_units_1_io_dis_uops_0_frs3_en;
  wire  issue_units_1_io_dis_uops_0_fp_val;
  wire  issue_units_1_io_dis_uops_0_fp_single;
  wire  issue_units_1_io_dis_uops_0_xcpt_pf_if;
  wire  issue_units_1_io_dis_uops_0_xcpt_ae_if;
  wire  issue_units_1_io_dis_uops_0_replay_if;
  wire  issue_units_1_io_dis_uops_0_xcpt_ma_if;
  wire [63:0] issue_units_1_io_dis_uops_0_debug_wdata;
  wire [31:0] issue_units_1_io_dis_uops_0_debug_events_fetch_seq;
  wire  issue_units_1_io_dis_uops_1_valid;
  wire [8:0] issue_units_1_io_dis_uops_1_uopc;
  wire [31:0] issue_units_1_io_dis_uops_1_inst;
  wire [39:0] issue_units_1_io_dis_uops_1_pc;
  wire [1:0] issue_units_1_io_dis_uops_1_iqtype;
  wire [9:0] issue_units_1_io_dis_uops_1_fu_code;
  wire  issue_units_1_io_dis_uops_1_allocate_brtag;
  wire  issue_units_1_io_dis_uops_1_is_br_or_jmp;
  wire  issue_units_1_io_dis_uops_1_is_jump;
  wire  issue_units_1_io_dis_uops_1_is_jal;
  wire  issue_units_1_io_dis_uops_1_is_ret;
  wire  issue_units_1_io_dis_uops_1_is_call;
  wire [7:0] issue_units_1_io_dis_uops_1_br_mask;
  wire [2:0] issue_units_1_io_dis_uops_1_br_tag;
  wire  issue_units_1_io_dis_uops_1_br_prediction_btb_blame;
  wire  issue_units_1_io_dis_uops_1_br_prediction_btb_hit;
  wire  issue_units_1_io_dis_uops_1_br_prediction_btb_taken;
  wire  issue_units_1_io_dis_uops_1_br_prediction_bpd_blame;
  wire  issue_units_1_io_dis_uops_1_br_prediction_bpd_hit;
  wire  issue_units_1_io_dis_uops_1_br_prediction_bpd_taken;
  wire [1:0] issue_units_1_io_dis_uops_1_br_prediction_bim_resp_value;
  wire [5:0] issue_units_1_io_dis_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_1_io_dis_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_info;
  wire  issue_units_1_io_dis_uops_1_stat_brjmp_mispredicted;
  wire  issue_units_1_io_dis_uops_1_stat_btb_made_pred;
  wire  issue_units_1_io_dis_uops_1_stat_btb_mispredicted;
  wire  issue_units_1_io_dis_uops_1_stat_bpd_made_pred;
  wire  issue_units_1_io_dis_uops_1_stat_bpd_mispredicted;
  wire [2:0] issue_units_1_io_dis_uops_1_fetch_pc_lob;
  wire [19:0] issue_units_1_io_dis_uops_1_imm_packed;
  wire [11:0] issue_units_1_io_dis_uops_1_csr_addr;
  wire [6:0] issue_units_1_io_dis_uops_1_rob_idx;
  wire [3:0] issue_units_1_io_dis_uops_1_ldq_idx;
  wire [3:0] issue_units_1_io_dis_uops_1_stq_idx;
  wire [5:0] issue_units_1_io_dis_uops_1_brob_idx;
  wire [6:0] issue_units_1_io_dis_uops_1_pdst;
  wire [6:0] issue_units_1_io_dis_uops_1_pop1;
  wire [6:0] issue_units_1_io_dis_uops_1_pop2;
  wire [6:0] issue_units_1_io_dis_uops_1_pop3;
  wire  issue_units_1_io_dis_uops_1_prs1_busy;
  wire  issue_units_1_io_dis_uops_1_prs2_busy;
  wire  issue_units_1_io_dis_uops_1_prs3_busy;
  wire [6:0] issue_units_1_io_dis_uops_1_stale_pdst;
  wire  issue_units_1_io_dis_uops_1_exception;
  wire [63:0] issue_units_1_io_dis_uops_1_exc_cause;
  wire  issue_units_1_io_dis_uops_1_bypassable;
  wire [4:0] issue_units_1_io_dis_uops_1_mem_cmd;
  wire [2:0] issue_units_1_io_dis_uops_1_mem_typ;
  wire  issue_units_1_io_dis_uops_1_is_fence;
  wire  issue_units_1_io_dis_uops_1_is_fencei;
  wire  issue_units_1_io_dis_uops_1_is_store;
  wire  issue_units_1_io_dis_uops_1_is_amo;
  wire  issue_units_1_io_dis_uops_1_is_load;
  wire  issue_units_1_io_dis_uops_1_is_sys_pc2epc;
  wire  issue_units_1_io_dis_uops_1_is_unique;
  wire  issue_units_1_io_dis_uops_1_flush_on_commit;
  wire [5:0] issue_units_1_io_dis_uops_1_ldst;
  wire [5:0] issue_units_1_io_dis_uops_1_lrs1;
  wire [5:0] issue_units_1_io_dis_uops_1_lrs2;
  wire [5:0] issue_units_1_io_dis_uops_1_lrs3;
  wire  issue_units_1_io_dis_uops_1_ldst_val;
  wire [1:0] issue_units_1_io_dis_uops_1_dst_rtype;
  wire [1:0] issue_units_1_io_dis_uops_1_lrs1_rtype;
  wire [1:0] issue_units_1_io_dis_uops_1_lrs2_rtype;
  wire  issue_units_1_io_dis_uops_1_frs3_en;
  wire  issue_units_1_io_dis_uops_1_fp_val;
  wire  issue_units_1_io_dis_uops_1_fp_single;
  wire  issue_units_1_io_dis_uops_1_xcpt_pf_if;
  wire  issue_units_1_io_dis_uops_1_xcpt_ae_if;
  wire  issue_units_1_io_dis_uops_1_replay_if;
  wire  issue_units_1_io_dis_uops_1_xcpt_ma_if;
  wire [63:0] issue_units_1_io_dis_uops_1_debug_wdata;
  wire [31:0] issue_units_1_io_dis_uops_1_debug_events_fetch_seq;
  wire  issue_units_1_io_dis_readys_0;
  wire  issue_units_1_io_dis_readys_1;
  wire  issue_units_1_io_iss_valids_0;
  wire  issue_units_1_io_iss_valids_1;
  wire  issue_units_1_io_iss_uops_0_valid;
  wire [1:0] issue_units_1_io_iss_uops_0_iw_state;
  wire [8:0] issue_units_1_io_iss_uops_0_uopc;
  wire [31:0] issue_units_1_io_iss_uops_0_inst;
  wire [39:0] issue_units_1_io_iss_uops_0_pc;
  wire [1:0] issue_units_1_io_iss_uops_0_iqtype;
  wire [9:0] issue_units_1_io_iss_uops_0_fu_code;
  wire  issue_units_1_io_iss_uops_0_allocate_brtag;
  wire  issue_units_1_io_iss_uops_0_is_br_or_jmp;
  wire  issue_units_1_io_iss_uops_0_is_jump;
  wire  issue_units_1_io_iss_uops_0_is_jal;
  wire  issue_units_1_io_iss_uops_0_is_ret;
  wire  issue_units_1_io_iss_uops_0_is_call;
  wire [7:0] issue_units_1_io_iss_uops_0_br_mask;
  wire [2:0] issue_units_1_io_iss_uops_0_br_tag;
  wire  issue_units_1_io_iss_uops_0_br_prediction_btb_blame;
  wire  issue_units_1_io_iss_uops_0_br_prediction_btb_hit;
  wire  issue_units_1_io_iss_uops_0_br_prediction_btb_taken;
  wire  issue_units_1_io_iss_uops_0_br_prediction_bpd_blame;
  wire  issue_units_1_io_iss_uops_0_br_prediction_bpd_hit;
  wire  issue_units_1_io_iss_uops_0_br_prediction_bpd_taken;
  wire [1:0] issue_units_1_io_iss_uops_0_br_prediction_bim_resp_value;
  wire [5:0] issue_units_1_io_iss_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_1_io_iss_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_info;
  wire  issue_units_1_io_iss_uops_0_stat_brjmp_mispredicted;
  wire  issue_units_1_io_iss_uops_0_stat_btb_made_pred;
  wire  issue_units_1_io_iss_uops_0_stat_btb_mispredicted;
  wire  issue_units_1_io_iss_uops_0_stat_bpd_made_pred;
  wire  issue_units_1_io_iss_uops_0_stat_bpd_mispredicted;
  wire [2:0] issue_units_1_io_iss_uops_0_fetch_pc_lob;
  wire [19:0] issue_units_1_io_iss_uops_0_imm_packed;
  wire [11:0] issue_units_1_io_iss_uops_0_csr_addr;
  wire [6:0] issue_units_1_io_iss_uops_0_rob_idx;
  wire [3:0] issue_units_1_io_iss_uops_0_ldq_idx;
  wire [3:0] issue_units_1_io_iss_uops_0_stq_idx;
  wire [5:0] issue_units_1_io_iss_uops_0_brob_idx;
  wire [6:0] issue_units_1_io_iss_uops_0_pdst;
  wire [6:0] issue_units_1_io_iss_uops_0_pop1;
  wire [6:0] issue_units_1_io_iss_uops_0_pop2;
  wire [6:0] issue_units_1_io_iss_uops_0_pop3;
  wire  issue_units_1_io_iss_uops_0_prs1_busy;
  wire  issue_units_1_io_iss_uops_0_prs2_busy;
  wire  issue_units_1_io_iss_uops_0_prs3_busy;
  wire [6:0] issue_units_1_io_iss_uops_0_stale_pdst;
  wire  issue_units_1_io_iss_uops_0_exception;
  wire [63:0] issue_units_1_io_iss_uops_0_exc_cause;
  wire  issue_units_1_io_iss_uops_0_bypassable;
  wire [4:0] issue_units_1_io_iss_uops_0_mem_cmd;
  wire [2:0] issue_units_1_io_iss_uops_0_mem_typ;
  wire  issue_units_1_io_iss_uops_0_is_fence;
  wire  issue_units_1_io_iss_uops_0_is_fencei;
  wire  issue_units_1_io_iss_uops_0_is_store;
  wire  issue_units_1_io_iss_uops_0_is_amo;
  wire  issue_units_1_io_iss_uops_0_is_load;
  wire  issue_units_1_io_iss_uops_0_is_sys_pc2epc;
  wire  issue_units_1_io_iss_uops_0_is_unique;
  wire  issue_units_1_io_iss_uops_0_flush_on_commit;
  wire [5:0] issue_units_1_io_iss_uops_0_ldst;
  wire [5:0] issue_units_1_io_iss_uops_0_lrs1;
  wire [5:0] issue_units_1_io_iss_uops_0_lrs2;
  wire [5:0] issue_units_1_io_iss_uops_0_lrs3;
  wire  issue_units_1_io_iss_uops_0_ldst_val;
  wire [1:0] issue_units_1_io_iss_uops_0_dst_rtype;
  wire [1:0] issue_units_1_io_iss_uops_0_lrs1_rtype;
  wire [1:0] issue_units_1_io_iss_uops_0_lrs2_rtype;
  wire  issue_units_1_io_iss_uops_0_frs3_en;
  wire  issue_units_1_io_iss_uops_0_fp_val;
  wire  issue_units_1_io_iss_uops_0_fp_single;
  wire  issue_units_1_io_iss_uops_0_xcpt_pf_if;
  wire  issue_units_1_io_iss_uops_0_xcpt_ae_if;
  wire  issue_units_1_io_iss_uops_0_replay_if;
  wire  issue_units_1_io_iss_uops_0_xcpt_ma_if;
  wire [63:0] issue_units_1_io_iss_uops_0_debug_wdata;
  wire [31:0] issue_units_1_io_iss_uops_0_debug_events_fetch_seq;
  wire  issue_units_1_io_iss_uops_1_valid;
  wire [1:0] issue_units_1_io_iss_uops_1_iw_state;
  wire [8:0] issue_units_1_io_iss_uops_1_uopc;
  wire [31:0] issue_units_1_io_iss_uops_1_inst;
  wire [39:0] issue_units_1_io_iss_uops_1_pc;
  wire [1:0] issue_units_1_io_iss_uops_1_iqtype;
  wire [9:0] issue_units_1_io_iss_uops_1_fu_code;
  wire  issue_units_1_io_iss_uops_1_allocate_brtag;
  wire  issue_units_1_io_iss_uops_1_is_br_or_jmp;
  wire  issue_units_1_io_iss_uops_1_is_jump;
  wire  issue_units_1_io_iss_uops_1_is_jal;
  wire  issue_units_1_io_iss_uops_1_is_ret;
  wire  issue_units_1_io_iss_uops_1_is_call;
  wire [7:0] issue_units_1_io_iss_uops_1_br_mask;
  wire [2:0] issue_units_1_io_iss_uops_1_br_tag;
  wire  issue_units_1_io_iss_uops_1_br_prediction_btb_blame;
  wire  issue_units_1_io_iss_uops_1_br_prediction_btb_hit;
  wire  issue_units_1_io_iss_uops_1_br_prediction_btb_taken;
  wire  issue_units_1_io_iss_uops_1_br_prediction_bpd_blame;
  wire  issue_units_1_io_iss_uops_1_br_prediction_bpd_hit;
  wire  issue_units_1_io_iss_uops_1_br_prediction_bpd_taken;
  wire [1:0] issue_units_1_io_iss_uops_1_br_prediction_bim_resp_value;
  wire [5:0] issue_units_1_io_iss_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] issue_units_1_io_iss_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_info;
  wire  issue_units_1_io_iss_uops_1_stat_brjmp_mispredicted;
  wire  issue_units_1_io_iss_uops_1_stat_btb_made_pred;
  wire  issue_units_1_io_iss_uops_1_stat_btb_mispredicted;
  wire  issue_units_1_io_iss_uops_1_stat_bpd_made_pred;
  wire  issue_units_1_io_iss_uops_1_stat_bpd_mispredicted;
  wire [2:0] issue_units_1_io_iss_uops_1_fetch_pc_lob;
  wire [19:0] issue_units_1_io_iss_uops_1_imm_packed;
  wire [11:0] issue_units_1_io_iss_uops_1_csr_addr;
  wire [6:0] issue_units_1_io_iss_uops_1_rob_idx;
  wire [3:0] issue_units_1_io_iss_uops_1_ldq_idx;
  wire [3:0] issue_units_1_io_iss_uops_1_stq_idx;
  wire [5:0] issue_units_1_io_iss_uops_1_brob_idx;
  wire [6:0] issue_units_1_io_iss_uops_1_pdst;
  wire [6:0] issue_units_1_io_iss_uops_1_pop1;
  wire [6:0] issue_units_1_io_iss_uops_1_pop2;
  wire [6:0] issue_units_1_io_iss_uops_1_pop3;
  wire  issue_units_1_io_iss_uops_1_prs1_busy;
  wire  issue_units_1_io_iss_uops_1_prs2_busy;
  wire  issue_units_1_io_iss_uops_1_prs3_busy;
  wire [6:0] issue_units_1_io_iss_uops_1_stale_pdst;
  wire  issue_units_1_io_iss_uops_1_exception;
  wire [63:0] issue_units_1_io_iss_uops_1_exc_cause;
  wire  issue_units_1_io_iss_uops_1_bypassable;
  wire [4:0] issue_units_1_io_iss_uops_1_mem_cmd;
  wire [2:0] issue_units_1_io_iss_uops_1_mem_typ;
  wire  issue_units_1_io_iss_uops_1_is_fence;
  wire  issue_units_1_io_iss_uops_1_is_fencei;
  wire  issue_units_1_io_iss_uops_1_is_store;
  wire  issue_units_1_io_iss_uops_1_is_amo;
  wire  issue_units_1_io_iss_uops_1_is_load;
  wire  issue_units_1_io_iss_uops_1_is_sys_pc2epc;
  wire  issue_units_1_io_iss_uops_1_is_unique;
  wire  issue_units_1_io_iss_uops_1_flush_on_commit;
  wire [5:0] issue_units_1_io_iss_uops_1_ldst;
  wire [5:0] issue_units_1_io_iss_uops_1_lrs1;
  wire [5:0] issue_units_1_io_iss_uops_1_lrs2;
  wire [5:0] issue_units_1_io_iss_uops_1_lrs3;
  wire  issue_units_1_io_iss_uops_1_ldst_val;
  wire [1:0] issue_units_1_io_iss_uops_1_dst_rtype;
  wire [1:0] issue_units_1_io_iss_uops_1_lrs1_rtype;
  wire [1:0] issue_units_1_io_iss_uops_1_lrs2_rtype;
  wire  issue_units_1_io_iss_uops_1_frs3_en;
  wire  issue_units_1_io_iss_uops_1_fp_val;
  wire  issue_units_1_io_iss_uops_1_fp_single;
  wire  issue_units_1_io_iss_uops_1_xcpt_pf_if;
  wire  issue_units_1_io_iss_uops_1_xcpt_ae_if;
  wire  issue_units_1_io_iss_uops_1_replay_if;
  wire  issue_units_1_io_iss_uops_1_xcpt_ma_if;
  wire [63:0] issue_units_1_io_iss_uops_1_debug_wdata;
  wire [31:0] issue_units_1_io_iss_uops_1_debug_events_fetch_seq;
  wire  issue_units_1_io_wakeup_pdsts_0_valid;
  wire [6:0] issue_units_1_io_wakeup_pdsts_0_bits;
  wire  issue_units_1_io_wakeup_pdsts_1_valid;
  wire [6:0] issue_units_1_io_wakeup_pdsts_1_bits;
  wire  issue_units_1_io_wakeup_pdsts_2_valid;
  wire [6:0] issue_units_1_io_wakeup_pdsts_2_bits;
  wire  issue_units_1_io_wakeup_pdsts_3_valid;
  wire [6:0] issue_units_1_io_wakeup_pdsts_3_bits;
  wire  issue_units_1_io_wakeup_pdsts_4_valid;
  wire [6:0] issue_units_1_io_wakeup_pdsts_4_bits;
  wire [9:0] issue_units_1_io_fu_types_0;
  wire  issue_units_1_io_brinfo_valid;
  wire  issue_units_1_io_brinfo_mispredict;
  wire [7:0] issue_units_1_io_brinfo_mask;
  wire  issue_units_1_io_flush_pipeline;
  wire  iregfile_clock;
  wire [6:0] iregfile_io_read_ports_0_addr;
  wire [63:0] iregfile_io_read_ports_0_data;
  wire [6:0] iregfile_io_read_ports_1_addr;
  wire [63:0] iregfile_io_read_ports_1_data;
  wire [6:0] iregfile_io_read_ports_2_addr;
  wire [63:0] iregfile_io_read_ports_2_data;
  wire [6:0] iregfile_io_read_ports_3_addr;
  wire [63:0] iregfile_io_read_ports_3_data;
  wire [6:0] iregfile_io_read_ports_4_addr;
  wire [63:0] iregfile_io_read_ports_4_data;
  wire [6:0] iregfile_io_read_ports_5_addr;
  wire [63:0] iregfile_io_read_ports_5_data;
  wire  iregfile_io_write_ports_0_valid;
  wire [6:0] iregfile_io_write_ports_0_bits_addr;
  wire [63:0] iregfile_io_write_ports_0_bits_data;
  wire  iregfile_io_write_ports_1_valid;
  wire [6:0] iregfile_io_write_ports_1_bits_addr;
  wire [63:0] iregfile_io_write_ports_1_bits_data;
  wire  iregfile_io_write_ports_2_valid;
  wire [6:0] iregfile_io_write_ports_2_bits_addr;
  wire [63:0] iregfile_io_write_ports_2_bits_data;
  wire  ll_wbarb_io_in_0_valid;
  wire [6:0] ll_wbarb_io_in_0_bits_uop_rob_idx;
  wire [6:0] ll_wbarb_io_in_0_bits_uop_pdst;
  wire  ll_wbarb_io_in_0_bits_uop_is_store;
  wire  ll_wbarb_io_in_0_bits_uop_is_amo;
  wire [1:0] ll_wbarb_io_in_0_bits_uop_dst_rtype;
  wire [63:0] ll_wbarb_io_in_0_bits_data;
  wire  ll_wbarb_io_in_1_ready;
  wire  ll_wbarb_io_in_1_valid;
  wire [6:0] ll_wbarb_io_in_1_bits_uop_rob_idx;
  wire [6:0] ll_wbarb_io_in_1_bits_uop_pdst;
  wire  ll_wbarb_io_in_1_bits_uop_is_store;
  wire  ll_wbarb_io_in_1_bits_uop_is_amo;
  wire [1:0] ll_wbarb_io_in_1_bits_uop_dst_rtype;
  wire [63:0] ll_wbarb_io_in_1_bits_data;
  wire  ll_wbarb_io_out_ready;
  wire  ll_wbarb_io_out_valid;
  wire [6:0] ll_wbarb_io_out_bits_uop_rob_idx;
  wire [6:0] ll_wbarb_io_out_bits_uop_pdst;
  wire  ll_wbarb_io_out_bits_uop_is_store;
  wire  ll_wbarb_io_out_bits_uop_is_amo;
  wire [1:0] ll_wbarb_io_out_bits_uop_dst_rtype;
  wire [63:0] ll_wbarb_io_out_bits_data;
  wire  iregister_read_clock;
  wire  iregister_read_reset;
  wire  iregister_read_io_iss_valids_0;
  wire  iregister_read_io_iss_valids_1;
  wire  iregister_read_io_iss_valids_2;
  wire [8:0] iregister_read_io_iss_uops_0_uopc;
  wire [7:0] iregister_read_io_iss_uops_0_br_mask;
  wire [19:0] iregister_read_io_iss_uops_0_imm_packed;
  wire [6:0] iregister_read_io_iss_uops_0_rob_idx;
  wire [3:0] iregister_read_io_iss_uops_0_ldq_idx;
  wire [3:0] iregister_read_io_iss_uops_0_stq_idx;
  wire [6:0] iregister_read_io_iss_uops_0_pdst;
  wire [6:0] iregister_read_io_iss_uops_0_pop1;
  wire [6:0] iregister_read_io_iss_uops_0_pop2;
  wire [4:0] iregister_read_io_iss_uops_0_mem_cmd;
  wire [2:0] iregister_read_io_iss_uops_0_mem_typ;
  wire  iregister_read_io_iss_uops_0_is_fence;
  wire  iregister_read_io_iss_uops_0_is_store;
  wire  iregister_read_io_iss_uops_0_is_amo;
  wire  iregister_read_io_iss_uops_0_is_load;
  wire [1:0] iregister_read_io_iss_uops_0_dst_rtype;
  wire [1:0] iregister_read_io_iss_uops_0_lrs1_rtype;
  wire [1:0] iregister_read_io_iss_uops_0_lrs2_rtype;
  wire  iregister_read_io_iss_uops_0_fp_val;
  wire  iregister_read_io_iss_uops_1_valid;
  wire [1:0] iregister_read_io_iss_uops_1_iw_state;
  wire [8:0] iregister_read_io_iss_uops_1_uopc;
  wire [31:0] iregister_read_io_iss_uops_1_inst;
  wire [39:0] iregister_read_io_iss_uops_1_pc;
  wire [1:0] iregister_read_io_iss_uops_1_iqtype;
  wire [9:0] iregister_read_io_iss_uops_1_fu_code;
  wire  iregister_read_io_iss_uops_1_allocate_brtag;
  wire  iregister_read_io_iss_uops_1_is_br_or_jmp;
  wire  iregister_read_io_iss_uops_1_is_jump;
  wire  iregister_read_io_iss_uops_1_is_jal;
  wire  iregister_read_io_iss_uops_1_is_ret;
  wire  iregister_read_io_iss_uops_1_is_call;
  wire [7:0] iregister_read_io_iss_uops_1_br_mask;
  wire [2:0] iregister_read_io_iss_uops_1_br_tag;
  wire  iregister_read_io_iss_uops_1_br_prediction_btb_blame;
  wire  iregister_read_io_iss_uops_1_br_prediction_btb_hit;
  wire  iregister_read_io_iss_uops_1_br_prediction_btb_taken;
  wire  iregister_read_io_iss_uops_1_br_prediction_bpd_blame;
  wire  iregister_read_io_iss_uops_1_br_prediction_bpd_hit;
  wire  iregister_read_io_iss_uops_1_br_prediction_bpd_taken;
  wire [1:0] iregister_read_io_iss_uops_1_br_prediction_bim_resp_value;
  wire [5:0] iregister_read_io_iss_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] iregister_read_io_iss_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] iregister_read_io_iss_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iregister_read_io_iss_uops_1_br_prediction_bpd_resp_info;
  wire  iregister_read_io_iss_uops_1_stat_brjmp_mispredicted;
  wire  iregister_read_io_iss_uops_1_stat_btb_made_pred;
  wire  iregister_read_io_iss_uops_1_stat_btb_mispredicted;
  wire  iregister_read_io_iss_uops_1_stat_bpd_made_pred;
  wire  iregister_read_io_iss_uops_1_stat_bpd_mispredicted;
  wire [2:0] iregister_read_io_iss_uops_1_fetch_pc_lob;
  wire [19:0] iregister_read_io_iss_uops_1_imm_packed;
  wire [11:0] iregister_read_io_iss_uops_1_csr_addr;
  wire [6:0] iregister_read_io_iss_uops_1_rob_idx;
  wire [3:0] iregister_read_io_iss_uops_1_ldq_idx;
  wire [3:0] iregister_read_io_iss_uops_1_stq_idx;
  wire [5:0] iregister_read_io_iss_uops_1_brob_idx;
  wire [6:0] iregister_read_io_iss_uops_1_pdst;
  wire [6:0] iregister_read_io_iss_uops_1_pop1;
  wire [6:0] iregister_read_io_iss_uops_1_pop2;
  wire [6:0] iregister_read_io_iss_uops_1_pop3;
  wire  iregister_read_io_iss_uops_1_prs1_busy;
  wire  iregister_read_io_iss_uops_1_prs2_busy;
  wire  iregister_read_io_iss_uops_1_prs3_busy;
  wire [6:0] iregister_read_io_iss_uops_1_stale_pdst;
  wire  iregister_read_io_iss_uops_1_exception;
  wire [63:0] iregister_read_io_iss_uops_1_exc_cause;
  wire  iregister_read_io_iss_uops_1_bypassable;
  wire [4:0] iregister_read_io_iss_uops_1_mem_cmd;
  wire [2:0] iregister_read_io_iss_uops_1_mem_typ;
  wire  iregister_read_io_iss_uops_1_is_fence;
  wire  iregister_read_io_iss_uops_1_is_fencei;
  wire  iregister_read_io_iss_uops_1_is_store;
  wire  iregister_read_io_iss_uops_1_is_amo;
  wire  iregister_read_io_iss_uops_1_is_load;
  wire  iregister_read_io_iss_uops_1_is_sys_pc2epc;
  wire  iregister_read_io_iss_uops_1_is_unique;
  wire  iregister_read_io_iss_uops_1_flush_on_commit;
  wire [5:0] iregister_read_io_iss_uops_1_ldst;
  wire [5:0] iregister_read_io_iss_uops_1_lrs1;
  wire [5:0] iregister_read_io_iss_uops_1_lrs2;
  wire [5:0] iregister_read_io_iss_uops_1_lrs3;
  wire  iregister_read_io_iss_uops_1_ldst_val;
  wire [1:0] iregister_read_io_iss_uops_1_dst_rtype;
  wire [1:0] iregister_read_io_iss_uops_1_lrs1_rtype;
  wire [1:0] iregister_read_io_iss_uops_1_lrs2_rtype;
  wire  iregister_read_io_iss_uops_1_frs3_en;
  wire  iregister_read_io_iss_uops_1_fp_val;
  wire  iregister_read_io_iss_uops_1_fp_single;
  wire  iregister_read_io_iss_uops_1_xcpt_pf_if;
  wire  iregister_read_io_iss_uops_1_xcpt_ae_if;
  wire  iregister_read_io_iss_uops_1_replay_if;
  wire  iregister_read_io_iss_uops_1_xcpt_ma_if;
  wire [63:0] iregister_read_io_iss_uops_1_debug_wdata;
  wire [31:0] iregister_read_io_iss_uops_1_debug_events_fetch_seq;
  wire  iregister_read_io_iss_uops_2_valid;
  wire [1:0] iregister_read_io_iss_uops_2_iw_state;
  wire [8:0] iregister_read_io_iss_uops_2_uopc;
  wire [31:0] iregister_read_io_iss_uops_2_inst;
  wire [39:0] iregister_read_io_iss_uops_2_pc;
  wire [1:0] iregister_read_io_iss_uops_2_iqtype;
  wire [9:0] iregister_read_io_iss_uops_2_fu_code;
  wire  iregister_read_io_iss_uops_2_allocate_brtag;
  wire  iregister_read_io_iss_uops_2_is_br_or_jmp;
  wire  iregister_read_io_iss_uops_2_is_jump;
  wire  iregister_read_io_iss_uops_2_is_jal;
  wire  iregister_read_io_iss_uops_2_is_ret;
  wire  iregister_read_io_iss_uops_2_is_call;
  wire [7:0] iregister_read_io_iss_uops_2_br_mask;
  wire [2:0] iregister_read_io_iss_uops_2_br_tag;
  wire  iregister_read_io_iss_uops_2_br_prediction_btb_blame;
  wire  iregister_read_io_iss_uops_2_br_prediction_btb_hit;
  wire  iregister_read_io_iss_uops_2_br_prediction_btb_taken;
  wire  iregister_read_io_iss_uops_2_br_prediction_bpd_blame;
  wire  iregister_read_io_iss_uops_2_br_prediction_bpd_hit;
  wire  iregister_read_io_iss_uops_2_br_prediction_bpd_taken;
  wire [1:0] iregister_read_io_iss_uops_2_br_prediction_bim_resp_value;
  wire [5:0] iregister_read_io_iss_uops_2_br_prediction_bim_resp_entry_idx;
  wire [1:0] iregister_read_io_iss_uops_2_br_prediction_bim_resp_way_idx;
  wire [1:0] iregister_read_io_iss_uops_2_br_prediction_bpd_resp_takens;
  wire [14:0] iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history;
  wire [14:0] iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_u;
  wire [7:0] iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iregister_read_io_iss_uops_2_br_prediction_bpd_resp_info;
  wire  iregister_read_io_iss_uops_2_stat_brjmp_mispredicted;
  wire  iregister_read_io_iss_uops_2_stat_btb_made_pred;
  wire  iregister_read_io_iss_uops_2_stat_btb_mispredicted;
  wire  iregister_read_io_iss_uops_2_stat_bpd_made_pred;
  wire  iregister_read_io_iss_uops_2_stat_bpd_mispredicted;
  wire [2:0] iregister_read_io_iss_uops_2_fetch_pc_lob;
  wire [19:0] iregister_read_io_iss_uops_2_imm_packed;
  wire [11:0] iregister_read_io_iss_uops_2_csr_addr;
  wire [6:0] iregister_read_io_iss_uops_2_rob_idx;
  wire [3:0] iregister_read_io_iss_uops_2_ldq_idx;
  wire [3:0] iregister_read_io_iss_uops_2_stq_idx;
  wire [5:0] iregister_read_io_iss_uops_2_brob_idx;
  wire [6:0] iregister_read_io_iss_uops_2_pdst;
  wire [6:0] iregister_read_io_iss_uops_2_pop1;
  wire [6:0] iregister_read_io_iss_uops_2_pop2;
  wire [6:0] iregister_read_io_iss_uops_2_pop3;
  wire  iregister_read_io_iss_uops_2_prs1_busy;
  wire  iregister_read_io_iss_uops_2_prs2_busy;
  wire  iregister_read_io_iss_uops_2_prs3_busy;
  wire [6:0] iregister_read_io_iss_uops_2_stale_pdst;
  wire  iregister_read_io_iss_uops_2_exception;
  wire [63:0] iregister_read_io_iss_uops_2_exc_cause;
  wire  iregister_read_io_iss_uops_2_bypassable;
  wire [4:0] iregister_read_io_iss_uops_2_mem_cmd;
  wire [2:0] iregister_read_io_iss_uops_2_mem_typ;
  wire  iregister_read_io_iss_uops_2_is_fence;
  wire  iregister_read_io_iss_uops_2_is_fencei;
  wire  iregister_read_io_iss_uops_2_is_store;
  wire  iregister_read_io_iss_uops_2_is_amo;
  wire  iregister_read_io_iss_uops_2_is_load;
  wire  iregister_read_io_iss_uops_2_is_sys_pc2epc;
  wire  iregister_read_io_iss_uops_2_is_unique;
  wire  iregister_read_io_iss_uops_2_flush_on_commit;
  wire [5:0] iregister_read_io_iss_uops_2_ldst;
  wire [5:0] iregister_read_io_iss_uops_2_lrs1;
  wire [5:0] iregister_read_io_iss_uops_2_lrs2;
  wire [5:0] iregister_read_io_iss_uops_2_lrs3;
  wire  iregister_read_io_iss_uops_2_ldst_val;
  wire [1:0] iregister_read_io_iss_uops_2_dst_rtype;
  wire [1:0] iregister_read_io_iss_uops_2_lrs1_rtype;
  wire [1:0] iregister_read_io_iss_uops_2_lrs2_rtype;
  wire  iregister_read_io_iss_uops_2_frs3_en;
  wire  iregister_read_io_iss_uops_2_fp_val;
  wire  iregister_read_io_iss_uops_2_fp_single;
  wire  iregister_read_io_iss_uops_2_xcpt_pf_if;
  wire  iregister_read_io_iss_uops_2_xcpt_ae_if;
  wire  iregister_read_io_iss_uops_2_replay_if;
  wire  iregister_read_io_iss_uops_2_xcpt_ma_if;
  wire [63:0] iregister_read_io_iss_uops_2_debug_wdata;
  wire [31:0] iregister_read_io_iss_uops_2_debug_events_fetch_seq;
  wire [6:0] iregister_read_io_rf_read_ports_0_addr;
  wire [63:0] iregister_read_io_rf_read_ports_0_data;
  wire [6:0] iregister_read_io_rf_read_ports_1_addr;
  wire [63:0] iregister_read_io_rf_read_ports_1_data;
  wire [6:0] iregister_read_io_rf_read_ports_2_addr;
  wire [63:0] iregister_read_io_rf_read_ports_2_data;
  wire [6:0] iregister_read_io_rf_read_ports_3_addr;
  wire [63:0] iregister_read_io_rf_read_ports_3_data;
  wire [6:0] iregister_read_io_rf_read_ports_4_addr;
  wire [63:0] iregister_read_io_rf_read_ports_4_data;
  wire [6:0] iregister_read_io_rf_read_ports_5_addr;
  wire [63:0] iregister_read_io_rf_read_ports_5_data;
  wire  iregister_read_io_bypass_valid_0;
  wire  iregister_read_io_bypass_valid_1;
  wire  iregister_read_io_bypass_valid_2;
  wire  iregister_read_io_bypass_valid_3;
  wire  iregister_read_io_bypass_uop_0_ctrl_rf_wen;
  wire [6:0] iregister_read_io_bypass_uop_0_pdst;
  wire [1:0] iregister_read_io_bypass_uop_0_dst_rtype;
  wire  iregister_read_io_bypass_uop_1_ctrl_rf_wen;
  wire [6:0] iregister_read_io_bypass_uop_1_pdst;
  wire [1:0] iregister_read_io_bypass_uop_1_dst_rtype;
  wire  iregister_read_io_bypass_uop_2_ctrl_rf_wen;
  wire [6:0] iregister_read_io_bypass_uop_2_pdst;
  wire [1:0] iregister_read_io_bypass_uop_2_dst_rtype;
  wire  iregister_read_io_bypass_uop_3_ctrl_rf_wen;
  wire [6:0] iregister_read_io_bypass_uop_3_pdst;
  wire [1:0] iregister_read_io_bypass_uop_3_dst_rtype;
  wire [63:0] iregister_read_io_bypass_data_0;
  wire [63:0] iregister_read_io_bypass_data_1;
  wire [63:0] iregister_read_io_bypass_data_2;
  wire [63:0] iregister_read_io_bypass_data_3;
  wire  iregister_read_io_exe_reqs_0_valid;
  wire [8:0] iregister_read_io_exe_reqs_0_bits_uop_uopc;
  wire  iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_load;
  wire  iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_sta;
  wire  iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_std;
  wire [7:0] iregister_read_io_exe_reqs_0_bits_uop_br_mask;
  wire [19:0] iregister_read_io_exe_reqs_0_bits_uop_imm_packed;
  wire [6:0] iregister_read_io_exe_reqs_0_bits_uop_rob_idx;
  wire [3:0] iregister_read_io_exe_reqs_0_bits_uop_ldq_idx;
  wire [3:0] iregister_read_io_exe_reqs_0_bits_uop_stq_idx;
  wire [6:0] iregister_read_io_exe_reqs_0_bits_uop_pdst;
  wire [4:0] iregister_read_io_exe_reqs_0_bits_uop_mem_cmd;
  wire [2:0] iregister_read_io_exe_reqs_0_bits_uop_mem_typ;
  wire  iregister_read_io_exe_reqs_0_bits_uop_is_fence;
  wire  iregister_read_io_exe_reqs_0_bits_uop_is_store;
  wire  iregister_read_io_exe_reqs_0_bits_uop_is_amo;
  wire  iregister_read_io_exe_reqs_0_bits_uop_is_load;
  wire [1:0] iregister_read_io_exe_reqs_0_bits_uop_dst_rtype;
  wire  iregister_read_io_exe_reqs_0_bits_uop_fp_val;
  wire [63:0] iregister_read_io_exe_reqs_0_bits_rs1_data;
  wire [63:0] iregister_read_io_exe_reqs_0_bits_rs2_data;
  wire  iregister_read_io_exe_reqs_1_valid;
  wire  iregister_read_io_exe_reqs_1_bits_uop_valid;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_iw_state;
  wire [8:0] iregister_read_io_exe_reqs_1_bits_uop_uopc;
  wire [31:0] iregister_read_io_exe_reqs_1_bits_uop_inst;
  wire [39:0] iregister_read_io_exe_reqs_1_bits_uop_pc;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_iqtype;
  wire [9:0] iregister_read_io_exe_reqs_1_bits_uop_fu_code;
  wire [3:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_br_type;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_op1_sel;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_op2_sel;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_imm_sel;
  wire [3:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_op_fcn;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ctrl_fcn_dw;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ctrl_rf_wen;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_ctrl_csr_cmd;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_load;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_sta;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_std;
  wire  iregister_read_io_exe_reqs_1_bits_uop_allocate_brtag;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_br_or_jmp;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_jump;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_jal;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_ret;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_call;
  wire [7:0] iregister_read_io_exe_reqs_1_bits_uop_br_mask;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_br_tag;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_blame;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_hit;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_taken;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_blame;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_hit;
  wire  iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_taken;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_value;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_takens;
  wire [14:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history;
  wire [14:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_info;
  wire  iregister_read_io_exe_reqs_1_bits_uop_stat_brjmp_mispredicted;
  wire  iregister_read_io_exe_reqs_1_bits_uop_stat_btb_made_pred;
  wire  iregister_read_io_exe_reqs_1_bits_uop_stat_btb_mispredicted;
  wire  iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_made_pred;
  wire  iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_mispredicted;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_fetch_pc_lob;
  wire [19:0] iregister_read_io_exe_reqs_1_bits_uop_imm_packed;
  wire [11:0] iregister_read_io_exe_reqs_1_bits_uop_csr_addr;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_rob_idx;
  wire [3:0] iregister_read_io_exe_reqs_1_bits_uop_ldq_idx;
  wire [3:0] iregister_read_io_exe_reqs_1_bits_uop_stq_idx;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_brob_idx;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_pdst;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_pop1;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_pop2;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_pop3;
  wire  iregister_read_io_exe_reqs_1_bits_uop_prs1_busy;
  wire  iregister_read_io_exe_reqs_1_bits_uop_prs2_busy;
  wire  iregister_read_io_exe_reqs_1_bits_uop_prs3_busy;
  wire [6:0] iregister_read_io_exe_reqs_1_bits_uop_stale_pdst;
  wire  iregister_read_io_exe_reqs_1_bits_uop_exception;
  wire [63:0] iregister_read_io_exe_reqs_1_bits_uop_exc_cause;
  wire  iregister_read_io_exe_reqs_1_bits_uop_bypassable;
  wire [4:0] iregister_read_io_exe_reqs_1_bits_uop_mem_cmd;
  wire [2:0] iregister_read_io_exe_reqs_1_bits_uop_mem_typ;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_fence;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_fencei;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_store;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_amo;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_load;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_sys_pc2epc;
  wire  iregister_read_io_exe_reqs_1_bits_uop_is_unique;
  wire  iregister_read_io_exe_reqs_1_bits_uop_flush_on_commit;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_ldst;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_lrs1;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_lrs2;
  wire [5:0] iregister_read_io_exe_reqs_1_bits_uop_lrs3;
  wire  iregister_read_io_exe_reqs_1_bits_uop_ldst_val;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_dst_rtype;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_lrs1_rtype;
  wire [1:0] iregister_read_io_exe_reqs_1_bits_uop_lrs2_rtype;
  wire  iregister_read_io_exe_reqs_1_bits_uop_frs3_en;
  wire  iregister_read_io_exe_reqs_1_bits_uop_fp_val;
  wire  iregister_read_io_exe_reqs_1_bits_uop_fp_single;
  wire  iregister_read_io_exe_reqs_1_bits_uop_xcpt_pf_if;
  wire  iregister_read_io_exe_reqs_1_bits_uop_xcpt_ae_if;
  wire  iregister_read_io_exe_reqs_1_bits_uop_replay_if;
  wire  iregister_read_io_exe_reqs_1_bits_uop_xcpt_ma_if;
  wire [63:0] iregister_read_io_exe_reqs_1_bits_uop_debug_wdata;
  wire [31:0] iregister_read_io_exe_reqs_1_bits_uop_debug_events_fetch_seq;
  wire [63:0] iregister_read_io_exe_reqs_1_bits_rs1_data;
  wire [63:0] iregister_read_io_exe_reqs_1_bits_rs2_data;
  wire  iregister_read_io_exe_reqs_2_valid;
  wire  iregister_read_io_exe_reqs_2_bits_uop_valid;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_iw_state;
  wire [8:0] iregister_read_io_exe_reqs_2_bits_uop_uopc;
  wire [31:0] iregister_read_io_exe_reqs_2_bits_uop_inst;
  wire [39:0] iregister_read_io_exe_reqs_2_bits_uop_pc;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_iqtype;
  wire [9:0] iregister_read_io_exe_reqs_2_bits_uop_fu_code;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_ctrl_op1_sel;
  wire [2:0] iregister_read_io_exe_reqs_2_bits_uop_ctrl_op2_sel;
  wire [2:0] iregister_read_io_exe_reqs_2_bits_uop_ctrl_imm_sel;
  wire [3:0] iregister_read_io_exe_reqs_2_bits_uop_ctrl_op_fcn;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ctrl_fcn_dw;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ctrl_rf_wen;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_load;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_sta;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_std;
  wire  iregister_read_io_exe_reqs_2_bits_uop_allocate_brtag;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_br_or_jmp;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_jump;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_jal;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_ret;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_call;
  wire [7:0] iregister_read_io_exe_reqs_2_bits_uop_br_mask;
  wire [2:0] iregister_read_io_exe_reqs_2_bits_uop_br_tag;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_blame;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_hit;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_taken;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_blame;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_hit;
  wire  iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_taken;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_value;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_entry_idx;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_way_idx;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_takens;
  wire [14:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history;
  wire [14:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_u;
  wire [7:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_info;
  wire  iregister_read_io_exe_reqs_2_bits_uop_stat_brjmp_mispredicted;
  wire  iregister_read_io_exe_reqs_2_bits_uop_stat_btb_made_pred;
  wire  iregister_read_io_exe_reqs_2_bits_uop_stat_btb_mispredicted;
  wire  iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_made_pred;
  wire  iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_mispredicted;
  wire [2:0] iregister_read_io_exe_reqs_2_bits_uop_fetch_pc_lob;
  wire [19:0] iregister_read_io_exe_reqs_2_bits_uop_imm_packed;
  wire [11:0] iregister_read_io_exe_reqs_2_bits_uop_csr_addr;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_rob_idx;
  wire [3:0] iregister_read_io_exe_reqs_2_bits_uop_ldq_idx;
  wire [3:0] iregister_read_io_exe_reqs_2_bits_uop_stq_idx;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_brob_idx;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_pdst;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_pop1;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_pop2;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_pop3;
  wire  iregister_read_io_exe_reqs_2_bits_uop_prs1_busy;
  wire  iregister_read_io_exe_reqs_2_bits_uop_prs2_busy;
  wire  iregister_read_io_exe_reqs_2_bits_uop_prs3_busy;
  wire [6:0] iregister_read_io_exe_reqs_2_bits_uop_stale_pdst;
  wire  iregister_read_io_exe_reqs_2_bits_uop_exception;
  wire [63:0] iregister_read_io_exe_reqs_2_bits_uop_exc_cause;
  wire  iregister_read_io_exe_reqs_2_bits_uop_bypassable;
  wire [4:0] iregister_read_io_exe_reqs_2_bits_uop_mem_cmd;
  wire [2:0] iregister_read_io_exe_reqs_2_bits_uop_mem_typ;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_fence;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_fencei;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_store;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_amo;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_load;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_sys_pc2epc;
  wire  iregister_read_io_exe_reqs_2_bits_uop_is_unique;
  wire  iregister_read_io_exe_reqs_2_bits_uop_flush_on_commit;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_ldst;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_lrs1;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_lrs2;
  wire [5:0] iregister_read_io_exe_reqs_2_bits_uop_lrs3;
  wire  iregister_read_io_exe_reqs_2_bits_uop_ldst_val;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_dst_rtype;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_lrs1_rtype;
  wire [1:0] iregister_read_io_exe_reqs_2_bits_uop_lrs2_rtype;
  wire  iregister_read_io_exe_reqs_2_bits_uop_frs3_en;
  wire  iregister_read_io_exe_reqs_2_bits_uop_fp_val;
  wire  iregister_read_io_exe_reqs_2_bits_uop_fp_single;
  wire  iregister_read_io_exe_reqs_2_bits_uop_xcpt_pf_if;
  wire  iregister_read_io_exe_reqs_2_bits_uop_xcpt_ae_if;
  wire  iregister_read_io_exe_reqs_2_bits_uop_replay_if;
  wire  iregister_read_io_exe_reqs_2_bits_uop_xcpt_ma_if;
  wire [63:0] iregister_read_io_exe_reqs_2_bits_uop_debug_wdata;
  wire [31:0] iregister_read_io_exe_reqs_2_bits_uop_debug_events_fetch_seq;
  wire [63:0] iregister_read_io_exe_reqs_2_bits_rs1_data;
  wire [63:0] iregister_read_io_exe_reqs_2_bits_rs2_data;
  wire  iregister_read_io_kill;
  wire  iregister_read_io_brinfo_valid;
  wire  iregister_read_io_brinfo_mispredict;
  wire [7:0] iregister_read_io_brinfo_mask;
  wire  dc_shim_clock;
  wire  dc_shim_reset;
  wire  dc_shim_io_core_req_valid;
  wire [39:0] dc_shim_io_core_req_bits_addr;
  wire [8:0] dc_shim_io_core_req_bits_uop_uopc;
  wire [7:0] dc_shim_io_core_req_bits_uop_br_mask;
  wire [6:0] dc_shim_io_core_req_bits_uop_rob_idx;
  wire [3:0] dc_shim_io_core_req_bits_uop_ldq_idx;
  wire [3:0] dc_shim_io_core_req_bits_uop_stq_idx;
  wire [6:0] dc_shim_io_core_req_bits_uop_pdst;
  wire [4:0] dc_shim_io_core_req_bits_uop_mem_cmd;
  wire [2:0] dc_shim_io_core_req_bits_uop_mem_typ;
  wire  dc_shim_io_core_req_bits_uop_is_store;
  wire  dc_shim_io_core_req_bits_uop_is_amo;
  wire  dc_shim_io_core_req_bits_uop_is_load;
  wire [1:0] dc_shim_io_core_req_bits_uop_dst_rtype;
  wire  dc_shim_io_core_req_bits_uop_fp_val;
  wire [63:0] dc_shim_io_core_req_bits_data;
  wire  dc_shim_io_core_req_bits_kill;
  wire  dc_shim_io_core_resp_valid;
  wire [63:0] dc_shim_io_core_resp_bits_data_subword;
  wire [8:0] dc_shim_io_core_resp_bits_uop_uopc;
  wire [6:0] dc_shim_io_core_resp_bits_uop_rob_idx;
  wire [3:0] dc_shim_io_core_resp_bits_uop_ldq_idx;
  wire [3:0] dc_shim_io_core_resp_bits_uop_stq_idx;
  wire [6:0] dc_shim_io_core_resp_bits_uop_pdst;
  wire [4:0] dc_shim_io_core_resp_bits_uop_mem_cmd;
  wire [2:0] dc_shim_io_core_resp_bits_uop_mem_typ;
  wire  dc_shim_io_core_resp_bits_uop_is_store;
  wire  dc_shim_io_core_resp_bits_uop_is_amo;
  wire  dc_shim_io_core_resp_bits_uop_is_load;
  wire [1:0] dc_shim_io_core_resp_bits_uop_dst_rtype;
  wire  dc_shim_io_core_resp_bits_uop_fp_val;
  wire  dc_shim_io_core_brinfo_valid;
  wire  dc_shim_io_core_brinfo_mispredict;
  wire [7:0] dc_shim_io_core_brinfo_mask;
  wire  dc_shim_io_core_nack_valid;
  wire [3:0] dc_shim_io_core_nack_lsu_idx;
  wire  dc_shim_io_core_nack_isload;
  wire  dc_shim_io_core_nack_cache_nack;
  wire  dc_shim_io_core_flush_pipe;
  wire  dc_shim_io_core_invalidate_lr;
  wire  dc_shim_io_core_ordered;
  wire  dc_shim_io_dmem_req_ready;
  wire  dc_shim_io_dmem_req_valid;
  wire [39:0] dc_shim_io_dmem_req_bits_addr;
  wire [6:0] dc_shim_io_dmem_req_bits_tag;
  wire [4:0] dc_shim_io_dmem_req_bits_cmd;
  wire [2:0] dc_shim_io_dmem_req_bits_typ;
  wire  dc_shim_io_dmem_s1_kill;
  wire [63:0] dc_shim_io_dmem_s1_data_data;
  wire  dc_shim_io_dmem_s2_nack;
  wire  dc_shim_io_dmem_resp_valid;
  wire [6:0] dc_shim_io_dmem_resp_bits_tag;
  wire [63:0] dc_shim_io_dmem_resp_bits_data;
  wire  dc_shim_io_dmem_resp_bits_has_data;
  wire  dc_shim_io_dmem_s2_xcpt_ma_ld;
  wire  dc_shim_io_dmem_s2_xcpt_ma_st;
  wire  dc_shim_io_dmem_s2_xcpt_pf_ld;
  wire  dc_shim_io_dmem_s2_xcpt_pf_st;
  wire  dc_shim_io_dmem_invalidate_lr;
  wire  dc_shim_io_dmem_ordered;
  wire  lsu_clock;
  wire  lsu_reset;
  wire  lsu_io_dec_st_vals_0;
  wire  lsu_io_dec_st_vals_1;
  wire  lsu_io_dec_ld_vals_0;
  wire  lsu_io_dec_ld_vals_1;
  wire [8:0] lsu_io_dec_uops_0_uopc;
  wire [7:0] lsu_io_dec_uops_0_br_mask;
  wire [6:0] lsu_io_dec_uops_0_rob_idx;
  wire [3:0] lsu_io_dec_uops_0_ldq_idx;
  wire [3:0] lsu_io_dec_uops_0_stq_idx;
  wire [4:0] lsu_io_dec_uops_0_mem_cmd;
  wire [2:0] lsu_io_dec_uops_0_mem_typ;
  wire  lsu_io_dec_uops_0_is_fence;
  wire  lsu_io_dec_uops_0_is_store;
  wire  lsu_io_dec_uops_0_is_amo;
  wire  lsu_io_dec_uops_0_is_load;
  wire [1:0] lsu_io_dec_uops_0_dst_rtype;
  wire  lsu_io_dec_uops_0_fp_val;
  wire [8:0] lsu_io_dec_uops_1_uopc;
  wire [7:0] lsu_io_dec_uops_1_br_mask;
  wire [6:0] lsu_io_dec_uops_1_rob_idx;
  wire [3:0] lsu_io_dec_uops_1_ldq_idx;
  wire [3:0] lsu_io_dec_uops_1_stq_idx;
  wire [4:0] lsu_io_dec_uops_1_mem_cmd;
  wire [2:0] lsu_io_dec_uops_1_mem_typ;
  wire  lsu_io_dec_uops_1_is_fence;
  wire  lsu_io_dec_uops_1_is_store;
  wire  lsu_io_dec_uops_1_is_amo;
  wire  lsu_io_dec_uops_1_is_load;
  wire [1:0] lsu_io_dec_uops_1_dst_rtype;
  wire  lsu_io_dec_uops_1_fp_val;
  wire [3:0] lsu_io_new_ldq_idx;
  wire [3:0] lsu_io_new_stq_idx;
  wire  lsu_io_exe_resp_valid;
  wire [8:0] lsu_io_exe_resp_bits_uop_uopc;
  wire  lsu_io_exe_resp_bits_uop_ctrl_is_load;
  wire  lsu_io_exe_resp_bits_uop_ctrl_is_sta;
  wire  lsu_io_exe_resp_bits_uop_ctrl_is_std;
  wire [7:0] lsu_io_exe_resp_bits_uop_br_mask;
  wire [6:0] lsu_io_exe_resp_bits_uop_rob_idx;
  wire [3:0] lsu_io_exe_resp_bits_uop_ldq_idx;
  wire [3:0] lsu_io_exe_resp_bits_uop_stq_idx;
  wire [6:0] lsu_io_exe_resp_bits_uop_pdst;
  wire [4:0] lsu_io_exe_resp_bits_uop_mem_cmd;
  wire [2:0] lsu_io_exe_resp_bits_uop_mem_typ;
  wire  lsu_io_exe_resp_bits_uop_is_fence;
  wire  lsu_io_exe_resp_bits_uop_is_store;
  wire  lsu_io_exe_resp_bits_uop_is_amo;
  wire  lsu_io_exe_resp_bits_uop_is_load;
  wire [1:0] lsu_io_exe_resp_bits_uop_dst_rtype;
  wire  lsu_io_exe_resp_bits_uop_fp_val;
  wire [63:0] lsu_io_exe_resp_bits_data;
  wire [39:0] lsu_io_exe_resp_bits_addr;
  wire  lsu_io_exe_resp_bits_mxcpt_valid;
  wire [16:0] lsu_io_exe_resp_bits_mxcpt_bits;
  wire  lsu_io_exe_resp_bits_sfence_valid;
  wire  lsu_io_exe_resp_bits_sfence_bits_rs1;
  wire  lsu_io_exe_resp_bits_sfence_bits_rs2;
  wire [38:0] lsu_io_exe_resp_bits_sfence_bits_addr;
  wire  lsu_io_fp_stdata_valid;
  wire [7:0] lsu_io_fp_stdata_bits_uop_br_mask;
  wire [6:0] lsu_io_fp_stdata_bits_uop_rob_idx;
  wire [3:0] lsu_io_fp_stdata_bits_uop_stq_idx;
  wire  lsu_io_fp_stdata_bits_uop_is_amo;
  wire [63:0] lsu_io_fp_stdata_bits_data;
  wire  lsu_io_commit_store_mask_0;
  wire  lsu_io_commit_store_mask_1;
  wire  lsu_io_commit_load_mask_0;
  wire  lsu_io_commit_load_mask_1;
  wire  lsu_io_commit_load_at_rob_head;
  wire  lsu_io_memreq_val;
  wire [31:0] lsu_io_memreq_addr;
  wire [63:0] lsu_io_memreq_wdata;
  wire [8:0] lsu_io_memreq_uop_uopc;
  wire [7:0] lsu_io_memreq_uop_br_mask;
  wire [6:0] lsu_io_memreq_uop_rob_idx;
  wire [3:0] lsu_io_memreq_uop_ldq_idx;
  wire [3:0] lsu_io_memreq_uop_stq_idx;
  wire [6:0] lsu_io_memreq_uop_pdst;
  wire [4:0] lsu_io_memreq_uop_mem_cmd;
  wire [2:0] lsu_io_memreq_uop_mem_typ;
  wire  lsu_io_memreq_uop_is_store;
  wire  lsu_io_memreq_uop_is_amo;
  wire  lsu_io_memreq_uop_is_load;
  wire [1:0] lsu_io_memreq_uop_dst_rtype;
  wire  lsu_io_memreq_uop_fp_val;
  wire  lsu_io_memreq_kill;
  wire  lsu_io_forward_val;
  wire [63:0] lsu_io_forward_data;
  wire [8:0] lsu_io_forward_uop_uopc;
  wire [6:0] lsu_io_forward_uop_rob_idx;
  wire [3:0] lsu_io_forward_uop_ldq_idx;
  wire [3:0] lsu_io_forward_uop_stq_idx;
  wire [6:0] lsu_io_forward_uop_pdst;
  wire [2:0] lsu_io_forward_uop_mem_typ;
  wire  lsu_io_forward_uop_is_store;
  wire  lsu_io_forward_uop_is_amo;
  wire  lsu_io_forward_uop_is_load;
  wire [1:0] lsu_io_forward_uop_dst_rtype;
  wire  lsu_io_forward_uop_fp_val;
  wire  lsu_io_memresp_valid;
  wire [3:0] lsu_io_memresp_bits_ldq_idx;
  wire [3:0] lsu_io_memresp_bits_stq_idx;
  wire  lsu_io_memresp_bits_is_load;
  wire  lsu_io_brinfo_valid;
  wire  lsu_io_brinfo_mispredict;
  wire [7:0] lsu_io_brinfo_mask;
  wire [3:0] lsu_io_brinfo_ldq_idx;
  wire [3:0] lsu_io_brinfo_stq_idx;
  wire  lsu_io_laq_full;
  wire  lsu_io_stq_full;
  wire  lsu_io_exception;
  wire  lsu_io_lsu_clr_bsy_valid_0;
  wire  lsu_io_lsu_clr_bsy_valid_1;
  wire [6:0] lsu_io_lsu_clr_bsy_rob_idx_0;
  wire [6:0] lsu_io_lsu_clr_bsy_rob_idx_1;
  wire  lsu_io_lsu_fencei_rdy;
  wire  lsu_io_xcpt_valid;
  wire [7:0] lsu_io_xcpt_bits_uop_br_mask;
  wire [6:0] lsu_io_xcpt_bits_uop_rob_idx;
  wire [4:0] lsu_io_xcpt_bits_cause;
  wire [39:0] lsu_io_xcpt_bits_badvaddr;
  wire  lsu_io_nack_valid;
  wire [3:0] lsu_io_nack_lsu_idx;
  wire  lsu_io_nack_isload;
  wire  lsu_io_nack_cache_nack;
  wire  lsu_io_dmem_is_ordered;
  wire  lsu_io_ptw_req_ready;
  wire  lsu_io_ptw_req_valid;
  wire [26:0] lsu_io_ptw_req_bits_addr;
  wire  lsu_io_ptw_resp_valid;
  wire  lsu_io_ptw_resp_bits_ae;
  wire [53:0] lsu_io_ptw_resp_bits_pte_ppn;
  wire  lsu_io_ptw_resp_bits_pte_d;
  wire  lsu_io_ptw_resp_bits_pte_a;
  wire  lsu_io_ptw_resp_bits_pte_g;
  wire  lsu_io_ptw_resp_bits_pte_u;
  wire  lsu_io_ptw_resp_bits_pte_x;
  wire  lsu_io_ptw_resp_bits_pte_w;
  wire  lsu_io_ptw_resp_bits_pte_r;
  wire  lsu_io_ptw_resp_bits_pte_v;
  wire [1:0] lsu_io_ptw_resp_bits_level;
  wire  lsu_io_ptw_resp_bits_homogeneous;
  wire [3:0] lsu_io_ptw_ptbr_mode;
  wire [1:0] lsu_io_ptw_status_dprv;
  wire  lsu_io_ptw_status_mxr;
  wire  lsu_io_ptw_status_sum;
  wire  rob_clock;
  wire  rob_reset;
  wire  rob_io_enq_valids_0;
  wire  rob_io_enq_valids_1;
  wire [39:0] rob_io_enq_uops_0_pc;
  wire [7:0] rob_io_enq_uops_0_br_mask;
  wire [6:0] rob_io_enq_uops_0_rob_idx;
  wire [5:0] rob_io_enq_uops_0_brob_idx;
  wire [6:0] rob_io_enq_uops_0_pdst;
  wire [6:0] rob_io_enq_uops_0_stale_pdst;
  wire  rob_io_enq_uops_0_exception;
  wire [63:0] rob_io_enq_uops_0_exc_cause;
  wire  rob_io_enq_uops_0_is_fence;
  wire  rob_io_enq_uops_0_is_fencei;
  wire  rob_io_enq_uops_0_is_store;
  wire  rob_io_enq_uops_0_is_load;
  wire  rob_io_enq_uops_0_is_sys_pc2epc;
  wire  rob_io_enq_uops_0_is_unique;
  wire  rob_io_enq_uops_0_flush_on_commit;
  wire [5:0] rob_io_enq_uops_0_ldst;
  wire  rob_io_enq_uops_0_ldst_val;
  wire [1:0] rob_io_enq_uops_0_dst_rtype;
  wire  rob_io_enq_uops_0_fp_val;
  wire [7:0] rob_io_enq_uops_1_br_mask;
  wire [6:0] rob_io_enq_uops_1_rob_idx;
  wire [6:0] rob_io_enq_uops_1_pdst;
  wire [6:0] rob_io_enq_uops_1_stale_pdst;
  wire  rob_io_enq_uops_1_exception;
  wire [63:0] rob_io_enq_uops_1_exc_cause;
  wire  rob_io_enq_uops_1_is_fence;
  wire  rob_io_enq_uops_1_is_fencei;
  wire  rob_io_enq_uops_1_is_store;
  wire  rob_io_enq_uops_1_is_load;
  wire  rob_io_enq_uops_1_is_sys_pc2epc;
  wire  rob_io_enq_uops_1_is_unique;
  wire  rob_io_enq_uops_1_flush_on_commit;
  wire [5:0] rob_io_enq_uops_1_ldst;
  wire  rob_io_enq_uops_1_ldst_val;
  wire [1:0] rob_io_enq_uops_1_dst_rtype;
  wire  rob_io_enq_uops_1_fp_val;
  wire  rob_io_enq_has_br_or_jalr_in_packet;
  wire  rob_io_enq_partial_stall;
  wire  rob_io_enq_new_packet;
  wire [6:0] rob_io_curr_rob_tail;
  wire  rob_io_brinfo_valid;
  wire  rob_io_brinfo_mispredict;
  wire [7:0] rob_io_brinfo_mask;
  wire [6:0] rob_io_brinfo_rob_idx;
  wire [6:0] rob_io_get_pc_rob_idx;
  wire [39:0] rob_io_get_pc_curr_pc;
  wire [5:0] rob_io_get_pc_curr_brob_idx;
  wire  rob_io_get_pc_next_val;
  wire [39:0] rob_io_get_pc_next_pc;
  wire  rob_io_wb_resps_0_valid;
  wire [6:0] rob_io_wb_resps_0_bits_uop_rob_idx;
  wire [6:0] rob_io_wb_resps_0_bits_uop_pdst;
  wire  rob_io_wb_resps_1_valid;
  wire [6:0] rob_io_wb_resps_1_bits_uop_rob_idx;
  wire [6:0] rob_io_wb_resps_1_bits_uop_pdst;
  wire  rob_io_wb_resps_2_valid;
  wire [6:0] rob_io_wb_resps_2_bits_uop_rob_idx;
  wire [6:0] rob_io_wb_resps_2_bits_uop_pdst;
  wire  rob_io_wb_resps_3_valid;
  wire [6:0] rob_io_wb_resps_3_bits_uop_rob_idx;
  wire [6:0] rob_io_wb_resps_3_bits_uop_pdst;
  wire  rob_io_wb_resps_4_valid;
  wire [6:0] rob_io_wb_resps_4_bits_uop_rob_idx;
  wire [6:0] rob_io_wb_resps_4_bits_uop_pdst;
  wire  rob_io_lsu_clr_bsy_valid_0;
  wire  rob_io_lsu_clr_bsy_valid_1;
  wire [6:0] rob_io_lsu_clr_bsy_rob_idx_0;
  wire [6:0] rob_io_lsu_clr_bsy_rob_idx_1;
  wire  rob_io_fflags_0_valid;
  wire [6:0] rob_io_fflags_0_bits_uop_rob_idx;
  wire [4:0] rob_io_fflags_0_bits_flags;
  wire  rob_io_fflags_1_valid;
  wire [6:0] rob_io_fflags_1_bits_uop_rob_idx;
  wire [4:0] rob_io_fflags_1_bits_flags;
  wire  rob_io_lxcpt_valid;
  wire [7:0] rob_io_lxcpt_bits_uop_br_mask;
  wire [6:0] rob_io_lxcpt_bits_uop_rob_idx;
  wire [4:0] rob_io_lxcpt_bits_cause;
  wire [39:0] rob_io_lxcpt_bits_badvaddr;
  wire  rob_io_bxcpt_valid;
  wire [7:0] rob_io_bxcpt_bits_uop_br_mask;
  wire [6:0] rob_io_bxcpt_bits_uop_rob_idx;
  wire [39:0] rob_io_bxcpt_bits_badvaddr;
  wire  rob_io_commit_valids_0;
  wire  rob_io_commit_valids_1;
  wire [6:0] rob_io_commit_uops_0_pdst;
  wire [6:0] rob_io_commit_uops_0_stale_pdst;
  wire  rob_io_commit_uops_0_is_fencei;
  wire  rob_io_commit_uops_0_is_store;
  wire  rob_io_commit_uops_0_is_load;
  wire  rob_io_commit_uops_0_is_sys_pc2epc;
  wire  rob_io_commit_uops_0_flush_on_commit;
  wire [5:0] rob_io_commit_uops_0_ldst;
  wire [1:0] rob_io_commit_uops_0_dst_rtype;
  wire  rob_io_commit_uops_0_fp_val;
  wire [6:0] rob_io_commit_uops_1_pdst;
  wire [6:0] rob_io_commit_uops_1_stale_pdst;
  wire  rob_io_commit_uops_1_is_fencei;
  wire  rob_io_commit_uops_1_is_store;
  wire  rob_io_commit_uops_1_is_load;
  wire  rob_io_commit_uops_1_is_sys_pc2epc;
  wire  rob_io_commit_uops_1_flush_on_commit;
  wire [5:0] rob_io_commit_uops_1_ldst;
  wire [1:0] rob_io_commit_uops_1_dst_rtype;
  wire  rob_io_commit_uops_1_fp_val;
  wire  rob_io_commit_fflags_valid;
  wire [4:0] rob_io_commit_fflags_bits;
  wire  rob_io_commit_rbk_valids_0;
  wire  rob_io_commit_rbk_valids_1;
  wire  rob_io_commit_st_mask_0;
  wire  rob_io_commit_st_mask_1;
  wire  rob_io_commit_ld_mask_0;
  wire  rob_io_commit_ld_mask_1;
  wire  rob_io_com_load_is_at_rob_head;
  wire  rob_io_com_xcpt_valid;
  wire [63:0] rob_io_com_xcpt_bits_pc;
  wire [63:0] rob_io_com_xcpt_bits_cause;
  wire [63:0] rob_io_com_xcpt_bits_badvaddr;
  wire  rob_io_csr_eret;
  wire [39:0] rob_io_csr_evec;
  wire  rob_io_csr_stall;
  wire  rob_io_flush_valid;
  wire [63:0] rob_io_flush_bits_pc;
  wire  rob_io_clear_brob;
  wire  rob_io_empty;
  wire  rob_io_ready;
  wire  rob_io_brob_deallocate_valid;
  wire [5:0] rob_io_brob_deallocate_bits_brob_idx;
  wire  int_wakeups_0_valid;
  wire [6:0] int_wakeups_0_bits_uop_pdst;
  wire [1:0] int_wakeups_0_bits_uop_dst_rtype;
  wire  int_wakeups_1_valid;
  wire [6:0] int_wakeups_1_bits_uop_pdst;
  wire [1:0] int_wakeups_1_bits_uop_dst_rtype;
  wire  int_wakeups_2_valid;
  wire [6:0] int_wakeups_2_bits_uop_pdst;
  wire [1:0] int_wakeups_2_bits_uop_dst_rtype;
  wire  int_wakeups_3_valid;
  wire [6:0] int_wakeups_3_bits_uop_pdst;
  wire [1:0] int_wakeups_3_bits_uop_dst_rtype;
  wire  int_wakeups_4_valid;
  wire [6:0] int_wakeups_4_bits_uop_pdst;
  wire [1:0] int_wakeups_4_bits_uop_dst_rtype;
  wire  dec_valids_0;
  wire  dec_valids_1;
  wire  dec_uops_0_valid;
  wire [8:0] dec_uops_0_uopc;
  wire [31:0] dec_uops_0_inst;
  wire [39:0] dec_uops_0_pc;
  wire [1:0] dec_uops_0_iqtype;
  wire [9:0] dec_uops_0_fu_code;
  wire  dec_uops_0_allocate_brtag;
  wire  dec_uops_0_is_br_or_jmp;
  wire  dec_uops_0_is_jump;
  wire  dec_uops_0_is_jal;
  wire  dec_uops_0_is_ret;
  wire  dec_uops_0_is_call;
  wire [7:0] dec_uops_0_br_mask;
  wire [2:0] dec_uops_0_br_tag;
  wire  dec_uops_0_br_prediction_btb_blame;
  wire  dec_uops_0_br_prediction_btb_hit;
  wire  dec_uops_0_br_prediction_btb_taken;
  wire  dec_uops_0_br_prediction_bpd_blame;
  wire  dec_uops_0_br_prediction_bpd_hit;
  wire  dec_uops_0_br_prediction_bpd_taken;
  wire [1:0] dec_uops_0_br_prediction_bim_resp_value;
  wire [5:0] dec_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] dec_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] dec_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] dec_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] dec_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] dec_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dec_uops_0_br_prediction_bpd_resp_info;
  wire [2:0] dec_uops_0_fetch_pc_lob;
  wire [19:0] dec_uops_0_imm_packed;
  wire [6:0] dec_uops_0_rob_idx;
  wire [3:0] dec_uops_0_ldq_idx;
  wire [3:0] dec_uops_0_stq_idx;
  wire [5:0] dec_uops_0_brob_idx;
  wire  dec_uops_0_exception;
  wire [63:0] dec_uops_0_exc_cause;
  wire  dec_uops_0_bypassable;
  wire [4:0] dec_uops_0_mem_cmd;
  wire [2:0] dec_uops_0_mem_typ;
  wire  dec_uops_0_is_fence;
  wire  dec_uops_0_is_fencei;
  wire  dec_uops_0_is_store;
  wire  dec_uops_0_is_amo;
  wire  dec_uops_0_is_load;
  wire  dec_uops_0_is_sys_pc2epc;
  wire  dec_uops_0_is_unique;
  wire  dec_uops_0_flush_on_commit;
  wire [5:0] dec_uops_0_ldst;
  wire [5:0] dec_uops_0_lrs1;
  wire [5:0] dec_uops_0_lrs2;
  wire [5:0] dec_uops_0_lrs3;
  wire  dec_uops_0_ldst_val;
  wire [1:0] dec_uops_0_dst_rtype;
  wire [1:0] dec_uops_0_lrs1_rtype;
  wire [1:0] dec_uops_0_lrs2_rtype;
  wire  dec_uops_0_frs3_en;
  wire  dec_uops_0_fp_val;
  wire  dec_uops_0_fp_single;
  wire  dec_uops_0_xcpt_pf_if;
  wire  dec_uops_0_xcpt_ae_if;
  wire  dec_uops_0_replay_if;
  wire  dec_uops_0_xcpt_ma_if;
  wire [31:0] dec_uops_0_debug_events_fetch_seq;
  wire  dec_uops_1_valid;
  wire [8:0] dec_uops_1_uopc;
  wire [31:0] dec_uops_1_inst;
  wire [39:0] dec_uops_1_pc;
  wire [1:0] dec_uops_1_iqtype;
  wire [9:0] dec_uops_1_fu_code;
  wire  dec_uops_1_allocate_brtag;
  wire  dec_uops_1_is_br_or_jmp;
  wire  dec_uops_1_is_jump;
  wire  dec_uops_1_is_jal;
  wire  dec_uops_1_is_ret;
  wire  dec_uops_1_is_call;
  wire [7:0] dec_uops_1_br_mask;
  wire [2:0] dec_uops_1_br_tag;
  wire  dec_uops_1_br_prediction_btb_blame;
  wire  dec_uops_1_br_prediction_btb_hit;
  wire  dec_uops_1_br_prediction_btb_taken;
  wire  dec_uops_1_br_prediction_bpd_blame;
  wire  dec_uops_1_br_prediction_bpd_hit;
  wire  dec_uops_1_br_prediction_bpd_taken;
  wire [1:0] dec_uops_1_br_prediction_bim_resp_value;
  wire [5:0] dec_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] dec_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] dec_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] dec_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] dec_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] dec_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dec_uops_1_br_prediction_bpd_resp_info;
  wire [2:0] dec_uops_1_fetch_pc_lob;
  wire [19:0] dec_uops_1_imm_packed;
  wire [6:0] dec_uops_1_rob_idx;
  wire [3:0] dec_uops_1_ldq_idx;
  wire [3:0] dec_uops_1_stq_idx;
  wire [5:0] dec_uops_1_brob_idx;
  wire  dec_uops_1_exception;
  wire [63:0] dec_uops_1_exc_cause;
  wire  dec_uops_1_bypassable;
  wire [4:0] dec_uops_1_mem_cmd;
  wire [2:0] dec_uops_1_mem_typ;
  wire  dec_uops_1_is_fence;
  wire  dec_uops_1_is_fencei;
  wire  dec_uops_1_is_store;
  wire  dec_uops_1_is_amo;
  wire  dec_uops_1_is_load;
  wire  dec_uops_1_is_sys_pc2epc;
  wire  dec_uops_1_is_unique;
  wire  dec_uops_1_flush_on_commit;
  wire [5:0] dec_uops_1_ldst;
  wire [5:0] dec_uops_1_lrs1;
  wire [5:0] dec_uops_1_lrs2;
  wire [5:0] dec_uops_1_lrs3;
  wire  dec_uops_1_ldst_val;
  wire [1:0] dec_uops_1_dst_rtype;
  wire [1:0] dec_uops_1_lrs1_rtype;
  wire [1:0] dec_uops_1_lrs2_rtype;
  wire  dec_uops_1_frs3_en;
  wire  dec_uops_1_fp_val;
  wire  dec_uops_1_fp_single;
  wire  dec_uops_1_xcpt_pf_if;
  wire  dec_uops_1_xcpt_ae_if;
  wire  dec_uops_1_replay_if;
  wire  dec_uops_1_xcpt_ma_if;
  wire [31:0] dec_uops_1_debug_events_fetch_seq;
  wire  dec_will_fire_0;
  wire  dec_will_fire_1;
  wire  dec_rdy;
  wire  dis_valids_0;
  wire  dis_valids_1;
  wire  dis_uops_0_valid;
  wire [8:0] dis_uops_0_uopc;
  wire [31:0] dis_uops_0_inst;
  wire [39:0] dis_uops_0_pc;
  wire [1:0] dis_uops_0_iqtype;
  wire [9:0] dis_uops_0_fu_code;
  wire  dis_uops_0_allocate_brtag;
  wire  dis_uops_0_is_br_or_jmp;
  wire  dis_uops_0_is_jump;
  wire  dis_uops_0_is_jal;
  wire  dis_uops_0_is_ret;
  wire  dis_uops_0_is_call;
  wire [7:0] dis_uops_0_br_mask;
  wire [2:0] dis_uops_0_br_tag;
  wire  dis_uops_0_br_prediction_btb_blame;
  wire  dis_uops_0_br_prediction_btb_hit;
  wire  dis_uops_0_br_prediction_btb_taken;
  wire  dis_uops_0_br_prediction_bpd_blame;
  wire  dis_uops_0_br_prediction_bpd_hit;
  wire  dis_uops_0_br_prediction_bpd_taken;
  wire [1:0] dis_uops_0_br_prediction_bim_resp_value;
  wire [5:0] dis_uops_0_br_prediction_bim_resp_entry_idx;
  wire [1:0] dis_uops_0_br_prediction_bim_resp_way_idx;
  wire [1:0] dis_uops_0_br_prediction_bpd_resp_takens;
  wire [14:0] dis_uops_0_br_prediction_bpd_resp_history;
  wire [14:0] dis_uops_0_br_prediction_bpd_resp_history_u;
  wire [7:0] dis_uops_0_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dis_uops_0_br_prediction_bpd_resp_info;
  wire  dis_uops_0_stat_brjmp_mispredicted;
  wire  dis_uops_0_stat_btb_made_pred;
  wire  dis_uops_0_stat_btb_mispredicted;
  wire  dis_uops_0_stat_bpd_made_pred;
  wire  dis_uops_0_stat_bpd_mispredicted;
  wire [2:0] dis_uops_0_fetch_pc_lob;
  wire [19:0] dis_uops_0_imm_packed;
  wire [11:0] dis_uops_0_csr_addr;
  wire [6:0] dis_uops_0_rob_idx;
  wire [3:0] dis_uops_0_ldq_idx;
  wire [3:0] dis_uops_0_stq_idx;
  wire [5:0] dis_uops_0_brob_idx;
  wire [6:0] dis_uops_0_pdst;
  wire [6:0] dis_uops_0_pop1;
  wire [6:0] dis_uops_0_pop2;
  wire [6:0] dis_uops_0_pop3;
  wire  dis_uops_0_prs1_busy;
  wire  dis_uops_0_prs2_busy;
  wire  dis_uops_0_prs3_busy;
  wire [6:0] dis_uops_0_stale_pdst;
  wire  dis_uops_0_exception;
  wire [63:0] dis_uops_0_exc_cause;
  wire  dis_uops_0_bypassable;
  wire [4:0] dis_uops_0_mem_cmd;
  wire [2:0] dis_uops_0_mem_typ;
  wire  dis_uops_0_is_fence;
  wire  dis_uops_0_is_fencei;
  wire  dis_uops_0_is_store;
  wire  dis_uops_0_is_amo;
  wire  dis_uops_0_is_load;
  wire  dis_uops_0_is_sys_pc2epc;
  wire  dis_uops_0_is_unique;
  wire  dis_uops_0_flush_on_commit;
  wire [5:0] dis_uops_0_ldst;
  wire [5:0] dis_uops_0_lrs1;
  wire [5:0] dis_uops_0_lrs2;
  wire [5:0] dis_uops_0_lrs3;
  wire  dis_uops_0_ldst_val;
  wire [1:0] dis_uops_0_dst_rtype;
  wire [1:0] dis_uops_0_lrs1_rtype;
  wire [1:0] dis_uops_0_lrs2_rtype;
  wire  dis_uops_0_frs3_en;
  wire  dis_uops_0_fp_val;
  wire  dis_uops_0_fp_single;
  wire  dis_uops_0_xcpt_pf_if;
  wire  dis_uops_0_xcpt_ae_if;
  wire  dis_uops_0_replay_if;
  wire  dis_uops_0_xcpt_ma_if;
  wire [63:0] dis_uops_0_debug_wdata;
  wire [31:0] dis_uops_0_debug_events_fetch_seq;
  wire  dis_uops_1_valid;
  wire [8:0] dis_uops_1_uopc;
  wire [31:0] dis_uops_1_inst;
  wire [39:0] dis_uops_1_pc;
  wire [1:0] dis_uops_1_iqtype;
  wire [9:0] dis_uops_1_fu_code;
  wire  dis_uops_1_allocate_brtag;
  wire  dis_uops_1_is_br_or_jmp;
  wire  dis_uops_1_is_jump;
  wire  dis_uops_1_is_jal;
  wire  dis_uops_1_is_ret;
  wire  dis_uops_1_is_call;
  wire [7:0] dis_uops_1_br_mask;
  wire [2:0] dis_uops_1_br_tag;
  wire  dis_uops_1_br_prediction_btb_blame;
  wire  dis_uops_1_br_prediction_btb_hit;
  wire  dis_uops_1_br_prediction_btb_taken;
  wire  dis_uops_1_br_prediction_bpd_blame;
  wire  dis_uops_1_br_prediction_bpd_hit;
  wire  dis_uops_1_br_prediction_bpd_taken;
  wire [1:0] dis_uops_1_br_prediction_bim_resp_value;
  wire [5:0] dis_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] dis_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] dis_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] dis_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] dis_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] dis_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] dis_uops_1_br_prediction_bpd_resp_info;
  wire  dis_uops_1_stat_brjmp_mispredicted;
  wire  dis_uops_1_stat_btb_made_pred;
  wire  dis_uops_1_stat_btb_mispredicted;
  wire  dis_uops_1_stat_bpd_made_pred;
  wire  dis_uops_1_stat_bpd_mispredicted;
  wire [2:0] dis_uops_1_fetch_pc_lob;
  wire [19:0] dis_uops_1_imm_packed;
  wire [11:0] dis_uops_1_csr_addr;
  wire [6:0] dis_uops_1_rob_idx;
  wire [3:0] dis_uops_1_ldq_idx;
  wire [3:0] dis_uops_1_stq_idx;
  wire [5:0] dis_uops_1_brob_idx;
  wire [6:0] dis_uops_1_pdst;
  wire [6:0] dis_uops_1_pop1;
  wire [6:0] dis_uops_1_pop2;
  wire [6:0] dis_uops_1_pop3;
  wire  dis_uops_1_prs1_busy;
  wire  dis_uops_1_prs2_busy;
  wire  dis_uops_1_prs3_busy;
  wire [6:0] dis_uops_1_stale_pdst;
  wire  dis_uops_1_exception;
  wire [63:0] dis_uops_1_exc_cause;
  wire  dis_uops_1_bypassable;
  wire [4:0] dis_uops_1_mem_cmd;
  wire [2:0] dis_uops_1_mem_typ;
  wire  dis_uops_1_is_fence;
  wire  dis_uops_1_is_fencei;
  wire  dis_uops_1_is_store;
  wire  dis_uops_1_is_amo;
  wire  dis_uops_1_is_load;
  wire  dis_uops_1_is_sys_pc2epc;
  wire  dis_uops_1_is_unique;
  wire  dis_uops_1_flush_on_commit;
  wire [5:0] dis_uops_1_ldst;
  wire [5:0] dis_uops_1_lrs1;
  wire [5:0] dis_uops_1_lrs2;
  wire [5:0] dis_uops_1_lrs3;
  wire  dis_uops_1_ldst_val;
  wire [1:0] dis_uops_1_dst_rtype;
  wire [1:0] dis_uops_1_lrs1_rtype;
  wire [1:0] dis_uops_1_lrs2_rtype;
  wire  dis_uops_1_frs3_en;
  wire  dis_uops_1_fp_val;
  wire  dis_uops_1_fp_single;
  wire  dis_uops_1_xcpt_pf_if;
  wire  dis_uops_1_xcpt_ae_if;
  wire  dis_uops_1_replay_if;
  wire  dis_uops_1_xcpt_ma_if;
  wire [63:0] dis_uops_1_debug_wdata;
  wire [31:0] dis_uops_1_debug_events_fetch_seq;
  wire  iss_valids_0;
  wire  iss_valids_1;
  wire  iss_valids_2;
  wire [8:0] iss_uops_0_uopc;
  wire [7:0] iss_uops_0_br_mask;
  wire [19:0] iss_uops_0_imm_packed;
  wire [6:0] iss_uops_0_rob_idx;
  wire [3:0] iss_uops_0_ldq_idx;
  wire [3:0] iss_uops_0_stq_idx;
  wire [6:0] iss_uops_0_pdst;
  wire [6:0] iss_uops_0_pop1;
  wire [6:0] iss_uops_0_pop2;
  wire [4:0] iss_uops_0_mem_cmd;
  wire [2:0] iss_uops_0_mem_typ;
  wire  iss_uops_0_is_fence;
  wire  iss_uops_0_is_store;
  wire  iss_uops_0_is_amo;
  wire  iss_uops_0_is_load;
  wire [1:0] iss_uops_0_dst_rtype;
  wire [1:0] iss_uops_0_lrs1_rtype;
  wire [1:0] iss_uops_0_lrs2_rtype;
  wire  iss_uops_0_fp_val;
  wire  iss_uops_1_valid;
  wire [1:0] iss_uops_1_iw_state;
  wire [8:0] iss_uops_1_uopc;
  wire [31:0] iss_uops_1_inst;
  wire [39:0] iss_uops_1_pc;
  wire [1:0] iss_uops_1_iqtype;
  wire [9:0] iss_uops_1_fu_code;
  wire  iss_uops_1_allocate_brtag;
  wire  iss_uops_1_is_br_or_jmp;
  wire  iss_uops_1_is_jump;
  wire  iss_uops_1_is_jal;
  wire  iss_uops_1_is_ret;
  wire  iss_uops_1_is_call;
  wire [7:0] iss_uops_1_br_mask;
  wire [2:0] iss_uops_1_br_tag;
  wire  iss_uops_1_br_prediction_btb_blame;
  wire  iss_uops_1_br_prediction_btb_hit;
  wire  iss_uops_1_br_prediction_btb_taken;
  wire  iss_uops_1_br_prediction_bpd_blame;
  wire  iss_uops_1_br_prediction_bpd_hit;
  wire  iss_uops_1_br_prediction_bpd_taken;
  wire [1:0] iss_uops_1_br_prediction_bim_resp_value;
  wire [5:0] iss_uops_1_br_prediction_bim_resp_entry_idx;
  wire [1:0] iss_uops_1_br_prediction_bim_resp_way_idx;
  wire [1:0] iss_uops_1_br_prediction_bpd_resp_takens;
  wire [14:0] iss_uops_1_br_prediction_bpd_resp_history;
  wire [14:0] iss_uops_1_br_prediction_bpd_resp_history_u;
  wire [7:0] iss_uops_1_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iss_uops_1_br_prediction_bpd_resp_info;
  wire  iss_uops_1_stat_brjmp_mispredicted;
  wire  iss_uops_1_stat_btb_made_pred;
  wire  iss_uops_1_stat_btb_mispredicted;
  wire  iss_uops_1_stat_bpd_made_pred;
  wire  iss_uops_1_stat_bpd_mispredicted;
  wire [2:0] iss_uops_1_fetch_pc_lob;
  wire [19:0] iss_uops_1_imm_packed;
  wire [11:0] iss_uops_1_csr_addr;
  wire [6:0] iss_uops_1_rob_idx;
  wire [3:0] iss_uops_1_ldq_idx;
  wire [3:0] iss_uops_1_stq_idx;
  wire [5:0] iss_uops_1_brob_idx;
  wire [6:0] iss_uops_1_pdst;
  wire [6:0] iss_uops_1_pop1;
  wire [6:0] iss_uops_1_pop2;
  wire [6:0] iss_uops_1_pop3;
  wire  iss_uops_1_prs1_busy;
  wire  iss_uops_1_prs2_busy;
  wire  iss_uops_1_prs3_busy;
  wire [6:0] iss_uops_1_stale_pdst;
  wire  iss_uops_1_exception;
  wire [63:0] iss_uops_1_exc_cause;
  wire  iss_uops_1_bypassable;
  wire [4:0] iss_uops_1_mem_cmd;
  wire [2:0] iss_uops_1_mem_typ;
  wire  iss_uops_1_is_fence;
  wire  iss_uops_1_is_fencei;
  wire  iss_uops_1_is_store;
  wire  iss_uops_1_is_amo;
  wire  iss_uops_1_is_load;
  wire  iss_uops_1_is_sys_pc2epc;
  wire  iss_uops_1_is_unique;
  wire  iss_uops_1_flush_on_commit;
  wire [5:0] iss_uops_1_ldst;
  wire [5:0] iss_uops_1_lrs1;
  wire [5:0] iss_uops_1_lrs2;
  wire [5:0] iss_uops_1_lrs3;
  wire  iss_uops_1_ldst_val;
  wire [1:0] iss_uops_1_dst_rtype;
  wire [1:0] iss_uops_1_lrs1_rtype;
  wire [1:0] iss_uops_1_lrs2_rtype;
  wire  iss_uops_1_frs3_en;
  wire  iss_uops_1_fp_val;
  wire  iss_uops_1_fp_single;
  wire  iss_uops_1_xcpt_pf_if;
  wire  iss_uops_1_xcpt_ae_if;
  wire  iss_uops_1_replay_if;
  wire  iss_uops_1_xcpt_ma_if;
  wire [63:0] iss_uops_1_debug_wdata;
  wire [31:0] iss_uops_1_debug_events_fetch_seq;
  wire  iss_uops_2_valid;
  wire [1:0] iss_uops_2_iw_state;
  wire [8:0] iss_uops_2_uopc;
  wire [31:0] iss_uops_2_inst;
  wire [39:0] iss_uops_2_pc;
  wire [1:0] iss_uops_2_iqtype;
  wire [9:0] iss_uops_2_fu_code;
  wire  iss_uops_2_allocate_brtag;
  wire  iss_uops_2_is_br_or_jmp;
  wire  iss_uops_2_is_jump;
  wire  iss_uops_2_is_jal;
  wire  iss_uops_2_is_ret;
  wire  iss_uops_2_is_call;
  wire [7:0] iss_uops_2_br_mask;
  wire [2:0] iss_uops_2_br_tag;
  wire  iss_uops_2_br_prediction_btb_blame;
  wire  iss_uops_2_br_prediction_btb_hit;
  wire  iss_uops_2_br_prediction_btb_taken;
  wire  iss_uops_2_br_prediction_bpd_blame;
  wire  iss_uops_2_br_prediction_bpd_hit;
  wire  iss_uops_2_br_prediction_bpd_taken;
  wire [1:0] iss_uops_2_br_prediction_bim_resp_value;
  wire [5:0] iss_uops_2_br_prediction_bim_resp_entry_idx;
  wire [1:0] iss_uops_2_br_prediction_bim_resp_way_idx;
  wire [1:0] iss_uops_2_br_prediction_bpd_resp_takens;
  wire [14:0] iss_uops_2_br_prediction_bpd_resp_history;
  wire [14:0] iss_uops_2_br_prediction_bpd_resp_history_u;
  wire [7:0] iss_uops_2_br_prediction_bpd_resp_history_ptr;
  wire [14:0] iss_uops_2_br_prediction_bpd_resp_info;
  wire  iss_uops_2_stat_brjmp_mispredicted;
  wire  iss_uops_2_stat_btb_made_pred;
  wire  iss_uops_2_stat_btb_mispredicted;
  wire  iss_uops_2_stat_bpd_made_pred;
  wire  iss_uops_2_stat_bpd_mispredicted;
  wire [2:0] iss_uops_2_fetch_pc_lob;
  wire [19:0] iss_uops_2_imm_packed;
  wire [11:0] iss_uops_2_csr_addr;
  wire [6:0] iss_uops_2_rob_idx;
  wire [3:0] iss_uops_2_ldq_idx;
  wire [3:0] iss_uops_2_stq_idx;
  wire [5:0] iss_uops_2_brob_idx;
  wire [6:0] iss_uops_2_pdst;
  wire [6:0] iss_uops_2_pop1;
  wire [6:0] iss_uops_2_pop2;
  wire [6:0] iss_uops_2_pop3;
  wire  iss_uops_2_prs1_busy;
  wire  iss_uops_2_prs2_busy;
  wire  iss_uops_2_prs3_busy;
  wire [6:0] iss_uops_2_stale_pdst;
  wire  iss_uops_2_exception;
  wire [63:0] iss_uops_2_exc_cause;
  wire  iss_uops_2_bypassable;
  wire [4:0] iss_uops_2_mem_cmd;
  wire [2:0] iss_uops_2_mem_typ;
  wire  iss_uops_2_is_fence;
  wire  iss_uops_2_is_fencei;
  wire  iss_uops_2_is_store;
  wire  iss_uops_2_is_amo;
  wire  iss_uops_2_is_load;
  wire  iss_uops_2_is_sys_pc2epc;
  wire  iss_uops_2_is_unique;
  wire  iss_uops_2_flush_on_commit;
  wire [5:0] iss_uops_2_ldst;
  wire [5:0] iss_uops_2_lrs1;
  wire [5:0] iss_uops_2_lrs2;
  wire [5:0] iss_uops_2_lrs3;
  wire  iss_uops_2_ldst_val;
  wire [1:0] iss_uops_2_dst_rtype;
  wire [1:0] iss_uops_2_lrs1_rtype;
  wire [1:0] iss_uops_2_lrs2_rtype;
  wire  iss_uops_2_frs3_en;
  wire  iss_uops_2_fp_val;
  wire  iss_uops_2_fp_single;
  wire  iss_uops_2_xcpt_pf_if;
  wire  iss_uops_2_xcpt_ae_if;
  wire  iss_uops_2_replay_if;
  wire  iss_uops_2_xcpt_ma_if;
  wire [63:0] iss_uops_2_debug_wdata;
  wire [31:0] iss_uops_2_debug_events_fetch_seq;
  wire  bypasses_valid_0;
  wire  bypasses_valid_1;
  wire  bypasses_valid_2;
  wire  bypasses_valid_3;
  wire  bypasses_uop_0_ctrl_rf_wen;
  wire [6:0] bypasses_uop_0_pdst;
  wire [1:0] bypasses_uop_0_dst_rtype;
  wire  bypasses_uop_1_ctrl_rf_wen;
  wire [6:0] bypasses_uop_1_pdst;
  wire [1:0] bypasses_uop_1_dst_rtype;
  wire  bypasses_uop_2_ctrl_rf_wen;
  wire [6:0] bypasses_uop_2_pdst;
  wire [1:0] bypasses_uop_2_dst_rtype;
  wire  bypasses_uop_3_ctrl_rf_wen;
  wire [6:0] bypasses_uop_3_pdst;
  wire [1:0] bypasses_uop_3_dst_rtype;
  wire [63:0] bypasses_data_0;
  wire [63:0] bypasses_data_1;
  wire [63:0] bypasses_data_2;
  wire [63:0] bypasses_data_3;
  wire  br_unit_take_pc;
  wire [39:0] br_unit_target;
  wire  br_unit_brinfo_valid;
  wire  br_unit_brinfo_mispredict;
  wire [7:0] br_unit_brinfo_mask;
  wire [2:0] br_unit_brinfo_tag;
  wire [7:0] br_unit_brinfo_exe_mask;
  wire [6:0] br_unit_brinfo_rob_idx;
  wire [3:0] br_unit_brinfo_ldq_idx;
  wire [3:0] br_unit_brinfo_stq_idx;
  wire  br_unit_brinfo_is_jr;
  wire  br_unit_btb_update_valid;
  wire [38:0] br_unit_btb_update_bits_pc;
  wire [38:0] br_unit_btb_update_bits_target;
  wire [38:0] br_unit_btb_update_bits_cfi_pc;
  wire [2:0] br_unit_btb_update_bits_bpd_type;
  wire [2:0] br_unit_btb_update_bits_cfi_type;
  wire  br_unit_bim_update_valid;
  wire  br_unit_bim_update_bits_taken;
  wire [1:0] br_unit_bim_update_bits_bim_resp_value;
  wire [5:0] br_unit_bim_update_bits_bim_resp_entry_idx;
  wire [1:0] br_unit_bim_update_bits_bim_resp_way_idx;
  wire  br_unit_bpd_update_valid;
  wire [2:0] br_unit_bpd_update_bits_br_pc;
  wire [5:0] br_unit_bpd_update_bits_brob_idx;
  wire  br_unit_bpd_update_bits_mispredict;
  wire [14:0] br_unit_bpd_update_bits_history;
  wire [7:0] br_unit_bpd_update_bits_history_ptr;
  wire  br_unit_bpd_update_bits_bpd_predict_val;
  wire  br_unit_bpd_update_bits_bpd_mispredict;
  wire  br_unit_bpd_update_bits_taken;
  wire  br_unit_bpd_update_bits_is_br;
  wire  br_unit_bpd_update_bits_new_pc_same_packet;
  wire  br_unit_xcpt_valid;
  wire [7:0] br_unit_xcpt_bits_uop_br_mask;
  wire [6:0] br_unit_xcpt_bits_uop_rob_idx;
  wire [39:0] br_unit_xcpt_bits_badvaddr;
  wire  csr_clock;
  wire  csr_reset;
  wire  csr_io_interrupts_debug;
  wire  csr_io_interrupts_mtip;
  wire  csr_io_interrupts_msip;
  wire  csr_io_interrupts_meip;
  wire  csr_io_interrupts_seip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [63:0] csr_io_rw_rdata;
  wire [63:0] csr_io_rw_wdata;
  wire [11:0] csr_io_decode_0_csr;
  wire  csr_io_decode_0_fp_illegal;
  wire  csr_io_decode_0_read_illegal;
  wire  csr_io_decode_0_write_illegal;
  wire  csr_io_decode_0_write_flush;
  wire  csr_io_decode_0_system_illegal;
  wire [11:0] csr_io_decode_1_csr;
  wire  csr_io_decode_1_fp_illegal;
  wire  csr_io_decode_1_read_illegal;
  wire  csr_io_decode_1_write_illegal;
  wire  csr_io_decode_1_write_flush;
  wire  csr_io_decode_1_system_illegal;
  wire  csr_io_csr_stall;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [31:0] csr_io_status_isa;
  wire [1:0] csr_io_status_dprv;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [26:0] csr_io_status_zero2;
  wire [1:0] csr_io_status_sxl;
  wire [1:0] csr_io_status_uxl;
  wire  csr_io_status_sd_rv32;
  wire [7:0] csr_io_status_zero1;
  wire  csr_io_status_tsr;
  wire  csr_io_status_tw;
  wire  csr_io_status_tvm;
  wire  csr_io_status_mxr;
  wire  csr_io_status_sum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [3:0] csr_io_ptbr_mode;
  wire [43:0] csr_io_ptbr_ppn;
  wire [39:0] csr_io_evec;
  wire  csr_io_exception;
  wire [1:0] csr_io_retire;
  wire [63:0] csr_io_cause;
  wire [39:0] csr_io_pc;
  wire [39:0] csr_io_badaddr;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_interrupt;
  wire [63:0] csr_io_interrupt_cause;
  wire [63:0] csr_io_counters_0_eventSel;
  wire [1:0] csr_io_counters_0_inc;
  wire [63:0] csr_io_counters_1_eventSel;
  wire [1:0] csr_io_counters_1_inc;
  wire [63:0] csr_io_counters_2_eventSel;
  wire [1:0] csr_io_counters_2_inc;
  wire [63:0] csr_io_counters_3_eventSel;
  wire [1:0] csr_io_counters_3_inc;
  wire [63:0] csr_io_counters_4_eventSel;
  wire [1:0] csr_io_counters_4_inc;
  wire [63:0] csr_io_counters_5_eventSel;
  wire [1:0] csr_io_counters_5_inc;
  wire [63:0] csr_io_counters_6_eventSel;
  wire [1:0] csr_io_counters_6_inc;
  wire [63:0] csr_io_counters_7_eventSel;
  wire [1:0] csr_io_counters_7_inc;
  wire [63:0] csr_io_counters_8_eventSel;
  wire [1:0] csr_io_counters_8_inc;
  wire [63:0] csr_io_counters_9_eventSel;
  wire [1:0] csr_io_counters_9_inc;
  wire [63:0] csr_io_counters_10_eventSel;
  wire [1:0] csr_io_counters_10_inc;
  wire [63:0] csr_io_counters_11_eventSel;
  wire [1:0] csr_io_counters_11_inc;
  wire [63:0] csr_io_counters_12_eventSel;
  wire [1:0] csr_io_counters_12_inc;
  wire [63:0] csr_io_counters_13_eventSel;
  wire [1:0] csr_io_counters_13_inc;
  wire [63:0] csr_io_counters_14_eventSel;
  wire [1:0] csr_io_counters_14_inc;
  wire [63:0] csr_io_counters_15_eventSel;
  wire [1:0] csr_io_counters_15_inc;
  wire [63:0] csr_io_counters_16_eventSel;
  wire [1:0] csr_io_counters_16_inc;
  wire [63:0] csr_io_counters_17_eventSel;
  wire [1:0] csr_io_counters_17_inc;
  wire [63:0] csr_io_counters_18_eventSel;
  wire [1:0] csr_io_counters_18_inc;
  wire [63:0] csr_io_counters_19_eventSel;
  wire [1:0] csr_io_counters_19_inc;
  wire [63:0] csr_io_counters_20_eventSel;
  wire [1:0] csr_io_counters_20_inc;
  wire [63:0] csr_io_counters_21_eventSel;
  wire [1:0] csr_io_counters_21_inc;
  wire [63:0] csr_io_counters_22_eventSel;
  wire [1:0] csr_io_counters_22_inc;
  wire [63:0] csr_io_counters_23_eventSel;
  wire [1:0] csr_io_counters_23_inc;
  wire [63:0] csr_io_counters_24_eventSel;
  wire [1:0] csr_io_counters_24_inc;
  wire [63:0] csr_io_counters_25_eventSel;
  wire [1:0] csr_io_counters_25_inc;
  wire [63:0] csr_io_counters_26_eventSel;
  wire [1:0] csr_io_counters_26_inc;
  wire [63:0] csr_io_counters_27_eventSel;
  wire [1:0] csr_io_counters_27_inc;
  wire [63:0] csr_io_counters_28_eventSel;
  wire [1:0] csr_io_counters_28_inc;
  reg  _T_1522;
  reg [31:0] _RAND_0;
  wire  _T_1523;
  wire  icache_blocked;
  wire [1:0] _T_1525;
  wire [55:0] _T_1526;
  wire [1:0] _T_1530;
  wire [3:0] _T_1532;
  wire [55:0] _GEN_13;
  wire [55:0] _T_1533;
  wire  _T_1535;
  wire  _T_1537;
  wire [1:0] _T_1538;
  wire [2:0] _T_1539;
  wire [1:0] _T_1540;
  wire [2:0] _T_1541;
  wire [5:0] _T_1542;
  wire [55:0] _GEN_14;
  wire [55:0] _T_1543;
  wire  _T_1545;
  wire [1:0] _T_1546;
  wire [2:0] _T_1547;
  wire [1:0] _T_1548;
  wire [2:0] _T_1549;
  wire [5:0] _T_1550;
  wire [55:0] _GEN_15;
  wire [55:0] _T_1551;
  wire  _T_1553;
  wire  _T_1555;
  wire  _T_1556;
  wire  _T_1558;
  wire  _T_1559;
  wire  _T_1561;
  wire  _T_1562;
  reg  _T_1564;
  reg [31:0] _RAND_1;
  wire [1:0] _T_1565;
  wire [55:0] _T_1566;
  wire [55:0] _T_1573;
  wire  _T_1575;
  wire [55:0] _T_1583;
  wire  _T_1585;
  wire [55:0] _T_1591;
  wire  _T_1593;
  wire  _T_1595;
  wire  _T_1596;
  wire  _T_1598;
  wire  _T_1599;
  wire  _T_1601;
  wire  _T_1602;
  reg  _T_1604;
  reg [31:0] _RAND_2;
  wire [1:0] _T_1605;
  wire [55:0] _T_1606;
  wire [55:0] _T_1613;
  wire  _T_1615;
  wire [55:0] _T_1623;
  wire  _T_1625;
  wire [55:0] _T_1631;
  wire  _T_1633;
  wire  _T_1635;
  wire  _T_1636;
  wire  _T_1638;
  wire  _T_1639;
  wire  _T_1641;
  wire  _T_1642;
  reg  _T_1644;
  reg [31:0] _RAND_3;
  wire [1:0] _T_1645;
  wire [55:0] _T_1646;
  wire [55:0] _T_1653;
  wire  _T_1655;
  wire [55:0] _T_1663;
  wire  _T_1665;
  wire [55:0] _T_1671;
  wire  _T_1673;
  wire  _T_1675;
  wire  _T_1676;
  wire  _T_1678;
  wire  _T_1679;
  wire  _T_1681;
  wire  _T_1682;
  reg  _T_1684;
  reg [31:0] _RAND_4;
  wire [1:0] _T_1685;
  wire [55:0] _T_1686;
  wire [55:0] _T_1693;
  wire  _T_1695;
  wire [55:0] _T_1703;
  wire  _T_1705;
  wire [55:0] _T_1711;
  wire  _T_1713;
  wire  _T_1715;
  wire  _T_1716;
  wire  _T_1718;
  wire  _T_1719;
  wire  _T_1721;
  wire  _T_1722;
  reg  _T_1724;
  reg [31:0] _RAND_5;
  wire [1:0] _T_1725;
  wire [55:0] _T_1726;
  wire [55:0] _T_1733;
  wire  _T_1735;
  wire [55:0] _T_1743;
  wire  _T_1745;
  wire [55:0] _T_1751;
  wire  _T_1753;
  wire  _T_1755;
  wire  _T_1756;
  wire  _T_1758;
  wire  _T_1759;
  wire  _T_1761;
  wire  _T_1762;
  reg  _T_1764;
  reg [31:0] _RAND_6;
  wire [1:0] _T_1765;
  wire [55:0] _T_1766;
  wire [55:0] _T_1773;
  wire  _T_1775;
  wire [55:0] _T_1783;
  wire  _T_1785;
  wire [55:0] _T_1791;
  wire  _T_1793;
  wire  _T_1795;
  wire  _T_1796;
  wire  _T_1798;
  wire  _T_1799;
  wire  _T_1801;
  wire  _T_1802;
  reg  _T_1804;
  reg [31:0] _RAND_7;
  wire [1:0] _T_1805;
  wire [55:0] _T_1806;
  wire [55:0] _T_1813;
  wire  _T_1815;
  wire [55:0] _T_1823;
  wire  _T_1825;
  wire [55:0] _T_1831;
  wire  _T_1833;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1838;
  wire  _T_1839;
  wire  _T_1841;
  wire  _T_1842;
  reg  _T_1844;
  reg [31:0] _RAND_8;
  wire [1:0] _T_1845;
  wire [55:0] _T_1846;
  wire [55:0] _T_1853;
  wire  _T_1855;
  wire [55:0] _T_1863;
  wire  _T_1865;
  wire [55:0] _T_1871;
  wire  _T_1873;
  wire  _T_1875;
  wire  _T_1876;
  wire  _T_1878;
  wire  _T_1879;
  wire  _T_1881;
  wire  _T_1882;
  reg  _T_1884;
  reg [31:0] _RAND_9;
  wire [1:0] _T_1885;
  wire [55:0] _T_1886;
  wire [55:0] _T_1893;
  wire  _T_1895;
  wire [55:0] _T_1903;
  wire  _T_1905;
  wire [55:0] _T_1911;
  wire  _T_1913;
  wire  _T_1915;
  wire  _T_1916;
  wire  _T_1918;
  wire  _T_1919;
  wire  _T_1921;
  wire  _T_1922;
  reg  _T_1924;
  reg [31:0] _RAND_10;
  wire [1:0] _T_1925;
  wire [55:0] _T_1926;
  wire [55:0] _T_1933;
  wire  _T_1935;
  wire [55:0] _T_1943;
  wire  _T_1945;
  wire [55:0] _T_1951;
  wire  _T_1953;
  wire  _T_1955;
  wire  _T_1956;
  wire  _T_1958;
  wire  _T_1959;
  wire  _T_1961;
  wire  _T_1962;
  reg  _T_1964;
  reg [31:0] _RAND_11;
  wire [1:0] _T_1965;
  wire [55:0] _T_1966;
  wire [55:0] _T_1973;
  wire  _T_1975;
  wire [55:0] _T_1983;
  wire  _T_1985;
  wire [55:0] _T_1991;
  wire  _T_1993;
  wire  _T_1995;
  wire  _T_1996;
  wire  _T_1998;
  wire  _T_1999;
  wire  _T_2001;
  wire  _T_2002;
  reg  _T_2004;
  reg [31:0] _RAND_12;
  wire [1:0] _T_2005;
  wire [55:0] _T_2006;
  wire [55:0] _T_2013;
  wire  _T_2015;
  wire [55:0] _T_2023;
  wire  _T_2025;
  wire [55:0] _T_2031;
  wire  _T_2033;
  wire  _T_2035;
  wire  _T_2036;
  wire  _T_2038;
  wire  _T_2039;
  wire  _T_2041;
  wire  _T_2042;
  reg  _T_2044;
  reg [31:0] _RAND_13;
  wire [1:0] _T_2045;
  wire [55:0] _T_2046;
  wire [55:0] _T_2053;
  wire  _T_2055;
  wire [55:0] _T_2063;
  wire  _T_2065;
  wire [55:0] _T_2071;
  wire  _T_2073;
  wire  _T_2075;
  wire  _T_2076;
  wire  _T_2078;
  wire  _T_2079;
  wire  _T_2081;
  wire  _T_2082;
  reg  _T_2084;
  reg [31:0] _RAND_14;
  wire [1:0] _T_2085;
  wire [55:0] _T_2086;
  wire [55:0] _T_2093;
  wire  _T_2095;
  wire [55:0] _T_2103;
  wire  _T_2105;
  wire [55:0] _T_2111;
  wire  _T_2113;
  wire  _T_2115;
  wire  _T_2116;
  wire  _T_2118;
  wire  _T_2119;
  wire  _T_2121;
  wire  _T_2122;
  reg  _T_2124;
  reg [31:0] _RAND_15;
  wire [1:0] _T_2125;
  wire [55:0] _T_2126;
  wire [55:0] _T_2133;
  wire  _T_2135;
  wire [55:0] _T_2143;
  wire  _T_2145;
  wire [55:0] _T_2151;
  wire  _T_2153;
  wire  _T_2155;
  wire  _T_2156;
  wire  _T_2158;
  wire  _T_2159;
  wire  _T_2161;
  wire  _T_2162;
  reg  _T_2164;
  reg [31:0] _RAND_16;
  wire [1:0] _T_2165;
  wire [55:0] _T_2166;
  wire [55:0] _T_2173;
  wire  _T_2175;
  wire [55:0] _T_2183;
  wire  _T_2185;
  wire [55:0] _T_2191;
  wire  _T_2193;
  wire  _T_2195;
  wire  _T_2196;
  wire  _T_2198;
  wire  _T_2199;
  wire  _T_2201;
  wire  _T_2202;
  reg  _T_2204;
  reg [31:0] _RAND_17;
  wire [1:0] _T_2205;
  wire [55:0] _T_2206;
  wire [55:0] _T_2213;
  wire  _T_2215;
  wire [55:0] _T_2223;
  wire  _T_2225;
  wire [55:0] _T_2231;
  wire  _T_2233;
  wire  _T_2235;
  wire  _T_2236;
  wire  _T_2238;
  wire  _T_2239;
  wire  _T_2241;
  wire  _T_2242;
  reg  _T_2244;
  reg [31:0] _RAND_18;
  wire [1:0] _T_2245;
  wire [55:0] _T_2246;
  wire [55:0] _T_2253;
  wire  _T_2255;
  wire [55:0] _T_2263;
  wire  _T_2265;
  wire [55:0] _T_2271;
  wire  _T_2273;
  wire  _T_2275;
  wire  _T_2276;
  wire  _T_2278;
  wire  _T_2279;
  wire  _T_2281;
  wire  _T_2282;
  reg  _T_2284;
  reg [31:0] _RAND_19;
  wire [1:0] _T_2285;
  wire [55:0] _T_2286;
  wire [55:0] _T_2293;
  wire  _T_2295;
  wire [55:0] _T_2303;
  wire  _T_2305;
  wire [55:0] _T_2311;
  wire  _T_2313;
  wire  _T_2315;
  wire  _T_2316;
  wire  _T_2318;
  wire  _T_2319;
  wire  _T_2321;
  wire  _T_2322;
  reg  _T_2324;
  reg [31:0] _RAND_20;
  wire [1:0] _T_2325;
  wire [55:0] _T_2326;
  wire [55:0] _T_2333;
  wire  _T_2335;
  wire [55:0] _T_2343;
  wire  _T_2345;
  wire [55:0] _T_2351;
  wire  _T_2353;
  wire  _T_2355;
  wire  _T_2356;
  wire  _T_2358;
  wire  _T_2359;
  wire  _T_2361;
  wire  _T_2362;
  reg  _T_2364;
  reg [31:0] _RAND_21;
  wire [1:0] _T_2365;
  wire [55:0] _T_2366;
  wire [55:0] _T_2373;
  wire  _T_2375;
  wire [55:0] _T_2383;
  wire  _T_2385;
  wire [55:0] _T_2391;
  wire  _T_2393;
  wire  _T_2395;
  wire  _T_2396;
  wire  _T_2398;
  wire  _T_2399;
  wire  _T_2401;
  wire  _T_2402;
  reg  _T_2404;
  reg [31:0] _RAND_22;
  wire [1:0] _T_2405;
  wire [55:0] _T_2406;
  wire [55:0] _T_2413;
  wire  _T_2415;
  wire [55:0] _T_2423;
  wire  _T_2425;
  wire [55:0] _T_2431;
  wire  _T_2433;
  wire  _T_2435;
  wire  _T_2436;
  wire  _T_2438;
  wire  _T_2439;
  wire  _T_2441;
  wire  _T_2442;
  reg  _T_2444;
  reg [31:0] _RAND_23;
  wire [1:0] _T_2445;
  wire [55:0] _T_2446;
  wire [55:0] _T_2453;
  wire  _T_2455;
  wire [55:0] _T_2463;
  wire  _T_2465;
  wire [55:0] _T_2471;
  wire  _T_2473;
  wire  _T_2475;
  wire  _T_2476;
  wire  _T_2478;
  wire  _T_2479;
  wire  _T_2481;
  wire  _T_2482;
  reg  _T_2484;
  reg [31:0] _RAND_24;
  wire [1:0] _T_2485;
  wire [55:0] _T_2486;
  wire [55:0] _T_2493;
  wire  _T_2495;
  wire [55:0] _T_2503;
  wire  _T_2505;
  wire [55:0] _T_2511;
  wire  _T_2513;
  wire  _T_2515;
  wire  _T_2516;
  wire  _T_2518;
  wire  _T_2519;
  wire  _T_2521;
  wire  _T_2522;
  reg  _T_2524;
  reg [31:0] _RAND_25;
  wire [1:0] _T_2525;
  wire [55:0] _T_2526;
  wire [55:0] _T_2533;
  wire  _T_2535;
  wire [55:0] _T_2543;
  wire  _T_2545;
  wire [55:0] _T_2551;
  wire  _T_2553;
  wire  _T_2555;
  wire  _T_2556;
  wire  _T_2558;
  wire  _T_2559;
  wire  _T_2561;
  wire  _T_2562;
  reg  _T_2564;
  reg [31:0] _RAND_26;
  wire [1:0] _T_2565;
  wire [55:0] _T_2566;
  wire [55:0] _T_2573;
  wire  _T_2575;
  wire [55:0] _T_2583;
  wire  _T_2585;
  wire [55:0] _T_2591;
  wire  _T_2593;
  wire  _T_2595;
  wire  _T_2596;
  wire  _T_2598;
  wire  _T_2599;
  wire  _T_2601;
  wire  _T_2602;
  reg  _T_2604;
  reg [31:0] _RAND_27;
  wire [1:0] _T_2605;
  wire [55:0] _T_2606;
  wire [55:0] _T_2613;
  wire  _T_2615;
  wire [55:0] _T_2623;
  wire  _T_2625;
  wire [55:0] _T_2631;
  wire  _T_2633;
  wire  _T_2635;
  wire  _T_2636;
  wire  _T_2638;
  wire  _T_2639;
  wire  _T_2641;
  wire  _T_2642;
  reg  _T_2644;
  reg [31:0] _RAND_28;
  wire [1:0] _T_2645;
  wire [55:0] _T_2646;
  wire [55:0] _T_2653;
  wire  _T_2655;
  wire [55:0] _T_2663;
  wire  _T_2665;
  wire [55:0] _T_2671;
  wire  _T_2673;
  wire  _T_2675;
  wire  _T_2676;
  wire  _T_2678;
  wire  _T_2679;
  wire  _T_2681;
  wire  _T_2682;
  reg  _T_2684;
  reg [31:0] _RAND_29;
  reg [63:0] debug_tsc_reg;
  reg [63:0] _RAND_30;
  reg [63:0] debug_irt_reg;
  reg [63:0] _RAND_31;
  wire [64:0] _T_2693;
  wire [63:0] _T_2694;
  wire [1:0] _T_2695;
  wire  _T_2696;
  wire  _T_2697;
  wire [1:0] _T_2698;
  wire [63:0] _GEN_100;
  wire [64:0] _T_2699;
  wire [63:0] _T_2700;
  wire  _T_2701;
  wire  _T_2702;
  reg  _T_2704;
  reg [31:0] _RAND_32;
  wire  _T_2705;
  wire  _T_2706;
  wire  _T_2707;
  wire  _T_2708;
  wire  _T_2710;
  wire  _T_2711;
  reg  _T_2715_valid;
  reg [31:0] _RAND_33;
  reg  _T_2715_bits_rs1;
  reg [31:0] _RAND_34;
  reg  _T_2715_bits_rs2;
  reg [31:0] _RAND_35;
  reg [38:0] _T_2715_bits_addr;
  reg [63:0] _RAND_36;
  reg [1:0] dec_finished_mask;
  reg [31:0] _RAND_37;
  wire  branch_mask_full_0;
  wire  branch_mask_full_1;
  wire  _T_2731;
  wire  _T_2732;
  wire  _T_2734;
  wire  _T_2735;
  wire  _T_2738;
  wire  _T_2739;
  wire  _T_2741;
  wire  _T_2743;
  wire  _T_2744;
  wire  _T_2746;
  wire  _T_2747;
  wire  _T_2749;
  wire  _T_2750;
  wire  _T_2751;
  wire  _T_2752;
  wire  _T_2753;
  wire  _T_2754;
  wire  _T_2755;
  wire  _T_2758;
  wire  _T_2759;
  wire  _T_2760;
  wire  _T_2763;
  wire  _T_2764;
  wire  _T_2765;
  wire  _T_2768;
  wire  _T_2770;
  wire  _T_2771;
  wire  _T_2773;
  wire  _T_2774;
  wire  _T_2775;
  wire  _T_2776;
  wire  _T_2778;
  wire  _T_2779;
  wire  _T_2783;
  wire  _T_2784;
  wire  _T_2790;
  wire  _T_2791;
  wire  _T_2792;
  wire  _T_2795;
  wire  _T_2796;
  wire  _T_2797;
  wire  _T_2798;
  wire  _T_2799;
  wire  _T_2800;
  wire  _T_2801;
  wire  _T_2804;
  wire  _T_2805;
  wire  _T_2808;
  wire  _T_2809;
  wire  _T_2810;
  wire  dec_last_inst_was_stalled;
  wire  dec_stall_next_inst;
  wire  _T_2813;
  wire  _T_2814;
  wire  _T_2817;
  wire  _T_2819;
  wire  _T_2820;
  wire [1:0] _T_2822;
  wire [1:0] _T_2823;
  wire [1:0] _GEN_0;
  wire  _T_2827;
  wire  _T_2828;
  wire  _T_2832;
  wire  _T_2833;
  wire [3:0] new_ldq_idx;
  wire [3:0] new_stq_idx;
  wire  _T_2836;
  wire [4:0] _T_2838;
  wire [3:0] _T_2839;
  wire [3:0] _T_2841;
  wire  _T_2842;
  wire [4:0] _T_2844;
  wire [3:0] _T_2845;
  wire [3:0] _T_2847;
  wire [7:0] _T_2859;
  wire [7:0] _T_2861;
  wire  _T_2862;
  wire  _T_2864;
  wire  _T_2865;
  wire  _T_2866;
  wire  _T_2868;
  wire  _T_2869;
  wire  dec_has_br_or_jalr_in_packet;
  wire  _T_2870;
  wire  _T_2872;
  wire  _T_2873;
  wire  _T_2874;
  wire [1:0] _T_2882;
  wire [1:0] _T_2883;
  wire [1:0] _T_2884;
  wire [1:0] _T_2885;
  wire [1:0] dis_readys;
  wire  _T_2886;
  wire  _T_2887;
  wire [1:0] _T_2899_0_bim_resp_value;
  wire [5:0] _T_2899_0_bim_resp_entry_idx;
  wire [1:0] _T_2899_0_bim_resp_way_idx;
  wire [14:0] _T_2899_0_bpd_resp_history;
  wire [7:0] _T_2899_0_bpd_resp_history_ptr;
  wire [1:0] _T_2899_1_bim_resp_value;
  wire [5:0] _T_2899_1_bim_resp_entry_idx;
  wire [1:0] _T_2899_1_bim_resp_way_idx;
  wire [14:0] _T_2899_1_bpd_resp_history;
  wire [7:0] _T_2899_1_bpd_resp_history_ptr;
  reg [2:0] _T_2923;
  reg [31:0] _RAND_38;
  reg [1:0] _T_2928_bim_resp_value;
  reg [31:0] _RAND_39;
  reg [5:0] _T_2928_bim_resp_entry_idx;
  reg [31:0] _RAND_40;
  reg [1:0] _T_2928_bim_resp_way_idx;
  reg [31:0] _RAND_41;
  reg [14:0] _T_2928_bpd_resp_history;
  reg [31:0] _RAND_42;
  reg [7:0] _T_2928_bpd_resp_history_ptr;
  reg [31:0] _RAND_43;
  wire  _T_2932;
  wire  _T_2933;
  wire  _T_2934;
  wire  _T_2935;
  wire  _T_2936;
  wire  _T_2937;
  wire  _T_2938;
  wire  _T_2940;
  wire  _T_2942;
  wire  _T_2944;
  wire  _T_2945;
  wire  _T_2947;
  wire  _T_2948;
  wire  _T_2949;
  wire  _T_2950;
  wire  _T_2951;
  wire  _T_2952;
  wire  _T_2953;
  wire  _T_2954;
  wire  _T_2955;
  wire  _T_2956;
  wire  _T_2958;
  wire  _T_2960;
  wire  _T_2962;
  wire  _T_2963;
  wire  _T_2965;
  wire  _T_2966;
  wire  _T_2967;
  wire  _T_2968;
  wire  _T_2974_valid;
  wire [8:0] _T_2974_uopc;
  wire [31:0] _T_2974_inst;
  wire [39:0] _T_2974_pc;
  wire [1:0] _T_2974_iqtype;
  wire [9:0] _T_2974_fu_code;
  wire  _T_2974_allocate_brtag;
  wire  _T_2974_is_br_or_jmp;
  wire  _T_2974_is_jump;
  wire  _T_2974_is_jal;
  wire  _T_2974_is_ret;
  wire  _T_2974_is_call;
  wire [7:0] _T_2974_br_mask;
  wire [2:0] _T_2974_br_tag;
  wire  _T_2974_br_prediction_btb_blame;
  wire  _T_2974_br_prediction_btb_hit;
  wire  _T_2974_br_prediction_btb_taken;
  wire  _T_2974_br_prediction_bpd_blame;
  wire  _T_2974_br_prediction_bpd_hit;
  wire  _T_2974_br_prediction_bpd_taken;
  wire [1:0] _T_2974_br_prediction_bim_resp_value;
  wire [5:0] _T_2974_br_prediction_bim_resp_entry_idx;
  wire [1:0] _T_2974_br_prediction_bim_resp_way_idx;
  wire [1:0] _T_2974_br_prediction_bpd_resp_takens;
  wire [14:0] _T_2974_br_prediction_bpd_resp_history;
  wire [14:0] _T_2974_br_prediction_bpd_resp_history_u;
  wire [7:0] _T_2974_br_prediction_bpd_resp_history_ptr;
  wire [14:0] _T_2974_br_prediction_bpd_resp_info;
  wire  _T_2974_stat_brjmp_mispredicted;
  wire  _T_2974_stat_btb_made_pred;
  wire  _T_2974_stat_btb_mispredicted;
  wire  _T_2974_stat_bpd_made_pred;
  wire  _T_2974_stat_bpd_mispredicted;
  wire [2:0] _T_2974_fetch_pc_lob;
  wire [19:0] _T_2974_imm_packed;
  wire [11:0] _T_2974_csr_addr;
  wire [6:0] _T_2974_rob_idx;
  wire [3:0] _T_2974_ldq_idx;
  wire [3:0] _T_2974_stq_idx;
  wire [5:0] _T_2974_brob_idx;
  wire [6:0] _T_2974_pdst;
  wire [6:0] _T_2974_pop1;
  wire [6:0] _T_2974_pop2;
  wire [6:0] _T_2974_pop3;
  wire  _T_2974_prs1_busy;
  wire  _T_2974_prs2_busy;
  wire  _T_2974_prs3_busy;
  wire [6:0] _T_2974_stale_pdst;
  wire  _T_2974_exception;
  wire [63:0] _T_2974_exc_cause;
  wire  _T_2974_bypassable;
  wire [4:0] _T_2974_mem_cmd;
  wire [2:0] _T_2974_mem_typ;
  wire  _T_2974_is_fence;
  wire  _T_2974_is_fencei;
  wire  _T_2974_is_store;
  wire  _T_2974_is_amo;
  wire  _T_2974_is_load;
  wire  _T_2974_is_sys_pc2epc;
  wire  _T_2974_is_unique;
  wire  _T_2974_flush_on_commit;
  wire [5:0] _T_2974_ldst;
  wire [5:0] _T_2974_lrs1;
  wire [5:0] _T_2974_lrs2;
  wire [5:0] _T_2974_lrs3;
  wire  _T_2974_ldst_val;
  wire [1:0] _T_2974_dst_rtype;
  wire [1:0] _T_2974_lrs1_rtype;
  wire [1:0] _T_2974_lrs2_rtype;
  wire  _T_2974_frs3_en;
  wire  _T_2974_fp_val;
  wire  _T_2974_fp_single;
  wire  _T_2974_xcpt_pf_if;
  wire  _T_2974_xcpt_ae_if;
  wire  _T_2974_replay_if;
  wire  _T_2974_xcpt_ma_if;
  wire [63:0] _T_2974_debug_wdata;
  wire [31:0] _T_2974_debug_events_fetch_seq;
  wire [7:0] _T_2979;
  wire [7:0] _T_2980;
  wire [7:0] _T_2981;
  wire  _T_2987_valid;
  wire [8:0] _T_2987_uopc;
  wire [31:0] _T_2987_inst;
  wire [39:0] _T_2987_pc;
  wire [1:0] _T_2987_iqtype;
  wire [9:0] _T_2987_fu_code;
  wire  _T_2987_allocate_brtag;
  wire  _T_2987_is_br_or_jmp;
  wire  _T_2987_is_jump;
  wire  _T_2987_is_jal;
  wire  _T_2987_is_ret;
  wire  _T_2987_is_call;
  wire [7:0] _T_2987_br_mask;
  wire [2:0] _T_2987_br_tag;
  wire  _T_2987_br_prediction_btb_blame;
  wire  _T_2987_br_prediction_btb_hit;
  wire  _T_2987_br_prediction_btb_taken;
  wire  _T_2987_br_prediction_bpd_blame;
  wire  _T_2987_br_prediction_bpd_hit;
  wire  _T_2987_br_prediction_bpd_taken;
  wire [1:0] _T_2987_br_prediction_bim_resp_value;
  wire [5:0] _T_2987_br_prediction_bim_resp_entry_idx;
  wire [1:0] _T_2987_br_prediction_bim_resp_way_idx;
  wire [1:0] _T_2987_br_prediction_bpd_resp_takens;
  wire [14:0] _T_2987_br_prediction_bpd_resp_history;
  wire [14:0] _T_2987_br_prediction_bpd_resp_history_u;
  wire [7:0] _T_2987_br_prediction_bpd_resp_history_ptr;
  wire [14:0] _T_2987_br_prediction_bpd_resp_info;
  wire  _T_2987_stat_brjmp_mispredicted;
  wire  _T_2987_stat_btb_made_pred;
  wire  _T_2987_stat_btb_mispredicted;
  wire  _T_2987_stat_bpd_made_pred;
  wire  _T_2987_stat_bpd_mispredicted;
  wire [2:0] _T_2987_fetch_pc_lob;
  wire [19:0] _T_2987_imm_packed;
  wire [11:0] _T_2987_csr_addr;
  wire [6:0] _T_2987_rob_idx;
  wire [3:0] _T_2987_ldq_idx;
  wire [3:0] _T_2987_stq_idx;
  wire [5:0] _T_2987_brob_idx;
  wire [6:0] _T_2987_pdst;
  wire [6:0] _T_2987_pop1;
  wire [6:0] _T_2987_pop2;
  wire [6:0] _T_2987_pop3;
  wire  _T_2987_prs1_busy;
  wire  _T_2987_prs2_busy;
  wire  _T_2987_prs3_busy;
  wire [6:0] _T_2987_stale_pdst;
  wire  _T_2987_exception;
  wire [63:0] _T_2987_exc_cause;
  wire  _T_2987_bypassable;
  wire [4:0] _T_2987_mem_cmd;
  wire [2:0] _T_2987_mem_typ;
  wire  _T_2987_is_fence;
  wire  _T_2987_is_fencei;
  wire  _T_2987_is_store;
  wire  _T_2987_is_amo;
  wire  _T_2987_is_load;
  wire  _T_2987_is_sys_pc2epc;
  wire  _T_2987_is_unique;
  wire  _T_2987_flush_on_commit;
  wire [5:0] _T_2987_ldst;
  wire [5:0] _T_2987_lrs1;
  wire [5:0] _T_2987_lrs2;
  wire [5:0] _T_2987_lrs3;
  wire  _T_2987_ldst_val;
  wire [1:0] _T_2987_dst_rtype;
  wire [1:0] _T_2987_lrs1_rtype;
  wire [1:0] _T_2987_lrs2_rtype;
  wire  _T_2987_frs3_en;
  wire  _T_2987_fp_val;
  wire  _T_2987_fp_single;
  wire  _T_2987_xcpt_pf_if;
  wire  _T_2987_xcpt_ae_if;
  wire  _T_2987_replay_if;
  wire  _T_2987_xcpt_ma_if;
  wire [63:0] _T_2987_debug_wdata;
  wire [31:0] _T_2987_debug_events_fetch_seq;
  wire [7:0] _T_2993;
  wire [7:0] _T_2994;
  wire  _T_2996;
  wire  _T_2997;
  wire  _T_2998;
  wire  _T_2999;
  wire  _T_3000;
  wire [1:0] _GEN_1;
  wire  _GEN_2;
  wire  _T_3003;
  wire  _T_3004;
  wire  _T_3005;
  wire  _T_3006;
  wire  _T_3007;
  wire [1:0] _GEN_3;
  wire  _GEN_4;
  wire  _T_3010;
  wire  _T_3011;
  wire  _T_3017;
  wire  _T_3018;
  wire  _T_3023;
  wire  _T_3024;
  wire [9:0] _T_3026;
  wire [9:0] _T_3027;
  reg [9:0] _T_3029;
  reg [31:0] _RAND_44;
  wire [9:0] _T_3030;
  wire [2:0] _T_3033;
  wire  _T_3038;
  wire  _GEN_9;
  wire  _T_3041;
  wire  _T_3042;
  wire  _T_3044;
  wire  _T_3045;
  wire  _T_3046;
  wire  _T_3051;
  wire  _T_3052;
  wire  _T_3055;
  wire  _T_3056;
  wire  _T_3061;
  wire  _T_3064;
  wire  _T_3065;
  wire  _T_3066;
  wire  _T_3067;
  wire  _T_3069;
  wire  _T_3071;
  wire  _T_3073;
  wire  _T_3075;
  wire  _T_3077;
  wire  _T_3078;
  wire  _T_3081;
  wire  _T_3082;
  wire  _T_3084;
  wire  _T_3086;
  wire  _T_3088;
  wire  _T_3090;
  wire  _T_3092;
  wire  _T_3095;
  wire [63:0] _T_3096;
  wire  _T_3098;
  wire  _T_3099;
  wire  _T_3101;
  wire  _T_3103;
  wire  _T_3105;
  wire  _T_3107;
  wire  _T_3108;
  wire  _T_3110;
  wire  _T_3112;
  wire  _T_3114;
  wire  _T_3116;
  wire  _T_3118;
  wire  _T_3119;
  wire  _T_3121;
  wire  _T_3123;
  wire  _T_3125;
  wire  _T_3130;
  wire  _T_3132;
  wire  _T_3133;
  wire  _T_3135;
  wire  _T_3137;
  wire  _T_3139;
  wire  _T_3141;
  wire  _T_3142;
  wire  _T_3144;
  wire  _T_3146;
  wire  _T_3148;
  wire  _T_3150;
  wire  _T_3152;
  wire  _T_3153;
  wire  _T_3155;
  wire  _T_3157;
  wire  _T_3159;
  wire  _T_3175_valid;
  wire [6:0] _T_3175_bits_addr;
  wire [63:0] _T_3175_bits_data;
  wire  _T_3182;
  wire  _T_3184;
  wire  _T_3185;
  wire  _T_3188;
  wire  _T_3189;
  wire  _T_3190;
  wire  _T_3192;
  wire  _T_3194;
  wire  _T_3196;
  wire  _T_3197;
  wire  _T_3199;
  wire  _T_3200;
  wire  _T_3204;
  wire  _T_3206;
  wire  _T_3207;
  wire  _T_3208;
  wire  _T_3210;
  wire  _T_3212;
  wire  _T_3214;
  wire  _T_3216;
  wire  _T_3217;
  wire  _T_3219;
  wire  _T_3220;
  wire  _T_3228;
  wire  _T_3229;
  wire  _T_3231;
  wire  _T_3232;
  wire  _T_3353;
  wire  _T_3354;
  wire  _T_3356;
  wire  _T_3358;
  wire  _T_3360;
  wire  _T_3362;
  wire  _T_3363;
  wire  _T_3365;
  wire  _T_3367;
  wire  _T_3369;
  wire  _T_3487;
  wire  _T_3488;
  wire  _T_3490;
  wire  _T_3492;
  wire  _T_3494;
  wire  _T_3496;
  wire  _T_3497;
  wire  _T_3499;
  wire  _T_3501;
  wire  _T_3503;
  reg [6:0] _T_3505;
  reg [31:0] _RAND_45;
  reg [39:0] _T_3507;
  reg [63:0] _RAND_46;
  reg [5:0] _T_3509;
  reg [31:0] _RAND_47;
  reg  _T_3511;
  reg [31:0] _RAND_48;
  reg [39:0] _T_3513;
  reg [63:0] _RAND_49;
  wire  _T_3516;
  wire  _T_3518;
  wire  _T_3520;
  wire  _T_3521;
  reg  _T_3523;
  reg [31:0] _RAND_50;
  wire  _T_3526;
  wire  _T_3528;
  wire  _T_3530;
  wire  _T_3532;
  reg [4:0] _T_3536;
  reg [31:0] _RAND_51;
  wire [5:0] _T_3537;
  reg [26:0] _T_3540;
  reg [31:0] _RAND_52;
  wire  _T_3541;
  wire [27:0] _T_3543;
  wire [26:0] _T_3544;
  wire [26:0] _GEN_10;
  wire [31:0] _T_3545;
  wire  _T_3548;
  wire  _T_3549;
  wire  _T_3551;
  wire [5:0] _GEN_11;
  wire [26:0] _GEN_12;
  wire  _T_3554;
  wire  _T_3556;
  wire  _T_3558;
  wire  _T_3560;
  MemExeUnit mem_unit (
    .clock(mem_unit_clock),
    .reset(mem_unit_reset),
    .io_req_valid(mem_unit_io_req_valid),
    .io_req_bits_uop_uopc(mem_unit_io_req_bits_uop_uopc),
    .io_req_bits_uop_ctrl_is_load(mem_unit_io_req_bits_uop_ctrl_is_load),
    .io_req_bits_uop_ctrl_is_sta(mem_unit_io_req_bits_uop_ctrl_is_sta),
    .io_req_bits_uop_ctrl_is_std(mem_unit_io_req_bits_uop_ctrl_is_std),
    .io_req_bits_uop_br_mask(mem_unit_io_req_bits_uop_br_mask),
    .io_req_bits_uop_imm_packed(mem_unit_io_req_bits_uop_imm_packed),
    .io_req_bits_uop_rob_idx(mem_unit_io_req_bits_uop_rob_idx),
    .io_req_bits_uop_ldq_idx(mem_unit_io_req_bits_uop_ldq_idx),
    .io_req_bits_uop_stq_idx(mem_unit_io_req_bits_uop_stq_idx),
    .io_req_bits_uop_pdst(mem_unit_io_req_bits_uop_pdst),
    .io_req_bits_uop_mem_cmd(mem_unit_io_req_bits_uop_mem_cmd),
    .io_req_bits_uop_mem_typ(mem_unit_io_req_bits_uop_mem_typ),
    .io_req_bits_uop_is_fence(mem_unit_io_req_bits_uop_is_fence),
    .io_req_bits_uop_is_store(mem_unit_io_req_bits_uop_is_store),
    .io_req_bits_uop_is_amo(mem_unit_io_req_bits_uop_is_amo),
    .io_req_bits_uop_is_load(mem_unit_io_req_bits_uop_is_load),
    .io_req_bits_uop_dst_rtype(mem_unit_io_req_bits_uop_dst_rtype),
    .io_req_bits_uop_fp_val(mem_unit_io_req_bits_uop_fp_val),
    .io_req_bits_rs1_data(mem_unit_io_req_bits_rs1_data),
    .io_req_bits_rs2_data(mem_unit_io_req_bits_rs2_data),
    .io_resp_0_valid(mem_unit_io_resp_0_valid),
    .io_resp_0_bits_uop_uopc(mem_unit_io_resp_0_bits_uop_uopc),
    .io_resp_0_bits_uop_ctrl_rf_wen(mem_unit_io_resp_0_bits_uop_ctrl_rf_wen),
    .io_resp_0_bits_uop_rob_idx(mem_unit_io_resp_0_bits_uop_rob_idx),
    .io_resp_0_bits_uop_pdst(mem_unit_io_resp_0_bits_uop_pdst),
    .io_resp_0_bits_uop_mem_typ(mem_unit_io_resp_0_bits_uop_mem_typ),
    .io_resp_0_bits_uop_is_store(mem_unit_io_resp_0_bits_uop_is_store),
    .io_resp_0_bits_uop_is_amo(mem_unit_io_resp_0_bits_uop_is_amo),
    .io_resp_0_bits_uop_dst_rtype(mem_unit_io_resp_0_bits_uop_dst_rtype),
    .io_resp_0_bits_uop_fp_val(mem_unit_io_resp_0_bits_uop_fp_val),
    .io_resp_0_bits_data(mem_unit_io_resp_0_bits_data),
    .io_brinfo_valid(mem_unit_io_brinfo_valid),
    .io_brinfo_mispredict(mem_unit_io_brinfo_mispredict),
    .io_brinfo_mask(mem_unit_io_brinfo_mask),
    .io_lsu_io_exe_resp_valid(mem_unit_io_lsu_io_exe_resp_valid),
    .io_lsu_io_exe_resp_bits_uop_uopc(mem_unit_io_lsu_io_exe_resp_bits_uop_uopc),
    .io_lsu_io_exe_resp_bits_uop_ctrl_is_load(mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_load),
    .io_lsu_io_exe_resp_bits_uop_ctrl_is_sta(mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_sta),
    .io_lsu_io_exe_resp_bits_uop_ctrl_is_std(mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_std),
    .io_lsu_io_exe_resp_bits_uop_br_mask(mem_unit_io_lsu_io_exe_resp_bits_uop_br_mask),
    .io_lsu_io_exe_resp_bits_uop_rob_idx(mem_unit_io_lsu_io_exe_resp_bits_uop_rob_idx),
    .io_lsu_io_exe_resp_bits_uop_ldq_idx(mem_unit_io_lsu_io_exe_resp_bits_uop_ldq_idx),
    .io_lsu_io_exe_resp_bits_uop_stq_idx(mem_unit_io_lsu_io_exe_resp_bits_uop_stq_idx),
    .io_lsu_io_exe_resp_bits_uop_pdst(mem_unit_io_lsu_io_exe_resp_bits_uop_pdst),
    .io_lsu_io_exe_resp_bits_uop_mem_cmd(mem_unit_io_lsu_io_exe_resp_bits_uop_mem_cmd),
    .io_lsu_io_exe_resp_bits_uop_mem_typ(mem_unit_io_lsu_io_exe_resp_bits_uop_mem_typ),
    .io_lsu_io_exe_resp_bits_uop_is_fence(mem_unit_io_lsu_io_exe_resp_bits_uop_is_fence),
    .io_lsu_io_exe_resp_bits_uop_is_store(mem_unit_io_lsu_io_exe_resp_bits_uop_is_store),
    .io_lsu_io_exe_resp_bits_uop_is_amo(mem_unit_io_lsu_io_exe_resp_bits_uop_is_amo),
    .io_lsu_io_exe_resp_bits_uop_is_load(mem_unit_io_lsu_io_exe_resp_bits_uop_is_load),
    .io_lsu_io_exe_resp_bits_uop_dst_rtype(mem_unit_io_lsu_io_exe_resp_bits_uop_dst_rtype),
    .io_lsu_io_exe_resp_bits_uop_fp_val(mem_unit_io_lsu_io_exe_resp_bits_uop_fp_val),
    .io_lsu_io_exe_resp_bits_data(mem_unit_io_lsu_io_exe_resp_bits_data),
    .io_lsu_io_exe_resp_bits_addr(mem_unit_io_lsu_io_exe_resp_bits_addr),
    .io_lsu_io_exe_resp_bits_mxcpt_valid(mem_unit_io_lsu_io_exe_resp_bits_mxcpt_valid),
    .io_lsu_io_exe_resp_bits_mxcpt_bits(mem_unit_io_lsu_io_exe_resp_bits_mxcpt_bits),
    .io_lsu_io_exe_resp_bits_sfence_valid(mem_unit_io_lsu_io_exe_resp_bits_sfence_valid),
    .io_lsu_io_exe_resp_bits_sfence_bits_rs1(mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs1),
    .io_lsu_io_exe_resp_bits_sfence_bits_rs2(mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs2),
    .io_lsu_io_exe_resp_bits_sfence_bits_addr(mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_addr),
    .io_lsu_io_memreq_val(mem_unit_io_lsu_io_memreq_val),
    .io_lsu_io_memreq_addr(mem_unit_io_lsu_io_memreq_addr),
    .io_lsu_io_memreq_wdata(mem_unit_io_lsu_io_memreq_wdata),
    .io_lsu_io_memreq_uop_uopc(mem_unit_io_lsu_io_memreq_uop_uopc),
    .io_lsu_io_memreq_uop_br_mask(mem_unit_io_lsu_io_memreq_uop_br_mask),
    .io_lsu_io_memreq_uop_rob_idx(mem_unit_io_lsu_io_memreq_uop_rob_idx),
    .io_lsu_io_memreq_uop_ldq_idx(mem_unit_io_lsu_io_memreq_uop_ldq_idx),
    .io_lsu_io_memreq_uop_stq_idx(mem_unit_io_lsu_io_memreq_uop_stq_idx),
    .io_lsu_io_memreq_uop_pdst(mem_unit_io_lsu_io_memreq_uop_pdst),
    .io_lsu_io_memreq_uop_mem_cmd(mem_unit_io_lsu_io_memreq_uop_mem_cmd),
    .io_lsu_io_memreq_uop_mem_typ(mem_unit_io_lsu_io_memreq_uop_mem_typ),
    .io_lsu_io_memreq_uop_is_store(mem_unit_io_lsu_io_memreq_uop_is_store),
    .io_lsu_io_memreq_uop_is_amo(mem_unit_io_lsu_io_memreq_uop_is_amo),
    .io_lsu_io_memreq_uop_is_load(mem_unit_io_lsu_io_memreq_uop_is_load),
    .io_lsu_io_memreq_uop_dst_rtype(mem_unit_io_lsu_io_memreq_uop_dst_rtype),
    .io_lsu_io_memreq_uop_fp_val(mem_unit_io_lsu_io_memreq_uop_fp_val),
    .io_lsu_io_memreq_kill(mem_unit_io_lsu_io_memreq_kill),
    .io_lsu_io_forward_val(mem_unit_io_lsu_io_forward_val),
    .io_lsu_io_forward_data(mem_unit_io_lsu_io_forward_data),
    .io_lsu_io_forward_uop_uopc(mem_unit_io_lsu_io_forward_uop_uopc),
    .io_lsu_io_forward_uop_rob_idx(mem_unit_io_lsu_io_forward_uop_rob_idx),
    .io_lsu_io_forward_uop_ldq_idx(mem_unit_io_lsu_io_forward_uop_ldq_idx),
    .io_lsu_io_forward_uop_stq_idx(mem_unit_io_lsu_io_forward_uop_stq_idx),
    .io_lsu_io_forward_uop_pdst(mem_unit_io_lsu_io_forward_uop_pdst),
    .io_lsu_io_forward_uop_mem_typ(mem_unit_io_lsu_io_forward_uop_mem_typ),
    .io_lsu_io_forward_uop_is_store(mem_unit_io_lsu_io_forward_uop_is_store),
    .io_lsu_io_forward_uop_is_amo(mem_unit_io_lsu_io_forward_uop_is_amo),
    .io_lsu_io_forward_uop_is_load(mem_unit_io_lsu_io_forward_uop_is_load),
    .io_lsu_io_forward_uop_dst_rtype(mem_unit_io_lsu_io_forward_uop_dst_rtype),
    .io_lsu_io_forward_uop_fp_val(mem_unit_io_lsu_io_forward_uop_fp_val),
    .io_lsu_io_memresp_valid(mem_unit_io_lsu_io_memresp_valid),
    .io_lsu_io_memresp_bits_ldq_idx(mem_unit_io_lsu_io_memresp_bits_ldq_idx),
    .io_lsu_io_memresp_bits_stq_idx(mem_unit_io_lsu_io_memresp_bits_stq_idx),
    .io_lsu_io_memresp_bits_is_load(mem_unit_io_lsu_io_memresp_bits_is_load),
    .io_dmem_req_valid(mem_unit_io_dmem_req_valid),
    .io_dmem_req_bits_addr(mem_unit_io_dmem_req_bits_addr),
    .io_dmem_req_bits_uop_uopc(mem_unit_io_dmem_req_bits_uop_uopc),
    .io_dmem_req_bits_uop_br_mask(mem_unit_io_dmem_req_bits_uop_br_mask),
    .io_dmem_req_bits_uop_rob_idx(mem_unit_io_dmem_req_bits_uop_rob_idx),
    .io_dmem_req_bits_uop_ldq_idx(mem_unit_io_dmem_req_bits_uop_ldq_idx),
    .io_dmem_req_bits_uop_stq_idx(mem_unit_io_dmem_req_bits_uop_stq_idx),
    .io_dmem_req_bits_uop_pdst(mem_unit_io_dmem_req_bits_uop_pdst),
    .io_dmem_req_bits_uop_mem_cmd(mem_unit_io_dmem_req_bits_uop_mem_cmd),
    .io_dmem_req_bits_uop_mem_typ(mem_unit_io_dmem_req_bits_uop_mem_typ),
    .io_dmem_req_bits_uop_is_store(mem_unit_io_dmem_req_bits_uop_is_store),
    .io_dmem_req_bits_uop_is_amo(mem_unit_io_dmem_req_bits_uop_is_amo),
    .io_dmem_req_bits_uop_is_load(mem_unit_io_dmem_req_bits_uop_is_load),
    .io_dmem_req_bits_uop_dst_rtype(mem_unit_io_dmem_req_bits_uop_dst_rtype),
    .io_dmem_req_bits_uop_fp_val(mem_unit_io_dmem_req_bits_uop_fp_val),
    .io_dmem_req_bits_data(mem_unit_io_dmem_req_bits_data),
    .io_dmem_req_bits_kill(mem_unit_io_dmem_req_bits_kill),
    .io_dmem_resp_valid(mem_unit_io_dmem_resp_valid),
    .io_dmem_resp_bits_data_subword(mem_unit_io_dmem_resp_bits_data_subword),
    .io_dmem_resp_bits_uop_uopc(mem_unit_io_dmem_resp_bits_uop_uopc),
    .io_dmem_resp_bits_uop_rob_idx(mem_unit_io_dmem_resp_bits_uop_rob_idx),
    .io_dmem_resp_bits_uop_ldq_idx(mem_unit_io_dmem_resp_bits_uop_ldq_idx),
    .io_dmem_resp_bits_uop_stq_idx(mem_unit_io_dmem_resp_bits_uop_stq_idx),
    .io_dmem_resp_bits_uop_pdst(mem_unit_io_dmem_resp_bits_uop_pdst),
    .io_dmem_resp_bits_uop_mem_cmd(mem_unit_io_dmem_resp_bits_uop_mem_cmd),
    .io_dmem_resp_bits_uop_mem_typ(mem_unit_io_dmem_resp_bits_uop_mem_typ),
    .io_dmem_resp_bits_uop_is_store(mem_unit_io_dmem_resp_bits_uop_is_store),
    .io_dmem_resp_bits_uop_is_amo(mem_unit_io_dmem_resp_bits_uop_is_amo),
    .io_dmem_resp_bits_uop_is_load(mem_unit_io_dmem_resp_bits_uop_is_load),
    .io_dmem_resp_bits_uop_dst_rtype(mem_unit_io_dmem_resp_bits_uop_dst_rtype),
    .io_dmem_resp_bits_uop_fp_val(mem_unit_io_dmem_resp_bits_uop_fp_val),
    .io_com_exception(mem_unit_io_com_exception)
  );
  ALUExeUnit csr_exe_unit (
    .clock(csr_exe_unit_clock),
    .reset(csr_exe_unit_reset),
    .io_fu_types(csr_exe_unit_io_fu_types),
    .io_req_valid(csr_exe_unit_io_req_valid),
    .io_req_bits_uop_valid(csr_exe_unit_io_req_bits_uop_valid),
    .io_req_bits_uop_iw_state(csr_exe_unit_io_req_bits_uop_iw_state),
    .io_req_bits_uop_uopc(csr_exe_unit_io_req_bits_uop_uopc),
    .io_req_bits_uop_inst(csr_exe_unit_io_req_bits_uop_inst),
    .io_req_bits_uop_pc(csr_exe_unit_io_req_bits_uop_pc),
    .io_req_bits_uop_iqtype(csr_exe_unit_io_req_bits_uop_iqtype),
    .io_req_bits_uop_fu_code(csr_exe_unit_io_req_bits_uop_fu_code),
    .io_req_bits_uop_ctrl_br_type(csr_exe_unit_io_req_bits_uop_ctrl_br_type),
    .io_req_bits_uop_ctrl_op1_sel(csr_exe_unit_io_req_bits_uop_ctrl_op1_sel),
    .io_req_bits_uop_ctrl_op2_sel(csr_exe_unit_io_req_bits_uop_ctrl_op2_sel),
    .io_req_bits_uop_ctrl_imm_sel(csr_exe_unit_io_req_bits_uop_ctrl_imm_sel),
    .io_req_bits_uop_ctrl_op_fcn(csr_exe_unit_io_req_bits_uop_ctrl_op_fcn),
    .io_req_bits_uop_ctrl_fcn_dw(csr_exe_unit_io_req_bits_uop_ctrl_fcn_dw),
    .io_req_bits_uop_ctrl_rf_wen(csr_exe_unit_io_req_bits_uop_ctrl_rf_wen),
    .io_req_bits_uop_ctrl_csr_cmd(csr_exe_unit_io_req_bits_uop_ctrl_csr_cmd),
    .io_req_bits_uop_ctrl_is_load(csr_exe_unit_io_req_bits_uop_ctrl_is_load),
    .io_req_bits_uop_ctrl_is_sta(csr_exe_unit_io_req_bits_uop_ctrl_is_sta),
    .io_req_bits_uop_ctrl_is_std(csr_exe_unit_io_req_bits_uop_ctrl_is_std),
    .io_req_bits_uop_allocate_brtag(csr_exe_unit_io_req_bits_uop_allocate_brtag),
    .io_req_bits_uop_is_br_or_jmp(csr_exe_unit_io_req_bits_uop_is_br_or_jmp),
    .io_req_bits_uop_is_jump(csr_exe_unit_io_req_bits_uop_is_jump),
    .io_req_bits_uop_is_jal(csr_exe_unit_io_req_bits_uop_is_jal),
    .io_req_bits_uop_is_ret(csr_exe_unit_io_req_bits_uop_is_ret),
    .io_req_bits_uop_is_call(csr_exe_unit_io_req_bits_uop_is_call),
    .io_req_bits_uop_br_mask(csr_exe_unit_io_req_bits_uop_br_mask),
    .io_req_bits_uop_br_tag(csr_exe_unit_io_req_bits_uop_br_tag),
    .io_req_bits_uop_br_prediction_btb_blame(csr_exe_unit_io_req_bits_uop_br_prediction_btb_blame),
    .io_req_bits_uop_br_prediction_btb_hit(csr_exe_unit_io_req_bits_uop_br_prediction_btb_hit),
    .io_req_bits_uop_br_prediction_btb_taken(csr_exe_unit_io_req_bits_uop_br_prediction_btb_taken),
    .io_req_bits_uop_br_prediction_bpd_blame(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_blame),
    .io_req_bits_uop_br_prediction_bpd_hit(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_hit),
    .io_req_bits_uop_br_prediction_bpd_taken(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_taken),
    .io_req_bits_uop_br_prediction_bim_resp_value(csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_value),
    .io_req_bits_uop_br_prediction_bim_resp_entry_idx(csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_entry_idx),
    .io_req_bits_uop_br_prediction_bim_resp_way_idx(csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_way_idx),
    .io_req_bits_uop_br_prediction_bpd_resp_takens(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_takens),
    .io_req_bits_uop_br_prediction_bpd_resp_history(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history),
    .io_req_bits_uop_br_prediction_bpd_resp_history_u(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_u),
    .io_req_bits_uop_br_prediction_bpd_resp_history_ptr(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr),
    .io_req_bits_uop_br_prediction_bpd_resp_info(csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_info),
    .io_req_bits_uop_stat_brjmp_mispredicted(csr_exe_unit_io_req_bits_uop_stat_brjmp_mispredicted),
    .io_req_bits_uop_stat_btb_made_pred(csr_exe_unit_io_req_bits_uop_stat_btb_made_pred),
    .io_req_bits_uop_stat_btb_mispredicted(csr_exe_unit_io_req_bits_uop_stat_btb_mispredicted),
    .io_req_bits_uop_stat_bpd_made_pred(csr_exe_unit_io_req_bits_uop_stat_bpd_made_pred),
    .io_req_bits_uop_stat_bpd_mispredicted(csr_exe_unit_io_req_bits_uop_stat_bpd_mispredicted),
    .io_req_bits_uop_fetch_pc_lob(csr_exe_unit_io_req_bits_uop_fetch_pc_lob),
    .io_req_bits_uop_imm_packed(csr_exe_unit_io_req_bits_uop_imm_packed),
    .io_req_bits_uop_csr_addr(csr_exe_unit_io_req_bits_uop_csr_addr),
    .io_req_bits_uop_rob_idx(csr_exe_unit_io_req_bits_uop_rob_idx),
    .io_req_bits_uop_ldq_idx(csr_exe_unit_io_req_bits_uop_ldq_idx),
    .io_req_bits_uop_stq_idx(csr_exe_unit_io_req_bits_uop_stq_idx),
    .io_req_bits_uop_brob_idx(csr_exe_unit_io_req_bits_uop_brob_idx),
    .io_req_bits_uop_pdst(csr_exe_unit_io_req_bits_uop_pdst),
    .io_req_bits_uop_pop1(csr_exe_unit_io_req_bits_uop_pop1),
    .io_req_bits_uop_pop2(csr_exe_unit_io_req_bits_uop_pop2),
    .io_req_bits_uop_pop3(csr_exe_unit_io_req_bits_uop_pop3),
    .io_req_bits_uop_prs1_busy(csr_exe_unit_io_req_bits_uop_prs1_busy),
    .io_req_bits_uop_prs2_busy(csr_exe_unit_io_req_bits_uop_prs2_busy),
    .io_req_bits_uop_prs3_busy(csr_exe_unit_io_req_bits_uop_prs3_busy),
    .io_req_bits_uop_stale_pdst(csr_exe_unit_io_req_bits_uop_stale_pdst),
    .io_req_bits_uop_exception(csr_exe_unit_io_req_bits_uop_exception),
    .io_req_bits_uop_exc_cause(csr_exe_unit_io_req_bits_uop_exc_cause),
    .io_req_bits_uop_bypassable(csr_exe_unit_io_req_bits_uop_bypassable),
    .io_req_bits_uop_mem_cmd(csr_exe_unit_io_req_bits_uop_mem_cmd),
    .io_req_bits_uop_mem_typ(csr_exe_unit_io_req_bits_uop_mem_typ),
    .io_req_bits_uop_is_fence(csr_exe_unit_io_req_bits_uop_is_fence),
    .io_req_bits_uop_is_fencei(csr_exe_unit_io_req_bits_uop_is_fencei),
    .io_req_bits_uop_is_store(csr_exe_unit_io_req_bits_uop_is_store),
    .io_req_bits_uop_is_amo(csr_exe_unit_io_req_bits_uop_is_amo),
    .io_req_bits_uop_is_load(csr_exe_unit_io_req_bits_uop_is_load),
    .io_req_bits_uop_is_sys_pc2epc(csr_exe_unit_io_req_bits_uop_is_sys_pc2epc),
    .io_req_bits_uop_is_unique(csr_exe_unit_io_req_bits_uop_is_unique),
    .io_req_bits_uop_flush_on_commit(csr_exe_unit_io_req_bits_uop_flush_on_commit),
    .io_req_bits_uop_ldst(csr_exe_unit_io_req_bits_uop_ldst),
    .io_req_bits_uop_lrs1(csr_exe_unit_io_req_bits_uop_lrs1),
    .io_req_bits_uop_lrs2(csr_exe_unit_io_req_bits_uop_lrs2),
    .io_req_bits_uop_lrs3(csr_exe_unit_io_req_bits_uop_lrs3),
    .io_req_bits_uop_ldst_val(csr_exe_unit_io_req_bits_uop_ldst_val),
    .io_req_bits_uop_dst_rtype(csr_exe_unit_io_req_bits_uop_dst_rtype),
    .io_req_bits_uop_lrs1_rtype(csr_exe_unit_io_req_bits_uop_lrs1_rtype),
    .io_req_bits_uop_lrs2_rtype(csr_exe_unit_io_req_bits_uop_lrs2_rtype),
    .io_req_bits_uop_frs3_en(csr_exe_unit_io_req_bits_uop_frs3_en),
    .io_req_bits_uop_fp_val(csr_exe_unit_io_req_bits_uop_fp_val),
    .io_req_bits_uop_fp_single(csr_exe_unit_io_req_bits_uop_fp_single),
    .io_req_bits_uop_xcpt_pf_if(csr_exe_unit_io_req_bits_uop_xcpt_pf_if),
    .io_req_bits_uop_xcpt_ae_if(csr_exe_unit_io_req_bits_uop_xcpt_ae_if),
    .io_req_bits_uop_replay_if(csr_exe_unit_io_req_bits_uop_replay_if),
    .io_req_bits_uop_xcpt_ma_if(csr_exe_unit_io_req_bits_uop_xcpt_ma_if),
    .io_req_bits_uop_debug_wdata(csr_exe_unit_io_req_bits_uop_debug_wdata),
    .io_req_bits_uop_debug_events_fetch_seq(csr_exe_unit_io_req_bits_uop_debug_events_fetch_seq),
    .io_req_bits_rs1_data(csr_exe_unit_io_req_bits_rs1_data),
    .io_req_bits_rs2_data(csr_exe_unit_io_req_bits_rs2_data),
    .io_req_bits_kill(csr_exe_unit_io_req_bits_kill),
    .io_resp_0_valid(csr_exe_unit_io_resp_0_valid),
    .io_resp_0_bits_uop_ctrl_rf_wen(csr_exe_unit_io_resp_0_bits_uop_ctrl_rf_wen),
    .io_resp_0_bits_uop_ctrl_csr_cmd(csr_exe_unit_io_resp_0_bits_uop_ctrl_csr_cmd),
    .io_resp_0_bits_uop_csr_addr(csr_exe_unit_io_resp_0_bits_uop_csr_addr),
    .io_resp_0_bits_uop_rob_idx(csr_exe_unit_io_resp_0_bits_uop_rob_idx),
    .io_resp_0_bits_uop_pdst(csr_exe_unit_io_resp_0_bits_uop_pdst),
    .io_resp_0_bits_uop_bypassable(csr_exe_unit_io_resp_0_bits_uop_bypassable),
    .io_resp_0_bits_uop_is_store(csr_exe_unit_io_resp_0_bits_uop_is_store),
    .io_resp_0_bits_uop_is_amo(csr_exe_unit_io_resp_0_bits_uop_is_amo),
    .io_resp_0_bits_uop_dst_rtype(csr_exe_unit_io_resp_0_bits_uop_dst_rtype),
    .io_resp_0_bits_data(csr_exe_unit_io_resp_0_bits_data),
    .io_bypass_valid_0(csr_exe_unit_io_bypass_valid_0),
    .io_bypass_valid_1(csr_exe_unit_io_bypass_valid_1),
    .io_bypass_valid_2(csr_exe_unit_io_bypass_valid_2),
    .io_bypass_uop_0_ctrl_rf_wen(csr_exe_unit_io_bypass_uop_0_ctrl_rf_wen),
    .io_bypass_uop_0_pdst(csr_exe_unit_io_bypass_uop_0_pdst),
    .io_bypass_uop_0_dst_rtype(csr_exe_unit_io_bypass_uop_0_dst_rtype),
    .io_bypass_uop_1_ctrl_rf_wen(csr_exe_unit_io_bypass_uop_1_ctrl_rf_wen),
    .io_bypass_uop_1_pdst(csr_exe_unit_io_bypass_uop_1_pdst),
    .io_bypass_uop_1_dst_rtype(csr_exe_unit_io_bypass_uop_1_dst_rtype),
    .io_bypass_uop_2_ctrl_rf_wen(csr_exe_unit_io_bypass_uop_2_ctrl_rf_wen),
    .io_bypass_uop_2_pdst(csr_exe_unit_io_bypass_uop_2_pdst),
    .io_bypass_uop_2_dst_rtype(csr_exe_unit_io_bypass_uop_2_dst_rtype),
    .io_bypass_data_0(csr_exe_unit_io_bypass_data_0),
    .io_bypass_data_1(csr_exe_unit_io_bypass_data_1),
    .io_bypass_data_2(csr_exe_unit_io_bypass_data_2),
    .io_brinfo_valid(csr_exe_unit_io_brinfo_valid),
    .io_brinfo_mispredict(csr_exe_unit_io_brinfo_mispredict),
    .io_brinfo_mask(csr_exe_unit_io_brinfo_mask),
    .io_br_unit_take_pc(csr_exe_unit_io_br_unit_take_pc),
    .io_br_unit_target(csr_exe_unit_io_br_unit_target),
    .io_br_unit_brinfo_valid(csr_exe_unit_io_br_unit_brinfo_valid),
    .io_br_unit_brinfo_mispredict(csr_exe_unit_io_br_unit_brinfo_mispredict),
    .io_br_unit_brinfo_mask(csr_exe_unit_io_br_unit_brinfo_mask),
    .io_br_unit_brinfo_tag(csr_exe_unit_io_br_unit_brinfo_tag),
    .io_br_unit_brinfo_exe_mask(csr_exe_unit_io_br_unit_brinfo_exe_mask),
    .io_br_unit_brinfo_rob_idx(csr_exe_unit_io_br_unit_brinfo_rob_idx),
    .io_br_unit_brinfo_ldq_idx(csr_exe_unit_io_br_unit_brinfo_ldq_idx),
    .io_br_unit_brinfo_stq_idx(csr_exe_unit_io_br_unit_brinfo_stq_idx),
    .io_br_unit_brinfo_is_jr(csr_exe_unit_io_br_unit_brinfo_is_jr),
    .io_br_unit_btb_update_valid(csr_exe_unit_io_br_unit_btb_update_valid),
    .io_br_unit_btb_update_bits_pc(csr_exe_unit_io_br_unit_btb_update_bits_pc),
    .io_br_unit_btb_update_bits_target(csr_exe_unit_io_br_unit_btb_update_bits_target),
    .io_br_unit_btb_update_bits_cfi_pc(csr_exe_unit_io_br_unit_btb_update_bits_cfi_pc),
    .io_br_unit_btb_update_bits_bpd_type(csr_exe_unit_io_br_unit_btb_update_bits_bpd_type),
    .io_br_unit_btb_update_bits_cfi_type(csr_exe_unit_io_br_unit_btb_update_bits_cfi_type),
    .io_br_unit_bim_update_valid(csr_exe_unit_io_br_unit_bim_update_valid),
    .io_br_unit_bim_update_bits_taken(csr_exe_unit_io_br_unit_bim_update_bits_taken),
    .io_br_unit_bim_update_bits_bim_resp_value(csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_value),
    .io_br_unit_bim_update_bits_bim_resp_entry_idx(csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_entry_idx),
    .io_br_unit_bim_update_bits_bim_resp_way_idx(csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_way_idx),
    .io_br_unit_bpd_update_valid(csr_exe_unit_io_br_unit_bpd_update_valid),
    .io_br_unit_bpd_update_bits_br_pc(csr_exe_unit_io_br_unit_bpd_update_bits_br_pc),
    .io_br_unit_bpd_update_bits_brob_idx(csr_exe_unit_io_br_unit_bpd_update_bits_brob_idx),
    .io_br_unit_bpd_update_bits_mispredict(csr_exe_unit_io_br_unit_bpd_update_bits_mispredict),
    .io_br_unit_bpd_update_bits_history(csr_exe_unit_io_br_unit_bpd_update_bits_history),
    .io_br_unit_bpd_update_bits_history_ptr(csr_exe_unit_io_br_unit_bpd_update_bits_history_ptr),
    .io_br_unit_bpd_update_bits_bpd_predict_val(csr_exe_unit_io_br_unit_bpd_update_bits_bpd_predict_val),
    .io_br_unit_bpd_update_bits_bpd_mispredict(csr_exe_unit_io_br_unit_bpd_update_bits_bpd_mispredict),
    .io_br_unit_bpd_update_bits_taken(csr_exe_unit_io_br_unit_bpd_update_bits_taken),
    .io_br_unit_bpd_update_bits_is_br(csr_exe_unit_io_br_unit_bpd_update_bits_is_br),
    .io_br_unit_bpd_update_bits_new_pc_same_packet(csr_exe_unit_io_br_unit_bpd_update_bits_new_pc_same_packet),
    .io_br_unit_xcpt_valid(csr_exe_unit_io_br_unit_xcpt_valid),
    .io_br_unit_xcpt_bits_uop_br_mask(csr_exe_unit_io_br_unit_xcpt_bits_uop_br_mask),
    .io_br_unit_xcpt_bits_uop_rob_idx(csr_exe_unit_io_br_unit_xcpt_bits_uop_rob_idx),
    .io_br_unit_xcpt_bits_badvaddr(csr_exe_unit_io_br_unit_xcpt_bits_badvaddr),
    .io_get_rob_pc_curr_pc(csr_exe_unit_io_get_rob_pc_curr_pc),
    .io_get_rob_pc_curr_brob_idx(csr_exe_unit_io_get_rob_pc_curr_brob_idx),
    .io_get_rob_pc_next_val(csr_exe_unit_io_get_rob_pc_next_val),
    .io_get_rob_pc_next_pc(csr_exe_unit_io_get_rob_pc_next_pc),
    .io_get_pred_info_bim_resp_value(csr_exe_unit_io_get_pred_info_bim_resp_value),
    .io_get_pred_info_bim_resp_entry_idx(csr_exe_unit_io_get_pred_info_bim_resp_entry_idx),
    .io_get_pred_info_bim_resp_way_idx(csr_exe_unit_io_get_pred_info_bim_resp_way_idx),
    .io_get_pred_info_bpd_resp_history(csr_exe_unit_io_get_pred_info_bpd_resp_history),
    .io_get_pred_info_bpd_resp_history_ptr(csr_exe_unit_io_get_pred_info_bpd_resp_history_ptr),
    .io_status_debug(csr_exe_unit_io_status_debug)
  );
  ALUExeUnit_1 ALUExeUnit (
    .clock(ALUExeUnit_clock),
    .reset(ALUExeUnit_reset),
    .io_req_valid(ALUExeUnit_io_req_valid),
    .io_req_bits_uop_valid(ALUExeUnit_io_req_bits_uop_valid),
    .io_req_bits_uop_iw_state(ALUExeUnit_io_req_bits_uop_iw_state),
    .io_req_bits_uop_uopc(ALUExeUnit_io_req_bits_uop_uopc),
    .io_req_bits_uop_inst(ALUExeUnit_io_req_bits_uop_inst),
    .io_req_bits_uop_pc(ALUExeUnit_io_req_bits_uop_pc),
    .io_req_bits_uop_iqtype(ALUExeUnit_io_req_bits_uop_iqtype),
    .io_req_bits_uop_fu_code(ALUExeUnit_io_req_bits_uop_fu_code),
    .io_req_bits_uop_ctrl_op1_sel(ALUExeUnit_io_req_bits_uop_ctrl_op1_sel),
    .io_req_bits_uop_ctrl_op2_sel(ALUExeUnit_io_req_bits_uop_ctrl_op2_sel),
    .io_req_bits_uop_ctrl_imm_sel(ALUExeUnit_io_req_bits_uop_ctrl_imm_sel),
    .io_req_bits_uop_ctrl_op_fcn(ALUExeUnit_io_req_bits_uop_ctrl_op_fcn),
    .io_req_bits_uop_ctrl_fcn_dw(ALUExeUnit_io_req_bits_uop_ctrl_fcn_dw),
    .io_req_bits_uop_ctrl_rf_wen(ALUExeUnit_io_req_bits_uop_ctrl_rf_wen),
    .io_req_bits_uop_ctrl_is_load(ALUExeUnit_io_req_bits_uop_ctrl_is_load),
    .io_req_bits_uop_ctrl_is_sta(ALUExeUnit_io_req_bits_uop_ctrl_is_sta),
    .io_req_bits_uop_ctrl_is_std(ALUExeUnit_io_req_bits_uop_ctrl_is_std),
    .io_req_bits_uop_allocate_brtag(ALUExeUnit_io_req_bits_uop_allocate_brtag),
    .io_req_bits_uop_is_br_or_jmp(ALUExeUnit_io_req_bits_uop_is_br_or_jmp),
    .io_req_bits_uop_is_jump(ALUExeUnit_io_req_bits_uop_is_jump),
    .io_req_bits_uop_is_jal(ALUExeUnit_io_req_bits_uop_is_jal),
    .io_req_bits_uop_is_ret(ALUExeUnit_io_req_bits_uop_is_ret),
    .io_req_bits_uop_is_call(ALUExeUnit_io_req_bits_uop_is_call),
    .io_req_bits_uop_br_mask(ALUExeUnit_io_req_bits_uop_br_mask),
    .io_req_bits_uop_br_tag(ALUExeUnit_io_req_bits_uop_br_tag),
    .io_req_bits_uop_br_prediction_btb_blame(ALUExeUnit_io_req_bits_uop_br_prediction_btb_blame),
    .io_req_bits_uop_br_prediction_btb_hit(ALUExeUnit_io_req_bits_uop_br_prediction_btb_hit),
    .io_req_bits_uop_br_prediction_btb_taken(ALUExeUnit_io_req_bits_uop_br_prediction_btb_taken),
    .io_req_bits_uop_br_prediction_bpd_blame(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_blame),
    .io_req_bits_uop_br_prediction_bpd_hit(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_hit),
    .io_req_bits_uop_br_prediction_bpd_taken(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_taken),
    .io_req_bits_uop_br_prediction_bim_resp_value(ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_value),
    .io_req_bits_uop_br_prediction_bim_resp_entry_idx(ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_entry_idx),
    .io_req_bits_uop_br_prediction_bim_resp_way_idx(ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_way_idx),
    .io_req_bits_uop_br_prediction_bpd_resp_takens(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_takens),
    .io_req_bits_uop_br_prediction_bpd_resp_history(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history),
    .io_req_bits_uop_br_prediction_bpd_resp_history_u(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_u),
    .io_req_bits_uop_br_prediction_bpd_resp_history_ptr(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr),
    .io_req_bits_uop_br_prediction_bpd_resp_info(ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_info),
    .io_req_bits_uop_stat_brjmp_mispredicted(ALUExeUnit_io_req_bits_uop_stat_brjmp_mispredicted),
    .io_req_bits_uop_stat_btb_made_pred(ALUExeUnit_io_req_bits_uop_stat_btb_made_pred),
    .io_req_bits_uop_stat_btb_mispredicted(ALUExeUnit_io_req_bits_uop_stat_btb_mispredicted),
    .io_req_bits_uop_stat_bpd_made_pred(ALUExeUnit_io_req_bits_uop_stat_bpd_made_pred),
    .io_req_bits_uop_stat_bpd_mispredicted(ALUExeUnit_io_req_bits_uop_stat_bpd_mispredicted),
    .io_req_bits_uop_fetch_pc_lob(ALUExeUnit_io_req_bits_uop_fetch_pc_lob),
    .io_req_bits_uop_imm_packed(ALUExeUnit_io_req_bits_uop_imm_packed),
    .io_req_bits_uop_csr_addr(ALUExeUnit_io_req_bits_uop_csr_addr),
    .io_req_bits_uop_rob_idx(ALUExeUnit_io_req_bits_uop_rob_idx),
    .io_req_bits_uop_ldq_idx(ALUExeUnit_io_req_bits_uop_ldq_idx),
    .io_req_bits_uop_stq_idx(ALUExeUnit_io_req_bits_uop_stq_idx),
    .io_req_bits_uop_brob_idx(ALUExeUnit_io_req_bits_uop_brob_idx),
    .io_req_bits_uop_pdst(ALUExeUnit_io_req_bits_uop_pdst),
    .io_req_bits_uop_pop1(ALUExeUnit_io_req_bits_uop_pop1),
    .io_req_bits_uop_pop2(ALUExeUnit_io_req_bits_uop_pop2),
    .io_req_bits_uop_pop3(ALUExeUnit_io_req_bits_uop_pop3),
    .io_req_bits_uop_prs1_busy(ALUExeUnit_io_req_bits_uop_prs1_busy),
    .io_req_bits_uop_prs2_busy(ALUExeUnit_io_req_bits_uop_prs2_busy),
    .io_req_bits_uop_prs3_busy(ALUExeUnit_io_req_bits_uop_prs3_busy),
    .io_req_bits_uop_stale_pdst(ALUExeUnit_io_req_bits_uop_stale_pdst),
    .io_req_bits_uop_exception(ALUExeUnit_io_req_bits_uop_exception),
    .io_req_bits_uop_exc_cause(ALUExeUnit_io_req_bits_uop_exc_cause),
    .io_req_bits_uop_bypassable(ALUExeUnit_io_req_bits_uop_bypassable),
    .io_req_bits_uop_mem_cmd(ALUExeUnit_io_req_bits_uop_mem_cmd),
    .io_req_bits_uop_mem_typ(ALUExeUnit_io_req_bits_uop_mem_typ),
    .io_req_bits_uop_is_fence(ALUExeUnit_io_req_bits_uop_is_fence),
    .io_req_bits_uop_is_fencei(ALUExeUnit_io_req_bits_uop_is_fencei),
    .io_req_bits_uop_is_store(ALUExeUnit_io_req_bits_uop_is_store),
    .io_req_bits_uop_is_amo(ALUExeUnit_io_req_bits_uop_is_amo),
    .io_req_bits_uop_is_load(ALUExeUnit_io_req_bits_uop_is_load),
    .io_req_bits_uop_is_sys_pc2epc(ALUExeUnit_io_req_bits_uop_is_sys_pc2epc),
    .io_req_bits_uop_is_unique(ALUExeUnit_io_req_bits_uop_is_unique),
    .io_req_bits_uop_flush_on_commit(ALUExeUnit_io_req_bits_uop_flush_on_commit),
    .io_req_bits_uop_ldst(ALUExeUnit_io_req_bits_uop_ldst),
    .io_req_bits_uop_lrs1(ALUExeUnit_io_req_bits_uop_lrs1),
    .io_req_bits_uop_lrs2(ALUExeUnit_io_req_bits_uop_lrs2),
    .io_req_bits_uop_lrs3(ALUExeUnit_io_req_bits_uop_lrs3),
    .io_req_bits_uop_ldst_val(ALUExeUnit_io_req_bits_uop_ldst_val),
    .io_req_bits_uop_dst_rtype(ALUExeUnit_io_req_bits_uop_dst_rtype),
    .io_req_bits_uop_lrs1_rtype(ALUExeUnit_io_req_bits_uop_lrs1_rtype),
    .io_req_bits_uop_lrs2_rtype(ALUExeUnit_io_req_bits_uop_lrs2_rtype),
    .io_req_bits_uop_frs3_en(ALUExeUnit_io_req_bits_uop_frs3_en),
    .io_req_bits_uop_fp_val(ALUExeUnit_io_req_bits_uop_fp_val),
    .io_req_bits_uop_fp_single(ALUExeUnit_io_req_bits_uop_fp_single),
    .io_req_bits_uop_xcpt_pf_if(ALUExeUnit_io_req_bits_uop_xcpt_pf_if),
    .io_req_bits_uop_xcpt_ae_if(ALUExeUnit_io_req_bits_uop_xcpt_ae_if),
    .io_req_bits_uop_replay_if(ALUExeUnit_io_req_bits_uop_replay_if),
    .io_req_bits_uop_xcpt_ma_if(ALUExeUnit_io_req_bits_uop_xcpt_ma_if),
    .io_req_bits_uop_debug_wdata(ALUExeUnit_io_req_bits_uop_debug_wdata),
    .io_req_bits_uop_debug_events_fetch_seq(ALUExeUnit_io_req_bits_uop_debug_events_fetch_seq),
    .io_req_bits_rs1_data(ALUExeUnit_io_req_bits_rs1_data),
    .io_req_bits_rs2_data(ALUExeUnit_io_req_bits_rs2_data),
    .io_req_bits_kill(ALUExeUnit_io_req_bits_kill),
    .io_resp_0_valid(ALUExeUnit_io_resp_0_valid),
    .io_resp_0_bits_uop_ctrl_rf_wen(ALUExeUnit_io_resp_0_bits_uop_ctrl_rf_wen),
    .io_resp_0_bits_uop_rob_idx(ALUExeUnit_io_resp_0_bits_uop_rob_idx),
    .io_resp_0_bits_uop_pdst(ALUExeUnit_io_resp_0_bits_uop_pdst),
    .io_resp_0_bits_uop_bypassable(ALUExeUnit_io_resp_0_bits_uop_bypassable),
    .io_resp_0_bits_uop_is_store(ALUExeUnit_io_resp_0_bits_uop_is_store),
    .io_resp_0_bits_uop_is_amo(ALUExeUnit_io_resp_0_bits_uop_is_amo),
    .io_resp_0_bits_uop_dst_rtype(ALUExeUnit_io_resp_0_bits_uop_dst_rtype),
    .io_resp_0_bits_data(ALUExeUnit_io_resp_0_bits_data),
    .io_bypass_valid_0(ALUExeUnit_io_bypass_valid_0),
    .io_bypass_uop_0_ctrl_rf_wen(ALUExeUnit_io_bypass_uop_0_ctrl_rf_wen),
    .io_bypass_uop_0_pdst(ALUExeUnit_io_bypass_uop_0_pdst),
    .io_bypass_uop_0_dst_rtype(ALUExeUnit_io_bypass_uop_0_dst_rtype),
    .io_bypass_data_0(ALUExeUnit_io_bypass_data_0),
    .io_brinfo_valid(ALUExeUnit_io_brinfo_valid),
    .io_brinfo_mispredict(ALUExeUnit_io_brinfo_mispredict),
    .io_brinfo_mask(ALUExeUnit_io_brinfo_mask)
  );
  FpPipeline fp_pipeline (
    .clock(fp_pipeline_clock),
    .reset(fp_pipeline_reset),
    .io_brinfo_valid(fp_pipeline_io_brinfo_valid),
    .io_brinfo_mispredict(fp_pipeline_io_brinfo_mispredict),
    .io_brinfo_mask(fp_pipeline_io_brinfo_mask),
    .io_flush_pipeline(fp_pipeline_io_flush_pipeline),
    .io_fcsr_rm(fp_pipeline_io_fcsr_rm),
    .io_dis_valids_0(fp_pipeline_io_dis_valids_0),
    .io_dis_valids_1(fp_pipeline_io_dis_valids_1),
    .io_dis_uops_0_valid(fp_pipeline_io_dis_uops_0_valid),
    .io_dis_uops_0_uopc(fp_pipeline_io_dis_uops_0_uopc),
    .io_dis_uops_0_inst(fp_pipeline_io_dis_uops_0_inst),
    .io_dis_uops_0_pc(fp_pipeline_io_dis_uops_0_pc),
    .io_dis_uops_0_iqtype(fp_pipeline_io_dis_uops_0_iqtype),
    .io_dis_uops_0_fu_code(fp_pipeline_io_dis_uops_0_fu_code),
    .io_dis_uops_0_allocate_brtag(fp_pipeline_io_dis_uops_0_allocate_brtag),
    .io_dis_uops_0_is_br_or_jmp(fp_pipeline_io_dis_uops_0_is_br_or_jmp),
    .io_dis_uops_0_is_jump(fp_pipeline_io_dis_uops_0_is_jump),
    .io_dis_uops_0_is_jal(fp_pipeline_io_dis_uops_0_is_jal),
    .io_dis_uops_0_is_ret(fp_pipeline_io_dis_uops_0_is_ret),
    .io_dis_uops_0_is_call(fp_pipeline_io_dis_uops_0_is_call),
    .io_dis_uops_0_br_mask(fp_pipeline_io_dis_uops_0_br_mask),
    .io_dis_uops_0_br_tag(fp_pipeline_io_dis_uops_0_br_tag),
    .io_dis_uops_0_br_prediction_btb_blame(fp_pipeline_io_dis_uops_0_br_prediction_btb_blame),
    .io_dis_uops_0_br_prediction_btb_hit(fp_pipeline_io_dis_uops_0_br_prediction_btb_hit),
    .io_dis_uops_0_br_prediction_btb_taken(fp_pipeline_io_dis_uops_0_br_prediction_btb_taken),
    .io_dis_uops_0_br_prediction_bpd_blame(fp_pipeline_io_dis_uops_0_br_prediction_bpd_blame),
    .io_dis_uops_0_br_prediction_bpd_hit(fp_pipeline_io_dis_uops_0_br_prediction_bpd_hit),
    .io_dis_uops_0_br_prediction_bpd_taken(fp_pipeline_io_dis_uops_0_br_prediction_bpd_taken),
    .io_dis_uops_0_br_prediction_bim_resp_value(fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_value),
    .io_dis_uops_0_br_prediction_bim_resp_entry_idx(fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_0_br_prediction_bim_resp_way_idx(fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_way_idx),
    .io_dis_uops_0_br_prediction_bpd_resp_takens(fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_takens),
    .io_dis_uops_0_br_prediction_bpd_resp_history(fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history),
    .io_dis_uops_0_br_prediction_bpd_resp_history_u(fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_u),
    .io_dis_uops_0_br_prediction_bpd_resp_history_ptr(fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_0_br_prediction_bpd_resp_info(fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_info),
    .io_dis_uops_0_stat_brjmp_mispredicted(fp_pipeline_io_dis_uops_0_stat_brjmp_mispredicted),
    .io_dis_uops_0_stat_btb_made_pred(fp_pipeline_io_dis_uops_0_stat_btb_made_pred),
    .io_dis_uops_0_stat_btb_mispredicted(fp_pipeline_io_dis_uops_0_stat_btb_mispredicted),
    .io_dis_uops_0_stat_bpd_made_pred(fp_pipeline_io_dis_uops_0_stat_bpd_made_pred),
    .io_dis_uops_0_stat_bpd_mispredicted(fp_pipeline_io_dis_uops_0_stat_bpd_mispredicted),
    .io_dis_uops_0_fetch_pc_lob(fp_pipeline_io_dis_uops_0_fetch_pc_lob),
    .io_dis_uops_0_imm_packed(fp_pipeline_io_dis_uops_0_imm_packed),
    .io_dis_uops_0_csr_addr(fp_pipeline_io_dis_uops_0_csr_addr),
    .io_dis_uops_0_rob_idx(fp_pipeline_io_dis_uops_0_rob_idx),
    .io_dis_uops_0_ldq_idx(fp_pipeline_io_dis_uops_0_ldq_idx),
    .io_dis_uops_0_stq_idx(fp_pipeline_io_dis_uops_0_stq_idx),
    .io_dis_uops_0_brob_idx(fp_pipeline_io_dis_uops_0_brob_idx),
    .io_dis_uops_0_pdst(fp_pipeline_io_dis_uops_0_pdst),
    .io_dis_uops_0_pop1(fp_pipeline_io_dis_uops_0_pop1),
    .io_dis_uops_0_pop2(fp_pipeline_io_dis_uops_0_pop2),
    .io_dis_uops_0_pop3(fp_pipeline_io_dis_uops_0_pop3),
    .io_dis_uops_0_prs1_busy(fp_pipeline_io_dis_uops_0_prs1_busy),
    .io_dis_uops_0_prs2_busy(fp_pipeline_io_dis_uops_0_prs2_busy),
    .io_dis_uops_0_prs3_busy(fp_pipeline_io_dis_uops_0_prs3_busy),
    .io_dis_uops_0_stale_pdst(fp_pipeline_io_dis_uops_0_stale_pdst),
    .io_dis_uops_0_exception(fp_pipeline_io_dis_uops_0_exception),
    .io_dis_uops_0_exc_cause(fp_pipeline_io_dis_uops_0_exc_cause),
    .io_dis_uops_0_bypassable(fp_pipeline_io_dis_uops_0_bypassable),
    .io_dis_uops_0_mem_cmd(fp_pipeline_io_dis_uops_0_mem_cmd),
    .io_dis_uops_0_mem_typ(fp_pipeline_io_dis_uops_0_mem_typ),
    .io_dis_uops_0_is_fence(fp_pipeline_io_dis_uops_0_is_fence),
    .io_dis_uops_0_is_fencei(fp_pipeline_io_dis_uops_0_is_fencei),
    .io_dis_uops_0_is_store(fp_pipeline_io_dis_uops_0_is_store),
    .io_dis_uops_0_is_amo(fp_pipeline_io_dis_uops_0_is_amo),
    .io_dis_uops_0_is_load(fp_pipeline_io_dis_uops_0_is_load),
    .io_dis_uops_0_is_sys_pc2epc(fp_pipeline_io_dis_uops_0_is_sys_pc2epc),
    .io_dis_uops_0_is_unique(fp_pipeline_io_dis_uops_0_is_unique),
    .io_dis_uops_0_flush_on_commit(fp_pipeline_io_dis_uops_0_flush_on_commit),
    .io_dis_uops_0_ldst(fp_pipeline_io_dis_uops_0_ldst),
    .io_dis_uops_0_lrs1(fp_pipeline_io_dis_uops_0_lrs1),
    .io_dis_uops_0_lrs2(fp_pipeline_io_dis_uops_0_lrs2),
    .io_dis_uops_0_lrs3(fp_pipeline_io_dis_uops_0_lrs3),
    .io_dis_uops_0_ldst_val(fp_pipeline_io_dis_uops_0_ldst_val),
    .io_dis_uops_0_dst_rtype(fp_pipeline_io_dis_uops_0_dst_rtype),
    .io_dis_uops_0_lrs1_rtype(fp_pipeline_io_dis_uops_0_lrs1_rtype),
    .io_dis_uops_0_lrs2_rtype(fp_pipeline_io_dis_uops_0_lrs2_rtype),
    .io_dis_uops_0_frs3_en(fp_pipeline_io_dis_uops_0_frs3_en),
    .io_dis_uops_0_fp_val(fp_pipeline_io_dis_uops_0_fp_val),
    .io_dis_uops_0_fp_single(fp_pipeline_io_dis_uops_0_fp_single),
    .io_dis_uops_0_xcpt_pf_if(fp_pipeline_io_dis_uops_0_xcpt_pf_if),
    .io_dis_uops_0_xcpt_ae_if(fp_pipeline_io_dis_uops_0_xcpt_ae_if),
    .io_dis_uops_0_replay_if(fp_pipeline_io_dis_uops_0_replay_if),
    .io_dis_uops_0_xcpt_ma_if(fp_pipeline_io_dis_uops_0_xcpt_ma_if),
    .io_dis_uops_0_debug_wdata(fp_pipeline_io_dis_uops_0_debug_wdata),
    .io_dis_uops_0_debug_events_fetch_seq(fp_pipeline_io_dis_uops_0_debug_events_fetch_seq),
    .io_dis_uops_1_valid(fp_pipeline_io_dis_uops_1_valid),
    .io_dis_uops_1_uopc(fp_pipeline_io_dis_uops_1_uopc),
    .io_dis_uops_1_inst(fp_pipeline_io_dis_uops_1_inst),
    .io_dis_uops_1_pc(fp_pipeline_io_dis_uops_1_pc),
    .io_dis_uops_1_iqtype(fp_pipeline_io_dis_uops_1_iqtype),
    .io_dis_uops_1_fu_code(fp_pipeline_io_dis_uops_1_fu_code),
    .io_dis_uops_1_allocate_brtag(fp_pipeline_io_dis_uops_1_allocate_brtag),
    .io_dis_uops_1_is_br_or_jmp(fp_pipeline_io_dis_uops_1_is_br_or_jmp),
    .io_dis_uops_1_is_jump(fp_pipeline_io_dis_uops_1_is_jump),
    .io_dis_uops_1_is_jal(fp_pipeline_io_dis_uops_1_is_jal),
    .io_dis_uops_1_is_ret(fp_pipeline_io_dis_uops_1_is_ret),
    .io_dis_uops_1_is_call(fp_pipeline_io_dis_uops_1_is_call),
    .io_dis_uops_1_br_mask(fp_pipeline_io_dis_uops_1_br_mask),
    .io_dis_uops_1_br_tag(fp_pipeline_io_dis_uops_1_br_tag),
    .io_dis_uops_1_br_prediction_btb_blame(fp_pipeline_io_dis_uops_1_br_prediction_btb_blame),
    .io_dis_uops_1_br_prediction_btb_hit(fp_pipeline_io_dis_uops_1_br_prediction_btb_hit),
    .io_dis_uops_1_br_prediction_btb_taken(fp_pipeline_io_dis_uops_1_br_prediction_btb_taken),
    .io_dis_uops_1_br_prediction_bpd_blame(fp_pipeline_io_dis_uops_1_br_prediction_bpd_blame),
    .io_dis_uops_1_br_prediction_bpd_hit(fp_pipeline_io_dis_uops_1_br_prediction_bpd_hit),
    .io_dis_uops_1_br_prediction_bpd_taken(fp_pipeline_io_dis_uops_1_br_prediction_bpd_taken),
    .io_dis_uops_1_br_prediction_bim_resp_value(fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_value),
    .io_dis_uops_1_br_prediction_bim_resp_entry_idx(fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_1_br_prediction_bim_resp_way_idx(fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_way_idx),
    .io_dis_uops_1_br_prediction_bpd_resp_takens(fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_takens),
    .io_dis_uops_1_br_prediction_bpd_resp_history(fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history),
    .io_dis_uops_1_br_prediction_bpd_resp_history_u(fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_u),
    .io_dis_uops_1_br_prediction_bpd_resp_history_ptr(fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_1_br_prediction_bpd_resp_info(fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_info),
    .io_dis_uops_1_stat_brjmp_mispredicted(fp_pipeline_io_dis_uops_1_stat_brjmp_mispredicted),
    .io_dis_uops_1_stat_btb_made_pred(fp_pipeline_io_dis_uops_1_stat_btb_made_pred),
    .io_dis_uops_1_stat_btb_mispredicted(fp_pipeline_io_dis_uops_1_stat_btb_mispredicted),
    .io_dis_uops_1_stat_bpd_made_pred(fp_pipeline_io_dis_uops_1_stat_bpd_made_pred),
    .io_dis_uops_1_stat_bpd_mispredicted(fp_pipeline_io_dis_uops_1_stat_bpd_mispredicted),
    .io_dis_uops_1_fetch_pc_lob(fp_pipeline_io_dis_uops_1_fetch_pc_lob),
    .io_dis_uops_1_imm_packed(fp_pipeline_io_dis_uops_1_imm_packed),
    .io_dis_uops_1_csr_addr(fp_pipeline_io_dis_uops_1_csr_addr),
    .io_dis_uops_1_rob_idx(fp_pipeline_io_dis_uops_1_rob_idx),
    .io_dis_uops_1_ldq_idx(fp_pipeline_io_dis_uops_1_ldq_idx),
    .io_dis_uops_1_stq_idx(fp_pipeline_io_dis_uops_1_stq_idx),
    .io_dis_uops_1_brob_idx(fp_pipeline_io_dis_uops_1_brob_idx),
    .io_dis_uops_1_pdst(fp_pipeline_io_dis_uops_1_pdst),
    .io_dis_uops_1_pop1(fp_pipeline_io_dis_uops_1_pop1),
    .io_dis_uops_1_pop2(fp_pipeline_io_dis_uops_1_pop2),
    .io_dis_uops_1_pop3(fp_pipeline_io_dis_uops_1_pop3),
    .io_dis_uops_1_prs1_busy(fp_pipeline_io_dis_uops_1_prs1_busy),
    .io_dis_uops_1_prs2_busy(fp_pipeline_io_dis_uops_1_prs2_busy),
    .io_dis_uops_1_prs3_busy(fp_pipeline_io_dis_uops_1_prs3_busy),
    .io_dis_uops_1_stale_pdst(fp_pipeline_io_dis_uops_1_stale_pdst),
    .io_dis_uops_1_exception(fp_pipeline_io_dis_uops_1_exception),
    .io_dis_uops_1_exc_cause(fp_pipeline_io_dis_uops_1_exc_cause),
    .io_dis_uops_1_bypassable(fp_pipeline_io_dis_uops_1_bypassable),
    .io_dis_uops_1_mem_cmd(fp_pipeline_io_dis_uops_1_mem_cmd),
    .io_dis_uops_1_mem_typ(fp_pipeline_io_dis_uops_1_mem_typ),
    .io_dis_uops_1_is_fence(fp_pipeline_io_dis_uops_1_is_fence),
    .io_dis_uops_1_is_fencei(fp_pipeline_io_dis_uops_1_is_fencei),
    .io_dis_uops_1_is_store(fp_pipeline_io_dis_uops_1_is_store),
    .io_dis_uops_1_is_amo(fp_pipeline_io_dis_uops_1_is_amo),
    .io_dis_uops_1_is_load(fp_pipeline_io_dis_uops_1_is_load),
    .io_dis_uops_1_is_sys_pc2epc(fp_pipeline_io_dis_uops_1_is_sys_pc2epc),
    .io_dis_uops_1_is_unique(fp_pipeline_io_dis_uops_1_is_unique),
    .io_dis_uops_1_flush_on_commit(fp_pipeline_io_dis_uops_1_flush_on_commit),
    .io_dis_uops_1_ldst(fp_pipeline_io_dis_uops_1_ldst),
    .io_dis_uops_1_lrs1(fp_pipeline_io_dis_uops_1_lrs1),
    .io_dis_uops_1_lrs2(fp_pipeline_io_dis_uops_1_lrs2),
    .io_dis_uops_1_lrs3(fp_pipeline_io_dis_uops_1_lrs3),
    .io_dis_uops_1_ldst_val(fp_pipeline_io_dis_uops_1_ldst_val),
    .io_dis_uops_1_dst_rtype(fp_pipeline_io_dis_uops_1_dst_rtype),
    .io_dis_uops_1_lrs1_rtype(fp_pipeline_io_dis_uops_1_lrs1_rtype),
    .io_dis_uops_1_lrs2_rtype(fp_pipeline_io_dis_uops_1_lrs2_rtype),
    .io_dis_uops_1_frs3_en(fp_pipeline_io_dis_uops_1_frs3_en),
    .io_dis_uops_1_fp_val(fp_pipeline_io_dis_uops_1_fp_val),
    .io_dis_uops_1_fp_single(fp_pipeline_io_dis_uops_1_fp_single),
    .io_dis_uops_1_xcpt_pf_if(fp_pipeline_io_dis_uops_1_xcpt_pf_if),
    .io_dis_uops_1_xcpt_ae_if(fp_pipeline_io_dis_uops_1_xcpt_ae_if),
    .io_dis_uops_1_replay_if(fp_pipeline_io_dis_uops_1_replay_if),
    .io_dis_uops_1_xcpt_ma_if(fp_pipeline_io_dis_uops_1_xcpt_ma_if),
    .io_dis_uops_1_debug_wdata(fp_pipeline_io_dis_uops_1_debug_wdata),
    .io_dis_uops_1_debug_events_fetch_seq(fp_pipeline_io_dis_uops_1_debug_events_fetch_seq),
    .io_dis_readys_0(fp_pipeline_io_dis_readys_0),
    .io_dis_readys_1(fp_pipeline_io_dis_readys_1),
    .io_ll_wport_valid(fp_pipeline_io_ll_wport_valid),
    .io_ll_wport_bits_uop_rob_idx(fp_pipeline_io_ll_wport_bits_uop_rob_idx),
    .io_ll_wport_bits_uop_pdst(fp_pipeline_io_ll_wport_bits_uop_pdst),
    .io_ll_wport_bits_uop_mem_typ(fp_pipeline_io_ll_wport_bits_uop_mem_typ),
    .io_ll_wport_bits_uop_dst_rtype(fp_pipeline_io_ll_wport_bits_uop_dst_rtype),
    .io_ll_wport_bits_uop_fp_val(fp_pipeline_io_ll_wport_bits_uop_fp_val),
    .io_ll_wport_bits_data(fp_pipeline_io_ll_wport_bits_data),
    .io_fromint_valid(fp_pipeline_io_fromint_valid),
    .io_fromint_bits_uop_uopc(fp_pipeline_io_fromint_bits_uop_uopc),
    .io_fromint_bits_uop_ctrl_rf_wen(fp_pipeline_io_fromint_bits_uop_ctrl_rf_wen),
    .io_fromint_bits_uop_br_mask(fp_pipeline_io_fromint_bits_uop_br_mask),
    .io_fromint_bits_uop_imm_packed(fp_pipeline_io_fromint_bits_uop_imm_packed),
    .io_fromint_bits_uop_rob_idx(fp_pipeline_io_fromint_bits_uop_rob_idx),
    .io_fromint_bits_uop_pdst(fp_pipeline_io_fromint_bits_uop_pdst),
    .io_fromint_bits_uop_dst_rtype(fp_pipeline_io_fromint_bits_uop_dst_rtype),
    .io_fromint_bits_uop_fp_val(fp_pipeline_io_fromint_bits_uop_fp_val),
    .io_fromint_bits_rs1_data(fp_pipeline_io_fromint_bits_rs1_data),
    .io_tosdq_valid(fp_pipeline_io_tosdq_valid),
    .io_tosdq_bits_uop_br_mask(fp_pipeline_io_tosdq_bits_uop_br_mask),
    .io_tosdq_bits_uop_rob_idx(fp_pipeline_io_tosdq_bits_uop_rob_idx),
    .io_tosdq_bits_uop_stq_idx(fp_pipeline_io_tosdq_bits_uop_stq_idx),
    .io_tosdq_bits_uop_is_amo(fp_pipeline_io_tosdq_bits_uop_is_amo),
    .io_tosdq_bits_data(fp_pipeline_io_tosdq_bits_data),
    .io_toint_ready(fp_pipeline_io_toint_ready),
    .io_toint_valid(fp_pipeline_io_toint_valid),
    .io_toint_bits_uop_rob_idx(fp_pipeline_io_toint_bits_uop_rob_idx),
    .io_toint_bits_uop_pdst(fp_pipeline_io_toint_bits_uop_pdst),
    .io_toint_bits_uop_is_store(fp_pipeline_io_toint_bits_uop_is_store),
    .io_toint_bits_uop_is_amo(fp_pipeline_io_toint_bits_uop_is_amo),
    .io_toint_bits_uop_dst_rtype(fp_pipeline_io_toint_bits_uop_dst_rtype),
    .io_toint_bits_data(fp_pipeline_io_toint_bits_data),
    .io_wakeups_0_valid(fp_pipeline_io_wakeups_0_valid),
    .io_wakeups_0_bits_uop_rob_idx(fp_pipeline_io_wakeups_0_bits_uop_rob_idx),
    .io_wakeups_0_bits_uop_pdst(fp_pipeline_io_wakeups_0_bits_uop_pdst),
    .io_wakeups_0_bits_uop_dst_rtype(fp_pipeline_io_wakeups_0_bits_uop_dst_rtype),
    .io_wakeups_0_bits_uop_fp_val(fp_pipeline_io_wakeups_0_bits_uop_fp_val),
    .io_wakeups_0_bits_fflags_valid(fp_pipeline_io_wakeups_0_bits_fflags_valid),
    .io_wakeups_0_bits_fflags_bits_uop_rob_idx(fp_pipeline_io_wakeups_0_bits_fflags_bits_uop_rob_idx),
    .io_wakeups_0_bits_fflags_bits_flags(fp_pipeline_io_wakeups_0_bits_fflags_bits_flags),
    .io_wakeups_1_valid(fp_pipeline_io_wakeups_1_valid),
    .io_wakeups_1_bits_uop_rob_idx(fp_pipeline_io_wakeups_1_bits_uop_rob_idx),
    .io_wakeups_1_bits_uop_pdst(fp_pipeline_io_wakeups_1_bits_uop_pdst),
    .io_wakeups_1_bits_uop_dst_rtype(fp_pipeline_io_wakeups_1_bits_uop_dst_rtype),
    .io_wakeups_1_bits_uop_fp_val(fp_pipeline_io_wakeups_1_bits_uop_fp_val),
    .io_wakeups_1_bits_fflags_valid(fp_pipeline_io_wakeups_1_bits_fflags_valid),
    .io_wakeups_1_bits_fflags_bits_uop_rob_idx(fp_pipeline_io_wakeups_1_bits_fflags_bits_uop_rob_idx),
    .io_wakeups_1_bits_fflags_bits_flags(fp_pipeline_io_wakeups_1_bits_fflags_bits_flags)
  );
  FetchUnit fetch_unit (
    .clock(fetch_unit_clock),
    .reset(fetch_unit_reset),
    .io_imem_req_valid(fetch_unit_io_imem_req_valid),
    .io_imem_req_bits_pc(fetch_unit_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(fetch_unit_io_imem_req_bits_speculative),
    .io_imem_resp_ready(fetch_unit_io_imem_resp_ready),
    .io_imem_resp_valid(fetch_unit_io_imem_resp_valid),
    .io_imem_resp_bits_pc(fetch_unit_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(fetch_unit_io_imem_resp_bits_data),
    .io_imem_resp_bits_mask(fetch_unit_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_pf_inst(fetch_unit_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(fetch_unit_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(fetch_unit_io_imem_resp_bits_replay),
    .io_f2_btb_resp_bits_bim_resp_value(fetch_unit_io_f2_btb_resp_bits_bim_resp_value),
    .io_f2_btb_resp_bits_bim_resp_entry_idx(fetch_unit_io_f2_btb_resp_bits_bim_resp_entry_idx),
    .io_f2_btb_resp_bits_bim_resp_way_idx(fetch_unit_io_f2_btb_resp_bits_bim_resp_way_idx),
    .io_f2_bpd_resp_bits_takens(fetch_unit_io_f2_bpd_resp_bits_takens),
    .io_f2_bpd_resp_bits_info(fetch_unit_io_f2_bpd_resp_bits_info),
    .io_f3_bpd_resp_bits_history(fetch_unit_io_f3_bpd_resp_bits_history),
    .io_f3_bpd_resp_bits_history_ptr(fetch_unit_io_f3_bpd_resp_bits_history_ptr),
    .io_f3_btb_update_valid(fetch_unit_io_f3_btb_update_valid),
    .io_f3_btb_update_bits_pc(fetch_unit_io_f3_btb_update_bits_pc),
    .io_f3_btb_update_bits_target(fetch_unit_io_f3_btb_update_bits_target),
    .io_f3_btb_update_bits_cfi_pc(fetch_unit_io_f3_btb_update_bits_cfi_pc),
    .io_f3_btb_update_bits_bpd_type(fetch_unit_io_f3_btb_update_bits_bpd_type),
    .io_f3_btb_update_bits_cfi_type(fetch_unit_io_f3_btb_update_bits_cfi_type),
    .io_f3_hist_update_valid(fetch_unit_io_f3_hist_update_valid),
    .io_f3_hist_update_bits_taken(fetch_unit_io_f3_hist_update_bits_taken),
    .io_f3_bim_update_valid(fetch_unit_io_f3_bim_update_valid),
    .io_f3_bim_update_bits_taken(fetch_unit_io_f3_bim_update_bits_taken),
    .io_f3_bim_update_bits_bim_resp_value(fetch_unit_io_f3_bim_update_bits_bim_resp_value),
    .io_f3_bim_update_bits_bim_resp_entry_idx(fetch_unit_io_f3_bim_update_bits_bim_resp_entry_idx),
    .io_f3_bim_update_bits_bim_resp_way_idx(fetch_unit_io_f3_bim_update_bits_bim_resp_way_idx),
    .io_br_unit_take_pc(fetch_unit_io_br_unit_take_pc),
    .io_br_unit_target(fetch_unit_io_br_unit_target),
    .io_clear_fetchbuffer(fetch_unit_io_clear_fetchbuffer),
    .io_flush_take_pc(fetch_unit_io_flush_take_pc),
    .io_flush_pc(fetch_unit_io_flush_pc),
    .io_sfence_take_pc(fetch_unit_io_sfence_take_pc),
    .io_sfence_addr(fetch_unit_io_sfence_addr),
    .io_resp_ready(fetch_unit_io_resp_ready),
    .io_resp_valid(fetch_unit_io_resp_valid),
    .io_resp_bits_pc(fetch_unit_io_resp_bits_pc),
    .io_resp_bits_insts_0(fetch_unit_io_resp_bits_insts_0),
    .io_resp_bits_insts_1(fetch_unit_io_resp_bits_insts_1),
    .io_resp_bits_mask(fetch_unit_io_resp_bits_mask),
    .io_resp_bits_xcpt_pf_if(fetch_unit_io_resp_bits_xcpt_pf_if),
    .io_resp_bits_xcpt_ae_if(fetch_unit_io_resp_bits_xcpt_ae_if),
    .io_resp_bits_replay_if(fetch_unit_io_resp_bits_replay_if),
    .io_resp_bits_xcpt_ma_if_oh(fetch_unit_io_resp_bits_xcpt_ma_if_oh),
    .io_resp_bits_bpu_info_0_btb_blame(fetch_unit_io_resp_bits_bpu_info_0_btb_blame),
    .io_resp_bits_bpu_info_0_btb_hit(fetch_unit_io_resp_bits_bpu_info_0_btb_hit),
    .io_resp_bits_bpu_info_0_btb_taken(fetch_unit_io_resp_bits_bpu_info_0_btb_taken),
    .io_resp_bits_bpu_info_0_bpd_blame(fetch_unit_io_resp_bits_bpu_info_0_bpd_blame),
    .io_resp_bits_bpu_info_0_bpd_hit(fetch_unit_io_resp_bits_bpu_info_0_bpd_hit),
    .io_resp_bits_bpu_info_0_bpd_taken(fetch_unit_io_resp_bits_bpu_info_0_bpd_taken),
    .io_resp_bits_bpu_info_0_bim_resp_value(fetch_unit_io_resp_bits_bpu_info_0_bim_resp_value),
    .io_resp_bits_bpu_info_0_bim_resp_entry_idx(fetch_unit_io_resp_bits_bpu_info_0_bim_resp_entry_idx),
    .io_resp_bits_bpu_info_0_bim_resp_way_idx(fetch_unit_io_resp_bits_bpu_info_0_bim_resp_way_idx),
    .io_resp_bits_bpu_info_0_bpd_resp_takens(fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_takens),
    .io_resp_bits_bpu_info_0_bpd_resp_history(fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history),
    .io_resp_bits_bpu_info_0_bpd_resp_history_u(fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_u),
    .io_resp_bits_bpu_info_0_bpd_resp_history_ptr(fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_ptr),
    .io_resp_bits_bpu_info_0_bpd_resp_info(fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_info),
    .io_resp_bits_bpu_info_1_btb_blame(fetch_unit_io_resp_bits_bpu_info_1_btb_blame),
    .io_resp_bits_bpu_info_1_btb_hit(fetch_unit_io_resp_bits_bpu_info_1_btb_hit),
    .io_resp_bits_bpu_info_1_btb_taken(fetch_unit_io_resp_bits_bpu_info_1_btb_taken),
    .io_resp_bits_bpu_info_1_bpd_blame(fetch_unit_io_resp_bits_bpu_info_1_bpd_blame),
    .io_resp_bits_bpu_info_1_bpd_hit(fetch_unit_io_resp_bits_bpu_info_1_bpd_hit),
    .io_resp_bits_bpu_info_1_bpd_taken(fetch_unit_io_resp_bits_bpu_info_1_bpd_taken),
    .io_resp_bits_bpu_info_1_bim_resp_value(fetch_unit_io_resp_bits_bpu_info_1_bim_resp_value),
    .io_resp_bits_bpu_info_1_bim_resp_entry_idx(fetch_unit_io_resp_bits_bpu_info_1_bim_resp_entry_idx),
    .io_resp_bits_bpu_info_1_bim_resp_way_idx(fetch_unit_io_resp_bits_bpu_info_1_bim_resp_way_idx),
    .io_resp_bits_bpu_info_1_bpd_resp_takens(fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_takens),
    .io_resp_bits_bpu_info_1_bpd_resp_history(fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history),
    .io_resp_bits_bpu_info_1_bpd_resp_history_u(fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_u),
    .io_resp_bits_bpu_info_1_bpd_resp_history_ptr(fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_ptr),
    .io_resp_bits_bpu_info_1_bpd_resp_info(fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_info),
    .io_resp_bits_debug_events_0_fetch_seq(fetch_unit_io_resp_bits_debug_events_0_fetch_seq),
    .io_resp_bits_debug_events_1_fetch_seq(fetch_unit_io_resp_bits_debug_events_1_fetch_seq),
    .io_stalled(fetch_unit_io_stalled)
  );
  BranchPredictionStage bpd_stage (
    .clock(bpd_stage_clock),
    .reset(bpd_stage_reset),
    .io_fetch_stalled(bpd_stage_io_fetch_stalled),
    .io_f2_btb_resp_bits_bim_resp_value(bpd_stage_io_f2_btb_resp_bits_bim_resp_value),
    .io_f2_btb_resp_bits_bim_resp_entry_idx(bpd_stage_io_f2_btb_resp_bits_bim_resp_entry_idx),
    .io_f2_btb_resp_bits_bim_resp_way_idx(bpd_stage_io_f2_btb_resp_bits_bim_resp_way_idx),
    .io_f2_bpd_resp_bits_takens(bpd_stage_io_f2_bpd_resp_bits_takens),
    .io_f2_bpd_resp_bits_info(bpd_stage_io_f2_bpd_resp_bits_info),
    .io_f3_bpd_resp_bits_history(bpd_stage_io_f3_bpd_resp_bits_history),
    .io_f3_bpd_resp_bits_history_ptr(bpd_stage_io_f3_bpd_resp_bits_history_ptr),
    .io_f3_btb_update_valid(bpd_stage_io_f3_btb_update_valid),
    .io_f3_btb_update_bits_pc(bpd_stage_io_f3_btb_update_bits_pc),
    .io_f3_btb_update_bits_target(bpd_stage_io_f3_btb_update_bits_target),
    .io_f3_btb_update_bits_cfi_pc(bpd_stage_io_f3_btb_update_bits_cfi_pc),
    .io_f3_btb_update_bits_bpd_type(bpd_stage_io_f3_btb_update_bits_bpd_type),
    .io_f3_btb_update_bits_cfi_type(bpd_stage_io_f3_btb_update_bits_cfi_type),
    .io_f3_hist_update_valid(bpd_stage_io_f3_hist_update_valid),
    .io_f3_hist_update_bits_taken(bpd_stage_io_f3_hist_update_bits_taken),
    .io_f3_bim_update_valid(bpd_stage_io_f3_bim_update_valid),
    .io_f3_bim_update_bits_taken(bpd_stage_io_f3_bim_update_bits_taken),
    .io_f3_bim_update_bits_bim_resp_value(bpd_stage_io_f3_bim_update_bits_bim_resp_value),
    .io_f3_bim_update_bits_bim_resp_entry_idx(bpd_stage_io_f3_bim_update_bits_bim_resp_entry_idx),
    .io_f3_bim_update_bits_bim_resp_way_idx(bpd_stage_io_f3_bim_update_bits_bim_resp_way_idx),
    .io_br_unit_btb_update_valid(bpd_stage_io_br_unit_btb_update_valid),
    .io_br_unit_btb_update_bits_pc(bpd_stage_io_br_unit_btb_update_bits_pc),
    .io_br_unit_btb_update_bits_target(bpd_stage_io_br_unit_btb_update_bits_target),
    .io_br_unit_btb_update_bits_cfi_pc(bpd_stage_io_br_unit_btb_update_bits_cfi_pc),
    .io_br_unit_btb_update_bits_bpd_type(bpd_stage_io_br_unit_btb_update_bits_bpd_type),
    .io_br_unit_btb_update_bits_cfi_type(bpd_stage_io_br_unit_btb_update_bits_cfi_type),
    .io_br_unit_bim_update_valid(bpd_stage_io_br_unit_bim_update_valid),
    .io_br_unit_bim_update_bits_taken(bpd_stage_io_br_unit_bim_update_bits_taken),
    .io_br_unit_bim_update_bits_bim_resp_value(bpd_stage_io_br_unit_bim_update_bits_bim_resp_value),
    .io_br_unit_bim_update_bits_bim_resp_entry_idx(bpd_stage_io_br_unit_bim_update_bits_bim_resp_entry_idx),
    .io_br_unit_bim_update_bits_bim_resp_way_idx(bpd_stage_io_br_unit_bim_update_bits_bim_resp_way_idx),
    .io_br_unit_bpd_update_valid(bpd_stage_io_br_unit_bpd_update_valid),
    .io_br_unit_bpd_update_bits_mispredict(bpd_stage_io_br_unit_bpd_update_bits_mispredict),
    .io_br_unit_bpd_update_bits_history(bpd_stage_io_br_unit_bpd_update_bits_history),
    .io_br_unit_bpd_update_bits_history_ptr(bpd_stage_io_br_unit_bpd_update_bits_history_ptr),
    .io_br_unit_bpd_update_bits_bpd_mispredict(bpd_stage_io_br_unit_bpd_update_bits_bpd_mispredict),
    .io_br_unit_bpd_update_bits_taken(bpd_stage_io_br_unit_bpd_update_bits_taken),
    .io_br_unit_bpd_update_bits_new_pc_same_packet(bpd_stage_io_br_unit_bpd_update_bits_new_pc_same_packet),
    .io_brob_allocate_ready(bpd_stage_io_brob_allocate_ready),
    .io_brob_allocate_valid(bpd_stage_io_brob_allocate_valid),
    .io_brob_allocate_bits_ctrl_brob_idx(bpd_stage_io_brob_allocate_bits_ctrl_brob_idx),
    .io_brob_allocate_bits_info_info(bpd_stage_io_brob_allocate_bits_info_info),
    .io_brob_allocate_brob_tail(bpd_stage_io_brob_allocate_brob_tail),
    .io_brob_deallocate_valid(bpd_stage_io_brob_deallocate_valid),
    .io_brob_deallocate_bits_brob_idx(bpd_stage_io_brob_deallocate_bits_brob_idx),
    .io_brob_bpd_update_valid(bpd_stage_io_brob_bpd_update_valid),
    .io_brob_bpd_update_bits_br_pc(bpd_stage_io_brob_bpd_update_bits_br_pc),
    .io_brob_bpd_update_bits_brob_idx(bpd_stage_io_brob_bpd_update_bits_brob_idx),
    .io_brob_bpd_update_bits_mispredict(bpd_stage_io_brob_bpd_update_bits_mispredict),
    .io_brob_bpd_update_bits_bpd_predict_val(bpd_stage_io_brob_bpd_update_bits_bpd_predict_val),
    .io_brob_bpd_update_bits_bpd_mispredict(bpd_stage_io_brob_bpd_update_bits_bpd_mispredict),
    .io_brob_bpd_update_bits_taken(bpd_stage_io_brob_bpd_update_bits_taken),
    .io_brob_bpd_update_bits_is_br(bpd_stage_io_brob_bpd_update_bits_is_br),
    .io_brob_flush(bpd_stage_io_brob_flush),
    .io_flush(bpd_stage_io_flush),
    .io_redirect(bpd_stage_io_redirect),
    .io_status_debug(bpd_stage_io_status_debug)
  );
  FetchSerializerNtoM dec_serializer (
    .io_enq_ready(dec_serializer_io_enq_ready),
    .io_enq_valid(dec_serializer_io_enq_valid),
    .io_enq_bits_pc(dec_serializer_io_enq_bits_pc),
    .io_enq_bits_insts_0(dec_serializer_io_enq_bits_insts_0),
    .io_enq_bits_insts_1(dec_serializer_io_enq_bits_insts_1),
    .io_enq_bits_mask(dec_serializer_io_enq_bits_mask),
    .io_enq_bits_xcpt_pf_if(dec_serializer_io_enq_bits_xcpt_pf_if),
    .io_enq_bits_xcpt_ae_if(dec_serializer_io_enq_bits_xcpt_ae_if),
    .io_enq_bits_replay_if(dec_serializer_io_enq_bits_replay_if),
    .io_enq_bits_xcpt_ma_if_oh(dec_serializer_io_enq_bits_xcpt_ma_if_oh),
    .io_enq_bits_bpu_info_0_btb_blame(dec_serializer_io_enq_bits_bpu_info_0_btb_blame),
    .io_enq_bits_bpu_info_0_btb_hit(dec_serializer_io_enq_bits_bpu_info_0_btb_hit),
    .io_enq_bits_bpu_info_0_btb_taken(dec_serializer_io_enq_bits_bpu_info_0_btb_taken),
    .io_enq_bits_bpu_info_0_bpd_blame(dec_serializer_io_enq_bits_bpu_info_0_bpd_blame),
    .io_enq_bits_bpu_info_0_bpd_hit(dec_serializer_io_enq_bits_bpu_info_0_bpd_hit),
    .io_enq_bits_bpu_info_0_bpd_taken(dec_serializer_io_enq_bits_bpu_info_0_bpd_taken),
    .io_enq_bits_bpu_info_0_bim_resp_value(dec_serializer_io_enq_bits_bpu_info_0_bim_resp_value),
    .io_enq_bits_bpu_info_0_bim_resp_entry_idx(dec_serializer_io_enq_bits_bpu_info_0_bim_resp_entry_idx),
    .io_enq_bits_bpu_info_0_bim_resp_way_idx(dec_serializer_io_enq_bits_bpu_info_0_bim_resp_way_idx),
    .io_enq_bits_bpu_info_0_bpd_resp_takens(dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_takens),
    .io_enq_bits_bpu_info_0_bpd_resp_history(dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history),
    .io_enq_bits_bpu_info_0_bpd_resp_history_u(dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_u),
    .io_enq_bits_bpu_info_0_bpd_resp_history_ptr(dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_ptr),
    .io_enq_bits_bpu_info_0_bpd_resp_info(dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_info),
    .io_enq_bits_bpu_info_1_btb_blame(dec_serializer_io_enq_bits_bpu_info_1_btb_blame),
    .io_enq_bits_bpu_info_1_btb_hit(dec_serializer_io_enq_bits_bpu_info_1_btb_hit),
    .io_enq_bits_bpu_info_1_btb_taken(dec_serializer_io_enq_bits_bpu_info_1_btb_taken),
    .io_enq_bits_bpu_info_1_bpd_blame(dec_serializer_io_enq_bits_bpu_info_1_bpd_blame),
    .io_enq_bits_bpu_info_1_bpd_hit(dec_serializer_io_enq_bits_bpu_info_1_bpd_hit),
    .io_enq_bits_bpu_info_1_bpd_taken(dec_serializer_io_enq_bits_bpu_info_1_bpd_taken),
    .io_enq_bits_bpu_info_1_bim_resp_value(dec_serializer_io_enq_bits_bpu_info_1_bim_resp_value),
    .io_enq_bits_bpu_info_1_bim_resp_entry_idx(dec_serializer_io_enq_bits_bpu_info_1_bim_resp_entry_idx),
    .io_enq_bits_bpu_info_1_bim_resp_way_idx(dec_serializer_io_enq_bits_bpu_info_1_bim_resp_way_idx),
    .io_enq_bits_bpu_info_1_bpd_resp_takens(dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_takens),
    .io_enq_bits_bpu_info_1_bpd_resp_history(dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history),
    .io_enq_bits_bpu_info_1_bpd_resp_history_u(dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_u),
    .io_enq_bits_bpu_info_1_bpd_resp_history_ptr(dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_ptr),
    .io_enq_bits_bpu_info_1_bpd_resp_info(dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_info),
    .io_enq_bits_debug_events_0_fetch_seq(dec_serializer_io_enq_bits_debug_events_0_fetch_seq),
    .io_enq_bits_debug_events_1_fetch_seq(dec_serializer_io_enq_bits_debug_events_1_fetch_seq),
    .io_deq_ready(dec_serializer_io_deq_ready),
    .io_deq_valid(dec_serializer_io_deq_valid),
    .io_deq_bits_uops_0_valid(dec_serializer_io_deq_bits_uops_0_valid),
    .io_deq_bits_uops_0_inst(dec_serializer_io_deq_bits_uops_0_inst),
    .io_deq_bits_uops_0_pc(dec_serializer_io_deq_bits_uops_0_pc),
    .io_deq_bits_uops_0_br_prediction_btb_blame(dec_serializer_io_deq_bits_uops_0_br_prediction_btb_blame),
    .io_deq_bits_uops_0_br_prediction_btb_hit(dec_serializer_io_deq_bits_uops_0_br_prediction_btb_hit),
    .io_deq_bits_uops_0_br_prediction_btb_taken(dec_serializer_io_deq_bits_uops_0_br_prediction_btb_taken),
    .io_deq_bits_uops_0_br_prediction_bpd_blame(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_blame),
    .io_deq_bits_uops_0_br_prediction_bpd_hit(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_hit),
    .io_deq_bits_uops_0_br_prediction_bpd_taken(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_taken),
    .io_deq_bits_uops_0_br_prediction_bim_resp_value(dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_value),
    .io_deq_bits_uops_0_br_prediction_bim_resp_entry_idx(dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_entry_idx),
    .io_deq_bits_uops_0_br_prediction_bim_resp_way_idx(dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_way_idx),
    .io_deq_bits_uops_0_br_prediction_bpd_resp_takens(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_takens),
    .io_deq_bits_uops_0_br_prediction_bpd_resp_history(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history),
    .io_deq_bits_uops_0_br_prediction_bpd_resp_history_u(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_u),
    .io_deq_bits_uops_0_br_prediction_bpd_resp_history_ptr(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_deq_bits_uops_0_br_prediction_bpd_resp_info(dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_info),
    .io_deq_bits_uops_0_fetch_pc_lob(dec_serializer_io_deq_bits_uops_0_fetch_pc_lob),
    .io_deq_bits_uops_0_xcpt_pf_if(dec_serializer_io_deq_bits_uops_0_xcpt_pf_if),
    .io_deq_bits_uops_0_xcpt_ae_if(dec_serializer_io_deq_bits_uops_0_xcpt_ae_if),
    .io_deq_bits_uops_0_replay_if(dec_serializer_io_deq_bits_uops_0_replay_if),
    .io_deq_bits_uops_0_xcpt_ma_if(dec_serializer_io_deq_bits_uops_0_xcpt_ma_if),
    .io_deq_bits_uops_0_debug_events_fetch_seq(dec_serializer_io_deq_bits_uops_0_debug_events_fetch_seq),
    .io_deq_bits_uops_1_valid(dec_serializer_io_deq_bits_uops_1_valid),
    .io_deq_bits_uops_1_inst(dec_serializer_io_deq_bits_uops_1_inst),
    .io_deq_bits_uops_1_pc(dec_serializer_io_deq_bits_uops_1_pc),
    .io_deq_bits_uops_1_br_prediction_btb_blame(dec_serializer_io_deq_bits_uops_1_br_prediction_btb_blame),
    .io_deq_bits_uops_1_br_prediction_btb_hit(dec_serializer_io_deq_bits_uops_1_br_prediction_btb_hit),
    .io_deq_bits_uops_1_br_prediction_btb_taken(dec_serializer_io_deq_bits_uops_1_br_prediction_btb_taken),
    .io_deq_bits_uops_1_br_prediction_bpd_blame(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_blame),
    .io_deq_bits_uops_1_br_prediction_bpd_hit(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_hit),
    .io_deq_bits_uops_1_br_prediction_bpd_taken(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_taken),
    .io_deq_bits_uops_1_br_prediction_bim_resp_value(dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_value),
    .io_deq_bits_uops_1_br_prediction_bim_resp_entry_idx(dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_entry_idx),
    .io_deq_bits_uops_1_br_prediction_bim_resp_way_idx(dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_way_idx),
    .io_deq_bits_uops_1_br_prediction_bpd_resp_takens(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_takens),
    .io_deq_bits_uops_1_br_prediction_bpd_resp_history(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history),
    .io_deq_bits_uops_1_br_prediction_bpd_resp_history_u(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_u),
    .io_deq_bits_uops_1_br_prediction_bpd_resp_history_ptr(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_deq_bits_uops_1_br_prediction_bpd_resp_info(dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_info),
    .io_deq_bits_uops_1_fetch_pc_lob(dec_serializer_io_deq_bits_uops_1_fetch_pc_lob),
    .io_deq_bits_uops_1_xcpt_pf_if(dec_serializer_io_deq_bits_uops_1_xcpt_pf_if),
    .io_deq_bits_uops_1_xcpt_ae_if(dec_serializer_io_deq_bits_uops_1_xcpt_ae_if),
    .io_deq_bits_uops_1_replay_if(dec_serializer_io_deq_bits_uops_1_replay_if),
    .io_deq_bits_uops_1_xcpt_ma_if(dec_serializer_io_deq_bits_uops_1_xcpt_ma_if),
    .io_deq_bits_uops_1_debug_events_fetch_seq(dec_serializer_io_deq_bits_uops_1_debug_events_fetch_seq),
    .io_deq_bits_bpd_resp_info(dec_serializer_io_deq_bits_bpd_resp_info)
  );
  DecodeUnit decode_units_0 (
    .io_enq_uop_valid(decode_units_0_io_enq_uop_valid),
    .io_enq_uop_inst(decode_units_0_io_enq_uop_inst),
    .io_enq_uop_pc(decode_units_0_io_enq_uop_pc),
    .io_enq_uop_br_prediction_btb_blame(decode_units_0_io_enq_uop_br_prediction_btb_blame),
    .io_enq_uop_br_prediction_btb_hit(decode_units_0_io_enq_uop_br_prediction_btb_hit),
    .io_enq_uop_br_prediction_btb_taken(decode_units_0_io_enq_uop_br_prediction_btb_taken),
    .io_enq_uop_br_prediction_bpd_blame(decode_units_0_io_enq_uop_br_prediction_bpd_blame),
    .io_enq_uop_br_prediction_bpd_hit(decode_units_0_io_enq_uop_br_prediction_bpd_hit),
    .io_enq_uop_br_prediction_bpd_taken(decode_units_0_io_enq_uop_br_prediction_bpd_taken),
    .io_enq_uop_br_prediction_bim_resp_value(decode_units_0_io_enq_uop_br_prediction_bim_resp_value),
    .io_enq_uop_br_prediction_bim_resp_entry_idx(decode_units_0_io_enq_uop_br_prediction_bim_resp_entry_idx),
    .io_enq_uop_br_prediction_bim_resp_way_idx(decode_units_0_io_enq_uop_br_prediction_bim_resp_way_idx),
    .io_enq_uop_br_prediction_bpd_resp_takens(decode_units_0_io_enq_uop_br_prediction_bpd_resp_takens),
    .io_enq_uop_br_prediction_bpd_resp_history(decode_units_0_io_enq_uop_br_prediction_bpd_resp_history),
    .io_enq_uop_br_prediction_bpd_resp_history_u(decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_u),
    .io_enq_uop_br_prediction_bpd_resp_history_ptr(decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_ptr),
    .io_enq_uop_br_prediction_bpd_resp_info(decode_units_0_io_enq_uop_br_prediction_bpd_resp_info),
    .io_enq_uop_fetch_pc_lob(decode_units_0_io_enq_uop_fetch_pc_lob),
    .io_enq_uop_xcpt_pf_if(decode_units_0_io_enq_uop_xcpt_pf_if),
    .io_enq_uop_xcpt_ae_if(decode_units_0_io_enq_uop_xcpt_ae_if),
    .io_enq_uop_replay_if(decode_units_0_io_enq_uop_replay_if),
    .io_enq_uop_xcpt_ma_if(decode_units_0_io_enq_uop_xcpt_ma_if),
    .io_enq_uop_debug_events_fetch_seq(decode_units_0_io_enq_uop_debug_events_fetch_seq),
    .io_deq_uop_valid(decode_units_0_io_deq_uop_valid),
    .io_deq_uop_uopc(decode_units_0_io_deq_uop_uopc),
    .io_deq_uop_inst(decode_units_0_io_deq_uop_inst),
    .io_deq_uop_pc(decode_units_0_io_deq_uop_pc),
    .io_deq_uop_iqtype(decode_units_0_io_deq_uop_iqtype),
    .io_deq_uop_fu_code(decode_units_0_io_deq_uop_fu_code),
    .io_deq_uop_allocate_brtag(decode_units_0_io_deq_uop_allocate_brtag),
    .io_deq_uop_is_br_or_jmp(decode_units_0_io_deq_uop_is_br_or_jmp),
    .io_deq_uop_is_jump(decode_units_0_io_deq_uop_is_jump),
    .io_deq_uop_is_jal(decode_units_0_io_deq_uop_is_jal),
    .io_deq_uop_is_ret(decode_units_0_io_deq_uop_is_ret),
    .io_deq_uop_is_call(decode_units_0_io_deq_uop_is_call),
    .io_deq_uop_br_prediction_btb_blame(decode_units_0_io_deq_uop_br_prediction_btb_blame),
    .io_deq_uop_br_prediction_btb_hit(decode_units_0_io_deq_uop_br_prediction_btb_hit),
    .io_deq_uop_br_prediction_btb_taken(decode_units_0_io_deq_uop_br_prediction_btb_taken),
    .io_deq_uop_br_prediction_bpd_blame(decode_units_0_io_deq_uop_br_prediction_bpd_blame),
    .io_deq_uop_br_prediction_bpd_hit(decode_units_0_io_deq_uop_br_prediction_bpd_hit),
    .io_deq_uop_br_prediction_bpd_taken(decode_units_0_io_deq_uop_br_prediction_bpd_taken),
    .io_deq_uop_br_prediction_bim_resp_value(decode_units_0_io_deq_uop_br_prediction_bim_resp_value),
    .io_deq_uop_br_prediction_bim_resp_entry_idx(decode_units_0_io_deq_uop_br_prediction_bim_resp_entry_idx),
    .io_deq_uop_br_prediction_bim_resp_way_idx(decode_units_0_io_deq_uop_br_prediction_bim_resp_way_idx),
    .io_deq_uop_br_prediction_bpd_resp_takens(decode_units_0_io_deq_uop_br_prediction_bpd_resp_takens),
    .io_deq_uop_br_prediction_bpd_resp_history(decode_units_0_io_deq_uop_br_prediction_bpd_resp_history),
    .io_deq_uop_br_prediction_bpd_resp_history_u(decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_u),
    .io_deq_uop_br_prediction_bpd_resp_history_ptr(decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_ptr),
    .io_deq_uop_br_prediction_bpd_resp_info(decode_units_0_io_deq_uop_br_prediction_bpd_resp_info),
    .io_deq_uop_fetch_pc_lob(decode_units_0_io_deq_uop_fetch_pc_lob),
    .io_deq_uop_imm_packed(decode_units_0_io_deq_uop_imm_packed),
    .io_deq_uop_exception(decode_units_0_io_deq_uop_exception),
    .io_deq_uop_exc_cause(decode_units_0_io_deq_uop_exc_cause),
    .io_deq_uop_bypassable(decode_units_0_io_deq_uop_bypassable),
    .io_deq_uop_mem_cmd(decode_units_0_io_deq_uop_mem_cmd),
    .io_deq_uop_mem_typ(decode_units_0_io_deq_uop_mem_typ),
    .io_deq_uop_is_fence(decode_units_0_io_deq_uop_is_fence),
    .io_deq_uop_is_fencei(decode_units_0_io_deq_uop_is_fencei),
    .io_deq_uop_is_store(decode_units_0_io_deq_uop_is_store),
    .io_deq_uop_is_amo(decode_units_0_io_deq_uop_is_amo),
    .io_deq_uop_is_load(decode_units_0_io_deq_uop_is_load),
    .io_deq_uop_is_sys_pc2epc(decode_units_0_io_deq_uop_is_sys_pc2epc),
    .io_deq_uop_is_unique(decode_units_0_io_deq_uop_is_unique),
    .io_deq_uop_flush_on_commit(decode_units_0_io_deq_uop_flush_on_commit),
    .io_deq_uop_ldst(decode_units_0_io_deq_uop_ldst),
    .io_deq_uop_lrs1(decode_units_0_io_deq_uop_lrs1),
    .io_deq_uop_lrs2(decode_units_0_io_deq_uop_lrs2),
    .io_deq_uop_lrs3(decode_units_0_io_deq_uop_lrs3),
    .io_deq_uop_ldst_val(decode_units_0_io_deq_uop_ldst_val),
    .io_deq_uop_dst_rtype(decode_units_0_io_deq_uop_dst_rtype),
    .io_deq_uop_lrs1_rtype(decode_units_0_io_deq_uop_lrs1_rtype),
    .io_deq_uop_lrs2_rtype(decode_units_0_io_deq_uop_lrs2_rtype),
    .io_deq_uop_frs3_en(decode_units_0_io_deq_uop_frs3_en),
    .io_deq_uop_fp_val(decode_units_0_io_deq_uop_fp_val),
    .io_deq_uop_fp_single(decode_units_0_io_deq_uop_fp_single),
    .io_deq_uop_xcpt_pf_if(decode_units_0_io_deq_uop_xcpt_pf_if),
    .io_deq_uop_xcpt_ae_if(decode_units_0_io_deq_uop_xcpt_ae_if),
    .io_deq_uop_replay_if(decode_units_0_io_deq_uop_replay_if),
    .io_deq_uop_xcpt_ma_if(decode_units_0_io_deq_uop_xcpt_ma_if),
    .io_deq_uop_debug_events_fetch_seq(decode_units_0_io_deq_uop_debug_events_fetch_seq),
    .io_status_isa(decode_units_0_io_status_isa),
    .io_csr_decode_csr(decode_units_0_io_csr_decode_csr),
    .io_csr_decode_fp_illegal(decode_units_0_io_csr_decode_fp_illegal),
    .io_csr_decode_read_illegal(decode_units_0_io_csr_decode_read_illegal),
    .io_csr_decode_write_illegal(decode_units_0_io_csr_decode_write_illegal),
    .io_csr_decode_write_flush(decode_units_0_io_csr_decode_write_flush),
    .io_csr_decode_system_illegal(decode_units_0_io_csr_decode_system_illegal),
    .io_interrupt(decode_units_0_io_interrupt),
    .io_interrupt_cause(decode_units_0_io_interrupt_cause)
  );
  DecodeUnit_1 decode_units_1 (
    .io_enq_uop_valid(decode_units_1_io_enq_uop_valid),
    .io_enq_uop_inst(decode_units_1_io_enq_uop_inst),
    .io_enq_uop_pc(decode_units_1_io_enq_uop_pc),
    .io_enq_uop_br_prediction_btb_blame(decode_units_1_io_enq_uop_br_prediction_btb_blame),
    .io_enq_uop_br_prediction_btb_hit(decode_units_1_io_enq_uop_br_prediction_btb_hit),
    .io_enq_uop_br_prediction_btb_taken(decode_units_1_io_enq_uop_br_prediction_btb_taken),
    .io_enq_uop_br_prediction_bpd_blame(decode_units_1_io_enq_uop_br_prediction_bpd_blame),
    .io_enq_uop_br_prediction_bpd_hit(decode_units_1_io_enq_uop_br_prediction_bpd_hit),
    .io_enq_uop_br_prediction_bpd_taken(decode_units_1_io_enq_uop_br_prediction_bpd_taken),
    .io_enq_uop_br_prediction_bim_resp_value(decode_units_1_io_enq_uop_br_prediction_bim_resp_value),
    .io_enq_uop_br_prediction_bim_resp_entry_idx(decode_units_1_io_enq_uop_br_prediction_bim_resp_entry_idx),
    .io_enq_uop_br_prediction_bim_resp_way_idx(decode_units_1_io_enq_uop_br_prediction_bim_resp_way_idx),
    .io_enq_uop_br_prediction_bpd_resp_takens(decode_units_1_io_enq_uop_br_prediction_bpd_resp_takens),
    .io_enq_uop_br_prediction_bpd_resp_history(decode_units_1_io_enq_uop_br_prediction_bpd_resp_history),
    .io_enq_uop_br_prediction_bpd_resp_history_u(decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_u),
    .io_enq_uop_br_prediction_bpd_resp_history_ptr(decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_ptr),
    .io_enq_uop_br_prediction_bpd_resp_info(decode_units_1_io_enq_uop_br_prediction_bpd_resp_info),
    .io_enq_uop_fetch_pc_lob(decode_units_1_io_enq_uop_fetch_pc_lob),
    .io_enq_uop_xcpt_pf_if(decode_units_1_io_enq_uop_xcpt_pf_if),
    .io_enq_uop_xcpt_ae_if(decode_units_1_io_enq_uop_xcpt_ae_if),
    .io_enq_uop_replay_if(decode_units_1_io_enq_uop_replay_if),
    .io_enq_uop_xcpt_ma_if(decode_units_1_io_enq_uop_xcpt_ma_if),
    .io_enq_uop_debug_events_fetch_seq(decode_units_1_io_enq_uop_debug_events_fetch_seq),
    .io_deq_uop_valid(decode_units_1_io_deq_uop_valid),
    .io_deq_uop_uopc(decode_units_1_io_deq_uop_uopc),
    .io_deq_uop_inst(decode_units_1_io_deq_uop_inst),
    .io_deq_uop_pc(decode_units_1_io_deq_uop_pc),
    .io_deq_uop_iqtype(decode_units_1_io_deq_uop_iqtype),
    .io_deq_uop_fu_code(decode_units_1_io_deq_uop_fu_code),
    .io_deq_uop_allocate_brtag(decode_units_1_io_deq_uop_allocate_brtag),
    .io_deq_uop_is_br_or_jmp(decode_units_1_io_deq_uop_is_br_or_jmp),
    .io_deq_uop_is_jump(decode_units_1_io_deq_uop_is_jump),
    .io_deq_uop_is_jal(decode_units_1_io_deq_uop_is_jal),
    .io_deq_uop_is_ret(decode_units_1_io_deq_uop_is_ret),
    .io_deq_uop_is_call(decode_units_1_io_deq_uop_is_call),
    .io_deq_uop_br_prediction_btb_blame(decode_units_1_io_deq_uop_br_prediction_btb_blame),
    .io_deq_uop_br_prediction_btb_hit(decode_units_1_io_deq_uop_br_prediction_btb_hit),
    .io_deq_uop_br_prediction_btb_taken(decode_units_1_io_deq_uop_br_prediction_btb_taken),
    .io_deq_uop_br_prediction_bpd_blame(decode_units_1_io_deq_uop_br_prediction_bpd_blame),
    .io_deq_uop_br_prediction_bpd_hit(decode_units_1_io_deq_uop_br_prediction_bpd_hit),
    .io_deq_uop_br_prediction_bpd_taken(decode_units_1_io_deq_uop_br_prediction_bpd_taken),
    .io_deq_uop_br_prediction_bim_resp_value(decode_units_1_io_deq_uop_br_prediction_bim_resp_value),
    .io_deq_uop_br_prediction_bim_resp_entry_idx(decode_units_1_io_deq_uop_br_prediction_bim_resp_entry_idx),
    .io_deq_uop_br_prediction_bim_resp_way_idx(decode_units_1_io_deq_uop_br_prediction_bim_resp_way_idx),
    .io_deq_uop_br_prediction_bpd_resp_takens(decode_units_1_io_deq_uop_br_prediction_bpd_resp_takens),
    .io_deq_uop_br_prediction_bpd_resp_history(decode_units_1_io_deq_uop_br_prediction_bpd_resp_history),
    .io_deq_uop_br_prediction_bpd_resp_history_u(decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_u),
    .io_deq_uop_br_prediction_bpd_resp_history_ptr(decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_ptr),
    .io_deq_uop_br_prediction_bpd_resp_info(decode_units_1_io_deq_uop_br_prediction_bpd_resp_info),
    .io_deq_uop_fetch_pc_lob(decode_units_1_io_deq_uop_fetch_pc_lob),
    .io_deq_uop_imm_packed(decode_units_1_io_deq_uop_imm_packed),
    .io_deq_uop_exception(decode_units_1_io_deq_uop_exception),
    .io_deq_uop_exc_cause(decode_units_1_io_deq_uop_exc_cause),
    .io_deq_uop_bypassable(decode_units_1_io_deq_uop_bypassable),
    .io_deq_uop_mem_cmd(decode_units_1_io_deq_uop_mem_cmd),
    .io_deq_uop_mem_typ(decode_units_1_io_deq_uop_mem_typ),
    .io_deq_uop_is_fence(decode_units_1_io_deq_uop_is_fence),
    .io_deq_uop_is_fencei(decode_units_1_io_deq_uop_is_fencei),
    .io_deq_uop_is_store(decode_units_1_io_deq_uop_is_store),
    .io_deq_uop_is_amo(decode_units_1_io_deq_uop_is_amo),
    .io_deq_uop_is_load(decode_units_1_io_deq_uop_is_load),
    .io_deq_uop_is_sys_pc2epc(decode_units_1_io_deq_uop_is_sys_pc2epc),
    .io_deq_uop_is_unique(decode_units_1_io_deq_uop_is_unique),
    .io_deq_uop_flush_on_commit(decode_units_1_io_deq_uop_flush_on_commit),
    .io_deq_uop_ldst(decode_units_1_io_deq_uop_ldst),
    .io_deq_uop_lrs1(decode_units_1_io_deq_uop_lrs1),
    .io_deq_uop_lrs2(decode_units_1_io_deq_uop_lrs2),
    .io_deq_uop_lrs3(decode_units_1_io_deq_uop_lrs3),
    .io_deq_uop_ldst_val(decode_units_1_io_deq_uop_ldst_val),
    .io_deq_uop_dst_rtype(decode_units_1_io_deq_uop_dst_rtype),
    .io_deq_uop_lrs1_rtype(decode_units_1_io_deq_uop_lrs1_rtype),
    .io_deq_uop_lrs2_rtype(decode_units_1_io_deq_uop_lrs2_rtype),
    .io_deq_uop_frs3_en(decode_units_1_io_deq_uop_frs3_en),
    .io_deq_uop_fp_val(decode_units_1_io_deq_uop_fp_val),
    .io_deq_uop_fp_single(decode_units_1_io_deq_uop_fp_single),
    .io_deq_uop_xcpt_pf_if(decode_units_1_io_deq_uop_xcpt_pf_if),
    .io_deq_uop_xcpt_ae_if(decode_units_1_io_deq_uop_xcpt_ae_if),
    .io_deq_uop_replay_if(decode_units_1_io_deq_uop_replay_if),
    .io_deq_uop_xcpt_ma_if(decode_units_1_io_deq_uop_xcpt_ma_if),
    .io_deq_uop_debug_events_fetch_seq(decode_units_1_io_deq_uop_debug_events_fetch_seq),
    .io_status_isa(decode_units_1_io_status_isa),
    .io_csr_decode_csr(decode_units_1_io_csr_decode_csr),
    .io_csr_decode_fp_illegal(decode_units_1_io_csr_decode_fp_illegal),
    .io_csr_decode_read_illegal(decode_units_1_io_csr_decode_read_illegal),
    .io_csr_decode_write_illegal(decode_units_1_io_csr_decode_write_illegal),
    .io_csr_decode_write_flush(decode_units_1_io_csr_decode_write_flush),
    .io_csr_decode_system_illegal(decode_units_1_io_csr_decode_system_illegal),
    .io_interrupt(decode_units_1_io_interrupt),
    .io_interrupt_cause(decode_units_1_io_interrupt_cause)
  );
  BranchMaskGenerationLogic dec_brmask_logic (
    .clock(dec_brmask_logic_clock),
    .reset(dec_brmask_logic_reset),
    .io_is_branch_0(dec_brmask_logic_io_is_branch_0),
    .io_is_branch_1(dec_brmask_logic_io_is_branch_1),
    .io_will_fire_0(dec_brmask_logic_io_will_fire_0),
    .io_will_fire_1(dec_brmask_logic_io_will_fire_1),
    .io_br_tag_0(dec_brmask_logic_io_br_tag_0),
    .io_br_tag_1(dec_brmask_logic_io_br_tag_1),
    .io_br_mask_0(dec_brmask_logic_io_br_mask_0),
    .io_br_mask_1(dec_brmask_logic_io_br_mask_1),
    .io_is_full_0(dec_brmask_logic_io_is_full_0),
    .io_is_full_1(dec_brmask_logic_io_is_full_1),
    .io_brinfo_valid(dec_brmask_logic_io_brinfo_valid),
    .io_brinfo_mispredict(dec_brmask_logic_io_brinfo_mispredict),
    .io_brinfo_mask(dec_brmask_logic_io_brinfo_mask),
    .io_brinfo_exe_mask(dec_brmask_logic_io_brinfo_exe_mask),
    .io_flush_pipeline(dec_brmask_logic_io_flush_pipeline)
  );
  RenameStage rename_stage (
    .clock(rename_stage_clock),
    .reset(rename_stage_reset),
    .io_inst_can_proceed_0(rename_stage_io_inst_can_proceed_0),
    .io_inst_can_proceed_1(rename_stage_io_inst_can_proceed_1),
    .io_kill(rename_stage_io_kill),
    .io_dec_will_fire_0(rename_stage_io_dec_will_fire_0),
    .io_dec_will_fire_1(rename_stage_io_dec_will_fire_1),
    .io_dec_uops_0_valid(rename_stage_io_dec_uops_0_valid),
    .io_dec_uops_0_uopc(rename_stage_io_dec_uops_0_uopc),
    .io_dec_uops_0_inst(rename_stage_io_dec_uops_0_inst),
    .io_dec_uops_0_pc(rename_stage_io_dec_uops_0_pc),
    .io_dec_uops_0_iqtype(rename_stage_io_dec_uops_0_iqtype),
    .io_dec_uops_0_fu_code(rename_stage_io_dec_uops_0_fu_code),
    .io_dec_uops_0_allocate_brtag(rename_stage_io_dec_uops_0_allocate_brtag),
    .io_dec_uops_0_is_br_or_jmp(rename_stage_io_dec_uops_0_is_br_or_jmp),
    .io_dec_uops_0_is_jump(rename_stage_io_dec_uops_0_is_jump),
    .io_dec_uops_0_is_jal(rename_stage_io_dec_uops_0_is_jal),
    .io_dec_uops_0_is_ret(rename_stage_io_dec_uops_0_is_ret),
    .io_dec_uops_0_is_call(rename_stage_io_dec_uops_0_is_call),
    .io_dec_uops_0_br_mask(rename_stage_io_dec_uops_0_br_mask),
    .io_dec_uops_0_br_tag(rename_stage_io_dec_uops_0_br_tag),
    .io_dec_uops_0_br_prediction_btb_blame(rename_stage_io_dec_uops_0_br_prediction_btb_blame),
    .io_dec_uops_0_br_prediction_btb_hit(rename_stage_io_dec_uops_0_br_prediction_btb_hit),
    .io_dec_uops_0_br_prediction_btb_taken(rename_stage_io_dec_uops_0_br_prediction_btb_taken),
    .io_dec_uops_0_br_prediction_bpd_blame(rename_stage_io_dec_uops_0_br_prediction_bpd_blame),
    .io_dec_uops_0_br_prediction_bpd_hit(rename_stage_io_dec_uops_0_br_prediction_bpd_hit),
    .io_dec_uops_0_br_prediction_bpd_taken(rename_stage_io_dec_uops_0_br_prediction_bpd_taken),
    .io_dec_uops_0_br_prediction_bim_resp_value(rename_stage_io_dec_uops_0_br_prediction_bim_resp_value),
    .io_dec_uops_0_br_prediction_bim_resp_entry_idx(rename_stage_io_dec_uops_0_br_prediction_bim_resp_entry_idx),
    .io_dec_uops_0_br_prediction_bim_resp_way_idx(rename_stage_io_dec_uops_0_br_prediction_bim_resp_way_idx),
    .io_dec_uops_0_br_prediction_bpd_resp_takens(rename_stage_io_dec_uops_0_br_prediction_bpd_resp_takens),
    .io_dec_uops_0_br_prediction_bpd_resp_history(rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history),
    .io_dec_uops_0_br_prediction_bpd_resp_history_u(rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_u),
    .io_dec_uops_0_br_prediction_bpd_resp_history_ptr(rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_dec_uops_0_br_prediction_bpd_resp_info(rename_stage_io_dec_uops_0_br_prediction_bpd_resp_info),
    .io_dec_uops_0_fetch_pc_lob(rename_stage_io_dec_uops_0_fetch_pc_lob),
    .io_dec_uops_0_imm_packed(rename_stage_io_dec_uops_0_imm_packed),
    .io_dec_uops_0_rob_idx(rename_stage_io_dec_uops_0_rob_idx),
    .io_dec_uops_0_ldq_idx(rename_stage_io_dec_uops_0_ldq_idx),
    .io_dec_uops_0_stq_idx(rename_stage_io_dec_uops_0_stq_idx),
    .io_dec_uops_0_brob_idx(rename_stage_io_dec_uops_0_brob_idx),
    .io_dec_uops_0_exception(rename_stage_io_dec_uops_0_exception),
    .io_dec_uops_0_exc_cause(rename_stage_io_dec_uops_0_exc_cause),
    .io_dec_uops_0_bypassable(rename_stage_io_dec_uops_0_bypassable),
    .io_dec_uops_0_mem_cmd(rename_stage_io_dec_uops_0_mem_cmd),
    .io_dec_uops_0_mem_typ(rename_stage_io_dec_uops_0_mem_typ),
    .io_dec_uops_0_is_fence(rename_stage_io_dec_uops_0_is_fence),
    .io_dec_uops_0_is_fencei(rename_stage_io_dec_uops_0_is_fencei),
    .io_dec_uops_0_is_store(rename_stage_io_dec_uops_0_is_store),
    .io_dec_uops_0_is_amo(rename_stage_io_dec_uops_0_is_amo),
    .io_dec_uops_0_is_load(rename_stage_io_dec_uops_0_is_load),
    .io_dec_uops_0_is_sys_pc2epc(rename_stage_io_dec_uops_0_is_sys_pc2epc),
    .io_dec_uops_0_is_unique(rename_stage_io_dec_uops_0_is_unique),
    .io_dec_uops_0_flush_on_commit(rename_stage_io_dec_uops_0_flush_on_commit),
    .io_dec_uops_0_ldst(rename_stage_io_dec_uops_0_ldst),
    .io_dec_uops_0_lrs1(rename_stage_io_dec_uops_0_lrs1),
    .io_dec_uops_0_lrs2(rename_stage_io_dec_uops_0_lrs2),
    .io_dec_uops_0_lrs3(rename_stage_io_dec_uops_0_lrs3),
    .io_dec_uops_0_ldst_val(rename_stage_io_dec_uops_0_ldst_val),
    .io_dec_uops_0_dst_rtype(rename_stage_io_dec_uops_0_dst_rtype),
    .io_dec_uops_0_lrs1_rtype(rename_stage_io_dec_uops_0_lrs1_rtype),
    .io_dec_uops_0_lrs2_rtype(rename_stage_io_dec_uops_0_lrs2_rtype),
    .io_dec_uops_0_frs3_en(rename_stage_io_dec_uops_0_frs3_en),
    .io_dec_uops_0_fp_val(rename_stage_io_dec_uops_0_fp_val),
    .io_dec_uops_0_fp_single(rename_stage_io_dec_uops_0_fp_single),
    .io_dec_uops_0_xcpt_pf_if(rename_stage_io_dec_uops_0_xcpt_pf_if),
    .io_dec_uops_0_xcpt_ae_if(rename_stage_io_dec_uops_0_xcpt_ae_if),
    .io_dec_uops_0_replay_if(rename_stage_io_dec_uops_0_replay_if),
    .io_dec_uops_0_xcpt_ma_if(rename_stage_io_dec_uops_0_xcpt_ma_if),
    .io_dec_uops_0_debug_events_fetch_seq(rename_stage_io_dec_uops_0_debug_events_fetch_seq),
    .io_dec_uops_1_valid(rename_stage_io_dec_uops_1_valid),
    .io_dec_uops_1_uopc(rename_stage_io_dec_uops_1_uopc),
    .io_dec_uops_1_inst(rename_stage_io_dec_uops_1_inst),
    .io_dec_uops_1_pc(rename_stage_io_dec_uops_1_pc),
    .io_dec_uops_1_iqtype(rename_stage_io_dec_uops_1_iqtype),
    .io_dec_uops_1_fu_code(rename_stage_io_dec_uops_1_fu_code),
    .io_dec_uops_1_allocate_brtag(rename_stage_io_dec_uops_1_allocate_brtag),
    .io_dec_uops_1_is_br_or_jmp(rename_stage_io_dec_uops_1_is_br_or_jmp),
    .io_dec_uops_1_is_jump(rename_stage_io_dec_uops_1_is_jump),
    .io_dec_uops_1_is_jal(rename_stage_io_dec_uops_1_is_jal),
    .io_dec_uops_1_is_ret(rename_stage_io_dec_uops_1_is_ret),
    .io_dec_uops_1_is_call(rename_stage_io_dec_uops_1_is_call),
    .io_dec_uops_1_br_mask(rename_stage_io_dec_uops_1_br_mask),
    .io_dec_uops_1_br_tag(rename_stage_io_dec_uops_1_br_tag),
    .io_dec_uops_1_br_prediction_btb_blame(rename_stage_io_dec_uops_1_br_prediction_btb_blame),
    .io_dec_uops_1_br_prediction_btb_hit(rename_stage_io_dec_uops_1_br_prediction_btb_hit),
    .io_dec_uops_1_br_prediction_btb_taken(rename_stage_io_dec_uops_1_br_prediction_btb_taken),
    .io_dec_uops_1_br_prediction_bpd_blame(rename_stage_io_dec_uops_1_br_prediction_bpd_blame),
    .io_dec_uops_1_br_prediction_bpd_hit(rename_stage_io_dec_uops_1_br_prediction_bpd_hit),
    .io_dec_uops_1_br_prediction_bpd_taken(rename_stage_io_dec_uops_1_br_prediction_bpd_taken),
    .io_dec_uops_1_br_prediction_bim_resp_value(rename_stage_io_dec_uops_1_br_prediction_bim_resp_value),
    .io_dec_uops_1_br_prediction_bim_resp_entry_idx(rename_stage_io_dec_uops_1_br_prediction_bim_resp_entry_idx),
    .io_dec_uops_1_br_prediction_bim_resp_way_idx(rename_stage_io_dec_uops_1_br_prediction_bim_resp_way_idx),
    .io_dec_uops_1_br_prediction_bpd_resp_takens(rename_stage_io_dec_uops_1_br_prediction_bpd_resp_takens),
    .io_dec_uops_1_br_prediction_bpd_resp_history(rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history),
    .io_dec_uops_1_br_prediction_bpd_resp_history_u(rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_u),
    .io_dec_uops_1_br_prediction_bpd_resp_history_ptr(rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_dec_uops_1_br_prediction_bpd_resp_info(rename_stage_io_dec_uops_1_br_prediction_bpd_resp_info),
    .io_dec_uops_1_fetch_pc_lob(rename_stage_io_dec_uops_1_fetch_pc_lob),
    .io_dec_uops_1_imm_packed(rename_stage_io_dec_uops_1_imm_packed),
    .io_dec_uops_1_rob_idx(rename_stage_io_dec_uops_1_rob_idx),
    .io_dec_uops_1_ldq_idx(rename_stage_io_dec_uops_1_ldq_idx),
    .io_dec_uops_1_stq_idx(rename_stage_io_dec_uops_1_stq_idx),
    .io_dec_uops_1_brob_idx(rename_stage_io_dec_uops_1_brob_idx),
    .io_dec_uops_1_exception(rename_stage_io_dec_uops_1_exception),
    .io_dec_uops_1_exc_cause(rename_stage_io_dec_uops_1_exc_cause),
    .io_dec_uops_1_bypassable(rename_stage_io_dec_uops_1_bypassable),
    .io_dec_uops_1_mem_cmd(rename_stage_io_dec_uops_1_mem_cmd),
    .io_dec_uops_1_mem_typ(rename_stage_io_dec_uops_1_mem_typ),
    .io_dec_uops_1_is_fence(rename_stage_io_dec_uops_1_is_fence),
    .io_dec_uops_1_is_fencei(rename_stage_io_dec_uops_1_is_fencei),
    .io_dec_uops_1_is_store(rename_stage_io_dec_uops_1_is_store),
    .io_dec_uops_1_is_amo(rename_stage_io_dec_uops_1_is_amo),
    .io_dec_uops_1_is_load(rename_stage_io_dec_uops_1_is_load),
    .io_dec_uops_1_is_sys_pc2epc(rename_stage_io_dec_uops_1_is_sys_pc2epc),
    .io_dec_uops_1_is_unique(rename_stage_io_dec_uops_1_is_unique),
    .io_dec_uops_1_flush_on_commit(rename_stage_io_dec_uops_1_flush_on_commit),
    .io_dec_uops_1_ldst(rename_stage_io_dec_uops_1_ldst),
    .io_dec_uops_1_lrs1(rename_stage_io_dec_uops_1_lrs1),
    .io_dec_uops_1_lrs2(rename_stage_io_dec_uops_1_lrs2),
    .io_dec_uops_1_lrs3(rename_stage_io_dec_uops_1_lrs3),
    .io_dec_uops_1_ldst_val(rename_stage_io_dec_uops_1_ldst_val),
    .io_dec_uops_1_dst_rtype(rename_stage_io_dec_uops_1_dst_rtype),
    .io_dec_uops_1_lrs1_rtype(rename_stage_io_dec_uops_1_lrs1_rtype),
    .io_dec_uops_1_lrs2_rtype(rename_stage_io_dec_uops_1_lrs2_rtype),
    .io_dec_uops_1_frs3_en(rename_stage_io_dec_uops_1_frs3_en),
    .io_dec_uops_1_fp_val(rename_stage_io_dec_uops_1_fp_val),
    .io_dec_uops_1_fp_single(rename_stage_io_dec_uops_1_fp_single),
    .io_dec_uops_1_xcpt_pf_if(rename_stage_io_dec_uops_1_xcpt_pf_if),
    .io_dec_uops_1_xcpt_ae_if(rename_stage_io_dec_uops_1_xcpt_ae_if),
    .io_dec_uops_1_replay_if(rename_stage_io_dec_uops_1_replay_if),
    .io_dec_uops_1_xcpt_ma_if(rename_stage_io_dec_uops_1_xcpt_ma_if),
    .io_dec_uops_1_debug_events_fetch_seq(rename_stage_io_dec_uops_1_debug_events_fetch_seq),
    .io_ren1_mask_0(rename_stage_io_ren1_mask_0),
    .io_ren1_mask_1(rename_stage_io_ren1_mask_1),
    .io_ren1_uops_0_pc(rename_stage_io_ren1_uops_0_pc),
    .io_ren1_uops_0_br_mask(rename_stage_io_ren1_uops_0_br_mask),
    .io_ren1_uops_0_rob_idx(rename_stage_io_ren1_uops_0_rob_idx),
    .io_ren1_uops_0_brob_idx(rename_stage_io_ren1_uops_0_brob_idx),
    .io_ren1_uops_0_pdst(rename_stage_io_ren1_uops_0_pdst),
    .io_ren1_uops_0_stale_pdst(rename_stage_io_ren1_uops_0_stale_pdst),
    .io_ren1_uops_0_exception(rename_stage_io_ren1_uops_0_exception),
    .io_ren1_uops_0_exc_cause(rename_stage_io_ren1_uops_0_exc_cause),
    .io_ren1_uops_0_is_fence(rename_stage_io_ren1_uops_0_is_fence),
    .io_ren1_uops_0_is_fencei(rename_stage_io_ren1_uops_0_is_fencei),
    .io_ren1_uops_0_is_store(rename_stage_io_ren1_uops_0_is_store),
    .io_ren1_uops_0_is_load(rename_stage_io_ren1_uops_0_is_load),
    .io_ren1_uops_0_is_sys_pc2epc(rename_stage_io_ren1_uops_0_is_sys_pc2epc),
    .io_ren1_uops_0_is_unique(rename_stage_io_ren1_uops_0_is_unique),
    .io_ren1_uops_0_flush_on_commit(rename_stage_io_ren1_uops_0_flush_on_commit),
    .io_ren1_uops_0_ldst(rename_stage_io_ren1_uops_0_ldst),
    .io_ren1_uops_0_ldst_val(rename_stage_io_ren1_uops_0_ldst_val),
    .io_ren1_uops_0_dst_rtype(rename_stage_io_ren1_uops_0_dst_rtype),
    .io_ren1_uops_0_fp_val(rename_stage_io_ren1_uops_0_fp_val),
    .io_ren1_uops_1_br_mask(rename_stage_io_ren1_uops_1_br_mask),
    .io_ren1_uops_1_rob_idx(rename_stage_io_ren1_uops_1_rob_idx),
    .io_ren1_uops_1_pdst(rename_stage_io_ren1_uops_1_pdst),
    .io_ren1_uops_1_stale_pdst(rename_stage_io_ren1_uops_1_stale_pdst),
    .io_ren1_uops_1_exception(rename_stage_io_ren1_uops_1_exception),
    .io_ren1_uops_1_exc_cause(rename_stage_io_ren1_uops_1_exc_cause),
    .io_ren1_uops_1_is_fence(rename_stage_io_ren1_uops_1_is_fence),
    .io_ren1_uops_1_is_fencei(rename_stage_io_ren1_uops_1_is_fencei),
    .io_ren1_uops_1_is_store(rename_stage_io_ren1_uops_1_is_store),
    .io_ren1_uops_1_is_load(rename_stage_io_ren1_uops_1_is_load),
    .io_ren1_uops_1_is_sys_pc2epc(rename_stage_io_ren1_uops_1_is_sys_pc2epc),
    .io_ren1_uops_1_is_unique(rename_stage_io_ren1_uops_1_is_unique),
    .io_ren1_uops_1_flush_on_commit(rename_stage_io_ren1_uops_1_flush_on_commit),
    .io_ren1_uops_1_ldst(rename_stage_io_ren1_uops_1_ldst),
    .io_ren1_uops_1_ldst_val(rename_stage_io_ren1_uops_1_ldst_val),
    .io_ren1_uops_1_dst_rtype(rename_stage_io_ren1_uops_1_dst_rtype),
    .io_ren1_uops_1_fp_val(rename_stage_io_ren1_uops_1_fp_val),
    .io_ren2_mask_0(rename_stage_io_ren2_mask_0),
    .io_ren2_mask_1(rename_stage_io_ren2_mask_1),
    .io_ren2_uops_0_valid(rename_stage_io_ren2_uops_0_valid),
    .io_ren2_uops_0_uopc(rename_stage_io_ren2_uops_0_uopc),
    .io_ren2_uops_0_inst(rename_stage_io_ren2_uops_0_inst),
    .io_ren2_uops_0_pc(rename_stage_io_ren2_uops_0_pc),
    .io_ren2_uops_0_iqtype(rename_stage_io_ren2_uops_0_iqtype),
    .io_ren2_uops_0_fu_code(rename_stage_io_ren2_uops_0_fu_code),
    .io_ren2_uops_0_allocate_brtag(rename_stage_io_ren2_uops_0_allocate_brtag),
    .io_ren2_uops_0_is_br_or_jmp(rename_stage_io_ren2_uops_0_is_br_or_jmp),
    .io_ren2_uops_0_is_jump(rename_stage_io_ren2_uops_0_is_jump),
    .io_ren2_uops_0_is_jal(rename_stage_io_ren2_uops_0_is_jal),
    .io_ren2_uops_0_is_ret(rename_stage_io_ren2_uops_0_is_ret),
    .io_ren2_uops_0_is_call(rename_stage_io_ren2_uops_0_is_call),
    .io_ren2_uops_0_br_mask(rename_stage_io_ren2_uops_0_br_mask),
    .io_ren2_uops_0_br_tag(rename_stage_io_ren2_uops_0_br_tag),
    .io_ren2_uops_0_br_prediction_btb_blame(rename_stage_io_ren2_uops_0_br_prediction_btb_blame),
    .io_ren2_uops_0_br_prediction_btb_hit(rename_stage_io_ren2_uops_0_br_prediction_btb_hit),
    .io_ren2_uops_0_br_prediction_btb_taken(rename_stage_io_ren2_uops_0_br_prediction_btb_taken),
    .io_ren2_uops_0_br_prediction_bpd_blame(rename_stage_io_ren2_uops_0_br_prediction_bpd_blame),
    .io_ren2_uops_0_br_prediction_bpd_hit(rename_stage_io_ren2_uops_0_br_prediction_bpd_hit),
    .io_ren2_uops_0_br_prediction_bpd_taken(rename_stage_io_ren2_uops_0_br_prediction_bpd_taken),
    .io_ren2_uops_0_br_prediction_bim_resp_value(rename_stage_io_ren2_uops_0_br_prediction_bim_resp_value),
    .io_ren2_uops_0_br_prediction_bim_resp_entry_idx(rename_stage_io_ren2_uops_0_br_prediction_bim_resp_entry_idx),
    .io_ren2_uops_0_br_prediction_bim_resp_way_idx(rename_stage_io_ren2_uops_0_br_prediction_bim_resp_way_idx),
    .io_ren2_uops_0_br_prediction_bpd_resp_takens(rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_takens),
    .io_ren2_uops_0_br_prediction_bpd_resp_history(rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history),
    .io_ren2_uops_0_br_prediction_bpd_resp_history_u(rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_u),
    .io_ren2_uops_0_br_prediction_bpd_resp_history_ptr(rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_ren2_uops_0_br_prediction_bpd_resp_info(rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_info),
    .io_ren2_uops_0_stat_brjmp_mispredicted(rename_stage_io_ren2_uops_0_stat_brjmp_mispredicted),
    .io_ren2_uops_0_stat_btb_made_pred(rename_stage_io_ren2_uops_0_stat_btb_made_pred),
    .io_ren2_uops_0_stat_btb_mispredicted(rename_stage_io_ren2_uops_0_stat_btb_mispredicted),
    .io_ren2_uops_0_stat_bpd_made_pred(rename_stage_io_ren2_uops_0_stat_bpd_made_pred),
    .io_ren2_uops_0_stat_bpd_mispredicted(rename_stage_io_ren2_uops_0_stat_bpd_mispredicted),
    .io_ren2_uops_0_fetch_pc_lob(rename_stage_io_ren2_uops_0_fetch_pc_lob),
    .io_ren2_uops_0_imm_packed(rename_stage_io_ren2_uops_0_imm_packed),
    .io_ren2_uops_0_csr_addr(rename_stage_io_ren2_uops_0_csr_addr),
    .io_ren2_uops_0_rob_idx(rename_stage_io_ren2_uops_0_rob_idx),
    .io_ren2_uops_0_ldq_idx(rename_stage_io_ren2_uops_0_ldq_idx),
    .io_ren2_uops_0_stq_idx(rename_stage_io_ren2_uops_0_stq_idx),
    .io_ren2_uops_0_brob_idx(rename_stage_io_ren2_uops_0_brob_idx),
    .io_ren2_uops_0_pdst(rename_stage_io_ren2_uops_0_pdst),
    .io_ren2_uops_0_pop1(rename_stage_io_ren2_uops_0_pop1),
    .io_ren2_uops_0_pop2(rename_stage_io_ren2_uops_0_pop2),
    .io_ren2_uops_0_pop3(rename_stage_io_ren2_uops_0_pop3),
    .io_ren2_uops_0_prs1_busy(rename_stage_io_ren2_uops_0_prs1_busy),
    .io_ren2_uops_0_prs2_busy(rename_stage_io_ren2_uops_0_prs2_busy),
    .io_ren2_uops_0_prs3_busy(rename_stage_io_ren2_uops_0_prs3_busy),
    .io_ren2_uops_0_stale_pdst(rename_stage_io_ren2_uops_0_stale_pdst),
    .io_ren2_uops_0_exception(rename_stage_io_ren2_uops_0_exception),
    .io_ren2_uops_0_exc_cause(rename_stage_io_ren2_uops_0_exc_cause),
    .io_ren2_uops_0_bypassable(rename_stage_io_ren2_uops_0_bypassable),
    .io_ren2_uops_0_mem_cmd(rename_stage_io_ren2_uops_0_mem_cmd),
    .io_ren2_uops_0_mem_typ(rename_stage_io_ren2_uops_0_mem_typ),
    .io_ren2_uops_0_is_fence(rename_stage_io_ren2_uops_0_is_fence),
    .io_ren2_uops_0_is_fencei(rename_stage_io_ren2_uops_0_is_fencei),
    .io_ren2_uops_0_is_store(rename_stage_io_ren2_uops_0_is_store),
    .io_ren2_uops_0_is_amo(rename_stage_io_ren2_uops_0_is_amo),
    .io_ren2_uops_0_is_load(rename_stage_io_ren2_uops_0_is_load),
    .io_ren2_uops_0_is_sys_pc2epc(rename_stage_io_ren2_uops_0_is_sys_pc2epc),
    .io_ren2_uops_0_is_unique(rename_stage_io_ren2_uops_0_is_unique),
    .io_ren2_uops_0_flush_on_commit(rename_stage_io_ren2_uops_0_flush_on_commit),
    .io_ren2_uops_0_ldst(rename_stage_io_ren2_uops_0_ldst),
    .io_ren2_uops_0_lrs1(rename_stage_io_ren2_uops_0_lrs1),
    .io_ren2_uops_0_lrs2(rename_stage_io_ren2_uops_0_lrs2),
    .io_ren2_uops_0_lrs3(rename_stage_io_ren2_uops_0_lrs3),
    .io_ren2_uops_0_ldst_val(rename_stage_io_ren2_uops_0_ldst_val),
    .io_ren2_uops_0_dst_rtype(rename_stage_io_ren2_uops_0_dst_rtype),
    .io_ren2_uops_0_lrs1_rtype(rename_stage_io_ren2_uops_0_lrs1_rtype),
    .io_ren2_uops_0_lrs2_rtype(rename_stage_io_ren2_uops_0_lrs2_rtype),
    .io_ren2_uops_0_frs3_en(rename_stage_io_ren2_uops_0_frs3_en),
    .io_ren2_uops_0_fp_val(rename_stage_io_ren2_uops_0_fp_val),
    .io_ren2_uops_0_fp_single(rename_stage_io_ren2_uops_0_fp_single),
    .io_ren2_uops_0_xcpt_pf_if(rename_stage_io_ren2_uops_0_xcpt_pf_if),
    .io_ren2_uops_0_xcpt_ae_if(rename_stage_io_ren2_uops_0_xcpt_ae_if),
    .io_ren2_uops_0_replay_if(rename_stage_io_ren2_uops_0_replay_if),
    .io_ren2_uops_0_xcpt_ma_if(rename_stage_io_ren2_uops_0_xcpt_ma_if),
    .io_ren2_uops_0_debug_wdata(rename_stage_io_ren2_uops_0_debug_wdata),
    .io_ren2_uops_0_debug_events_fetch_seq(rename_stage_io_ren2_uops_0_debug_events_fetch_seq),
    .io_ren2_uops_1_valid(rename_stage_io_ren2_uops_1_valid),
    .io_ren2_uops_1_uopc(rename_stage_io_ren2_uops_1_uopc),
    .io_ren2_uops_1_inst(rename_stage_io_ren2_uops_1_inst),
    .io_ren2_uops_1_pc(rename_stage_io_ren2_uops_1_pc),
    .io_ren2_uops_1_iqtype(rename_stage_io_ren2_uops_1_iqtype),
    .io_ren2_uops_1_fu_code(rename_stage_io_ren2_uops_1_fu_code),
    .io_ren2_uops_1_allocate_brtag(rename_stage_io_ren2_uops_1_allocate_brtag),
    .io_ren2_uops_1_is_br_or_jmp(rename_stage_io_ren2_uops_1_is_br_or_jmp),
    .io_ren2_uops_1_is_jump(rename_stage_io_ren2_uops_1_is_jump),
    .io_ren2_uops_1_is_jal(rename_stage_io_ren2_uops_1_is_jal),
    .io_ren2_uops_1_is_ret(rename_stage_io_ren2_uops_1_is_ret),
    .io_ren2_uops_1_is_call(rename_stage_io_ren2_uops_1_is_call),
    .io_ren2_uops_1_br_mask(rename_stage_io_ren2_uops_1_br_mask),
    .io_ren2_uops_1_br_tag(rename_stage_io_ren2_uops_1_br_tag),
    .io_ren2_uops_1_br_prediction_btb_blame(rename_stage_io_ren2_uops_1_br_prediction_btb_blame),
    .io_ren2_uops_1_br_prediction_btb_hit(rename_stage_io_ren2_uops_1_br_prediction_btb_hit),
    .io_ren2_uops_1_br_prediction_btb_taken(rename_stage_io_ren2_uops_1_br_prediction_btb_taken),
    .io_ren2_uops_1_br_prediction_bpd_blame(rename_stage_io_ren2_uops_1_br_prediction_bpd_blame),
    .io_ren2_uops_1_br_prediction_bpd_hit(rename_stage_io_ren2_uops_1_br_prediction_bpd_hit),
    .io_ren2_uops_1_br_prediction_bpd_taken(rename_stage_io_ren2_uops_1_br_prediction_bpd_taken),
    .io_ren2_uops_1_br_prediction_bim_resp_value(rename_stage_io_ren2_uops_1_br_prediction_bim_resp_value),
    .io_ren2_uops_1_br_prediction_bim_resp_entry_idx(rename_stage_io_ren2_uops_1_br_prediction_bim_resp_entry_idx),
    .io_ren2_uops_1_br_prediction_bim_resp_way_idx(rename_stage_io_ren2_uops_1_br_prediction_bim_resp_way_idx),
    .io_ren2_uops_1_br_prediction_bpd_resp_takens(rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_takens),
    .io_ren2_uops_1_br_prediction_bpd_resp_history(rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history),
    .io_ren2_uops_1_br_prediction_bpd_resp_history_u(rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_u),
    .io_ren2_uops_1_br_prediction_bpd_resp_history_ptr(rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_ren2_uops_1_br_prediction_bpd_resp_info(rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_info),
    .io_ren2_uops_1_stat_brjmp_mispredicted(rename_stage_io_ren2_uops_1_stat_brjmp_mispredicted),
    .io_ren2_uops_1_stat_btb_made_pred(rename_stage_io_ren2_uops_1_stat_btb_made_pred),
    .io_ren2_uops_1_stat_btb_mispredicted(rename_stage_io_ren2_uops_1_stat_btb_mispredicted),
    .io_ren2_uops_1_stat_bpd_made_pred(rename_stage_io_ren2_uops_1_stat_bpd_made_pred),
    .io_ren2_uops_1_stat_bpd_mispredicted(rename_stage_io_ren2_uops_1_stat_bpd_mispredicted),
    .io_ren2_uops_1_fetch_pc_lob(rename_stage_io_ren2_uops_1_fetch_pc_lob),
    .io_ren2_uops_1_imm_packed(rename_stage_io_ren2_uops_1_imm_packed),
    .io_ren2_uops_1_csr_addr(rename_stage_io_ren2_uops_1_csr_addr),
    .io_ren2_uops_1_rob_idx(rename_stage_io_ren2_uops_1_rob_idx),
    .io_ren2_uops_1_ldq_idx(rename_stage_io_ren2_uops_1_ldq_idx),
    .io_ren2_uops_1_stq_idx(rename_stage_io_ren2_uops_1_stq_idx),
    .io_ren2_uops_1_brob_idx(rename_stage_io_ren2_uops_1_brob_idx),
    .io_ren2_uops_1_pdst(rename_stage_io_ren2_uops_1_pdst),
    .io_ren2_uops_1_pop1(rename_stage_io_ren2_uops_1_pop1),
    .io_ren2_uops_1_pop2(rename_stage_io_ren2_uops_1_pop2),
    .io_ren2_uops_1_pop3(rename_stage_io_ren2_uops_1_pop3),
    .io_ren2_uops_1_prs1_busy(rename_stage_io_ren2_uops_1_prs1_busy),
    .io_ren2_uops_1_prs2_busy(rename_stage_io_ren2_uops_1_prs2_busy),
    .io_ren2_uops_1_prs3_busy(rename_stage_io_ren2_uops_1_prs3_busy),
    .io_ren2_uops_1_stale_pdst(rename_stage_io_ren2_uops_1_stale_pdst),
    .io_ren2_uops_1_exception(rename_stage_io_ren2_uops_1_exception),
    .io_ren2_uops_1_exc_cause(rename_stage_io_ren2_uops_1_exc_cause),
    .io_ren2_uops_1_bypassable(rename_stage_io_ren2_uops_1_bypassable),
    .io_ren2_uops_1_mem_cmd(rename_stage_io_ren2_uops_1_mem_cmd),
    .io_ren2_uops_1_mem_typ(rename_stage_io_ren2_uops_1_mem_typ),
    .io_ren2_uops_1_is_fence(rename_stage_io_ren2_uops_1_is_fence),
    .io_ren2_uops_1_is_fencei(rename_stage_io_ren2_uops_1_is_fencei),
    .io_ren2_uops_1_is_store(rename_stage_io_ren2_uops_1_is_store),
    .io_ren2_uops_1_is_amo(rename_stage_io_ren2_uops_1_is_amo),
    .io_ren2_uops_1_is_load(rename_stage_io_ren2_uops_1_is_load),
    .io_ren2_uops_1_is_sys_pc2epc(rename_stage_io_ren2_uops_1_is_sys_pc2epc),
    .io_ren2_uops_1_is_unique(rename_stage_io_ren2_uops_1_is_unique),
    .io_ren2_uops_1_flush_on_commit(rename_stage_io_ren2_uops_1_flush_on_commit),
    .io_ren2_uops_1_ldst(rename_stage_io_ren2_uops_1_ldst),
    .io_ren2_uops_1_lrs1(rename_stage_io_ren2_uops_1_lrs1),
    .io_ren2_uops_1_lrs2(rename_stage_io_ren2_uops_1_lrs2),
    .io_ren2_uops_1_lrs3(rename_stage_io_ren2_uops_1_lrs3),
    .io_ren2_uops_1_ldst_val(rename_stage_io_ren2_uops_1_ldst_val),
    .io_ren2_uops_1_dst_rtype(rename_stage_io_ren2_uops_1_dst_rtype),
    .io_ren2_uops_1_lrs1_rtype(rename_stage_io_ren2_uops_1_lrs1_rtype),
    .io_ren2_uops_1_lrs2_rtype(rename_stage_io_ren2_uops_1_lrs2_rtype),
    .io_ren2_uops_1_frs3_en(rename_stage_io_ren2_uops_1_frs3_en),
    .io_ren2_uops_1_fp_val(rename_stage_io_ren2_uops_1_fp_val),
    .io_ren2_uops_1_fp_single(rename_stage_io_ren2_uops_1_fp_single),
    .io_ren2_uops_1_xcpt_pf_if(rename_stage_io_ren2_uops_1_xcpt_pf_if),
    .io_ren2_uops_1_xcpt_ae_if(rename_stage_io_ren2_uops_1_xcpt_ae_if),
    .io_ren2_uops_1_replay_if(rename_stage_io_ren2_uops_1_replay_if),
    .io_ren2_uops_1_xcpt_ma_if(rename_stage_io_ren2_uops_1_xcpt_ma_if),
    .io_ren2_uops_1_debug_wdata(rename_stage_io_ren2_uops_1_debug_wdata),
    .io_ren2_uops_1_debug_events_fetch_seq(rename_stage_io_ren2_uops_1_debug_events_fetch_seq),
    .io_ren_pred_info_0_bim_resp_value(rename_stage_io_ren_pred_info_0_bim_resp_value),
    .io_ren_pred_info_0_bim_resp_entry_idx(rename_stage_io_ren_pred_info_0_bim_resp_entry_idx),
    .io_ren_pred_info_0_bim_resp_way_idx(rename_stage_io_ren_pred_info_0_bim_resp_way_idx),
    .io_ren_pred_info_0_bpd_resp_history(rename_stage_io_ren_pred_info_0_bpd_resp_history),
    .io_ren_pred_info_0_bpd_resp_history_ptr(rename_stage_io_ren_pred_info_0_bpd_resp_history_ptr),
    .io_ren_pred_info_1_bim_resp_value(rename_stage_io_ren_pred_info_1_bim_resp_value),
    .io_ren_pred_info_1_bim_resp_entry_idx(rename_stage_io_ren_pred_info_1_bim_resp_entry_idx),
    .io_ren_pred_info_1_bim_resp_way_idx(rename_stage_io_ren_pred_info_1_bim_resp_way_idx),
    .io_ren_pred_info_1_bpd_resp_history(rename_stage_io_ren_pred_info_1_bpd_resp_history),
    .io_ren_pred_info_1_bpd_resp_history_ptr(rename_stage_io_ren_pred_info_1_bpd_resp_history_ptr),
    .io_brinfo_valid(rename_stage_io_brinfo_valid),
    .io_brinfo_mispredict(rename_stage_io_brinfo_mispredict),
    .io_brinfo_mask(rename_stage_io_brinfo_mask),
    .io_brinfo_tag(rename_stage_io_brinfo_tag),
    .io_get_pred_br_tag(rename_stage_io_get_pred_br_tag),
    .io_get_pred_info_bim_resp_value(rename_stage_io_get_pred_info_bim_resp_value),
    .io_get_pred_info_bim_resp_entry_idx(rename_stage_io_get_pred_info_bim_resp_entry_idx),
    .io_get_pred_info_bim_resp_way_idx(rename_stage_io_get_pred_info_bim_resp_way_idx),
    .io_get_pred_info_bpd_resp_history(rename_stage_io_get_pred_info_bpd_resp_history),
    .io_get_pred_info_bpd_resp_history_ptr(rename_stage_io_get_pred_info_bpd_resp_history_ptr),
    .io_dis_inst_can_proceed_0(rename_stage_io_dis_inst_can_proceed_0),
    .io_dis_inst_can_proceed_1(rename_stage_io_dis_inst_can_proceed_1),
    .io_int_wakeups_0_valid(rename_stage_io_int_wakeups_0_valid),
    .io_int_wakeups_0_bits_uop_pdst(rename_stage_io_int_wakeups_0_bits_uop_pdst),
    .io_int_wakeups_0_bits_uop_dst_rtype(rename_stage_io_int_wakeups_0_bits_uop_dst_rtype),
    .io_int_wakeups_1_valid(rename_stage_io_int_wakeups_1_valid),
    .io_int_wakeups_1_bits_uop_pdst(rename_stage_io_int_wakeups_1_bits_uop_pdst),
    .io_int_wakeups_1_bits_uop_dst_rtype(rename_stage_io_int_wakeups_1_bits_uop_dst_rtype),
    .io_int_wakeups_2_valid(rename_stage_io_int_wakeups_2_valid),
    .io_int_wakeups_2_bits_uop_pdst(rename_stage_io_int_wakeups_2_bits_uop_pdst),
    .io_int_wakeups_2_bits_uop_dst_rtype(rename_stage_io_int_wakeups_2_bits_uop_dst_rtype),
    .io_int_wakeups_3_valid(rename_stage_io_int_wakeups_3_valid),
    .io_int_wakeups_3_bits_uop_pdst(rename_stage_io_int_wakeups_3_bits_uop_pdst),
    .io_int_wakeups_3_bits_uop_dst_rtype(rename_stage_io_int_wakeups_3_bits_uop_dst_rtype),
    .io_int_wakeups_4_valid(rename_stage_io_int_wakeups_4_valid),
    .io_int_wakeups_4_bits_uop_pdst(rename_stage_io_int_wakeups_4_bits_uop_pdst),
    .io_int_wakeups_4_bits_uop_dst_rtype(rename_stage_io_int_wakeups_4_bits_uop_dst_rtype),
    .io_fp_wakeups_0_valid(rename_stage_io_fp_wakeups_0_valid),
    .io_fp_wakeups_0_bits_uop_pdst(rename_stage_io_fp_wakeups_0_bits_uop_pdst),
    .io_fp_wakeups_0_bits_uop_dst_rtype(rename_stage_io_fp_wakeups_0_bits_uop_dst_rtype),
    .io_fp_wakeups_1_valid(rename_stage_io_fp_wakeups_1_valid),
    .io_fp_wakeups_1_bits_uop_pdst(rename_stage_io_fp_wakeups_1_bits_uop_pdst),
    .io_fp_wakeups_1_bits_uop_dst_rtype(rename_stage_io_fp_wakeups_1_bits_uop_dst_rtype),
    .io_com_valids_0(rename_stage_io_com_valids_0),
    .io_com_valids_1(rename_stage_io_com_valids_1),
    .io_com_uops_0_pdst(rename_stage_io_com_uops_0_pdst),
    .io_com_uops_0_stale_pdst(rename_stage_io_com_uops_0_stale_pdst),
    .io_com_uops_0_ldst(rename_stage_io_com_uops_0_ldst),
    .io_com_uops_0_dst_rtype(rename_stage_io_com_uops_0_dst_rtype),
    .io_com_uops_1_pdst(rename_stage_io_com_uops_1_pdst),
    .io_com_uops_1_stale_pdst(rename_stage_io_com_uops_1_stale_pdst),
    .io_com_uops_1_ldst(rename_stage_io_com_uops_1_ldst),
    .io_com_uops_1_dst_rtype(rename_stage_io_com_uops_1_dst_rtype),
    .io_com_rbk_valids_0(rename_stage_io_com_rbk_valids_0),
    .io_com_rbk_valids_1(rename_stage_io_com_rbk_valids_1),
    .io_debug_rob_empty(rename_stage_io_debug_rob_empty)
  );
  IssueUnitCollasping_1 issue_units_0 (
    .clock(issue_units_0_clock),
    .reset(issue_units_0_reset),
    .io_dis_valids_0(issue_units_0_io_dis_valids_0),
    .io_dis_valids_1(issue_units_0_io_dis_valids_1),
    .io_dis_uops_0_valid(issue_units_0_io_dis_uops_0_valid),
    .io_dis_uops_0_uopc(issue_units_0_io_dis_uops_0_uopc),
    .io_dis_uops_0_inst(issue_units_0_io_dis_uops_0_inst),
    .io_dis_uops_0_pc(issue_units_0_io_dis_uops_0_pc),
    .io_dis_uops_0_iqtype(issue_units_0_io_dis_uops_0_iqtype),
    .io_dis_uops_0_fu_code(issue_units_0_io_dis_uops_0_fu_code),
    .io_dis_uops_0_allocate_brtag(issue_units_0_io_dis_uops_0_allocate_brtag),
    .io_dis_uops_0_is_br_or_jmp(issue_units_0_io_dis_uops_0_is_br_or_jmp),
    .io_dis_uops_0_is_jump(issue_units_0_io_dis_uops_0_is_jump),
    .io_dis_uops_0_is_jal(issue_units_0_io_dis_uops_0_is_jal),
    .io_dis_uops_0_is_ret(issue_units_0_io_dis_uops_0_is_ret),
    .io_dis_uops_0_is_call(issue_units_0_io_dis_uops_0_is_call),
    .io_dis_uops_0_br_mask(issue_units_0_io_dis_uops_0_br_mask),
    .io_dis_uops_0_br_tag(issue_units_0_io_dis_uops_0_br_tag),
    .io_dis_uops_0_br_prediction_btb_blame(issue_units_0_io_dis_uops_0_br_prediction_btb_blame),
    .io_dis_uops_0_br_prediction_btb_hit(issue_units_0_io_dis_uops_0_br_prediction_btb_hit),
    .io_dis_uops_0_br_prediction_btb_taken(issue_units_0_io_dis_uops_0_br_prediction_btb_taken),
    .io_dis_uops_0_br_prediction_bpd_blame(issue_units_0_io_dis_uops_0_br_prediction_bpd_blame),
    .io_dis_uops_0_br_prediction_bpd_hit(issue_units_0_io_dis_uops_0_br_prediction_bpd_hit),
    .io_dis_uops_0_br_prediction_bpd_taken(issue_units_0_io_dis_uops_0_br_prediction_bpd_taken),
    .io_dis_uops_0_br_prediction_bim_resp_value(issue_units_0_io_dis_uops_0_br_prediction_bim_resp_value),
    .io_dis_uops_0_br_prediction_bim_resp_entry_idx(issue_units_0_io_dis_uops_0_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_0_br_prediction_bim_resp_way_idx(issue_units_0_io_dis_uops_0_br_prediction_bim_resp_way_idx),
    .io_dis_uops_0_br_prediction_bpd_resp_takens(issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_takens),
    .io_dis_uops_0_br_prediction_bpd_resp_history(issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history),
    .io_dis_uops_0_br_prediction_bpd_resp_history_u(issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_u),
    .io_dis_uops_0_br_prediction_bpd_resp_history_ptr(issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_0_br_prediction_bpd_resp_info(issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_info),
    .io_dis_uops_0_stat_brjmp_mispredicted(issue_units_0_io_dis_uops_0_stat_brjmp_mispredicted),
    .io_dis_uops_0_stat_btb_made_pred(issue_units_0_io_dis_uops_0_stat_btb_made_pred),
    .io_dis_uops_0_stat_btb_mispredicted(issue_units_0_io_dis_uops_0_stat_btb_mispredicted),
    .io_dis_uops_0_stat_bpd_made_pred(issue_units_0_io_dis_uops_0_stat_bpd_made_pred),
    .io_dis_uops_0_stat_bpd_mispredicted(issue_units_0_io_dis_uops_0_stat_bpd_mispredicted),
    .io_dis_uops_0_fetch_pc_lob(issue_units_0_io_dis_uops_0_fetch_pc_lob),
    .io_dis_uops_0_imm_packed(issue_units_0_io_dis_uops_0_imm_packed),
    .io_dis_uops_0_csr_addr(issue_units_0_io_dis_uops_0_csr_addr),
    .io_dis_uops_0_rob_idx(issue_units_0_io_dis_uops_0_rob_idx),
    .io_dis_uops_0_ldq_idx(issue_units_0_io_dis_uops_0_ldq_idx),
    .io_dis_uops_0_stq_idx(issue_units_0_io_dis_uops_0_stq_idx),
    .io_dis_uops_0_brob_idx(issue_units_0_io_dis_uops_0_brob_idx),
    .io_dis_uops_0_pdst(issue_units_0_io_dis_uops_0_pdst),
    .io_dis_uops_0_pop1(issue_units_0_io_dis_uops_0_pop1),
    .io_dis_uops_0_pop2(issue_units_0_io_dis_uops_0_pop2),
    .io_dis_uops_0_pop3(issue_units_0_io_dis_uops_0_pop3),
    .io_dis_uops_0_prs1_busy(issue_units_0_io_dis_uops_0_prs1_busy),
    .io_dis_uops_0_prs2_busy(issue_units_0_io_dis_uops_0_prs2_busy),
    .io_dis_uops_0_prs3_busy(issue_units_0_io_dis_uops_0_prs3_busy),
    .io_dis_uops_0_stale_pdst(issue_units_0_io_dis_uops_0_stale_pdst),
    .io_dis_uops_0_exception(issue_units_0_io_dis_uops_0_exception),
    .io_dis_uops_0_exc_cause(issue_units_0_io_dis_uops_0_exc_cause),
    .io_dis_uops_0_bypassable(issue_units_0_io_dis_uops_0_bypassable),
    .io_dis_uops_0_mem_cmd(issue_units_0_io_dis_uops_0_mem_cmd),
    .io_dis_uops_0_mem_typ(issue_units_0_io_dis_uops_0_mem_typ),
    .io_dis_uops_0_is_fence(issue_units_0_io_dis_uops_0_is_fence),
    .io_dis_uops_0_is_fencei(issue_units_0_io_dis_uops_0_is_fencei),
    .io_dis_uops_0_is_store(issue_units_0_io_dis_uops_0_is_store),
    .io_dis_uops_0_is_amo(issue_units_0_io_dis_uops_0_is_amo),
    .io_dis_uops_0_is_load(issue_units_0_io_dis_uops_0_is_load),
    .io_dis_uops_0_is_sys_pc2epc(issue_units_0_io_dis_uops_0_is_sys_pc2epc),
    .io_dis_uops_0_is_unique(issue_units_0_io_dis_uops_0_is_unique),
    .io_dis_uops_0_flush_on_commit(issue_units_0_io_dis_uops_0_flush_on_commit),
    .io_dis_uops_0_ldst(issue_units_0_io_dis_uops_0_ldst),
    .io_dis_uops_0_lrs1(issue_units_0_io_dis_uops_0_lrs1),
    .io_dis_uops_0_lrs2(issue_units_0_io_dis_uops_0_lrs2),
    .io_dis_uops_0_lrs3(issue_units_0_io_dis_uops_0_lrs3),
    .io_dis_uops_0_ldst_val(issue_units_0_io_dis_uops_0_ldst_val),
    .io_dis_uops_0_dst_rtype(issue_units_0_io_dis_uops_0_dst_rtype),
    .io_dis_uops_0_lrs1_rtype(issue_units_0_io_dis_uops_0_lrs1_rtype),
    .io_dis_uops_0_lrs2_rtype(issue_units_0_io_dis_uops_0_lrs2_rtype),
    .io_dis_uops_0_frs3_en(issue_units_0_io_dis_uops_0_frs3_en),
    .io_dis_uops_0_fp_val(issue_units_0_io_dis_uops_0_fp_val),
    .io_dis_uops_0_fp_single(issue_units_0_io_dis_uops_0_fp_single),
    .io_dis_uops_0_xcpt_pf_if(issue_units_0_io_dis_uops_0_xcpt_pf_if),
    .io_dis_uops_0_xcpt_ae_if(issue_units_0_io_dis_uops_0_xcpt_ae_if),
    .io_dis_uops_0_replay_if(issue_units_0_io_dis_uops_0_replay_if),
    .io_dis_uops_0_xcpt_ma_if(issue_units_0_io_dis_uops_0_xcpt_ma_if),
    .io_dis_uops_0_debug_wdata(issue_units_0_io_dis_uops_0_debug_wdata),
    .io_dis_uops_0_debug_events_fetch_seq(issue_units_0_io_dis_uops_0_debug_events_fetch_seq),
    .io_dis_uops_1_valid(issue_units_0_io_dis_uops_1_valid),
    .io_dis_uops_1_uopc(issue_units_0_io_dis_uops_1_uopc),
    .io_dis_uops_1_inst(issue_units_0_io_dis_uops_1_inst),
    .io_dis_uops_1_pc(issue_units_0_io_dis_uops_1_pc),
    .io_dis_uops_1_iqtype(issue_units_0_io_dis_uops_1_iqtype),
    .io_dis_uops_1_fu_code(issue_units_0_io_dis_uops_1_fu_code),
    .io_dis_uops_1_allocate_brtag(issue_units_0_io_dis_uops_1_allocate_brtag),
    .io_dis_uops_1_is_br_or_jmp(issue_units_0_io_dis_uops_1_is_br_or_jmp),
    .io_dis_uops_1_is_jump(issue_units_0_io_dis_uops_1_is_jump),
    .io_dis_uops_1_is_jal(issue_units_0_io_dis_uops_1_is_jal),
    .io_dis_uops_1_is_ret(issue_units_0_io_dis_uops_1_is_ret),
    .io_dis_uops_1_is_call(issue_units_0_io_dis_uops_1_is_call),
    .io_dis_uops_1_br_mask(issue_units_0_io_dis_uops_1_br_mask),
    .io_dis_uops_1_br_tag(issue_units_0_io_dis_uops_1_br_tag),
    .io_dis_uops_1_br_prediction_btb_blame(issue_units_0_io_dis_uops_1_br_prediction_btb_blame),
    .io_dis_uops_1_br_prediction_btb_hit(issue_units_0_io_dis_uops_1_br_prediction_btb_hit),
    .io_dis_uops_1_br_prediction_btb_taken(issue_units_0_io_dis_uops_1_br_prediction_btb_taken),
    .io_dis_uops_1_br_prediction_bpd_blame(issue_units_0_io_dis_uops_1_br_prediction_bpd_blame),
    .io_dis_uops_1_br_prediction_bpd_hit(issue_units_0_io_dis_uops_1_br_prediction_bpd_hit),
    .io_dis_uops_1_br_prediction_bpd_taken(issue_units_0_io_dis_uops_1_br_prediction_bpd_taken),
    .io_dis_uops_1_br_prediction_bim_resp_value(issue_units_0_io_dis_uops_1_br_prediction_bim_resp_value),
    .io_dis_uops_1_br_prediction_bim_resp_entry_idx(issue_units_0_io_dis_uops_1_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_1_br_prediction_bim_resp_way_idx(issue_units_0_io_dis_uops_1_br_prediction_bim_resp_way_idx),
    .io_dis_uops_1_br_prediction_bpd_resp_takens(issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_takens),
    .io_dis_uops_1_br_prediction_bpd_resp_history(issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history),
    .io_dis_uops_1_br_prediction_bpd_resp_history_u(issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_u),
    .io_dis_uops_1_br_prediction_bpd_resp_history_ptr(issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_1_br_prediction_bpd_resp_info(issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_info),
    .io_dis_uops_1_stat_brjmp_mispredicted(issue_units_0_io_dis_uops_1_stat_brjmp_mispredicted),
    .io_dis_uops_1_stat_btb_made_pred(issue_units_0_io_dis_uops_1_stat_btb_made_pred),
    .io_dis_uops_1_stat_btb_mispredicted(issue_units_0_io_dis_uops_1_stat_btb_mispredicted),
    .io_dis_uops_1_stat_bpd_made_pred(issue_units_0_io_dis_uops_1_stat_bpd_made_pred),
    .io_dis_uops_1_stat_bpd_mispredicted(issue_units_0_io_dis_uops_1_stat_bpd_mispredicted),
    .io_dis_uops_1_fetch_pc_lob(issue_units_0_io_dis_uops_1_fetch_pc_lob),
    .io_dis_uops_1_imm_packed(issue_units_0_io_dis_uops_1_imm_packed),
    .io_dis_uops_1_csr_addr(issue_units_0_io_dis_uops_1_csr_addr),
    .io_dis_uops_1_rob_idx(issue_units_0_io_dis_uops_1_rob_idx),
    .io_dis_uops_1_ldq_idx(issue_units_0_io_dis_uops_1_ldq_idx),
    .io_dis_uops_1_stq_idx(issue_units_0_io_dis_uops_1_stq_idx),
    .io_dis_uops_1_brob_idx(issue_units_0_io_dis_uops_1_brob_idx),
    .io_dis_uops_1_pdst(issue_units_0_io_dis_uops_1_pdst),
    .io_dis_uops_1_pop1(issue_units_0_io_dis_uops_1_pop1),
    .io_dis_uops_1_pop2(issue_units_0_io_dis_uops_1_pop2),
    .io_dis_uops_1_pop3(issue_units_0_io_dis_uops_1_pop3),
    .io_dis_uops_1_prs1_busy(issue_units_0_io_dis_uops_1_prs1_busy),
    .io_dis_uops_1_prs2_busy(issue_units_0_io_dis_uops_1_prs2_busy),
    .io_dis_uops_1_prs3_busy(issue_units_0_io_dis_uops_1_prs3_busy),
    .io_dis_uops_1_stale_pdst(issue_units_0_io_dis_uops_1_stale_pdst),
    .io_dis_uops_1_exception(issue_units_0_io_dis_uops_1_exception),
    .io_dis_uops_1_exc_cause(issue_units_0_io_dis_uops_1_exc_cause),
    .io_dis_uops_1_bypassable(issue_units_0_io_dis_uops_1_bypassable),
    .io_dis_uops_1_mem_cmd(issue_units_0_io_dis_uops_1_mem_cmd),
    .io_dis_uops_1_mem_typ(issue_units_0_io_dis_uops_1_mem_typ),
    .io_dis_uops_1_is_fence(issue_units_0_io_dis_uops_1_is_fence),
    .io_dis_uops_1_is_fencei(issue_units_0_io_dis_uops_1_is_fencei),
    .io_dis_uops_1_is_store(issue_units_0_io_dis_uops_1_is_store),
    .io_dis_uops_1_is_amo(issue_units_0_io_dis_uops_1_is_amo),
    .io_dis_uops_1_is_load(issue_units_0_io_dis_uops_1_is_load),
    .io_dis_uops_1_is_sys_pc2epc(issue_units_0_io_dis_uops_1_is_sys_pc2epc),
    .io_dis_uops_1_is_unique(issue_units_0_io_dis_uops_1_is_unique),
    .io_dis_uops_1_flush_on_commit(issue_units_0_io_dis_uops_1_flush_on_commit),
    .io_dis_uops_1_ldst(issue_units_0_io_dis_uops_1_ldst),
    .io_dis_uops_1_lrs1(issue_units_0_io_dis_uops_1_lrs1),
    .io_dis_uops_1_lrs2(issue_units_0_io_dis_uops_1_lrs2),
    .io_dis_uops_1_lrs3(issue_units_0_io_dis_uops_1_lrs3),
    .io_dis_uops_1_ldst_val(issue_units_0_io_dis_uops_1_ldst_val),
    .io_dis_uops_1_dst_rtype(issue_units_0_io_dis_uops_1_dst_rtype),
    .io_dis_uops_1_lrs1_rtype(issue_units_0_io_dis_uops_1_lrs1_rtype),
    .io_dis_uops_1_lrs2_rtype(issue_units_0_io_dis_uops_1_lrs2_rtype),
    .io_dis_uops_1_frs3_en(issue_units_0_io_dis_uops_1_frs3_en),
    .io_dis_uops_1_fp_val(issue_units_0_io_dis_uops_1_fp_val),
    .io_dis_uops_1_fp_single(issue_units_0_io_dis_uops_1_fp_single),
    .io_dis_uops_1_xcpt_pf_if(issue_units_0_io_dis_uops_1_xcpt_pf_if),
    .io_dis_uops_1_xcpt_ae_if(issue_units_0_io_dis_uops_1_xcpt_ae_if),
    .io_dis_uops_1_replay_if(issue_units_0_io_dis_uops_1_replay_if),
    .io_dis_uops_1_xcpt_ma_if(issue_units_0_io_dis_uops_1_xcpt_ma_if),
    .io_dis_uops_1_debug_wdata(issue_units_0_io_dis_uops_1_debug_wdata),
    .io_dis_uops_1_debug_events_fetch_seq(issue_units_0_io_dis_uops_1_debug_events_fetch_seq),
    .io_dis_readys_0(issue_units_0_io_dis_readys_0),
    .io_dis_readys_1(issue_units_0_io_dis_readys_1),
    .io_iss_valids_0(issue_units_0_io_iss_valids_0),
    .io_iss_uops_0_uopc(issue_units_0_io_iss_uops_0_uopc),
    .io_iss_uops_0_br_mask(issue_units_0_io_iss_uops_0_br_mask),
    .io_iss_uops_0_imm_packed(issue_units_0_io_iss_uops_0_imm_packed),
    .io_iss_uops_0_rob_idx(issue_units_0_io_iss_uops_0_rob_idx),
    .io_iss_uops_0_ldq_idx(issue_units_0_io_iss_uops_0_ldq_idx),
    .io_iss_uops_0_stq_idx(issue_units_0_io_iss_uops_0_stq_idx),
    .io_iss_uops_0_pdst(issue_units_0_io_iss_uops_0_pdst),
    .io_iss_uops_0_pop1(issue_units_0_io_iss_uops_0_pop1),
    .io_iss_uops_0_pop2(issue_units_0_io_iss_uops_0_pop2),
    .io_iss_uops_0_mem_cmd(issue_units_0_io_iss_uops_0_mem_cmd),
    .io_iss_uops_0_mem_typ(issue_units_0_io_iss_uops_0_mem_typ),
    .io_iss_uops_0_is_fence(issue_units_0_io_iss_uops_0_is_fence),
    .io_iss_uops_0_is_store(issue_units_0_io_iss_uops_0_is_store),
    .io_iss_uops_0_is_amo(issue_units_0_io_iss_uops_0_is_amo),
    .io_iss_uops_0_is_load(issue_units_0_io_iss_uops_0_is_load),
    .io_iss_uops_0_dst_rtype(issue_units_0_io_iss_uops_0_dst_rtype),
    .io_iss_uops_0_lrs1_rtype(issue_units_0_io_iss_uops_0_lrs1_rtype),
    .io_iss_uops_0_lrs2_rtype(issue_units_0_io_iss_uops_0_lrs2_rtype),
    .io_iss_uops_0_fp_val(issue_units_0_io_iss_uops_0_fp_val),
    .io_wakeup_pdsts_0_valid(issue_units_0_io_wakeup_pdsts_0_valid),
    .io_wakeup_pdsts_0_bits(issue_units_0_io_wakeup_pdsts_0_bits),
    .io_wakeup_pdsts_1_valid(issue_units_0_io_wakeup_pdsts_1_valid),
    .io_wakeup_pdsts_1_bits(issue_units_0_io_wakeup_pdsts_1_bits),
    .io_wakeup_pdsts_2_valid(issue_units_0_io_wakeup_pdsts_2_valid),
    .io_wakeup_pdsts_2_bits(issue_units_0_io_wakeup_pdsts_2_bits),
    .io_wakeup_pdsts_3_valid(issue_units_0_io_wakeup_pdsts_3_valid),
    .io_wakeup_pdsts_3_bits(issue_units_0_io_wakeup_pdsts_3_bits),
    .io_wakeup_pdsts_4_valid(issue_units_0_io_wakeup_pdsts_4_valid),
    .io_wakeup_pdsts_4_bits(issue_units_0_io_wakeup_pdsts_4_bits),
    .io_brinfo_valid(issue_units_0_io_brinfo_valid),
    .io_brinfo_mispredict(issue_units_0_io_brinfo_mispredict),
    .io_brinfo_mask(issue_units_0_io_brinfo_mask),
    .io_flush_pipeline(issue_units_0_io_flush_pipeline)
  );
  IssueUnitCollasping_2 issue_units_1 (
    .clock(issue_units_1_clock),
    .reset(issue_units_1_reset),
    .io_dis_valids_0(issue_units_1_io_dis_valids_0),
    .io_dis_valids_1(issue_units_1_io_dis_valids_1),
    .io_dis_uops_0_valid(issue_units_1_io_dis_uops_0_valid),
    .io_dis_uops_0_uopc(issue_units_1_io_dis_uops_0_uopc),
    .io_dis_uops_0_inst(issue_units_1_io_dis_uops_0_inst),
    .io_dis_uops_0_pc(issue_units_1_io_dis_uops_0_pc),
    .io_dis_uops_0_iqtype(issue_units_1_io_dis_uops_0_iqtype),
    .io_dis_uops_0_fu_code(issue_units_1_io_dis_uops_0_fu_code),
    .io_dis_uops_0_allocate_brtag(issue_units_1_io_dis_uops_0_allocate_brtag),
    .io_dis_uops_0_is_br_or_jmp(issue_units_1_io_dis_uops_0_is_br_or_jmp),
    .io_dis_uops_0_is_jump(issue_units_1_io_dis_uops_0_is_jump),
    .io_dis_uops_0_is_jal(issue_units_1_io_dis_uops_0_is_jal),
    .io_dis_uops_0_is_ret(issue_units_1_io_dis_uops_0_is_ret),
    .io_dis_uops_0_is_call(issue_units_1_io_dis_uops_0_is_call),
    .io_dis_uops_0_br_mask(issue_units_1_io_dis_uops_0_br_mask),
    .io_dis_uops_0_br_tag(issue_units_1_io_dis_uops_0_br_tag),
    .io_dis_uops_0_br_prediction_btb_blame(issue_units_1_io_dis_uops_0_br_prediction_btb_blame),
    .io_dis_uops_0_br_prediction_btb_hit(issue_units_1_io_dis_uops_0_br_prediction_btb_hit),
    .io_dis_uops_0_br_prediction_btb_taken(issue_units_1_io_dis_uops_0_br_prediction_btb_taken),
    .io_dis_uops_0_br_prediction_bpd_blame(issue_units_1_io_dis_uops_0_br_prediction_bpd_blame),
    .io_dis_uops_0_br_prediction_bpd_hit(issue_units_1_io_dis_uops_0_br_prediction_bpd_hit),
    .io_dis_uops_0_br_prediction_bpd_taken(issue_units_1_io_dis_uops_0_br_prediction_bpd_taken),
    .io_dis_uops_0_br_prediction_bim_resp_value(issue_units_1_io_dis_uops_0_br_prediction_bim_resp_value),
    .io_dis_uops_0_br_prediction_bim_resp_entry_idx(issue_units_1_io_dis_uops_0_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_0_br_prediction_bim_resp_way_idx(issue_units_1_io_dis_uops_0_br_prediction_bim_resp_way_idx),
    .io_dis_uops_0_br_prediction_bpd_resp_takens(issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_takens),
    .io_dis_uops_0_br_prediction_bpd_resp_history(issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history),
    .io_dis_uops_0_br_prediction_bpd_resp_history_u(issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_u),
    .io_dis_uops_0_br_prediction_bpd_resp_history_ptr(issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_0_br_prediction_bpd_resp_info(issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_info),
    .io_dis_uops_0_stat_brjmp_mispredicted(issue_units_1_io_dis_uops_0_stat_brjmp_mispredicted),
    .io_dis_uops_0_stat_btb_made_pred(issue_units_1_io_dis_uops_0_stat_btb_made_pred),
    .io_dis_uops_0_stat_btb_mispredicted(issue_units_1_io_dis_uops_0_stat_btb_mispredicted),
    .io_dis_uops_0_stat_bpd_made_pred(issue_units_1_io_dis_uops_0_stat_bpd_made_pred),
    .io_dis_uops_0_stat_bpd_mispredicted(issue_units_1_io_dis_uops_0_stat_bpd_mispredicted),
    .io_dis_uops_0_fetch_pc_lob(issue_units_1_io_dis_uops_0_fetch_pc_lob),
    .io_dis_uops_0_imm_packed(issue_units_1_io_dis_uops_0_imm_packed),
    .io_dis_uops_0_csr_addr(issue_units_1_io_dis_uops_0_csr_addr),
    .io_dis_uops_0_rob_idx(issue_units_1_io_dis_uops_0_rob_idx),
    .io_dis_uops_0_ldq_idx(issue_units_1_io_dis_uops_0_ldq_idx),
    .io_dis_uops_0_stq_idx(issue_units_1_io_dis_uops_0_stq_idx),
    .io_dis_uops_0_brob_idx(issue_units_1_io_dis_uops_0_brob_idx),
    .io_dis_uops_0_pdst(issue_units_1_io_dis_uops_0_pdst),
    .io_dis_uops_0_pop1(issue_units_1_io_dis_uops_0_pop1),
    .io_dis_uops_0_pop2(issue_units_1_io_dis_uops_0_pop2),
    .io_dis_uops_0_pop3(issue_units_1_io_dis_uops_0_pop3),
    .io_dis_uops_0_prs1_busy(issue_units_1_io_dis_uops_0_prs1_busy),
    .io_dis_uops_0_prs2_busy(issue_units_1_io_dis_uops_0_prs2_busy),
    .io_dis_uops_0_prs3_busy(issue_units_1_io_dis_uops_0_prs3_busy),
    .io_dis_uops_0_stale_pdst(issue_units_1_io_dis_uops_0_stale_pdst),
    .io_dis_uops_0_exception(issue_units_1_io_dis_uops_0_exception),
    .io_dis_uops_0_exc_cause(issue_units_1_io_dis_uops_0_exc_cause),
    .io_dis_uops_0_bypassable(issue_units_1_io_dis_uops_0_bypassable),
    .io_dis_uops_0_mem_cmd(issue_units_1_io_dis_uops_0_mem_cmd),
    .io_dis_uops_0_mem_typ(issue_units_1_io_dis_uops_0_mem_typ),
    .io_dis_uops_0_is_fence(issue_units_1_io_dis_uops_0_is_fence),
    .io_dis_uops_0_is_fencei(issue_units_1_io_dis_uops_0_is_fencei),
    .io_dis_uops_0_is_store(issue_units_1_io_dis_uops_0_is_store),
    .io_dis_uops_0_is_amo(issue_units_1_io_dis_uops_0_is_amo),
    .io_dis_uops_0_is_load(issue_units_1_io_dis_uops_0_is_load),
    .io_dis_uops_0_is_sys_pc2epc(issue_units_1_io_dis_uops_0_is_sys_pc2epc),
    .io_dis_uops_0_is_unique(issue_units_1_io_dis_uops_0_is_unique),
    .io_dis_uops_0_flush_on_commit(issue_units_1_io_dis_uops_0_flush_on_commit),
    .io_dis_uops_0_ldst(issue_units_1_io_dis_uops_0_ldst),
    .io_dis_uops_0_lrs1(issue_units_1_io_dis_uops_0_lrs1),
    .io_dis_uops_0_lrs2(issue_units_1_io_dis_uops_0_lrs2),
    .io_dis_uops_0_lrs3(issue_units_1_io_dis_uops_0_lrs3),
    .io_dis_uops_0_ldst_val(issue_units_1_io_dis_uops_0_ldst_val),
    .io_dis_uops_0_dst_rtype(issue_units_1_io_dis_uops_0_dst_rtype),
    .io_dis_uops_0_lrs1_rtype(issue_units_1_io_dis_uops_0_lrs1_rtype),
    .io_dis_uops_0_lrs2_rtype(issue_units_1_io_dis_uops_0_lrs2_rtype),
    .io_dis_uops_0_frs3_en(issue_units_1_io_dis_uops_0_frs3_en),
    .io_dis_uops_0_fp_val(issue_units_1_io_dis_uops_0_fp_val),
    .io_dis_uops_0_fp_single(issue_units_1_io_dis_uops_0_fp_single),
    .io_dis_uops_0_xcpt_pf_if(issue_units_1_io_dis_uops_0_xcpt_pf_if),
    .io_dis_uops_0_xcpt_ae_if(issue_units_1_io_dis_uops_0_xcpt_ae_if),
    .io_dis_uops_0_replay_if(issue_units_1_io_dis_uops_0_replay_if),
    .io_dis_uops_0_xcpt_ma_if(issue_units_1_io_dis_uops_0_xcpt_ma_if),
    .io_dis_uops_0_debug_wdata(issue_units_1_io_dis_uops_0_debug_wdata),
    .io_dis_uops_0_debug_events_fetch_seq(issue_units_1_io_dis_uops_0_debug_events_fetch_seq),
    .io_dis_uops_1_valid(issue_units_1_io_dis_uops_1_valid),
    .io_dis_uops_1_uopc(issue_units_1_io_dis_uops_1_uopc),
    .io_dis_uops_1_inst(issue_units_1_io_dis_uops_1_inst),
    .io_dis_uops_1_pc(issue_units_1_io_dis_uops_1_pc),
    .io_dis_uops_1_iqtype(issue_units_1_io_dis_uops_1_iqtype),
    .io_dis_uops_1_fu_code(issue_units_1_io_dis_uops_1_fu_code),
    .io_dis_uops_1_allocate_brtag(issue_units_1_io_dis_uops_1_allocate_brtag),
    .io_dis_uops_1_is_br_or_jmp(issue_units_1_io_dis_uops_1_is_br_or_jmp),
    .io_dis_uops_1_is_jump(issue_units_1_io_dis_uops_1_is_jump),
    .io_dis_uops_1_is_jal(issue_units_1_io_dis_uops_1_is_jal),
    .io_dis_uops_1_is_ret(issue_units_1_io_dis_uops_1_is_ret),
    .io_dis_uops_1_is_call(issue_units_1_io_dis_uops_1_is_call),
    .io_dis_uops_1_br_mask(issue_units_1_io_dis_uops_1_br_mask),
    .io_dis_uops_1_br_tag(issue_units_1_io_dis_uops_1_br_tag),
    .io_dis_uops_1_br_prediction_btb_blame(issue_units_1_io_dis_uops_1_br_prediction_btb_blame),
    .io_dis_uops_1_br_prediction_btb_hit(issue_units_1_io_dis_uops_1_br_prediction_btb_hit),
    .io_dis_uops_1_br_prediction_btb_taken(issue_units_1_io_dis_uops_1_br_prediction_btb_taken),
    .io_dis_uops_1_br_prediction_bpd_blame(issue_units_1_io_dis_uops_1_br_prediction_bpd_blame),
    .io_dis_uops_1_br_prediction_bpd_hit(issue_units_1_io_dis_uops_1_br_prediction_bpd_hit),
    .io_dis_uops_1_br_prediction_bpd_taken(issue_units_1_io_dis_uops_1_br_prediction_bpd_taken),
    .io_dis_uops_1_br_prediction_bim_resp_value(issue_units_1_io_dis_uops_1_br_prediction_bim_resp_value),
    .io_dis_uops_1_br_prediction_bim_resp_entry_idx(issue_units_1_io_dis_uops_1_br_prediction_bim_resp_entry_idx),
    .io_dis_uops_1_br_prediction_bim_resp_way_idx(issue_units_1_io_dis_uops_1_br_prediction_bim_resp_way_idx),
    .io_dis_uops_1_br_prediction_bpd_resp_takens(issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_takens),
    .io_dis_uops_1_br_prediction_bpd_resp_history(issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history),
    .io_dis_uops_1_br_prediction_bpd_resp_history_u(issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_u),
    .io_dis_uops_1_br_prediction_bpd_resp_history_ptr(issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_dis_uops_1_br_prediction_bpd_resp_info(issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_info),
    .io_dis_uops_1_stat_brjmp_mispredicted(issue_units_1_io_dis_uops_1_stat_brjmp_mispredicted),
    .io_dis_uops_1_stat_btb_made_pred(issue_units_1_io_dis_uops_1_stat_btb_made_pred),
    .io_dis_uops_1_stat_btb_mispredicted(issue_units_1_io_dis_uops_1_stat_btb_mispredicted),
    .io_dis_uops_1_stat_bpd_made_pred(issue_units_1_io_dis_uops_1_stat_bpd_made_pred),
    .io_dis_uops_1_stat_bpd_mispredicted(issue_units_1_io_dis_uops_1_stat_bpd_mispredicted),
    .io_dis_uops_1_fetch_pc_lob(issue_units_1_io_dis_uops_1_fetch_pc_lob),
    .io_dis_uops_1_imm_packed(issue_units_1_io_dis_uops_1_imm_packed),
    .io_dis_uops_1_csr_addr(issue_units_1_io_dis_uops_1_csr_addr),
    .io_dis_uops_1_rob_idx(issue_units_1_io_dis_uops_1_rob_idx),
    .io_dis_uops_1_ldq_idx(issue_units_1_io_dis_uops_1_ldq_idx),
    .io_dis_uops_1_stq_idx(issue_units_1_io_dis_uops_1_stq_idx),
    .io_dis_uops_1_brob_idx(issue_units_1_io_dis_uops_1_brob_idx),
    .io_dis_uops_1_pdst(issue_units_1_io_dis_uops_1_pdst),
    .io_dis_uops_1_pop1(issue_units_1_io_dis_uops_1_pop1),
    .io_dis_uops_1_pop2(issue_units_1_io_dis_uops_1_pop2),
    .io_dis_uops_1_pop3(issue_units_1_io_dis_uops_1_pop3),
    .io_dis_uops_1_prs1_busy(issue_units_1_io_dis_uops_1_prs1_busy),
    .io_dis_uops_1_prs2_busy(issue_units_1_io_dis_uops_1_prs2_busy),
    .io_dis_uops_1_prs3_busy(issue_units_1_io_dis_uops_1_prs3_busy),
    .io_dis_uops_1_stale_pdst(issue_units_1_io_dis_uops_1_stale_pdst),
    .io_dis_uops_1_exception(issue_units_1_io_dis_uops_1_exception),
    .io_dis_uops_1_exc_cause(issue_units_1_io_dis_uops_1_exc_cause),
    .io_dis_uops_1_bypassable(issue_units_1_io_dis_uops_1_bypassable),
    .io_dis_uops_1_mem_cmd(issue_units_1_io_dis_uops_1_mem_cmd),
    .io_dis_uops_1_mem_typ(issue_units_1_io_dis_uops_1_mem_typ),
    .io_dis_uops_1_is_fence(issue_units_1_io_dis_uops_1_is_fence),
    .io_dis_uops_1_is_fencei(issue_units_1_io_dis_uops_1_is_fencei),
    .io_dis_uops_1_is_store(issue_units_1_io_dis_uops_1_is_store),
    .io_dis_uops_1_is_amo(issue_units_1_io_dis_uops_1_is_amo),
    .io_dis_uops_1_is_load(issue_units_1_io_dis_uops_1_is_load),
    .io_dis_uops_1_is_sys_pc2epc(issue_units_1_io_dis_uops_1_is_sys_pc2epc),
    .io_dis_uops_1_is_unique(issue_units_1_io_dis_uops_1_is_unique),
    .io_dis_uops_1_flush_on_commit(issue_units_1_io_dis_uops_1_flush_on_commit),
    .io_dis_uops_1_ldst(issue_units_1_io_dis_uops_1_ldst),
    .io_dis_uops_1_lrs1(issue_units_1_io_dis_uops_1_lrs1),
    .io_dis_uops_1_lrs2(issue_units_1_io_dis_uops_1_lrs2),
    .io_dis_uops_1_lrs3(issue_units_1_io_dis_uops_1_lrs3),
    .io_dis_uops_1_ldst_val(issue_units_1_io_dis_uops_1_ldst_val),
    .io_dis_uops_1_dst_rtype(issue_units_1_io_dis_uops_1_dst_rtype),
    .io_dis_uops_1_lrs1_rtype(issue_units_1_io_dis_uops_1_lrs1_rtype),
    .io_dis_uops_1_lrs2_rtype(issue_units_1_io_dis_uops_1_lrs2_rtype),
    .io_dis_uops_1_frs3_en(issue_units_1_io_dis_uops_1_frs3_en),
    .io_dis_uops_1_fp_val(issue_units_1_io_dis_uops_1_fp_val),
    .io_dis_uops_1_fp_single(issue_units_1_io_dis_uops_1_fp_single),
    .io_dis_uops_1_xcpt_pf_if(issue_units_1_io_dis_uops_1_xcpt_pf_if),
    .io_dis_uops_1_xcpt_ae_if(issue_units_1_io_dis_uops_1_xcpt_ae_if),
    .io_dis_uops_1_replay_if(issue_units_1_io_dis_uops_1_replay_if),
    .io_dis_uops_1_xcpt_ma_if(issue_units_1_io_dis_uops_1_xcpt_ma_if),
    .io_dis_uops_1_debug_wdata(issue_units_1_io_dis_uops_1_debug_wdata),
    .io_dis_uops_1_debug_events_fetch_seq(issue_units_1_io_dis_uops_1_debug_events_fetch_seq),
    .io_dis_readys_0(issue_units_1_io_dis_readys_0),
    .io_dis_readys_1(issue_units_1_io_dis_readys_1),
    .io_iss_valids_0(issue_units_1_io_iss_valids_0),
    .io_iss_valids_1(issue_units_1_io_iss_valids_1),
    .io_iss_uops_0_valid(issue_units_1_io_iss_uops_0_valid),
    .io_iss_uops_0_iw_state(issue_units_1_io_iss_uops_0_iw_state),
    .io_iss_uops_0_uopc(issue_units_1_io_iss_uops_0_uopc),
    .io_iss_uops_0_inst(issue_units_1_io_iss_uops_0_inst),
    .io_iss_uops_0_pc(issue_units_1_io_iss_uops_0_pc),
    .io_iss_uops_0_iqtype(issue_units_1_io_iss_uops_0_iqtype),
    .io_iss_uops_0_fu_code(issue_units_1_io_iss_uops_0_fu_code),
    .io_iss_uops_0_allocate_brtag(issue_units_1_io_iss_uops_0_allocate_brtag),
    .io_iss_uops_0_is_br_or_jmp(issue_units_1_io_iss_uops_0_is_br_or_jmp),
    .io_iss_uops_0_is_jump(issue_units_1_io_iss_uops_0_is_jump),
    .io_iss_uops_0_is_jal(issue_units_1_io_iss_uops_0_is_jal),
    .io_iss_uops_0_is_ret(issue_units_1_io_iss_uops_0_is_ret),
    .io_iss_uops_0_is_call(issue_units_1_io_iss_uops_0_is_call),
    .io_iss_uops_0_br_mask(issue_units_1_io_iss_uops_0_br_mask),
    .io_iss_uops_0_br_tag(issue_units_1_io_iss_uops_0_br_tag),
    .io_iss_uops_0_br_prediction_btb_blame(issue_units_1_io_iss_uops_0_br_prediction_btb_blame),
    .io_iss_uops_0_br_prediction_btb_hit(issue_units_1_io_iss_uops_0_br_prediction_btb_hit),
    .io_iss_uops_0_br_prediction_btb_taken(issue_units_1_io_iss_uops_0_br_prediction_btb_taken),
    .io_iss_uops_0_br_prediction_bpd_blame(issue_units_1_io_iss_uops_0_br_prediction_bpd_blame),
    .io_iss_uops_0_br_prediction_bpd_hit(issue_units_1_io_iss_uops_0_br_prediction_bpd_hit),
    .io_iss_uops_0_br_prediction_bpd_taken(issue_units_1_io_iss_uops_0_br_prediction_bpd_taken),
    .io_iss_uops_0_br_prediction_bim_resp_value(issue_units_1_io_iss_uops_0_br_prediction_bim_resp_value),
    .io_iss_uops_0_br_prediction_bim_resp_entry_idx(issue_units_1_io_iss_uops_0_br_prediction_bim_resp_entry_idx),
    .io_iss_uops_0_br_prediction_bim_resp_way_idx(issue_units_1_io_iss_uops_0_br_prediction_bim_resp_way_idx),
    .io_iss_uops_0_br_prediction_bpd_resp_takens(issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_takens),
    .io_iss_uops_0_br_prediction_bpd_resp_history(issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history),
    .io_iss_uops_0_br_prediction_bpd_resp_history_u(issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_u),
    .io_iss_uops_0_br_prediction_bpd_resp_history_ptr(issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_ptr),
    .io_iss_uops_0_br_prediction_bpd_resp_info(issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_info),
    .io_iss_uops_0_stat_brjmp_mispredicted(issue_units_1_io_iss_uops_0_stat_brjmp_mispredicted),
    .io_iss_uops_0_stat_btb_made_pred(issue_units_1_io_iss_uops_0_stat_btb_made_pred),
    .io_iss_uops_0_stat_btb_mispredicted(issue_units_1_io_iss_uops_0_stat_btb_mispredicted),
    .io_iss_uops_0_stat_bpd_made_pred(issue_units_1_io_iss_uops_0_stat_bpd_made_pred),
    .io_iss_uops_0_stat_bpd_mispredicted(issue_units_1_io_iss_uops_0_stat_bpd_mispredicted),
    .io_iss_uops_0_fetch_pc_lob(issue_units_1_io_iss_uops_0_fetch_pc_lob),
    .io_iss_uops_0_imm_packed(issue_units_1_io_iss_uops_0_imm_packed),
    .io_iss_uops_0_csr_addr(issue_units_1_io_iss_uops_0_csr_addr),
    .io_iss_uops_0_rob_idx(issue_units_1_io_iss_uops_0_rob_idx),
    .io_iss_uops_0_ldq_idx(issue_units_1_io_iss_uops_0_ldq_idx),
    .io_iss_uops_0_stq_idx(issue_units_1_io_iss_uops_0_stq_idx),
    .io_iss_uops_0_brob_idx(issue_units_1_io_iss_uops_0_brob_idx),
    .io_iss_uops_0_pdst(issue_units_1_io_iss_uops_0_pdst),
    .io_iss_uops_0_pop1(issue_units_1_io_iss_uops_0_pop1),
    .io_iss_uops_0_pop2(issue_units_1_io_iss_uops_0_pop2),
    .io_iss_uops_0_pop3(issue_units_1_io_iss_uops_0_pop3),
    .io_iss_uops_0_prs1_busy(issue_units_1_io_iss_uops_0_prs1_busy),
    .io_iss_uops_0_prs2_busy(issue_units_1_io_iss_uops_0_prs2_busy),
    .io_iss_uops_0_prs3_busy(issue_units_1_io_iss_uops_0_prs3_busy),
    .io_iss_uops_0_stale_pdst(issue_units_1_io_iss_uops_0_stale_pdst),
    .io_iss_uops_0_exception(issue_units_1_io_iss_uops_0_exception),
    .io_iss_uops_0_exc_cause(issue_units_1_io_iss_uops_0_exc_cause),
    .io_iss_uops_0_bypassable(issue_units_1_io_iss_uops_0_bypassable),
    .io_iss_uops_0_mem_cmd(issue_units_1_io_iss_uops_0_mem_cmd),
    .io_iss_uops_0_mem_typ(issue_units_1_io_iss_uops_0_mem_typ),
    .io_iss_uops_0_is_fence(issue_units_1_io_iss_uops_0_is_fence),
    .io_iss_uops_0_is_fencei(issue_units_1_io_iss_uops_0_is_fencei),
    .io_iss_uops_0_is_store(issue_units_1_io_iss_uops_0_is_store),
    .io_iss_uops_0_is_amo(issue_units_1_io_iss_uops_0_is_amo),
    .io_iss_uops_0_is_load(issue_units_1_io_iss_uops_0_is_load),
    .io_iss_uops_0_is_sys_pc2epc(issue_units_1_io_iss_uops_0_is_sys_pc2epc),
    .io_iss_uops_0_is_unique(issue_units_1_io_iss_uops_0_is_unique),
    .io_iss_uops_0_flush_on_commit(issue_units_1_io_iss_uops_0_flush_on_commit),
    .io_iss_uops_0_ldst(issue_units_1_io_iss_uops_0_ldst),
    .io_iss_uops_0_lrs1(issue_units_1_io_iss_uops_0_lrs1),
    .io_iss_uops_0_lrs2(issue_units_1_io_iss_uops_0_lrs2),
    .io_iss_uops_0_lrs3(issue_units_1_io_iss_uops_0_lrs3),
    .io_iss_uops_0_ldst_val(issue_units_1_io_iss_uops_0_ldst_val),
    .io_iss_uops_0_dst_rtype(issue_units_1_io_iss_uops_0_dst_rtype),
    .io_iss_uops_0_lrs1_rtype(issue_units_1_io_iss_uops_0_lrs1_rtype),
    .io_iss_uops_0_lrs2_rtype(issue_units_1_io_iss_uops_0_lrs2_rtype),
    .io_iss_uops_0_frs3_en(issue_units_1_io_iss_uops_0_frs3_en),
    .io_iss_uops_0_fp_val(issue_units_1_io_iss_uops_0_fp_val),
    .io_iss_uops_0_fp_single(issue_units_1_io_iss_uops_0_fp_single),
    .io_iss_uops_0_xcpt_pf_if(issue_units_1_io_iss_uops_0_xcpt_pf_if),
    .io_iss_uops_0_xcpt_ae_if(issue_units_1_io_iss_uops_0_xcpt_ae_if),
    .io_iss_uops_0_replay_if(issue_units_1_io_iss_uops_0_replay_if),
    .io_iss_uops_0_xcpt_ma_if(issue_units_1_io_iss_uops_0_xcpt_ma_if),
    .io_iss_uops_0_debug_wdata(issue_units_1_io_iss_uops_0_debug_wdata),
    .io_iss_uops_0_debug_events_fetch_seq(issue_units_1_io_iss_uops_0_debug_events_fetch_seq),
    .io_iss_uops_1_valid(issue_units_1_io_iss_uops_1_valid),
    .io_iss_uops_1_iw_state(issue_units_1_io_iss_uops_1_iw_state),
    .io_iss_uops_1_uopc(issue_units_1_io_iss_uops_1_uopc),
    .io_iss_uops_1_inst(issue_units_1_io_iss_uops_1_inst),
    .io_iss_uops_1_pc(issue_units_1_io_iss_uops_1_pc),
    .io_iss_uops_1_iqtype(issue_units_1_io_iss_uops_1_iqtype),
    .io_iss_uops_1_fu_code(issue_units_1_io_iss_uops_1_fu_code),
    .io_iss_uops_1_allocate_brtag(issue_units_1_io_iss_uops_1_allocate_brtag),
    .io_iss_uops_1_is_br_or_jmp(issue_units_1_io_iss_uops_1_is_br_or_jmp),
    .io_iss_uops_1_is_jump(issue_units_1_io_iss_uops_1_is_jump),
    .io_iss_uops_1_is_jal(issue_units_1_io_iss_uops_1_is_jal),
    .io_iss_uops_1_is_ret(issue_units_1_io_iss_uops_1_is_ret),
    .io_iss_uops_1_is_call(issue_units_1_io_iss_uops_1_is_call),
    .io_iss_uops_1_br_mask(issue_units_1_io_iss_uops_1_br_mask),
    .io_iss_uops_1_br_tag(issue_units_1_io_iss_uops_1_br_tag),
    .io_iss_uops_1_br_prediction_btb_blame(issue_units_1_io_iss_uops_1_br_prediction_btb_blame),
    .io_iss_uops_1_br_prediction_btb_hit(issue_units_1_io_iss_uops_1_br_prediction_btb_hit),
    .io_iss_uops_1_br_prediction_btb_taken(issue_units_1_io_iss_uops_1_br_prediction_btb_taken),
    .io_iss_uops_1_br_prediction_bpd_blame(issue_units_1_io_iss_uops_1_br_prediction_bpd_blame),
    .io_iss_uops_1_br_prediction_bpd_hit(issue_units_1_io_iss_uops_1_br_prediction_bpd_hit),
    .io_iss_uops_1_br_prediction_bpd_taken(issue_units_1_io_iss_uops_1_br_prediction_bpd_taken),
    .io_iss_uops_1_br_prediction_bim_resp_value(issue_units_1_io_iss_uops_1_br_prediction_bim_resp_value),
    .io_iss_uops_1_br_prediction_bim_resp_entry_idx(issue_units_1_io_iss_uops_1_br_prediction_bim_resp_entry_idx),
    .io_iss_uops_1_br_prediction_bim_resp_way_idx(issue_units_1_io_iss_uops_1_br_prediction_bim_resp_way_idx),
    .io_iss_uops_1_br_prediction_bpd_resp_takens(issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_takens),
    .io_iss_uops_1_br_prediction_bpd_resp_history(issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history),
    .io_iss_uops_1_br_prediction_bpd_resp_history_u(issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_u),
    .io_iss_uops_1_br_prediction_bpd_resp_history_ptr(issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_iss_uops_1_br_prediction_bpd_resp_info(issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_info),
    .io_iss_uops_1_stat_brjmp_mispredicted(issue_units_1_io_iss_uops_1_stat_brjmp_mispredicted),
    .io_iss_uops_1_stat_btb_made_pred(issue_units_1_io_iss_uops_1_stat_btb_made_pred),
    .io_iss_uops_1_stat_btb_mispredicted(issue_units_1_io_iss_uops_1_stat_btb_mispredicted),
    .io_iss_uops_1_stat_bpd_made_pred(issue_units_1_io_iss_uops_1_stat_bpd_made_pred),
    .io_iss_uops_1_stat_bpd_mispredicted(issue_units_1_io_iss_uops_1_stat_bpd_mispredicted),
    .io_iss_uops_1_fetch_pc_lob(issue_units_1_io_iss_uops_1_fetch_pc_lob),
    .io_iss_uops_1_imm_packed(issue_units_1_io_iss_uops_1_imm_packed),
    .io_iss_uops_1_csr_addr(issue_units_1_io_iss_uops_1_csr_addr),
    .io_iss_uops_1_rob_idx(issue_units_1_io_iss_uops_1_rob_idx),
    .io_iss_uops_1_ldq_idx(issue_units_1_io_iss_uops_1_ldq_idx),
    .io_iss_uops_1_stq_idx(issue_units_1_io_iss_uops_1_stq_idx),
    .io_iss_uops_1_brob_idx(issue_units_1_io_iss_uops_1_brob_idx),
    .io_iss_uops_1_pdst(issue_units_1_io_iss_uops_1_pdst),
    .io_iss_uops_1_pop1(issue_units_1_io_iss_uops_1_pop1),
    .io_iss_uops_1_pop2(issue_units_1_io_iss_uops_1_pop2),
    .io_iss_uops_1_pop3(issue_units_1_io_iss_uops_1_pop3),
    .io_iss_uops_1_prs1_busy(issue_units_1_io_iss_uops_1_prs1_busy),
    .io_iss_uops_1_prs2_busy(issue_units_1_io_iss_uops_1_prs2_busy),
    .io_iss_uops_1_prs3_busy(issue_units_1_io_iss_uops_1_prs3_busy),
    .io_iss_uops_1_stale_pdst(issue_units_1_io_iss_uops_1_stale_pdst),
    .io_iss_uops_1_exception(issue_units_1_io_iss_uops_1_exception),
    .io_iss_uops_1_exc_cause(issue_units_1_io_iss_uops_1_exc_cause),
    .io_iss_uops_1_bypassable(issue_units_1_io_iss_uops_1_bypassable),
    .io_iss_uops_1_mem_cmd(issue_units_1_io_iss_uops_1_mem_cmd),
    .io_iss_uops_1_mem_typ(issue_units_1_io_iss_uops_1_mem_typ),
    .io_iss_uops_1_is_fence(issue_units_1_io_iss_uops_1_is_fence),
    .io_iss_uops_1_is_fencei(issue_units_1_io_iss_uops_1_is_fencei),
    .io_iss_uops_1_is_store(issue_units_1_io_iss_uops_1_is_store),
    .io_iss_uops_1_is_amo(issue_units_1_io_iss_uops_1_is_amo),
    .io_iss_uops_1_is_load(issue_units_1_io_iss_uops_1_is_load),
    .io_iss_uops_1_is_sys_pc2epc(issue_units_1_io_iss_uops_1_is_sys_pc2epc),
    .io_iss_uops_1_is_unique(issue_units_1_io_iss_uops_1_is_unique),
    .io_iss_uops_1_flush_on_commit(issue_units_1_io_iss_uops_1_flush_on_commit),
    .io_iss_uops_1_ldst(issue_units_1_io_iss_uops_1_ldst),
    .io_iss_uops_1_lrs1(issue_units_1_io_iss_uops_1_lrs1),
    .io_iss_uops_1_lrs2(issue_units_1_io_iss_uops_1_lrs2),
    .io_iss_uops_1_lrs3(issue_units_1_io_iss_uops_1_lrs3),
    .io_iss_uops_1_ldst_val(issue_units_1_io_iss_uops_1_ldst_val),
    .io_iss_uops_1_dst_rtype(issue_units_1_io_iss_uops_1_dst_rtype),
    .io_iss_uops_1_lrs1_rtype(issue_units_1_io_iss_uops_1_lrs1_rtype),
    .io_iss_uops_1_lrs2_rtype(issue_units_1_io_iss_uops_1_lrs2_rtype),
    .io_iss_uops_1_frs3_en(issue_units_1_io_iss_uops_1_frs3_en),
    .io_iss_uops_1_fp_val(issue_units_1_io_iss_uops_1_fp_val),
    .io_iss_uops_1_fp_single(issue_units_1_io_iss_uops_1_fp_single),
    .io_iss_uops_1_xcpt_pf_if(issue_units_1_io_iss_uops_1_xcpt_pf_if),
    .io_iss_uops_1_xcpt_ae_if(issue_units_1_io_iss_uops_1_xcpt_ae_if),
    .io_iss_uops_1_replay_if(issue_units_1_io_iss_uops_1_replay_if),
    .io_iss_uops_1_xcpt_ma_if(issue_units_1_io_iss_uops_1_xcpt_ma_if),
    .io_iss_uops_1_debug_wdata(issue_units_1_io_iss_uops_1_debug_wdata),
    .io_iss_uops_1_debug_events_fetch_seq(issue_units_1_io_iss_uops_1_debug_events_fetch_seq),
    .io_wakeup_pdsts_0_valid(issue_units_1_io_wakeup_pdsts_0_valid),
    .io_wakeup_pdsts_0_bits(issue_units_1_io_wakeup_pdsts_0_bits),
    .io_wakeup_pdsts_1_valid(issue_units_1_io_wakeup_pdsts_1_valid),
    .io_wakeup_pdsts_1_bits(issue_units_1_io_wakeup_pdsts_1_bits),
    .io_wakeup_pdsts_2_valid(issue_units_1_io_wakeup_pdsts_2_valid),
    .io_wakeup_pdsts_2_bits(issue_units_1_io_wakeup_pdsts_2_bits),
    .io_wakeup_pdsts_3_valid(issue_units_1_io_wakeup_pdsts_3_valid),
    .io_wakeup_pdsts_3_bits(issue_units_1_io_wakeup_pdsts_3_bits),
    .io_wakeup_pdsts_4_valid(issue_units_1_io_wakeup_pdsts_4_valid),
    .io_wakeup_pdsts_4_bits(issue_units_1_io_wakeup_pdsts_4_bits),
    .io_fu_types_0(issue_units_1_io_fu_types_0),
    .io_brinfo_valid(issue_units_1_io_brinfo_valid),
    .io_brinfo_mispredict(issue_units_1_io_brinfo_mispredict),
    .io_brinfo_mask(issue_units_1_io_brinfo_mask),
    .io_flush_pipeline(issue_units_1_io_flush_pipeline)
  );
  RegisterFileBehavorial_1 iregfile (
    .clock(iregfile_clock),
    .io_read_ports_0_addr(iregfile_io_read_ports_0_addr),
    .io_read_ports_0_data(iregfile_io_read_ports_0_data),
    .io_read_ports_1_addr(iregfile_io_read_ports_1_addr),
    .io_read_ports_1_data(iregfile_io_read_ports_1_data),
    .io_read_ports_2_addr(iregfile_io_read_ports_2_addr),
    .io_read_ports_2_data(iregfile_io_read_ports_2_data),
    .io_read_ports_3_addr(iregfile_io_read_ports_3_addr),
    .io_read_ports_3_data(iregfile_io_read_ports_3_data),
    .io_read_ports_4_addr(iregfile_io_read_ports_4_addr),
    .io_read_ports_4_data(iregfile_io_read_ports_4_data),
    .io_read_ports_5_addr(iregfile_io_read_ports_5_addr),
    .io_read_ports_5_data(iregfile_io_read_ports_5_data),
    .io_write_ports_0_valid(iregfile_io_write_ports_0_valid),
    .io_write_ports_0_bits_addr(iregfile_io_write_ports_0_bits_addr),
    .io_write_ports_0_bits_data(iregfile_io_write_ports_0_bits_data),
    .io_write_ports_1_valid(iregfile_io_write_ports_1_valid),
    .io_write_ports_1_bits_addr(iregfile_io_write_ports_1_bits_addr),
    .io_write_ports_1_bits_data(iregfile_io_write_ports_1_bits_data),
    .io_write_ports_2_valid(iregfile_io_write_ports_2_valid),
    .io_write_ports_2_bits_addr(iregfile_io_write_ports_2_bits_addr),
    .io_write_ports_2_bits_data(iregfile_io_write_ports_2_bits_data)
  );
  Arbiter_13 ll_wbarb (
    .io_in_0_valid(ll_wbarb_io_in_0_valid),
    .io_in_0_bits_uop_rob_idx(ll_wbarb_io_in_0_bits_uop_rob_idx),
    .io_in_0_bits_uop_pdst(ll_wbarb_io_in_0_bits_uop_pdst),
    .io_in_0_bits_uop_is_store(ll_wbarb_io_in_0_bits_uop_is_store),
    .io_in_0_bits_uop_is_amo(ll_wbarb_io_in_0_bits_uop_is_amo),
    .io_in_0_bits_uop_dst_rtype(ll_wbarb_io_in_0_bits_uop_dst_rtype),
    .io_in_0_bits_data(ll_wbarb_io_in_0_bits_data),
    .io_in_1_ready(ll_wbarb_io_in_1_ready),
    .io_in_1_valid(ll_wbarb_io_in_1_valid),
    .io_in_1_bits_uop_rob_idx(ll_wbarb_io_in_1_bits_uop_rob_idx),
    .io_in_1_bits_uop_pdst(ll_wbarb_io_in_1_bits_uop_pdst),
    .io_in_1_bits_uop_is_store(ll_wbarb_io_in_1_bits_uop_is_store),
    .io_in_1_bits_uop_is_amo(ll_wbarb_io_in_1_bits_uop_is_amo),
    .io_in_1_bits_uop_dst_rtype(ll_wbarb_io_in_1_bits_uop_dst_rtype),
    .io_in_1_bits_data(ll_wbarb_io_in_1_bits_data),
    .io_out_ready(ll_wbarb_io_out_ready),
    .io_out_valid(ll_wbarb_io_out_valid),
    .io_out_bits_uop_rob_idx(ll_wbarb_io_out_bits_uop_rob_idx),
    .io_out_bits_uop_pdst(ll_wbarb_io_out_bits_uop_pdst),
    .io_out_bits_uop_is_store(ll_wbarb_io_out_bits_uop_is_store),
    .io_out_bits_uop_is_amo(ll_wbarb_io_out_bits_uop_is_amo),
    .io_out_bits_uop_dst_rtype(ll_wbarb_io_out_bits_uop_dst_rtype),
    .io_out_bits_data(ll_wbarb_io_out_bits_data)
  );
  RegisterRead_1 iregister_read (
    .clock(iregister_read_clock),
    .reset(iregister_read_reset),
    .io_iss_valids_0(iregister_read_io_iss_valids_0),
    .io_iss_valids_1(iregister_read_io_iss_valids_1),
    .io_iss_valids_2(iregister_read_io_iss_valids_2),
    .io_iss_uops_0_uopc(iregister_read_io_iss_uops_0_uopc),
    .io_iss_uops_0_br_mask(iregister_read_io_iss_uops_0_br_mask),
    .io_iss_uops_0_imm_packed(iregister_read_io_iss_uops_0_imm_packed),
    .io_iss_uops_0_rob_idx(iregister_read_io_iss_uops_0_rob_idx),
    .io_iss_uops_0_ldq_idx(iregister_read_io_iss_uops_0_ldq_idx),
    .io_iss_uops_0_stq_idx(iregister_read_io_iss_uops_0_stq_idx),
    .io_iss_uops_0_pdst(iregister_read_io_iss_uops_0_pdst),
    .io_iss_uops_0_pop1(iregister_read_io_iss_uops_0_pop1),
    .io_iss_uops_0_pop2(iregister_read_io_iss_uops_0_pop2),
    .io_iss_uops_0_mem_cmd(iregister_read_io_iss_uops_0_mem_cmd),
    .io_iss_uops_0_mem_typ(iregister_read_io_iss_uops_0_mem_typ),
    .io_iss_uops_0_is_fence(iregister_read_io_iss_uops_0_is_fence),
    .io_iss_uops_0_is_store(iregister_read_io_iss_uops_0_is_store),
    .io_iss_uops_0_is_amo(iregister_read_io_iss_uops_0_is_amo),
    .io_iss_uops_0_is_load(iregister_read_io_iss_uops_0_is_load),
    .io_iss_uops_0_dst_rtype(iregister_read_io_iss_uops_0_dst_rtype),
    .io_iss_uops_0_lrs1_rtype(iregister_read_io_iss_uops_0_lrs1_rtype),
    .io_iss_uops_0_lrs2_rtype(iregister_read_io_iss_uops_0_lrs2_rtype),
    .io_iss_uops_0_fp_val(iregister_read_io_iss_uops_0_fp_val),
    .io_iss_uops_1_valid(iregister_read_io_iss_uops_1_valid),
    .io_iss_uops_1_iw_state(iregister_read_io_iss_uops_1_iw_state),
    .io_iss_uops_1_uopc(iregister_read_io_iss_uops_1_uopc),
    .io_iss_uops_1_inst(iregister_read_io_iss_uops_1_inst),
    .io_iss_uops_1_pc(iregister_read_io_iss_uops_1_pc),
    .io_iss_uops_1_iqtype(iregister_read_io_iss_uops_1_iqtype),
    .io_iss_uops_1_fu_code(iregister_read_io_iss_uops_1_fu_code),
    .io_iss_uops_1_allocate_brtag(iregister_read_io_iss_uops_1_allocate_brtag),
    .io_iss_uops_1_is_br_or_jmp(iregister_read_io_iss_uops_1_is_br_or_jmp),
    .io_iss_uops_1_is_jump(iregister_read_io_iss_uops_1_is_jump),
    .io_iss_uops_1_is_jal(iregister_read_io_iss_uops_1_is_jal),
    .io_iss_uops_1_is_ret(iregister_read_io_iss_uops_1_is_ret),
    .io_iss_uops_1_is_call(iregister_read_io_iss_uops_1_is_call),
    .io_iss_uops_1_br_mask(iregister_read_io_iss_uops_1_br_mask),
    .io_iss_uops_1_br_tag(iregister_read_io_iss_uops_1_br_tag),
    .io_iss_uops_1_br_prediction_btb_blame(iregister_read_io_iss_uops_1_br_prediction_btb_blame),
    .io_iss_uops_1_br_prediction_btb_hit(iregister_read_io_iss_uops_1_br_prediction_btb_hit),
    .io_iss_uops_1_br_prediction_btb_taken(iregister_read_io_iss_uops_1_br_prediction_btb_taken),
    .io_iss_uops_1_br_prediction_bpd_blame(iregister_read_io_iss_uops_1_br_prediction_bpd_blame),
    .io_iss_uops_1_br_prediction_bpd_hit(iregister_read_io_iss_uops_1_br_prediction_bpd_hit),
    .io_iss_uops_1_br_prediction_bpd_taken(iregister_read_io_iss_uops_1_br_prediction_bpd_taken),
    .io_iss_uops_1_br_prediction_bim_resp_value(iregister_read_io_iss_uops_1_br_prediction_bim_resp_value),
    .io_iss_uops_1_br_prediction_bim_resp_entry_idx(iregister_read_io_iss_uops_1_br_prediction_bim_resp_entry_idx),
    .io_iss_uops_1_br_prediction_bim_resp_way_idx(iregister_read_io_iss_uops_1_br_prediction_bim_resp_way_idx),
    .io_iss_uops_1_br_prediction_bpd_resp_takens(iregister_read_io_iss_uops_1_br_prediction_bpd_resp_takens),
    .io_iss_uops_1_br_prediction_bpd_resp_history(iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history),
    .io_iss_uops_1_br_prediction_bpd_resp_history_u(iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_u),
    .io_iss_uops_1_br_prediction_bpd_resp_history_ptr(iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_ptr),
    .io_iss_uops_1_br_prediction_bpd_resp_info(iregister_read_io_iss_uops_1_br_prediction_bpd_resp_info),
    .io_iss_uops_1_stat_brjmp_mispredicted(iregister_read_io_iss_uops_1_stat_brjmp_mispredicted),
    .io_iss_uops_1_stat_btb_made_pred(iregister_read_io_iss_uops_1_stat_btb_made_pred),
    .io_iss_uops_1_stat_btb_mispredicted(iregister_read_io_iss_uops_1_stat_btb_mispredicted),
    .io_iss_uops_1_stat_bpd_made_pred(iregister_read_io_iss_uops_1_stat_bpd_made_pred),
    .io_iss_uops_1_stat_bpd_mispredicted(iregister_read_io_iss_uops_1_stat_bpd_mispredicted),
    .io_iss_uops_1_fetch_pc_lob(iregister_read_io_iss_uops_1_fetch_pc_lob),
    .io_iss_uops_1_imm_packed(iregister_read_io_iss_uops_1_imm_packed),
    .io_iss_uops_1_csr_addr(iregister_read_io_iss_uops_1_csr_addr),
    .io_iss_uops_1_rob_idx(iregister_read_io_iss_uops_1_rob_idx),
    .io_iss_uops_1_ldq_idx(iregister_read_io_iss_uops_1_ldq_idx),
    .io_iss_uops_1_stq_idx(iregister_read_io_iss_uops_1_stq_idx),
    .io_iss_uops_1_brob_idx(iregister_read_io_iss_uops_1_brob_idx),
    .io_iss_uops_1_pdst(iregister_read_io_iss_uops_1_pdst),
    .io_iss_uops_1_pop1(iregister_read_io_iss_uops_1_pop1),
    .io_iss_uops_1_pop2(iregister_read_io_iss_uops_1_pop2),
    .io_iss_uops_1_pop3(iregister_read_io_iss_uops_1_pop3),
    .io_iss_uops_1_prs1_busy(iregister_read_io_iss_uops_1_prs1_busy),
    .io_iss_uops_1_prs2_busy(iregister_read_io_iss_uops_1_prs2_busy),
    .io_iss_uops_1_prs3_busy(iregister_read_io_iss_uops_1_prs3_busy),
    .io_iss_uops_1_stale_pdst(iregister_read_io_iss_uops_1_stale_pdst),
    .io_iss_uops_1_exception(iregister_read_io_iss_uops_1_exception),
    .io_iss_uops_1_exc_cause(iregister_read_io_iss_uops_1_exc_cause),
    .io_iss_uops_1_bypassable(iregister_read_io_iss_uops_1_bypassable),
    .io_iss_uops_1_mem_cmd(iregister_read_io_iss_uops_1_mem_cmd),
    .io_iss_uops_1_mem_typ(iregister_read_io_iss_uops_1_mem_typ),
    .io_iss_uops_1_is_fence(iregister_read_io_iss_uops_1_is_fence),
    .io_iss_uops_1_is_fencei(iregister_read_io_iss_uops_1_is_fencei),
    .io_iss_uops_1_is_store(iregister_read_io_iss_uops_1_is_store),
    .io_iss_uops_1_is_amo(iregister_read_io_iss_uops_1_is_amo),
    .io_iss_uops_1_is_load(iregister_read_io_iss_uops_1_is_load),
    .io_iss_uops_1_is_sys_pc2epc(iregister_read_io_iss_uops_1_is_sys_pc2epc),
    .io_iss_uops_1_is_unique(iregister_read_io_iss_uops_1_is_unique),
    .io_iss_uops_1_flush_on_commit(iregister_read_io_iss_uops_1_flush_on_commit),
    .io_iss_uops_1_ldst(iregister_read_io_iss_uops_1_ldst),
    .io_iss_uops_1_lrs1(iregister_read_io_iss_uops_1_lrs1),
    .io_iss_uops_1_lrs2(iregister_read_io_iss_uops_1_lrs2),
    .io_iss_uops_1_lrs3(iregister_read_io_iss_uops_1_lrs3),
    .io_iss_uops_1_ldst_val(iregister_read_io_iss_uops_1_ldst_val),
    .io_iss_uops_1_dst_rtype(iregister_read_io_iss_uops_1_dst_rtype),
    .io_iss_uops_1_lrs1_rtype(iregister_read_io_iss_uops_1_lrs1_rtype),
    .io_iss_uops_1_lrs2_rtype(iregister_read_io_iss_uops_1_lrs2_rtype),
    .io_iss_uops_1_frs3_en(iregister_read_io_iss_uops_1_frs3_en),
    .io_iss_uops_1_fp_val(iregister_read_io_iss_uops_1_fp_val),
    .io_iss_uops_1_fp_single(iregister_read_io_iss_uops_1_fp_single),
    .io_iss_uops_1_xcpt_pf_if(iregister_read_io_iss_uops_1_xcpt_pf_if),
    .io_iss_uops_1_xcpt_ae_if(iregister_read_io_iss_uops_1_xcpt_ae_if),
    .io_iss_uops_1_replay_if(iregister_read_io_iss_uops_1_replay_if),
    .io_iss_uops_1_xcpt_ma_if(iregister_read_io_iss_uops_1_xcpt_ma_if),
    .io_iss_uops_1_debug_wdata(iregister_read_io_iss_uops_1_debug_wdata),
    .io_iss_uops_1_debug_events_fetch_seq(iregister_read_io_iss_uops_1_debug_events_fetch_seq),
    .io_iss_uops_2_valid(iregister_read_io_iss_uops_2_valid),
    .io_iss_uops_2_iw_state(iregister_read_io_iss_uops_2_iw_state),
    .io_iss_uops_2_uopc(iregister_read_io_iss_uops_2_uopc),
    .io_iss_uops_2_inst(iregister_read_io_iss_uops_2_inst),
    .io_iss_uops_2_pc(iregister_read_io_iss_uops_2_pc),
    .io_iss_uops_2_iqtype(iregister_read_io_iss_uops_2_iqtype),
    .io_iss_uops_2_fu_code(iregister_read_io_iss_uops_2_fu_code),
    .io_iss_uops_2_allocate_brtag(iregister_read_io_iss_uops_2_allocate_brtag),
    .io_iss_uops_2_is_br_or_jmp(iregister_read_io_iss_uops_2_is_br_or_jmp),
    .io_iss_uops_2_is_jump(iregister_read_io_iss_uops_2_is_jump),
    .io_iss_uops_2_is_jal(iregister_read_io_iss_uops_2_is_jal),
    .io_iss_uops_2_is_ret(iregister_read_io_iss_uops_2_is_ret),
    .io_iss_uops_2_is_call(iregister_read_io_iss_uops_2_is_call),
    .io_iss_uops_2_br_mask(iregister_read_io_iss_uops_2_br_mask),
    .io_iss_uops_2_br_tag(iregister_read_io_iss_uops_2_br_tag),
    .io_iss_uops_2_br_prediction_btb_blame(iregister_read_io_iss_uops_2_br_prediction_btb_blame),
    .io_iss_uops_2_br_prediction_btb_hit(iregister_read_io_iss_uops_2_br_prediction_btb_hit),
    .io_iss_uops_2_br_prediction_btb_taken(iregister_read_io_iss_uops_2_br_prediction_btb_taken),
    .io_iss_uops_2_br_prediction_bpd_blame(iregister_read_io_iss_uops_2_br_prediction_bpd_blame),
    .io_iss_uops_2_br_prediction_bpd_hit(iregister_read_io_iss_uops_2_br_prediction_bpd_hit),
    .io_iss_uops_2_br_prediction_bpd_taken(iregister_read_io_iss_uops_2_br_prediction_bpd_taken),
    .io_iss_uops_2_br_prediction_bim_resp_value(iregister_read_io_iss_uops_2_br_prediction_bim_resp_value),
    .io_iss_uops_2_br_prediction_bim_resp_entry_idx(iregister_read_io_iss_uops_2_br_prediction_bim_resp_entry_idx),
    .io_iss_uops_2_br_prediction_bim_resp_way_idx(iregister_read_io_iss_uops_2_br_prediction_bim_resp_way_idx),
    .io_iss_uops_2_br_prediction_bpd_resp_takens(iregister_read_io_iss_uops_2_br_prediction_bpd_resp_takens),
    .io_iss_uops_2_br_prediction_bpd_resp_history(iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history),
    .io_iss_uops_2_br_prediction_bpd_resp_history_u(iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_u),
    .io_iss_uops_2_br_prediction_bpd_resp_history_ptr(iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_ptr),
    .io_iss_uops_2_br_prediction_bpd_resp_info(iregister_read_io_iss_uops_2_br_prediction_bpd_resp_info),
    .io_iss_uops_2_stat_brjmp_mispredicted(iregister_read_io_iss_uops_2_stat_brjmp_mispredicted),
    .io_iss_uops_2_stat_btb_made_pred(iregister_read_io_iss_uops_2_stat_btb_made_pred),
    .io_iss_uops_2_stat_btb_mispredicted(iregister_read_io_iss_uops_2_stat_btb_mispredicted),
    .io_iss_uops_2_stat_bpd_made_pred(iregister_read_io_iss_uops_2_stat_bpd_made_pred),
    .io_iss_uops_2_stat_bpd_mispredicted(iregister_read_io_iss_uops_2_stat_bpd_mispredicted),
    .io_iss_uops_2_fetch_pc_lob(iregister_read_io_iss_uops_2_fetch_pc_lob),
    .io_iss_uops_2_imm_packed(iregister_read_io_iss_uops_2_imm_packed),
    .io_iss_uops_2_csr_addr(iregister_read_io_iss_uops_2_csr_addr),
    .io_iss_uops_2_rob_idx(iregister_read_io_iss_uops_2_rob_idx),
    .io_iss_uops_2_ldq_idx(iregister_read_io_iss_uops_2_ldq_idx),
    .io_iss_uops_2_stq_idx(iregister_read_io_iss_uops_2_stq_idx),
    .io_iss_uops_2_brob_idx(iregister_read_io_iss_uops_2_brob_idx),
    .io_iss_uops_2_pdst(iregister_read_io_iss_uops_2_pdst),
    .io_iss_uops_2_pop1(iregister_read_io_iss_uops_2_pop1),
    .io_iss_uops_2_pop2(iregister_read_io_iss_uops_2_pop2),
    .io_iss_uops_2_pop3(iregister_read_io_iss_uops_2_pop3),
    .io_iss_uops_2_prs1_busy(iregister_read_io_iss_uops_2_prs1_busy),
    .io_iss_uops_2_prs2_busy(iregister_read_io_iss_uops_2_prs2_busy),
    .io_iss_uops_2_prs3_busy(iregister_read_io_iss_uops_2_prs3_busy),
    .io_iss_uops_2_stale_pdst(iregister_read_io_iss_uops_2_stale_pdst),
    .io_iss_uops_2_exception(iregister_read_io_iss_uops_2_exception),
    .io_iss_uops_2_exc_cause(iregister_read_io_iss_uops_2_exc_cause),
    .io_iss_uops_2_bypassable(iregister_read_io_iss_uops_2_bypassable),
    .io_iss_uops_2_mem_cmd(iregister_read_io_iss_uops_2_mem_cmd),
    .io_iss_uops_2_mem_typ(iregister_read_io_iss_uops_2_mem_typ),
    .io_iss_uops_2_is_fence(iregister_read_io_iss_uops_2_is_fence),
    .io_iss_uops_2_is_fencei(iregister_read_io_iss_uops_2_is_fencei),
    .io_iss_uops_2_is_store(iregister_read_io_iss_uops_2_is_store),
    .io_iss_uops_2_is_amo(iregister_read_io_iss_uops_2_is_amo),
    .io_iss_uops_2_is_load(iregister_read_io_iss_uops_2_is_load),
    .io_iss_uops_2_is_sys_pc2epc(iregister_read_io_iss_uops_2_is_sys_pc2epc),
    .io_iss_uops_2_is_unique(iregister_read_io_iss_uops_2_is_unique),
    .io_iss_uops_2_flush_on_commit(iregister_read_io_iss_uops_2_flush_on_commit),
    .io_iss_uops_2_ldst(iregister_read_io_iss_uops_2_ldst),
    .io_iss_uops_2_lrs1(iregister_read_io_iss_uops_2_lrs1),
    .io_iss_uops_2_lrs2(iregister_read_io_iss_uops_2_lrs2),
    .io_iss_uops_2_lrs3(iregister_read_io_iss_uops_2_lrs3),
    .io_iss_uops_2_ldst_val(iregister_read_io_iss_uops_2_ldst_val),
    .io_iss_uops_2_dst_rtype(iregister_read_io_iss_uops_2_dst_rtype),
    .io_iss_uops_2_lrs1_rtype(iregister_read_io_iss_uops_2_lrs1_rtype),
    .io_iss_uops_2_lrs2_rtype(iregister_read_io_iss_uops_2_lrs2_rtype),
    .io_iss_uops_2_frs3_en(iregister_read_io_iss_uops_2_frs3_en),
    .io_iss_uops_2_fp_val(iregister_read_io_iss_uops_2_fp_val),
    .io_iss_uops_2_fp_single(iregister_read_io_iss_uops_2_fp_single),
    .io_iss_uops_2_xcpt_pf_if(iregister_read_io_iss_uops_2_xcpt_pf_if),
    .io_iss_uops_2_xcpt_ae_if(iregister_read_io_iss_uops_2_xcpt_ae_if),
    .io_iss_uops_2_replay_if(iregister_read_io_iss_uops_2_replay_if),
    .io_iss_uops_2_xcpt_ma_if(iregister_read_io_iss_uops_2_xcpt_ma_if),
    .io_iss_uops_2_debug_wdata(iregister_read_io_iss_uops_2_debug_wdata),
    .io_iss_uops_2_debug_events_fetch_seq(iregister_read_io_iss_uops_2_debug_events_fetch_seq),
    .io_rf_read_ports_0_addr(iregister_read_io_rf_read_ports_0_addr),
    .io_rf_read_ports_0_data(iregister_read_io_rf_read_ports_0_data),
    .io_rf_read_ports_1_addr(iregister_read_io_rf_read_ports_1_addr),
    .io_rf_read_ports_1_data(iregister_read_io_rf_read_ports_1_data),
    .io_rf_read_ports_2_addr(iregister_read_io_rf_read_ports_2_addr),
    .io_rf_read_ports_2_data(iregister_read_io_rf_read_ports_2_data),
    .io_rf_read_ports_3_addr(iregister_read_io_rf_read_ports_3_addr),
    .io_rf_read_ports_3_data(iregister_read_io_rf_read_ports_3_data),
    .io_rf_read_ports_4_addr(iregister_read_io_rf_read_ports_4_addr),
    .io_rf_read_ports_4_data(iregister_read_io_rf_read_ports_4_data),
    .io_rf_read_ports_5_addr(iregister_read_io_rf_read_ports_5_addr),
    .io_rf_read_ports_5_data(iregister_read_io_rf_read_ports_5_data),
    .io_bypass_valid_0(iregister_read_io_bypass_valid_0),
    .io_bypass_valid_1(iregister_read_io_bypass_valid_1),
    .io_bypass_valid_2(iregister_read_io_bypass_valid_2),
    .io_bypass_valid_3(iregister_read_io_bypass_valid_3),
    .io_bypass_uop_0_ctrl_rf_wen(iregister_read_io_bypass_uop_0_ctrl_rf_wen),
    .io_bypass_uop_0_pdst(iregister_read_io_bypass_uop_0_pdst),
    .io_bypass_uop_0_dst_rtype(iregister_read_io_bypass_uop_0_dst_rtype),
    .io_bypass_uop_1_ctrl_rf_wen(iregister_read_io_bypass_uop_1_ctrl_rf_wen),
    .io_bypass_uop_1_pdst(iregister_read_io_bypass_uop_1_pdst),
    .io_bypass_uop_1_dst_rtype(iregister_read_io_bypass_uop_1_dst_rtype),
    .io_bypass_uop_2_ctrl_rf_wen(iregister_read_io_bypass_uop_2_ctrl_rf_wen),
    .io_bypass_uop_2_pdst(iregister_read_io_bypass_uop_2_pdst),
    .io_bypass_uop_2_dst_rtype(iregister_read_io_bypass_uop_2_dst_rtype),
    .io_bypass_uop_3_ctrl_rf_wen(iregister_read_io_bypass_uop_3_ctrl_rf_wen),
    .io_bypass_uop_3_pdst(iregister_read_io_bypass_uop_3_pdst),
    .io_bypass_uop_3_dst_rtype(iregister_read_io_bypass_uop_3_dst_rtype),
    .io_bypass_data_0(iregister_read_io_bypass_data_0),
    .io_bypass_data_1(iregister_read_io_bypass_data_1),
    .io_bypass_data_2(iregister_read_io_bypass_data_2),
    .io_bypass_data_3(iregister_read_io_bypass_data_3),
    .io_exe_reqs_0_valid(iregister_read_io_exe_reqs_0_valid),
    .io_exe_reqs_0_bits_uop_uopc(iregister_read_io_exe_reqs_0_bits_uop_uopc),
    .io_exe_reqs_0_bits_uop_ctrl_is_load(iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_load),
    .io_exe_reqs_0_bits_uop_ctrl_is_sta(iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_sta),
    .io_exe_reqs_0_bits_uop_ctrl_is_std(iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_std),
    .io_exe_reqs_0_bits_uop_br_mask(iregister_read_io_exe_reqs_0_bits_uop_br_mask),
    .io_exe_reqs_0_bits_uop_imm_packed(iregister_read_io_exe_reqs_0_bits_uop_imm_packed),
    .io_exe_reqs_0_bits_uop_rob_idx(iregister_read_io_exe_reqs_0_bits_uop_rob_idx),
    .io_exe_reqs_0_bits_uop_ldq_idx(iregister_read_io_exe_reqs_0_bits_uop_ldq_idx),
    .io_exe_reqs_0_bits_uop_stq_idx(iregister_read_io_exe_reqs_0_bits_uop_stq_idx),
    .io_exe_reqs_0_bits_uop_pdst(iregister_read_io_exe_reqs_0_bits_uop_pdst),
    .io_exe_reqs_0_bits_uop_mem_cmd(iregister_read_io_exe_reqs_0_bits_uop_mem_cmd),
    .io_exe_reqs_0_bits_uop_mem_typ(iregister_read_io_exe_reqs_0_bits_uop_mem_typ),
    .io_exe_reqs_0_bits_uop_is_fence(iregister_read_io_exe_reqs_0_bits_uop_is_fence),
    .io_exe_reqs_0_bits_uop_is_store(iregister_read_io_exe_reqs_0_bits_uop_is_store),
    .io_exe_reqs_0_bits_uop_is_amo(iregister_read_io_exe_reqs_0_bits_uop_is_amo),
    .io_exe_reqs_0_bits_uop_is_load(iregister_read_io_exe_reqs_0_bits_uop_is_load),
    .io_exe_reqs_0_bits_uop_dst_rtype(iregister_read_io_exe_reqs_0_bits_uop_dst_rtype),
    .io_exe_reqs_0_bits_uop_fp_val(iregister_read_io_exe_reqs_0_bits_uop_fp_val),
    .io_exe_reqs_0_bits_rs1_data(iregister_read_io_exe_reqs_0_bits_rs1_data),
    .io_exe_reqs_0_bits_rs2_data(iregister_read_io_exe_reqs_0_bits_rs2_data),
    .io_exe_reqs_1_valid(iregister_read_io_exe_reqs_1_valid),
    .io_exe_reqs_1_bits_uop_valid(iregister_read_io_exe_reqs_1_bits_uop_valid),
    .io_exe_reqs_1_bits_uop_iw_state(iregister_read_io_exe_reqs_1_bits_uop_iw_state),
    .io_exe_reqs_1_bits_uop_uopc(iregister_read_io_exe_reqs_1_bits_uop_uopc),
    .io_exe_reqs_1_bits_uop_inst(iregister_read_io_exe_reqs_1_bits_uop_inst),
    .io_exe_reqs_1_bits_uop_pc(iregister_read_io_exe_reqs_1_bits_uop_pc),
    .io_exe_reqs_1_bits_uop_iqtype(iregister_read_io_exe_reqs_1_bits_uop_iqtype),
    .io_exe_reqs_1_bits_uop_fu_code(iregister_read_io_exe_reqs_1_bits_uop_fu_code),
    .io_exe_reqs_1_bits_uop_ctrl_br_type(iregister_read_io_exe_reqs_1_bits_uop_ctrl_br_type),
    .io_exe_reqs_1_bits_uop_ctrl_op1_sel(iregister_read_io_exe_reqs_1_bits_uop_ctrl_op1_sel),
    .io_exe_reqs_1_bits_uop_ctrl_op2_sel(iregister_read_io_exe_reqs_1_bits_uop_ctrl_op2_sel),
    .io_exe_reqs_1_bits_uop_ctrl_imm_sel(iregister_read_io_exe_reqs_1_bits_uop_ctrl_imm_sel),
    .io_exe_reqs_1_bits_uop_ctrl_op_fcn(iregister_read_io_exe_reqs_1_bits_uop_ctrl_op_fcn),
    .io_exe_reqs_1_bits_uop_ctrl_fcn_dw(iregister_read_io_exe_reqs_1_bits_uop_ctrl_fcn_dw),
    .io_exe_reqs_1_bits_uop_ctrl_rf_wen(iregister_read_io_exe_reqs_1_bits_uop_ctrl_rf_wen),
    .io_exe_reqs_1_bits_uop_ctrl_csr_cmd(iregister_read_io_exe_reqs_1_bits_uop_ctrl_csr_cmd),
    .io_exe_reqs_1_bits_uop_ctrl_is_load(iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_load),
    .io_exe_reqs_1_bits_uop_ctrl_is_sta(iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_sta),
    .io_exe_reqs_1_bits_uop_ctrl_is_std(iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_std),
    .io_exe_reqs_1_bits_uop_allocate_brtag(iregister_read_io_exe_reqs_1_bits_uop_allocate_brtag),
    .io_exe_reqs_1_bits_uop_is_br_or_jmp(iregister_read_io_exe_reqs_1_bits_uop_is_br_or_jmp),
    .io_exe_reqs_1_bits_uop_is_jump(iregister_read_io_exe_reqs_1_bits_uop_is_jump),
    .io_exe_reqs_1_bits_uop_is_jal(iregister_read_io_exe_reqs_1_bits_uop_is_jal),
    .io_exe_reqs_1_bits_uop_is_ret(iregister_read_io_exe_reqs_1_bits_uop_is_ret),
    .io_exe_reqs_1_bits_uop_is_call(iregister_read_io_exe_reqs_1_bits_uop_is_call),
    .io_exe_reqs_1_bits_uop_br_mask(iregister_read_io_exe_reqs_1_bits_uop_br_mask),
    .io_exe_reqs_1_bits_uop_br_tag(iregister_read_io_exe_reqs_1_bits_uop_br_tag),
    .io_exe_reqs_1_bits_uop_br_prediction_btb_blame(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_blame),
    .io_exe_reqs_1_bits_uop_br_prediction_btb_hit(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_hit),
    .io_exe_reqs_1_bits_uop_br_prediction_btb_taken(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_taken),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_blame(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_blame),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_hit(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_hit),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_taken(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_taken),
    .io_exe_reqs_1_bits_uop_br_prediction_bim_resp_value(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_value),
    .io_exe_reqs_1_bits_uop_br_prediction_bim_resp_entry_idx(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_entry_idx),
    .io_exe_reqs_1_bits_uop_br_prediction_bim_resp_way_idx(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_way_idx),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_takens(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_takens),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_u(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_u),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_ptr(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_ptr),
    .io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_info(iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_info),
    .io_exe_reqs_1_bits_uop_stat_brjmp_mispredicted(iregister_read_io_exe_reqs_1_bits_uop_stat_brjmp_mispredicted),
    .io_exe_reqs_1_bits_uop_stat_btb_made_pred(iregister_read_io_exe_reqs_1_bits_uop_stat_btb_made_pred),
    .io_exe_reqs_1_bits_uop_stat_btb_mispredicted(iregister_read_io_exe_reqs_1_bits_uop_stat_btb_mispredicted),
    .io_exe_reqs_1_bits_uop_stat_bpd_made_pred(iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_made_pred),
    .io_exe_reqs_1_bits_uop_stat_bpd_mispredicted(iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_mispredicted),
    .io_exe_reqs_1_bits_uop_fetch_pc_lob(iregister_read_io_exe_reqs_1_bits_uop_fetch_pc_lob),
    .io_exe_reqs_1_bits_uop_imm_packed(iregister_read_io_exe_reqs_1_bits_uop_imm_packed),
    .io_exe_reqs_1_bits_uop_csr_addr(iregister_read_io_exe_reqs_1_bits_uop_csr_addr),
    .io_exe_reqs_1_bits_uop_rob_idx(iregister_read_io_exe_reqs_1_bits_uop_rob_idx),
    .io_exe_reqs_1_bits_uop_ldq_idx(iregister_read_io_exe_reqs_1_bits_uop_ldq_idx),
    .io_exe_reqs_1_bits_uop_stq_idx(iregister_read_io_exe_reqs_1_bits_uop_stq_idx),
    .io_exe_reqs_1_bits_uop_brob_idx(iregister_read_io_exe_reqs_1_bits_uop_brob_idx),
    .io_exe_reqs_1_bits_uop_pdst(iregister_read_io_exe_reqs_1_bits_uop_pdst),
    .io_exe_reqs_1_bits_uop_pop1(iregister_read_io_exe_reqs_1_bits_uop_pop1),
    .io_exe_reqs_1_bits_uop_pop2(iregister_read_io_exe_reqs_1_bits_uop_pop2),
    .io_exe_reqs_1_bits_uop_pop3(iregister_read_io_exe_reqs_1_bits_uop_pop3),
    .io_exe_reqs_1_bits_uop_prs1_busy(iregister_read_io_exe_reqs_1_bits_uop_prs1_busy),
    .io_exe_reqs_1_bits_uop_prs2_busy(iregister_read_io_exe_reqs_1_bits_uop_prs2_busy),
    .io_exe_reqs_1_bits_uop_prs3_busy(iregister_read_io_exe_reqs_1_bits_uop_prs3_busy),
    .io_exe_reqs_1_bits_uop_stale_pdst(iregister_read_io_exe_reqs_1_bits_uop_stale_pdst),
    .io_exe_reqs_1_bits_uop_exception(iregister_read_io_exe_reqs_1_bits_uop_exception),
    .io_exe_reqs_1_bits_uop_exc_cause(iregister_read_io_exe_reqs_1_bits_uop_exc_cause),
    .io_exe_reqs_1_bits_uop_bypassable(iregister_read_io_exe_reqs_1_bits_uop_bypassable),
    .io_exe_reqs_1_bits_uop_mem_cmd(iregister_read_io_exe_reqs_1_bits_uop_mem_cmd),
    .io_exe_reqs_1_bits_uop_mem_typ(iregister_read_io_exe_reqs_1_bits_uop_mem_typ),
    .io_exe_reqs_1_bits_uop_is_fence(iregister_read_io_exe_reqs_1_bits_uop_is_fence),
    .io_exe_reqs_1_bits_uop_is_fencei(iregister_read_io_exe_reqs_1_bits_uop_is_fencei),
    .io_exe_reqs_1_bits_uop_is_store(iregister_read_io_exe_reqs_1_bits_uop_is_store),
    .io_exe_reqs_1_bits_uop_is_amo(iregister_read_io_exe_reqs_1_bits_uop_is_amo),
    .io_exe_reqs_1_bits_uop_is_load(iregister_read_io_exe_reqs_1_bits_uop_is_load),
    .io_exe_reqs_1_bits_uop_is_sys_pc2epc(iregister_read_io_exe_reqs_1_bits_uop_is_sys_pc2epc),
    .io_exe_reqs_1_bits_uop_is_unique(iregister_read_io_exe_reqs_1_bits_uop_is_unique),
    .io_exe_reqs_1_bits_uop_flush_on_commit(iregister_read_io_exe_reqs_1_bits_uop_flush_on_commit),
    .io_exe_reqs_1_bits_uop_ldst(iregister_read_io_exe_reqs_1_bits_uop_ldst),
    .io_exe_reqs_1_bits_uop_lrs1(iregister_read_io_exe_reqs_1_bits_uop_lrs1),
    .io_exe_reqs_1_bits_uop_lrs2(iregister_read_io_exe_reqs_1_bits_uop_lrs2),
    .io_exe_reqs_1_bits_uop_lrs3(iregister_read_io_exe_reqs_1_bits_uop_lrs3),
    .io_exe_reqs_1_bits_uop_ldst_val(iregister_read_io_exe_reqs_1_bits_uop_ldst_val),
    .io_exe_reqs_1_bits_uop_dst_rtype(iregister_read_io_exe_reqs_1_bits_uop_dst_rtype),
    .io_exe_reqs_1_bits_uop_lrs1_rtype(iregister_read_io_exe_reqs_1_bits_uop_lrs1_rtype),
    .io_exe_reqs_1_bits_uop_lrs2_rtype(iregister_read_io_exe_reqs_1_bits_uop_lrs2_rtype),
    .io_exe_reqs_1_bits_uop_frs3_en(iregister_read_io_exe_reqs_1_bits_uop_frs3_en),
    .io_exe_reqs_1_bits_uop_fp_val(iregister_read_io_exe_reqs_1_bits_uop_fp_val),
    .io_exe_reqs_1_bits_uop_fp_single(iregister_read_io_exe_reqs_1_bits_uop_fp_single),
    .io_exe_reqs_1_bits_uop_xcpt_pf_if(iregister_read_io_exe_reqs_1_bits_uop_xcpt_pf_if),
    .io_exe_reqs_1_bits_uop_xcpt_ae_if(iregister_read_io_exe_reqs_1_bits_uop_xcpt_ae_if),
    .io_exe_reqs_1_bits_uop_replay_if(iregister_read_io_exe_reqs_1_bits_uop_replay_if),
    .io_exe_reqs_1_bits_uop_xcpt_ma_if(iregister_read_io_exe_reqs_1_bits_uop_xcpt_ma_if),
    .io_exe_reqs_1_bits_uop_debug_wdata(iregister_read_io_exe_reqs_1_bits_uop_debug_wdata),
    .io_exe_reqs_1_bits_uop_debug_events_fetch_seq(iregister_read_io_exe_reqs_1_bits_uop_debug_events_fetch_seq),
    .io_exe_reqs_1_bits_rs1_data(iregister_read_io_exe_reqs_1_bits_rs1_data),
    .io_exe_reqs_1_bits_rs2_data(iregister_read_io_exe_reqs_1_bits_rs2_data),
    .io_exe_reqs_2_valid(iregister_read_io_exe_reqs_2_valid),
    .io_exe_reqs_2_bits_uop_valid(iregister_read_io_exe_reqs_2_bits_uop_valid),
    .io_exe_reqs_2_bits_uop_iw_state(iregister_read_io_exe_reqs_2_bits_uop_iw_state),
    .io_exe_reqs_2_bits_uop_uopc(iregister_read_io_exe_reqs_2_bits_uop_uopc),
    .io_exe_reqs_2_bits_uop_inst(iregister_read_io_exe_reqs_2_bits_uop_inst),
    .io_exe_reqs_2_bits_uop_pc(iregister_read_io_exe_reqs_2_bits_uop_pc),
    .io_exe_reqs_2_bits_uop_iqtype(iregister_read_io_exe_reqs_2_bits_uop_iqtype),
    .io_exe_reqs_2_bits_uop_fu_code(iregister_read_io_exe_reqs_2_bits_uop_fu_code),
    .io_exe_reqs_2_bits_uop_ctrl_op1_sel(iregister_read_io_exe_reqs_2_bits_uop_ctrl_op1_sel),
    .io_exe_reqs_2_bits_uop_ctrl_op2_sel(iregister_read_io_exe_reqs_2_bits_uop_ctrl_op2_sel),
    .io_exe_reqs_2_bits_uop_ctrl_imm_sel(iregister_read_io_exe_reqs_2_bits_uop_ctrl_imm_sel),
    .io_exe_reqs_2_bits_uop_ctrl_op_fcn(iregister_read_io_exe_reqs_2_bits_uop_ctrl_op_fcn),
    .io_exe_reqs_2_bits_uop_ctrl_fcn_dw(iregister_read_io_exe_reqs_2_bits_uop_ctrl_fcn_dw),
    .io_exe_reqs_2_bits_uop_ctrl_rf_wen(iregister_read_io_exe_reqs_2_bits_uop_ctrl_rf_wen),
    .io_exe_reqs_2_bits_uop_ctrl_is_load(iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_load),
    .io_exe_reqs_2_bits_uop_ctrl_is_sta(iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_sta),
    .io_exe_reqs_2_bits_uop_ctrl_is_std(iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_std),
    .io_exe_reqs_2_bits_uop_allocate_brtag(iregister_read_io_exe_reqs_2_bits_uop_allocate_brtag),
    .io_exe_reqs_2_bits_uop_is_br_or_jmp(iregister_read_io_exe_reqs_2_bits_uop_is_br_or_jmp),
    .io_exe_reqs_2_bits_uop_is_jump(iregister_read_io_exe_reqs_2_bits_uop_is_jump),
    .io_exe_reqs_2_bits_uop_is_jal(iregister_read_io_exe_reqs_2_bits_uop_is_jal),
    .io_exe_reqs_2_bits_uop_is_ret(iregister_read_io_exe_reqs_2_bits_uop_is_ret),
    .io_exe_reqs_2_bits_uop_is_call(iregister_read_io_exe_reqs_2_bits_uop_is_call),
    .io_exe_reqs_2_bits_uop_br_mask(iregister_read_io_exe_reqs_2_bits_uop_br_mask),
    .io_exe_reqs_2_bits_uop_br_tag(iregister_read_io_exe_reqs_2_bits_uop_br_tag),
    .io_exe_reqs_2_bits_uop_br_prediction_btb_blame(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_blame),
    .io_exe_reqs_2_bits_uop_br_prediction_btb_hit(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_hit),
    .io_exe_reqs_2_bits_uop_br_prediction_btb_taken(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_taken),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_blame(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_blame),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_hit(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_hit),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_taken(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_taken),
    .io_exe_reqs_2_bits_uop_br_prediction_bim_resp_value(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_value),
    .io_exe_reqs_2_bits_uop_br_prediction_bim_resp_entry_idx(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_entry_idx),
    .io_exe_reqs_2_bits_uop_br_prediction_bim_resp_way_idx(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_way_idx),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_takens(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_takens),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_u(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_u),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_ptr(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_ptr),
    .io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_info(iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_info),
    .io_exe_reqs_2_bits_uop_stat_brjmp_mispredicted(iregister_read_io_exe_reqs_2_bits_uop_stat_brjmp_mispredicted),
    .io_exe_reqs_2_bits_uop_stat_btb_made_pred(iregister_read_io_exe_reqs_2_bits_uop_stat_btb_made_pred),
    .io_exe_reqs_2_bits_uop_stat_btb_mispredicted(iregister_read_io_exe_reqs_2_bits_uop_stat_btb_mispredicted),
    .io_exe_reqs_2_bits_uop_stat_bpd_made_pred(iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_made_pred),
    .io_exe_reqs_2_bits_uop_stat_bpd_mispredicted(iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_mispredicted),
    .io_exe_reqs_2_bits_uop_fetch_pc_lob(iregister_read_io_exe_reqs_2_bits_uop_fetch_pc_lob),
    .io_exe_reqs_2_bits_uop_imm_packed(iregister_read_io_exe_reqs_2_bits_uop_imm_packed),
    .io_exe_reqs_2_bits_uop_csr_addr(iregister_read_io_exe_reqs_2_bits_uop_csr_addr),
    .io_exe_reqs_2_bits_uop_rob_idx(iregister_read_io_exe_reqs_2_bits_uop_rob_idx),
    .io_exe_reqs_2_bits_uop_ldq_idx(iregister_read_io_exe_reqs_2_bits_uop_ldq_idx),
    .io_exe_reqs_2_bits_uop_stq_idx(iregister_read_io_exe_reqs_2_bits_uop_stq_idx),
    .io_exe_reqs_2_bits_uop_brob_idx(iregister_read_io_exe_reqs_2_bits_uop_brob_idx),
    .io_exe_reqs_2_bits_uop_pdst(iregister_read_io_exe_reqs_2_bits_uop_pdst),
    .io_exe_reqs_2_bits_uop_pop1(iregister_read_io_exe_reqs_2_bits_uop_pop1),
    .io_exe_reqs_2_bits_uop_pop2(iregister_read_io_exe_reqs_2_bits_uop_pop2),
    .io_exe_reqs_2_bits_uop_pop3(iregister_read_io_exe_reqs_2_bits_uop_pop3),
    .io_exe_reqs_2_bits_uop_prs1_busy(iregister_read_io_exe_reqs_2_bits_uop_prs1_busy),
    .io_exe_reqs_2_bits_uop_prs2_busy(iregister_read_io_exe_reqs_2_bits_uop_prs2_busy),
    .io_exe_reqs_2_bits_uop_prs3_busy(iregister_read_io_exe_reqs_2_bits_uop_prs3_busy),
    .io_exe_reqs_2_bits_uop_stale_pdst(iregister_read_io_exe_reqs_2_bits_uop_stale_pdst),
    .io_exe_reqs_2_bits_uop_exception(iregister_read_io_exe_reqs_2_bits_uop_exception),
    .io_exe_reqs_2_bits_uop_exc_cause(iregister_read_io_exe_reqs_2_bits_uop_exc_cause),
    .io_exe_reqs_2_bits_uop_bypassable(iregister_read_io_exe_reqs_2_bits_uop_bypassable),
    .io_exe_reqs_2_bits_uop_mem_cmd(iregister_read_io_exe_reqs_2_bits_uop_mem_cmd),
    .io_exe_reqs_2_bits_uop_mem_typ(iregister_read_io_exe_reqs_2_bits_uop_mem_typ),
    .io_exe_reqs_2_bits_uop_is_fence(iregister_read_io_exe_reqs_2_bits_uop_is_fence),
    .io_exe_reqs_2_bits_uop_is_fencei(iregister_read_io_exe_reqs_2_bits_uop_is_fencei),
    .io_exe_reqs_2_bits_uop_is_store(iregister_read_io_exe_reqs_2_bits_uop_is_store),
    .io_exe_reqs_2_bits_uop_is_amo(iregister_read_io_exe_reqs_2_bits_uop_is_amo),
    .io_exe_reqs_2_bits_uop_is_load(iregister_read_io_exe_reqs_2_bits_uop_is_load),
    .io_exe_reqs_2_bits_uop_is_sys_pc2epc(iregister_read_io_exe_reqs_2_bits_uop_is_sys_pc2epc),
    .io_exe_reqs_2_bits_uop_is_unique(iregister_read_io_exe_reqs_2_bits_uop_is_unique),
    .io_exe_reqs_2_bits_uop_flush_on_commit(iregister_read_io_exe_reqs_2_bits_uop_flush_on_commit),
    .io_exe_reqs_2_bits_uop_ldst(iregister_read_io_exe_reqs_2_bits_uop_ldst),
    .io_exe_reqs_2_bits_uop_lrs1(iregister_read_io_exe_reqs_2_bits_uop_lrs1),
    .io_exe_reqs_2_bits_uop_lrs2(iregister_read_io_exe_reqs_2_bits_uop_lrs2),
    .io_exe_reqs_2_bits_uop_lrs3(iregister_read_io_exe_reqs_2_bits_uop_lrs3),
    .io_exe_reqs_2_bits_uop_ldst_val(iregister_read_io_exe_reqs_2_bits_uop_ldst_val),
    .io_exe_reqs_2_bits_uop_dst_rtype(iregister_read_io_exe_reqs_2_bits_uop_dst_rtype),
    .io_exe_reqs_2_bits_uop_lrs1_rtype(iregister_read_io_exe_reqs_2_bits_uop_lrs1_rtype),
    .io_exe_reqs_2_bits_uop_lrs2_rtype(iregister_read_io_exe_reqs_2_bits_uop_lrs2_rtype),
    .io_exe_reqs_2_bits_uop_frs3_en(iregister_read_io_exe_reqs_2_bits_uop_frs3_en),
    .io_exe_reqs_2_bits_uop_fp_val(iregister_read_io_exe_reqs_2_bits_uop_fp_val),
    .io_exe_reqs_2_bits_uop_fp_single(iregister_read_io_exe_reqs_2_bits_uop_fp_single),
    .io_exe_reqs_2_bits_uop_xcpt_pf_if(iregister_read_io_exe_reqs_2_bits_uop_xcpt_pf_if),
    .io_exe_reqs_2_bits_uop_xcpt_ae_if(iregister_read_io_exe_reqs_2_bits_uop_xcpt_ae_if),
    .io_exe_reqs_2_bits_uop_replay_if(iregister_read_io_exe_reqs_2_bits_uop_replay_if),
    .io_exe_reqs_2_bits_uop_xcpt_ma_if(iregister_read_io_exe_reqs_2_bits_uop_xcpt_ma_if),
    .io_exe_reqs_2_bits_uop_debug_wdata(iregister_read_io_exe_reqs_2_bits_uop_debug_wdata),
    .io_exe_reqs_2_bits_uop_debug_events_fetch_seq(iregister_read_io_exe_reqs_2_bits_uop_debug_events_fetch_seq),
    .io_exe_reqs_2_bits_rs1_data(iregister_read_io_exe_reqs_2_bits_rs1_data),
    .io_exe_reqs_2_bits_rs2_data(iregister_read_io_exe_reqs_2_bits_rs2_data),
    .io_kill(iregister_read_io_kill),
    .io_brinfo_valid(iregister_read_io_brinfo_valid),
    .io_brinfo_mispredict(iregister_read_io_brinfo_mispredict),
    .io_brinfo_mask(iregister_read_io_brinfo_mask)
  );
  DCacheShim dc_shim (
    .clock(dc_shim_clock),
    .reset(dc_shim_reset),
    .io_core_req_valid(dc_shim_io_core_req_valid),
    .io_core_req_bits_addr(dc_shim_io_core_req_bits_addr),
    .io_core_req_bits_uop_uopc(dc_shim_io_core_req_bits_uop_uopc),
    .io_core_req_bits_uop_br_mask(dc_shim_io_core_req_bits_uop_br_mask),
    .io_core_req_bits_uop_rob_idx(dc_shim_io_core_req_bits_uop_rob_idx),
    .io_core_req_bits_uop_ldq_idx(dc_shim_io_core_req_bits_uop_ldq_idx),
    .io_core_req_bits_uop_stq_idx(dc_shim_io_core_req_bits_uop_stq_idx),
    .io_core_req_bits_uop_pdst(dc_shim_io_core_req_bits_uop_pdst),
    .io_core_req_bits_uop_mem_cmd(dc_shim_io_core_req_bits_uop_mem_cmd),
    .io_core_req_bits_uop_mem_typ(dc_shim_io_core_req_bits_uop_mem_typ),
    .io_core_req_bits_uop_is_store(dc_shim_io_core_req_bits_uop_is_store),
    .io_core_req_bits_uop_is_amo(dc_shim_io_core_req_bits_uop_is_amo),
    .io_core_req_bits_uop_is_load(dc_shim_io_core_req_bits_uop_is_load),
    .io_core_req_bits_uop_dst_rtype(dc_shim_io_core_req_bits_uop_dst_rtype),
    .io_core_req_bits_uop_fp_val(dc_shim_io_core_req_bits_uop_fp_val),
    .io_core_req_bits_data(dc_shim_io_core_req_bits_data),
    .io_core_req_bits_kill(dc_shim_io_core_req_bits_kill),
    .io_core_resp_valid(dc_shim_io_core_resp_valid),
    .io_core_resp_bits_data_subword(dc_shim_io_core_resp_bits_data_subword),
    .io_core_resp_bits_uop_uopc(dc_shim_io_core_resp_bits_uop_uopc),
    .io_core_resp_bits_uop_rob_idx(dc_shim_io_core_resp_bits_uop_rob_idx),
    .io_core_resp_bits_uop_ldq_idx(dc_shim_io_core_resp_bits_uop_ldq_idx),
    .io_core_resp_bits_uop_stq_idx(dc_shim_io_core_resp_bits_uop_stq_idx),
    .io_core_resp_bits_uop_pdst(dc_shim_io_core_resp_bits_uop_pdst),
    .io_core_resp_bits_uop_mem_cmd(dc_shim_io_core_resp_bits_uop_mem_cmd),
    .io_core_resp_bits_uop_mem_typ(dc_shim_io_core_resp_bits_uop_mem_typ),
    .io_core_resp_bits_uop_is_store(dc_shim_io_core_resp_bits_uop_is_store),
    .io_core_resp_bits_uop_is_amo(dc_shim_io_core_resp_bits_uop_is_amo),
    .io_core_resp_bits_uop_is_load(dc_shim_io_core_resp_bits_uop_is_load),
    .io_core_resp_bits_uop_dst_rtype(dc_shim_io_core_resp_bits_uop_dst_rtype),
    .io_core_resp_bits_uop_fp_val(dc_shim_io_core_resp_bits_uop_fp_val),
    .io_core_brinfo_valid(dc_shim_io_core_brinfo_valid),
    .io_core_brinfo_mispredict(dc_shim_io_core_brinfo_mispredict),
    .io_core_brinfo_mask(dc_shim_io_core_brinfo_mask),
    .io_core_nack_valid(dc_shim_io_core_nack_valid),
    .io_core_nack_lsu_idx(dc_shim_io_core_nack_lsu_idx),
    .io_core_nack_isload(dc_shim_io_core_nack_isload),
    .io_core_nack_cache_nack(dc_shim_io_core_nack_cache_nack),
    .io_core_flush_pipe(dc_shim_io_core_flush_pipe),
    .io_core_invalidate_lr(dc_shim_io_core_invalidate_lr),
    .io_core_ordered(dc_shim_io_core_ordered),
    .io_dmem_req_ready(dc_shim_io_dmem_req_ready),
    .io_dmem_req_valid(dc_shim_io_dmem_req_valid),
    .io_dmem_req_bits_addr(dc_shim_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(dc_shim_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(dc_shim_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(dc_shim_io_dmem_req_bits_typ),
    .io_dmem_s1_kill(dc_shim_io_dmem_s1_kill),
    .io_dmem_s1_data_data(dc_shim_io_dmem_s1_data_data),
    .io_dmem_s2_nack(dc_shim_io_dmem_s2_nack),
    .io_dmem_resp_valid(dc_shim_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(dc_shim_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_data(dc_shim_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_has_data(dc_shim_io_dmem_resp_bits_has_data),
    .io_dmem_s2_xcpt_ma_ld(dc_shim_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(dc_shim_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(dc_shim_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(dc_shim_io_dmem_s2_xcpt_pf_st),
    .io_dmem_invalidate_lr(dc_shim_io_dmem_invalidate_lr),
    .io_dmem_ordered(dc_shim_io_dmem_ordered)
  );
  LoadStoreUnit lsu (
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_dec_st_vals_0(lsu_io_dec_st_vals_0),
    .io_dec_st_vals_1(lsu_io_dec_st_vals_1),
    .io_dec_ld_vals_0(lsu_io_dec_ld_vals_0),
    .io_dec_ld_vals_1(lsu_io_dec_ld_vals_1),
    .io_dec_uops_0_uopc(lsu_io_dec_uops_0_uopc),
    .io_dec_uops_0_br_mask(lsu_io_dec_uops_0_br_mask),
    .io_dec_uops_0_rob_idx(lsu_io_dec_uops_0_rob_idx),
    .io_dec_uops_0_ldq_idx(lsu_io_dec_uops_0_ldq_idx),
    .io_dec_uops_0_stq_idx(lsu_io_dec_uops_0_stq_idx),
    .io_dec_uops_0_mem_cmd(lsu_io_dec_uops_0_mem_cmd),
    .io_dec_uops_0_mem_typ(lsu_io_dec_uops_0_mem_typ),
    .io_dec_uops_0_is_fence(lsu_io_dec_uops_0_is_fence),
    .io_dec_uops_0_is_store(lsu_io_dec_uops_0_is_store),
    .io_dec_uops_0_is_amo(lsu_io_dec_uops_0_is_amo),
    .io_dec_uops_0_is_load(lsu_io_dec_uops_0_is_load),
    .io_dec_uops_0_dst_rtype(lsu_io_dec_uops_0_dst_rtype),
    .io_dec_uops_0_fp_val(lsu_io_dec_uops_0_fp_val),
    .io_dec_uops_1_uopc(lsu_io_dec_uops_1_uopc),
    .io_dec_uops_1_br_mask(lsu_io_dec_uops_1_br_mask),
    .io_dec_uops_1_rob_idx(lsu_io_dec_uops_1_rob_idx),
    .io_dec_uops_1_ldq_idx(lsu_io_dec_uops_1_ldq_idx),
    .io_dec_uops_1_stq_idx(lsu_io_dec_uops_1_stq_idx),
    .io_dec_uops_1_mem_cmd(lsu_io_dec_uops_1_mem_cmd),
    .io_dec_uops_1_mem_typ(lsu_io_dec_uops_1_mem_typ),
    .io_dec_uops_1_is_fence(lsu_io_dec_uops_1_is_fence),
    .io_dec_uops_1_is_store(lsu_io_dec_uops_1_is_store),
    .io_dec_uops_1_is_amo(lsu_io_dec_uops_1_is_amo),
    .io_dec_uops_1_is_load(lsu_io_dec_uops_1_is_load),
    .io_dec_uops_1_dst_rtype(lsu_io_dec_uops_1_dst_rtype),
    .io_dec_uops_1_fp_val(lsu_io_dec_uops_1_fp_val),
    .io_new_ldq_idx(lsu_io_new_ldq_idx),
    .io_new_stq_idx(lsu_io_new_stq_idx),
    .io_exe_resp_valid(lsu_io_exe_resp_valid),
    .io_exe_resp_bits_uop_uopc(lsu_io_exe_resp_bits_uop_uopc),
    .io_exe_resp_bits_uop_ctrl_is_load(lsu_io_exe_resp_bits_uop_ctrl_is_load),
    .io_exe_resp_bits_uop_ctrl_is_sta(lsu_io_exe_resp_bits_uop_ctrl_is_sta),
    .io_exe_resp_bits_uop_ctrl_is_std(lsu_io_exe_resp_bits_uop_ctrl_is_std),
    .io_exe_resp_bits_uop_br_mask(lsu_io_exe_resp_bits_uop_br_mask),
    .io_exe_resp_bits_uop_rob_idx(lsu_io_exe_resp_bits_uop_rob_idx),
    .io_exe_resp_bits_uop_ldq_idx(lsu_io_exe_resp_bits_uop_ldq_idx),
    .io_exe_resp_bits_uop_stq_idx(lsu_io_exe_resp_bits_uop_stq_idx),
    .io_exe_resp_bits_uop_pdst(lsu_io_exe_resp_bits_uop_pdst),
    .io_exe_resp_bits_uop_mem_cmd(lsu_io_exe_resp_bits_uop_mem_cmd),
    .io_exe_resp_bits_uop_mem_typ(lsu_io_exe_resp_bits_uop_mem_typ),
    .io_exe_resp_bits_uop_is_fence(lsu_io_exe_resp_bits_uop_is_fence),
    .io_exe_resp_bits_uop_is_store(lsu_io_exe_resp_bits_uop_is_store),
    .io_exe_resp_bits_uop_is_amo(lsu_io_exe_resp_bits_uop_is_amo),
    .io_exe_resp_bits_uop_is_load(lsu_io_exe_resp_bits_uop_is_load),
    .io_exe_resp_bits_uop_dst_rtype(lsu_io_exe_resp_bits_uop_dst_rtype),
    .io_exe_resp_bits_uop_fp_val(lsu_io_exe_resp_bits_uop_fp_val),
    .io_exe_resp_bits_data(lsu_io_exe_resp_bits_data),
    .io_exe_resp_bits_addr(lsu_io_exe_resp_bits_addr),
    .io_exe_resp_bits_mxcpt_valid(lsu_io_exe_resp_bits_mxcpt_valid),
    .io_exe_resp_bits_mxcpt_bits(lsu_io_exe_resp_bits_mxcpt_bits),
    .io_exe_resp_bits_sfence_valid(lsu_io_exe_resp_bits_sfence_valid),
    .io_exe_resp_bits_sfence_bits_rs1(lsu_io_exe_resp_bits_sfence_bits_rs1),
    .io_exe_resp_bits_sfence_bits_rs2(lsu_io_exe_resp_bits_sfence_bits_rs2),
    .io_exe_resp_bits_sfence_bits_addr(lsu_io_exe_resp_bits_sfence_bits_addr),
    .io_fp_stdata_valid(lsu_io_fp_stdata_valid),
    .io_fp_stdata_bits_uop_br_mask(lsu_io_fp_stdata_bits_uop_br_mask),
    .io_fp_stdata_bits_uop_rob_idx(lsu_io_fp_stdata_bits_uop_rob_idx),
    .io_fp_stdata_bits_uop_stq_idx(lsu_io_fp_stdata_bits_uop_stq_idx),
    .io_fp_stdata_bits_uop_is_amo(lsu_io_fp_stdata_bits_uop_is_amo),
    .io_fp_stdata_bits_data(lsu_io_fp_stdata_bits_data),
    .io_commit_store_mask_0(lsu_io_commit_store_mask_0),
    .io_commit_store_mask_1(lsu_io_commit_store_mask_1),
    .io_commit_load_mask_0(lsu_io_commit_load_mask_0),
    .io_commit_load_mask_1(lsu_io_commit_load_mask_1),
    .io_commit_load_at_rob_head(lsu_io_commit_load_at_rob_head),
    .io_memreq_val(lsu_io_memreq_val),
    .io_memreq_addr(lsu_io_memreq_addr),
    .io_memreq_wdata(lsu_io_memreq_wdata),
    .io_memreq_uop_uopc(lsu_io_memreq_uop_uopc),
    .io_memreq_uop_br_mask(lsu_io_memreq_uop_br_mask),
    .io_memreq_uop_rob_idx(lsu_io_memreq_uop_rob_idx),
    .io_memreq_uop_ldq_idx(lsu_io_memreq_uop_ldq_idx),
    .io_memreq_uop_stq_idx(lsu_io_memreq_uop_stq_idx),
    .io_memreq_uop_pdst(lsu_io_memreq_uop_pdst),
    .io_memreq_uop_mem_cmd(lsu_io_memreq_uop_mem_cmd),
    .io_memreq_uop_mem_typ(lsu_io_memreq_uop_mem_typ),
    .io_memreq_uop_is_store(lsu_io_memreq_uop_is_store),
    .io_memreq_uop_is_amo(lsu_io_memreq_uop_is_amo),
    .io_memreq_uop_is_load(lsu_io_memreq_uop_is_load),
    .io_memreq_uop_dst_rtype(lsu_io_memreq_uop_dst_rtype),
    .io_memreq_uop_fp_val(lsu_io_memreq_uop_fp_val),
    .io_memreq_kill(lsu_io_memreq_kill),
    .io_forward_val(lsu_io_forward_val),
    .io_forward_data(lsu_io_forward_data),
    .io_forward_uop_uopc(lsu_io_forward_uop_uopc),
    .io_forward_uop_rob_idx(lsu_io_forward_uop_rob_idx),
    .io_forward_uop_ldq_idx(lsu_io_forward_uop_ldq_idx),
    .io_forward_uop_stq_idx(lsu_io_forward_uop_stq_idx),
    .io_forward_uop_pdst(lsu_io_forward_uop_pdst),
    .io_forward_uop_mem_typ(lsu_io_forward_uop_mem_typ),
    .io_forward_uop_is_store(lsu_io_forward_uop_is_store),
    .io_forward_uop_is_amo(lsu_io_forward_uop_is_amo),
    .io_forward_uop_is_load(lsu_io_forward_uop_is_load),
    .io_forward_uop_dst_rtype(lsu_io_forward_uop_dst_rtype),
    .io_forward_uop_fp_val(lsu_io_forward_uop_fp_val),
    .io_memresp_valid(lsu_io_memresp_valid),
    .io_memresp_bits_ldq_idx(lsu_io_memresp_bits_ldq_idx),
    .io_memresp_bits_stq_idx(lsu_io_memresp_bits_stq_idx),
    .io_memresp_bits_is_load(lsu_io_memresp_bits_is_load),
    .io_brinfo_valid(lsu_io_brinfo_valid),
    .io_brinfo_mispredict(lsu_io_brinfo_mispredict),
    .io_brinfo_mask(lsu_io_brinfo_mask),
    .io_brinfo_ldq_idx(lsu_io_brinfo_ldq_idx),
    .io_brinfo_stq_idx(lsu_io_brinfo_stq_idx),
    .io_laq_full(lsu_io_laq_full),
    .io_stq_full(lsu_io_stq_full),
    .io_exception(lsu_io_exception),
    .io_lsu_clr_bsy_valid_0(lsu_io_lsu_clr_bsy_valid_0),
    .io_lsu_clr_bsy_valid_1(lsu_io_lsu_clr_bsy_valid_1),
    .io_lsu_clr_bsy_rob_idx_0(lsu_io_lsu_clr_bsy_rob_idx_0),
    .io_lsu_clr_bsy_rob_idx_1(lsu_io_lsu_clr_bsy_rob_idx_1),
    .io_lsu_fencei_rdy(lsu_io_lsu_fencei_rdy),
    .io_xcpt_valid(lsu_io_xcpt_valid),
    .io_xcpt_bits_uop_br_mask(lsu_io_xcpt_bits_uop_br_mask),
    .io_xcpt_bits_uop_rob_idx(lsu_io_xcpt_bits_uop_rob_idx),
    .io_xcpt_bits_cause(lsu_io_xcpt_bits_cause),
    .io_xcpt_bits_badvaddr(lsu_io_xcpt_bits_badvaddr),
    .io_nack_valid(lsu_io_nack_valid),
    .io_nack_lsu_idx(lsu_io_nack_lsu_idx),
    .io_nack_isload(lsu_io_nack_isload),
    .io_nack_cache_nack(lsu_io_nack_cache_nack),
    .io_dmem_is_ordered(lsu_io_dmem_is_ordered),
    .io_ptw_req_ready(lsu_io_ptw_req_ready),
    .io_ptw_req_valid(lsu_io_ptw_req_valid),
    .io_ptw_req_bits_addr(lsu_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(lsu_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(lsu_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(lsu_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(lsu_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(lsu_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(lsu_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(lsu_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(lsu_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(lsu_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(lsu_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(lsu_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(lsu_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(lsu_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(lsu_io_ptw_ptbr_mode),
    .io_ptw_status_dprv(lsu_io_ptw_status_dprv),
    .io_ptw_status_mxr(lsu_io_ptw_status_mxr),
    .io_ptw_status_sum(lsu_io_ptw_status_sum)
  );
  Rob rob (
    .clock(rob_clock),
    .reset(rob_reset),
    .io_enq_valids_0(rob_io_enq_valids_0),
    .io_enq_valids_1(rob_io_enq_valids_1),
    .io_enq_uops_0_pc(rob_io_enq_uops_0_pc),
    .io_enq_uops_0_br_mask(rob_io_enq_uops_0_br_mask),
    .io_enq_uops_0_rob_idx(rob_io_enq_uops_0_rob_idx),
    .io_enq_uops_0_brob_idx(rob_io_enq_uops_0_brob_idx),
    .io_enq_uops_0_pdst(rob_io_enq_uops_0_pdst),
    .io_enq_uops_0_stale_pdst(rob_io_enq_uops_0_stale_pdst),
    .io_enq_uops_0_exception(rob_io_enq_uops_0_exception),
    .io_enq_uops_0_exc_cause(rob_io_enq_uops_0_exc_cause),
    .io_enq_uops_0_is_fence(rob_io_enq_uops_0_is_fence),
    .io_enq_uops_0_is_fencei(rob_io_enq_uops_0_is_fencei),
    .io_enq_uops_0_is_store(rob_io_enq_uops_0_is_store),
    .io_enq_uops_0_is_load(rob_io_enq_uops_0_is_load),
    .io_enq_uops_0_is_sys_pc2epc(rob_io_enq_uops_0_is_sys_pc2epc),
    .io_enq_uops_0_is_unique(rob_io_enq_uops_0_is_unique),
    .io_enq_uops_0_flush_on_commit(rob_io_enq_uops_0_flush_on_commit),
    .io_enq_uops_0_ldst(rob_io_enq_uops_0_ldst),
    .io_enq_uops_0_ldst_val(rob_io_enq_uops_0_ldst_val),
    .io_enq_uops_0_dst_rtype(rob_io_enq_uops_0_dst_rtype),
    .io_enq_uops_0_fp_val(rob_io_enq_uops_0_fp_val),
    .io_enq_uops_1_br_mask(rob_io_enq_uops_1_br_mask),
    .io_enq_uops_1_rob_idx(rob_io_enq_uops_1_rob_idx),
    .io_enq_uops_1_pdst(rob_io_enq_uops_1_pdst),
    .io_enq_uops_1_stale_pdst(rob_io_enq_uops_1_stale_pdst),
    .io_enq_uops_1_exception(rob_io_enq_uops_1_exception),
    .io_enq_uops_1_exc_cause(rob_io_enq_uops_1_exc_cause),
    .io_enq_uops_1_is_fence(rob_io_enq_uops_1_is_fence),
    .io_enq_uops_1_is_fencei(rob_io_enq_uops_1_is_fencei),
    .io_enq_uops_1_is_store(rob_io_enq_uops_1_is_store),
    .io_enq_uops_1_is_load(rob_io_enq_uops_1_is_load),
    .io_enq_uops_1_is_sys_pc2epc(rob_io_enq_uops_1_is_sys_pc2epc),
    .io_enq_uops_1_is_unique(rob_io_enq_uops_1_is_unique),
    .io_enq_uops_1_flush_on_commit(rob_io_enq_uops_1_flush_on_commit),
    .io_enq_uops_1_ldst(rob_io_enq_uops_1_ldst),
    .io_enq_uops_1_ldst_val(rob_io_enq_uops_1_ldst_val),
    .io_enq_uops_1_dst_rtype(rob_io_enq_uops_1_dst_rtype),
    .io_enq_uops_1_fp_val(rob_io_enq_uops_1_fp_val),
    .io_enq_has_br_or_jalr_in_packet(rob_io_enq_has_br_or_jalr_in_packet),
    .io_enq_partial_stall(rob_io_enq_partial_stall),
    .io_enq_new_packet(rob_io_enq_new_packet),
    .io_curr_rob_tail(rob_io_curr_rob_tail),
    .io_brinfo_valid(rob_io_brinfo_valid),
    .io_brinfo_mispredict(rob_io_brinfo_mispredict),
    .io_brinfo_mask(rob_io_brinfo_mask),
    .io_brinfo_rob_idx(rob_io_brinfo_rob_idx),
    .io_get_pc_rob_idx(rob_io_get_pc_rob_idx),
    .io_get_pc_curr_pc(rob_io_get_pc_curr_pc),
    .io_get_pc_curr_brob_idx(rob_io_get_pc_curr_brob_idx),
    .io_get_pc_next_val(rob_io_get_pc_next_val),
    .io_get_pc_next_pc(rob_io_get_pc_next_pc),
    .io_wb_resps_0_valid(rob_io_wb_resps_0_valid),
    .io_wb_resps_0_bits_uop_rob_idx(rob_io_wb_resps_0_bits_uop_rob_idx),
    .io_wb_resps_0_bits_uop_pdst(rob_io_wb_resps_0_bits_uop_pdst),
    .io_wb_resps_1_valid(rob_io_wb_resps_1_valid),
    .io_wb_resps_1_bits_uop_rob_idx(rob_io_wb_resps_1_bits_uop_rob_idx),
    .io_wb_resps_1_bits_uop_pdst(rob_io_wb_resps_1_bits_uop_pdst),
    .io_wb_resps_2_valid(rob_io_wb_resps_2_valid),
    .io_wb_resps_2_bits_uop_rob_idx(rob_io_wb_resps_2_bits_uop_rob_idx),
    .io_wb_resps_2_bits_uop_pdst(rob_io_wb_resps_2_bits_uop_pdst),
    .io_wb_resps_3_valid(rob_io_wb_resps_3_valid),
    .io_wb_resps_3_bits_uop_rob_idx(rob_io_wb_resps_3_bits_uop_rob_idx),
    .io_wb_resps_3_bits_uop_pdst(rob_io_wb_resps_3_bits_uop_pdst),
    .io_wb_resps_4_valid(rob_io_wb_resps_4_valid),
    .io_wb_resps_4_bits_uop_rob_idx(rob_io_wb_resps_4_bits_uop_rob_idx),
    .io_wb_resps_4_bits_uop_pdst(rob_io_wb_resps_4_bits_uop_pdst),
    .io_lsu_clr_bsy_valid_0(rob_io_lsu_clr_bsy_valid_0),
    .io_lsu_clr_bsy_valid_1(rob_io_lsu_clr_bsy_valid_1),
    .io_lsu_clr_bsy_rob_idx_0(rob_io_lsu_clr_bsy_rob_idx_0),
    .io_lsu_clr_bsy_rob_idx_1(rob_io_lsu_clr_bsy_rob_idx_1),
    .io_fflags_0_valid(rob_io_fflags_0_valid),
    .io_fflags_0_bits_uop_rob_idx(rob_io_fflags_0_bits_uop_rob_idx),
    .io_fflags_0_bits_flags(rob_io_fflags_0_bits_flags),
    .io_fflags_1_valid(rob_io_fflags_1_valid),
    .io_fflags_1_bits_uop_rob_idx(rob_io_fflags_1_bits_uop_rob_idx),
    .io_fflags_1_bits_flags(rob_io_fflags_1_bits_flags),
    .io_lxcpt_valid(rob_io_lxcpt_valid),
    .io_lxcpt_bits_uop_br_mask(rob_io_lxcpt_bits_uop_br_mask),
    .io_lxcpt_bits_uop_rob_idx(rob_io_lxcpt_bits_uop_rob_idx),
    .io_lxcpt_bits_cause(rob_io_lxcpt_bits_cause),
    .io_lxcpt_bits_badvaddr(rob_io_lxcpt_bits_badvaddr),
    .io_bxcpt_valid(rob_io_bxcpt_valid),
    .io_bxcpt_bits_uop_br_mask(rob_io_bxcpt_bits_uop_br_mask),
    .io_bxcpt_bits_uop_rob_idx(rob_io_bxcpt_bits_uop_rob_idx),
    .io_bxcpt_bits_badvaddr(rob_io_bxcpt_bits_badvaddr),
    .io_commit_valids_0(rob_io_commit_valids_0),
    .io_commit_valids_1(rob_io_commit_valids_1),
    .io_commit_uops_0_pdst(rob_io_commit_uops_0_pdst),
    .io_commit_uops_0_stale_pdst(rob_io_commit_uops_0_stale_pdst),
    .io_commit_uops_0_is_fencei(rob_io_commit_uops_0_is_fencei),
    .io_commit_uops_0_is_store(rob_io_commit_uops_0_is_store),
    .io_commit_uops_0_is_load(rob_io_commit_uops_0_is_load),
    .io_commit_uops_0_is_sys_pc2epc(rob_io_commit_uops_0_is_sys_pc2epc),
    .io_commit_uops_0_flush_on_commit(rob_io_commit_uops_0_flush_on_commit),
    .io_commit_uops_0_ldst(rob_io_commit_uops_0_ldst),
    .io_commit_uops_0_dst_rtype(rob_io_commit_uops_0_dst_rtype),
    .io_commit_uops_0_fp_val(rob_io_commit_uops_0_fp_val),
    .io_commit_uops_1_pdst(rob_io_commit_uops_1_pdst),
    .io_commit_uops_1_stale_pdst(rob_io_commit_uops_1_stale_pdst),
    .io_commit_uops_1_is_fencei(rob_io_commit_uops_1_is_fencei),
    .io_commit_uops_1_is_store(rob_io_commit_uops_1_is_store),
    .io_commit_uops_1_is_load(rob_io_commit_uops_1_is_load),
    .io_commit_uops_1_is_sys_pc2epc(rob_io_commit_uops_1_is_sys_pc2epc),
    .io_commit_uops_1_flush_on_commit(rob_io_commit_uops_1_flush_on_commit),
    .io_commit_uops_1_ldst(rob_io_commit_uops_1_ldst),
    .io_commit_uops_1_dst_rtype(rob_io_commit_uops_1_dst_rtype),
    .io_commit_uops_1_fp_val(rob_io_commit_uops_1_fp_val),
    .io_commit_fflags_valid(rob_io_commit_fflags_valid),
    .io_commit_fflags_bits(rob_io_commit_fflags_bits),
    .io_commit_rbk_valids_0(rob_io_commit_rbk_valids_0),
    .io_commit_rbk_valids_1(rob_io_commit_rbk_valids_1),
    .io_commit_st_mask_0(rob_io_commit_st_mask_0),
    .io_commit_st_mask_1(rob_io_commit_st_mask_1),
    .io_commit_ld_mask_0(rob_io_commit_ld_mask_0),
    .io_commit_ld_mask_1(rob_io_commit_ld_mask_1),
    .io_com_load_is_at_rob_head(rob_io_com_load_is_at_rob_head),
    .io_com_xcpt_valid(rob_io_com_xcpt_valid),
    .io_com_xcpt_bits_pc(rob_io_com_xcpt_bits_pc),
    .io_com_xcpt_bits_cause(rob_io_com_xcpt_bits_cause),
    .io_com_xcpt_bits_badvaddr(rob_io_com_xcpt_bits_badvaddr),
    .io_csr_eret(rob_io_csr_eret),
    .io_csr_evec(rob_io_csr_evec),
    .io_csr_stall(rob_io_csr_stall),
    .io_flush_valid(rob_io_flush_valid),
    .io_flush_bits_pc(rob_io_flush_bits_pc),
    .io_clear_brob(rob_io_clear_brob),
    .io_empty(rob_io_empty),
    .io_ready(rob_io_ready),
    .io_brob_deallocate_valid(rob_io_brob_deallocate_valid),
    .io_brob_deallocate_bits_brob_idx(rob_io_brob_deallocate_bits_brob_idx)
  );
  CSRFile csr (
    .clock(csr_clock),
    .reset(csr_reset),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_interrupts_seip(csr_io_interrupts_seip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_0_csr(csr_io_decode_0_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_decode_1_csr(csr_io_decode_1_csr),
    .io_decode_1_fp_illegal(csr_io_decode_1_fp_illegal),
    .io_decode_1_read_illegal(csr_io_decode_1_read_illegal),
    .io_decode_1_write_illegal(csr_io_decode_1_write_illegal),
    .io_decode_1_write_flush(csr_io_decode_1_write_flush),
    .io_decode_1_system_illegal(csr_io_decode_1_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_counters_0_eventSel(csr_io_counters_0_eventSel),
    .io_counters_0_inc(csr_io_counters_0_inc),
    .io_counters_1_eventSel(csr_io_counters_1_eventSel),
    .io_counters_1_inc(csr_io_counters_1_inc),
    .io_counters_2_eventSel(csr_io_counters_2_eventSel),
    .io_counters_2_inc(csr_io_counters_2_inc),
    .io_counters_3_eventSel(csr_io_counters_3_eventSel),
    .io_counters_3_inc(csr_io_counters_3_inc),
    .io_counters_4_eventSel(csr_io_counters_4_eventSel),
    .io_counters_4_inc(csr_io_counters_4_inc),
    .io_counters_5_eventSel(csr_io_counters_5_eventSel),
    .io_counters_5_inc(csr_io_counters_5_inc),
    .io_counters_6_eventSel(csr_io_counters_6_eventSel),
    .io_counters_6_inc(csr_io_counters_6_inc),
    .io_counters_7_eventSel(csr_io_counters_7_eventSel),
    .io_counters_7_inc(csr_io_counters_7_inc),
    .io_counters_8_eventSel(csr_io_counters_8_eventSel),
    .io_counters_8_inc(csr_io_counters_8_inc),
    .io_counters_9_eventSel(csr_io_counters_9_eventSel),
    .io_counters_9_inc(csr_io_counters_9_inc),
    .io_counters_10_eventSel(csr_io_counters_10_eventSel),
    .io_counters_10_inc(csr_io_counters_10_inc),
    .io_counters_11_eventSel(csr_io_counters_11_eventSel),
    .io_counters_11_inc(csr_io_counters_11_inc),
    .io_counters_12_eventSel(csr_io_counters_12_eventSel),
    .io_counters_12_inc(csr_io_counters_12_inc),
    .io_counters_13_eventSel(csr_io_counters_13_eventSel),
    .io_counters_13_inc(csr_io_counters_13_inc),
    .io_counters_14_eventSel(csr_io_counters_14_eventSel),
    .io_counters_14_inc(csr_io_counters_14_inc),
    .io_counters_15_eventSel(csr_io_counters_15_eventSel),
    .io_counters_15_inc(csr_io_counters_15_inc),
    .io_counters_16_eventSel(csr_io_counters_16_eventSel),
    .io_counters_16_inc(csr_io_counters_16_inc),
    .io_counters_17_eventSel(csr_io_counters_17_eventSel),
    .io_counters_17_inc(csr_io_counters_17_inc),
    .io_counters_18_eventSel(csr_io_counters_18_eventSel),
    .io_counters_18_inc(csr_io_counters_18_inc),
    .io_counters_19_eventSel(csr_io_counters_19_eventSel),
    .io_counters_19_inc(csr_io_counters_19_inc),
    .io_counters_20_eventSel(csr_io_counters_20_eventSel),
    .io_counters_20_inc(csr_io_counters_20_inc),
    .io_counters_21_eventSel(csr_io_counters_21_eventSel),
    .io_counters_21_inc(csr_io_counters_21_inc),
    .io_counters_22_eventSel(csr_io_counters_22_eventSel),
    .io_counters_22_inc(csr_io_counters_22_inc),
    .io_counters_23_eventSel(csr_io_counters_23_eventSel),
    .io_counters_23_inc(csr_io_counters_23_inc),
    .io_counters_24_eventSel(csr_io_counters_24_eventSel),
    .io_counters_24_inc(csr_io_counters_24_inc),
    .io_counters_25_eventSel(csr_io_counters_25_eventSel),
    .io_counters_25_inc(csr_io_counters_25_inc),
    .io_counters_26_eventSel(csr_io_counters_26_eventSel),
    .io_counters_26_inc(csr_io_counters_26_inc),
    .io_counters_27_eventSel(csr_io_counters_27_eventSel),
    .io_counters_27_inc(csr_io_counters_27_inc),
    .io_counters_28_eventSel(csr_io_counters_28_eventSel),
    .io_counters_28_inc(csr_io_counters_28_inc)
  );
  assign _T_1523 = io_imem_resp_valid | _T_1522;
  assign icache_blocked = _T_1523 == 1'h0;
  assign _T_1525 = csr_io_counters_0_eventSel[1:0];
  assign _T_1526 = csr_io_counters_0_eventSel[63:8];
  assign _T_1530 = {1'h0,rob_io_com_xcpt_valid};
  assign _T_1532 = {2'h0,_T_1530};
  assign _GEN_13 = {{52'd0}, _T_1532};
  assign _T_1533 = _T_1526 & _GEN_13;
  assign _T_1535 = _T_1533 != 56'h0;
  assign _T_1537 = br_unit_brinfo_mispredict & br_unit_brinfo_is_jr;
  assign _T_1538 = {br_unit_brinfo_mispredict,1'h0};
  assign _T_1539 = {_T_1538,icache_blocked};
  assign _T_1540 = {br_unit_brinfo_valid,rob_io_flush_valid};
  assign _T_1541 = {_T_1540,_T_1537};
  assign _T_1542 = {_T_1541,_T_1539};
  assign _GEN_14 = {{50'd0}, _T_1542};
  assign _T_1543 = _T_1526 & _GEN_14;
  assign _T_1545 = _T_1543 != 56'h0;
  assign _T_1546 = {io_dmem_perf_release,io_dmem_perf_acquire};
  assign _T_1547 = {_T_1546,io_imem_perf_acquire};
  assign _T_1548 = {1'h0,io_dmem_perf_tlbMiss};
  assign _T_1549 = {_T_1548,io_imem_perf_tlbMiss};
  assign _T_1550 = {_T_1549,_T_1547};
  assign _GEN_15 = {{50'd0}, _T_1550};
  assign _T_1551 = _T_1526 & _GEN_15;
  assign _T_1553 = _T_1551 != 56'h0;
  assign _T_1555 = _T_1525 == 2'h1;
  assign _T_1556 = _T_1555 ? _T_1545 : _T_1535;
  assign _T_1558 = _T_1525 == 2'h2;
  assign _T_1559 = _T_1558 ? _T_1553 : _T_1556;
  assign _T_1561 = _T_1525 == 2'h3;
  assign _T_1562 = _T_1561 ? _T_1553 : _T_1559;
  assign _T_1565 = csr_io_counters_1_eventSel[1:0];
  assign _T_1566 = csr_io_counters_1_eventSel[63:8];
  assign _T_1573 = _T_1566 & _GEN_13;
  assign _T_1575 = _T_1573 != 56'h0;
  assign _T_1583 = _T_1566 & _GEN_14;
  assign _T_1585 = _T_1583 != 56'h0;
  assign _T_1591 = _T_1566 & _GEN_15;
  assign _T_1593 = _T_1591 != 56'h0;
  assign _T_1595 = _T_1565 == 2'h1;
  assign _T_1596 = _T_1595 ? _T_1585 : _T_1575;
  assign _T_1598 = _T_1565 == 2'h2;
  assign _T_1599 = _T_1598 ? _T_1593 : _T_1596;
  assign _T_1601 = _T_1565 == 2'h3;
  assign _T_1602 = _T_1601 ? _T_1593 : _T_1599;
  assign _T_1605 = csr_io_counters_2_eventSel[1:0];
  assign _T_1606 = csr_io_counters_2_eventSel[63:8];
  assign _T_1613 = _T_1606 & _GEN_13;
  assign _T_1615 = _T_1613 != 56'h0;
  assign _T_1623 = _T_1606 & _GEN_14;
  assign _T_1625 = _T_1623 != 56'h0;
  assign _T_1631 = _T_1606 & _GEN_15;
  assign _T_1633 = _T_1631 != 56'h0;
  assign _T_1635 = _T_1605 == 2'h1;
  assign _T_1636 = _T_1635 ? _T_1625 : _T_1615;
  assign _T_1638 = _T_1605 == 2'h2;
  assign _T_1639 = _T_1638 ? _T_1633 : _T_1636;
  assign _T_1641 = _T_1605 == 2'h3;
  assign _T_1642 = _T_1641 ? _T_1633 : _T_1639;
  assign _T_1645 = csr_io_counters_3_eventSel[1:0];
  assign _T_1646 = csr_io_counters_3_eventSel[63:8];
  assign _T_1653 = _T_1646 & _GEN_13;
  assign _T_1655 = _T_1653 != 56'h0;
  assign _T_1663 = _T_1646 & _GEN_14;
  assign _T_1665 = _T_1663 != 56'h0;
  assign _T_1671 = _T_1646 & _GEN_15;
  assign _T_1673 = _T_1671 != 56'h0;
  assign _T_1675 = _T_1645 == 2'h1;
  assign _T_1676 = _T_1675 ? _T_1665 : _T_1655;
  assign _T_1678 = _T_1645 == 2'h2;
  assign _T_1679 = _T_1678 ? _T_1673 : _T_1676;
  assign _T_1681 = _T_1645 == 2'h3;
  assign _T_1682 = _T_1681 ? _T_1673 : _T_1679;
  assign _T_1685 = csr_io_counters_4_eventSel[1:0];
  assign _T_1686 = csr_io_counters_4_eventSel[63:8];
  assign _T_1693 = _T_1686 & _GEN_13;
  assign _T_1695 = _T_1693 != 56'h0;
  assign _T_1703 = _T_1686 & _GEN_14;
  assign _T_1705 = _T_1703 != 56'h0;
  assign _T_1711 = _T_1686 & _GEN_15;
  assign _T_1713 = _T_1711 != 56'h0;
  assign _T_1715 = _T_1685 == 2'h1;
  assign _T_1716 = _T_1715 ? _T_1705 : _T_1695;
  assign _T_1718 = _T_1685 == 2'h2;
  assign _T_1719 = _T_1718 ? _T_1713 : _T_1716;
  assign _T_1721 = _T_1685 == 2'h3;
  assign _T_1722 = _T_1721 ? _T_1713 : _T_1719;
  assign _T_1725 = csr_io_counters_5_eventSel[1:0];
  assign _T_1726 = csr_io_counters_5_eventSel[63:8];
  assign _T_1733 = _T_1726 & _GEN_13;
  assign _T_1735 = _T_1733 != 56'h0;
  assign _T_1743 = _T_1726 & _GEN_14;
  assign _T_1745 = _T_1743 != 56'h0;
  assign _T_1751 = _T_1726 & _GEN_15;
  assign _T_1753 = _T_1751 != 56'h0;
  assign _T_1755 = _T_1725 == 2'h1;
  assign _T_1756 = _T_1755 ? _T_1745 : _T_1735;
  assign _T_1758 = _T_1725 == 2'h2;
  assign _T_1759 = _T_1758 ? _T_1753 : _T_1756;
  assign _T_1761 = _T_1725 == 2'h3;
  assign _T_1762 = _T_1761 ? _T_1753 : _T_1759;
  assign _T_1765 = csr_io_counters_6_eventSel[1:0];
  assign _T_1766 = csr_io_counters_6_eventSel[63:8];
  assign _T_1773 = _T_1766 & _GEN_13;
  assign _T_1775 = _T_1773 != 56'h0;
  assign _T_1783 = _T_1766 & _GEN_14;
  assign _T_1785 = _T_1783 != 56'h0;
  assign _T_1791 = _T_1766 & _GEN_15;
  assign _T_1793 = _T_1791 != 56'h0;
  assign _T_1795 = _T_1765 == 2'h1;
  assign _T_1796 = _T_1795 ? _T_1785 : _T_1775;
  assign _T_1798 = _T_1765 == 2'h2;
  assign _T_1799 = _T_1798 ? _T_1793 : _T_1796;
  assign _T_1801 = _T_1765 == 2'h3;
  assign _T_1802 = _T_1801 ? _T_1793 : _T_1799;
  assign _T_1805 = csr_io_counters_7_eventSel[1:0];
  assign _T_1806 = csr_io_counters_7_eventSel[63:8];
  assign _T_1813 = _T_1806 & _GEN_13;
  assign _T_1815 = _T_1813 != 56'h0;
  assign _T_1823 = _T_1806 & _GEN_14;
  assign _T_1825 = _T_1823 != 56'h0;
  assign _T_1831 = _T_1806 & _GEN_15;
  assign _T_1833 = _T_1831 != 56'h0;
  assign _T_1835 = _T_1805 == 2'h1;
  assign _T_1836 = _T_1835 ? _T_1825 : _T_1815;
  assign _T_1838 = _T_1805 == 2'h2;
  assign _T_1839 = _T_1838 ? _T_1833 : _T_1836;
  assign _T_1841 = _T_1805 == 2'h3;
  assign _T_1842 = _T_1841 ? _T_1833 : _T_1839;
  assign _T_1845 = csr_io_counters_8_eventSel[1:0];
  assign _T_1846 = csr_io_counters_8_eventSel[63:8];
  assign _T_1853 = _T_1846 & _GEN_13;
  assign _T_1855 = _T_1853 != 56'h0;
  assign _T_1863 = _T_1846 & _GEN_14;
  assign _T_1865 = _T_1863 != 56'h0;
  assign _T_1871 = _T_1846 & _GEN_15;
  assign _T_1873 = _T_1871 != 56'h0;
  assign _T_1875 = _T_1845 == 2'h1;
  assign _T_1876 = _T_1875 ? _T_1865 : _T_1855;
  assign _T_1878 = _T_1845 == 2'h2;
  assign _T_1879 = _T_1878 ? _T_1873 : _T_1876;
  assign _T_1881 = _T_1845 == 2'h3;
  assign _T_1882 = _T_1881 ? _T_1873 : _T_1879;
  assign _T_1885 = csr_io_counters_9_eventSel[1:0];
  assign _T_1886 = csr_io_counters_9_eventSel[63:8];
  assign _T_1893 = _T_1886 & _GEN_13;
  assign _T_1895 = _T_1893 != 56'h0;
  assign _T_1903 = _T_1886 & _GEN_14;
  assign _T_1905 = _T_1903 != 56'h0;
  assign _T_1911 = _T_1886 & _GEN_15;
  assign _T_1913 = _T_1911 != 56'h0;
  assign _T_1915 = _T_1885 == 2'h1;
  assign _T_1916 = _T_1915 ? _T_1905 : _T_1895;
  assign _T_1918 = _T_1885 == 2'h2;
  assign _T_1919 = _T_1918 ? _T_1913 : _T_1916;
  assign _T_1921 = _T_1885 == 2'h3;
  assign _T_1922 = _T_1921 ? _T_1913 : _T_1919;
  assign _T_1925 = csr_io_counters_10_eventSel[1:0];
  assign _T_1926 = csr_io_counters_10_eventSel[63:8];
  assign _T_1933 = _T_1926 & _GEN_13;
  assign _T_1935 = _T_1933 != 56'h0;
  assign _T_1943 = _T_1926 & _GEN_14;
  assign _T_1945 = _T_1943 != 56'h0;
  assign _T_1951 = _T_1926 & _GEN_15;
  assign _T_1953 = _T_1951 != 56'h0;
  assign _T_1955 = _T_1925 == 2'h1;
  assign _T_1956 = _T_1955 ? _T_1945 : _T_1935;
  assign _T_1958 = _T_1925 == 2'h2;
  assign _T_1959 = _T_1958 ? _T_1953 : _T_1956;
  assign _T_1961 = _T_1925 == 2'h3;
  assign _T_1962 = _T_1961 ? _T_1953 : _T_1959;
  assign _T_1965 = csr_io_counters_11_eventSel[1:0];
  assign _T_1966 = csr_io_counters_11_eventSel[63:8];
  assign _T_1973 = _T_1966 & _GEN_13;
  assign _T_1975 = _T_1973 != 56'h0;
  assign _T_1983 = _T_1966 & _GEN_14;
  assign _T_1985 = _T_1983 != 56'h0;
  assign _T_1991 = _T_1966 & _GEN_15;
  assign _T_1993 = _T_1991 != 56'h0;
  assign _T_1995 = _T_1965 == 2'h1;
  assign _T_1996 = _T_1995 ? _T_1985 : _T_1975;
  assign _T_1998 = _T_1965 == 2'h2;
  assign _T_1999 = _T_1998 ? _T_1993 : _T_1996;
  assign _T_2001 = _T_1965 == 2'h3;
  assign _T_2002 = _T_2001 ? _T_1993 : _T_1999;
  assign _T_2005 = csr_io_counters_12_eventSel[1:0];
  assign _T_2006 = csr_io_counters_12_eventSel[63:8];
  assign _T_2013 = _T_2006 & _GEN_13;
  assign _T_2015 = _T_2013 != 56'h0;
  assign _T_2023 = _T_2006 & _GEN_14;
  assign _T_2025 = _T_2023 != 56'h0;
  assign _T_2031 = _T_2006 & _GEN_15;
  assign _T_2033 = _T_2031 != 56'h0;
  assign _T_2035 = _T_2005 == 2'h1;
  assign _T_2036 = _T_2035 ? _T_2025 : _T_2015;
  assign _T_2038 = _T_2005 == 2'h2;
  assign _T_2039 = _T_2038 ? _T_2033 : _T_2036;
  assign _T_2041 = _T_2005 == 2'h3;
  assign _T_2042 = _T_2041 ? _T_2033 : _T_2039;
  assign _T_2045 = csr_io_counters_13_eventSel[1:0];
  assign _T_2046 = csr_io_counters_13_eventSel[63:8];
  assign _T_2053 = _T_2046 & _GEN_13;
  assign _T_2055 = _T_2053 != 56'h0;
  assign _T_2063 = _T_2046 & _GEN_14;
  assign _T_2065 = _T_2063 != 56'h0;
  assign _T_2071 = _T_2046 & _GEN_15;
  assign _T_2073 = _T_2071 != 56'h0;
  assign _T_2075 = _T_2045 == 2'h1;
  assign _T_2076 = _T_2075 ? _T_2065 : _T_2055;
  assign _T_2078 = _T_2045 == 2'h2;
  assign _T_2079 = _T_2078 ? _T_2073 : _T_2076;
  assign _T_2081 = _T_2045 == 2'h3;
  assign _T_2082 = _T_2081 ? _T_2073 : _T_2079;
  assign _T_2085 = csr_io_counters_14_eventSel[1:0];
  assign _T_2086 = csr_io_counters_14_eventSel[63:8];
  assign _T_2093 = _T_2086 & _GEN_13;
  assign _T_2095 = _T_2093 != 56'h0;
  assign _T_2103 = _T_2086 & _GEN_14;
  assign _T_2105 = _T_2103 != 56'h0;
  assign _T_2111 = _T_2086 & _GEN_15;
  assign _T_2113 = _T_2111 != 56'h0;
  assign _T_2115 = _T_2085 == 2'h1;
  assign _T_2116 = _T_2115 ? _T_2105 : _T_2095;
  assign _T_2118 = _T_2085 == 2'h2;
  assign _T_2119 = _T_2118 ? _T_2113 : _T_2116;
  assign _T_2121 = _T_2085 == 2'h3;
  assign _T_2122 = _T_2121 ? _T_2113 : _T_2119;
  assign _T_2125 = csr_io_counters_15_eventSel[1:0];
  assign _T_2126 = csr_io_counters_15_eventSel[63:8];
  assign _T_2133 = _T_2126 & _GEN_13;
  assign _T_2135 = _T_2133 != 56'h0;
  assign _T_2143 = _T_2126 & _GEN_14;
  assign _T_2145 = _T_2143 != 56'h0;
  assign _T_2151 = _T_2126 & _GEN_15;
  assign _T_2153 = _T_2151 != 56'h0;
  assign _T_2155 = _T_2125 == 2'h1;
  assign _T_2156 = _T_2155 ? _T_2145 : _T_2135;
  assign _T_2158 = _T_2125 == 2'h2;
  assign _T_2159 = _T_2158 ? _T_2153 : _T_2156;
  assign _T_2161 = _T_2125 == 2'h3;
  assign _T_2162 = _T_2161 ? _T_2153 : _T_2159;
  assign _T_2165 = csr_io_counters_16_eventSel[1:0];
  assign _T_2166 = csr_io_counters_16_eventSel[63:8];
  assign _T_2173 = _T_2166 & _GEN_13;
  assign _T_2175 = _T_2173 != 56'h0;
  assign _T_2183 = _T_2166 & _GEN_14;
  assign _T_2185 = _T_2183 != 56'h0;
  assign _T_2191 = _T_2166 & _GEN_15;
  assign _T_2193 = _T_2191 != 56'h0;
  assign _T_2195 = _T_2165 == 2'h1;
  assign _T_2196 = _T_2195 ? _T_2185 : _T_2175;
  assign _T_2198 = _T_2165 == 2'h2;
  assign _T_2199 = _T_2198 ? _T_2193 : _T_2196;
  assign _T_2201 = _T_2165 == 2'h3;
  assign _T_2202 = _T_2201 ? _T_2193 : _T_2199;
  assign _T_2205 = csr_io_counters_17_eventSel[1:0];
  assign _T_2206 = csr_io_counters_17_eventSel[63:8];
  assign _T_2213 = _T_2206 & _GEN_13;
  assign _T_2215 = _T_2213 != 56'h0;
  assign _T_2223 = _T_2206 & _GEN_14;
  assign _T_2225 = _T_2223 != 56'h0;
  assign _T_2231 = _T_2206 & _GEN_15;
  assign _T_2233 = _T_2231 != 56'h0;
  assign _T_2235 = _T_2205 == 2'h1;
  assign _T_2236 = _T_2235 ? _T_2225 : _T_2215;
  assign _T_2238 = _T_2205 == 2'h2;
  assign _T_2239 = _T_2238 ? _T_2233 : _T_2236;
  assign _T_2241 = _T_2205 == 2'h3;
  assign _T_2242 = _T_2241 ? _T_2233 : _T_2239;
  assign _T_2245 = csr_io_counters_18_eventSel[1:0];
  assign _T_2246 = csr_io_counters_18_eventSel[63:8];
  assign _T_2253 = _T_2246 & _GEN_13;
  assign _T_2255 = _T_2253 != 56'h0;
  assign _T_2263 = _T_2246 & _GEN_14;
  assign _T_2265 = _T_2263 != 56'h0;
  assign _T_2271 = _T_2246 & _GEN_15;
  assign _T_2273 = _T_2271 != 56'h0;
  assign _T_2275 = _T_2245 == 2'h1;
  assign _T_2276 = _T_2275 ? _T_2265 : _T_2255;
  assign _T_2278 = _T_2245 == 2'h2;
  assign _T_2279 = _T_2278 ? _T_2273 : _T_2276;
  assign _T_2281 = _T_2245 == 2'h3;
  assign _T_2282 = _T_2281 ? _T_2273 : _T_2279;
  assign _T_2285 = csr_io_counters_19_eventSel[1:0];
  assign _T_2286 = csr_io_counters_19_eventSel[63:8];
  assign _T_2293 = _T_2286 & _GEN_13;
  assign _T_2295 = _T_2293 != 56'h0;
  assign _T_2303 = _T_2286 & _GEN_14;
  assign _T_2305 = _T_2303 != 56'h0;
  assign _T_2311 = _T_2286 & _GEN_15;
  assign _T_2313 = _T_2311 != 56'h0;
  assign _T_2315 = _T_2285 == 2'h1;
  assign _T_2316 = _T_2315 ? _T_2305 : _T_2295;
  assign _T_2318 = _T_2285 == 2'h2;
  assign _T_2319 = _T_2318 ? _T_2313 : _T_2316;
  assign _T_2321 = _T_2285 == 2'h3;
  assign _T_2322 = _T_2321 ? _T_2313 : _T_2319;
  assign _T_2325 = csr_io_counters_20_eventSel[1:0];
  assign _T_2326 = csr_io_counters_20_eventSel[63:8];
  assign _T_2333 = _T_2326 & _GEN_13;
  assign _T_2335 = _T_2333 != 56'h0;
  assign _T_2343 = _T_2326 & _GEN_14;
  assign _T_2345 = _T_2343 != 56'h0;
  assign _T_2351 = _T_2326 & _GEN_15;
  assign _T_2353 = _T_2351 != 56'h0;
  assign _T_2355 = _T_2325 == 2'h1;
  assign _T_2356 = _T_2355 ? _T_2345 : _T_2335;
  assign _T_2358 = _T_2325 == 2'h2;
  assign _T_2359 = _T_2358 ? _T_2353 : _T_2356;
  assign _T_2361 = _T_2325 == 2'h3;
  assign _T_2362 = _T_2361 ? _T_2353 : _T_2359;
  assign _T_2365 = csr_io_counters_21_eventSel[1:0];
  assign _T_2366 = csr_io_counters_21_eventSel[63:8];
  assign _T_2373 = _T_2366 & _GEN_13;
  assign _T_2375 = _T_2373 != 56'h0;
  assign _T_2383 = _T_2366 & _GEN_14;
  assign _T_2385 = _T_2383 != 56'h0;
  assign _T_2391 = _T_2366 & _GEN_15;
  assign _T_2393 = _T_2391 != 56'h0;
  assign _T_2395 = _T_2365 == 2'h1;
  assign _T_2396 = _T_2395 ? _T_2385 : _T_2375;
  assign _T_2398 = _T_2365 == 2'h2;
  assign _T_2399 = _T_2398 ? _T_2393 : _T_2396;
  assign _T_2401 = _T_2365 == 2'h3;
  assign _T_2402 = _T_2401 ? _T_2393 : _T_2399;
  assign _T_2405 = csr_io_counters_22_eventSel[1:0];
  assign _T_2406 = csr_io_counters_22_eventSel[63:8];
  assign _T_2413 = _T_2406 & _GEN_13;
  assign _T_2415 = _T_2413 != 56'h0;
  assign _T_2423 = _T_2406 & _GEN_14;
  assign _T_2425 = _T_2423 != 56'h0;
  assign _T_2431 = _T_2406 & _GEN_15;
  assign _T_2433 = _T_2431 != 56'h0;
  assign _T_2435 = _T_2405 == 2'h1;
  assign _T_2436 = _T_2435 ? _T_2425 : _T_2415;
  assign _T_2438 = _T_2405 == 2'h2;
  assign _T_2439 = _T_2438 ? _T_2433 : _T_2436;
  assign _T_2441 = _T_2405 == 2'h3;
  assign _T_2442 = _T_2441 ? _T_2433 : _T_2439;
  assign _T_2445 = csr_io_counters_23_eventSel[1:0];
  assign _T_2446 = csr_io_counters_23_eventSel[63:8];
  assign _T_2453 = _T_2446 & _GEN_13;
  assign _T_2455 = _T_2453 != 56'h0;
  assign _T_2463 = _T_2446 & _GEN_14;
  assign _T_2465 = _T_2463 != 56'h0;
  assign _T_2471 = _T_2446 & _GEN_15;
  assign _T_2473 = _T_2471 != 56'h0;
  assign _T_2475 = _T_2445 == 2'h1;
  assign _T_2476 = _T_2475 ? _T_2465 : _T_2455;
  assign _T_2478 = _T_2445 == 2'h2;
  assign _T_2479 = _T_2478 ? _T_2473 : _T_2476;
  assign _T_2481 = _T_2445 == 2'h3;
  assign _T_2482 = _T_2481 ? _T_2473 : _T_2479;
  assign _T_2485 = csr_io_counters_24_eventSel[1:0];
  assign _T_2486 = csr_io_counters_24_eventSel[63:8];
  assign _T_2493 = _T_2486 & _GEN_13;
  assign _T_2495 = _T_2493 != 56'h0;
  assign _T_2503 = _T_2486 & _GEN_14;
  assign _T_2505 = _T_2503 != 56'h0;
  assign _T_2511 = _T_2486 & _GEN_15;
  assign _T_2513 = _T_2511 != 56'h0;
  assign _T_2515 = _T_2485 == 2'h1;
  assign _T_2516 = _T_2515 ? _T_2505 : _T_2495;
  assign _T_2518 = _T_2485 == 2'h2;
  assign _T_2519 = _T_2518 ? _T_2513 : _T_2516;
  assign _T_2521 = _T_2485 == 2'h3;
  assign _T_2522 = _T_2521 ? _T_2513 : _T_2519;
  assign _T_2525 = csr_io_counters_25_eventSel[1:0];
  assign _T_2526 = csr_io_counters_25_eventSel[63:8];
  assign _T_2533 = _T_2526 & _GEN_13;
  assign _T_2535 = _T_2533 != 56'h0;
  assign _T_2543 = _T_2526 & _GEN_14;
  assign _T_2545 = _T_2543 != 56'h0;
  assign _T_2551 = _T_2526 & _GEN_15;
  assign _T_2553 = _T_2551 != 56'h0;
  assign _T_2555 = _T_2525 == 2'h1;
  assign _T_2556 = _T_2555 ? _T_2545 : _T_2535;
  assign _T_2558 = _T_2525 == 2'h2;
  assign _T_2559 = _T_2558 ? _T_2553 : _T_2556;
  assign _T_2561 = _T_2525 == 2'h3;
  assign _T_2562 = _T_2561 ? _T_2553 : _T_2559;
  assign _T_2565 = csr_io_counters_26_eventSel[1:0];
  assign _T_2566 = csr_io_counters_26_eventSel[63:8];
  assign _T_2573 = _T_2566 & _GEN_13;
  assign _T_2575 = _T_2573 != 56'h0;
  assign _T_2583 = _T_2566 & _GEN_14;
  assign _T_2585 = _T_2583 != 56'h0;
  assign _T_2591 = _T_2566 & _GEN_15;
  assign _T_2593 = _T_2591 != 56'h0;
  assign _T_2595 = _T_2565 == 2'h1;
  assign _T_2596 = _T_2595 ? _T_2585 : _T_2575;
  assign _T_2598 = _T_2565 == 2'h2;
  assign _T_2599 = _T_2598 ? _T_2593 : _T_2596;
  assign _T_2601 = _T_2565 == 2'h3;
  assign _T_2602 = _T_2601 ? _T_2593 : _T_2599;
  assign _T_2605 = csr_io_counters_27_eventSel[1:0];
  assign _T_2606 = csr_io_counters_27_eventSel[63:8];
  assign _T_2613 = _T_2606 & _GEN_13;
  assign _T_2615 = _T_2613 != 56'h0;
  assign _T_2623 = _T_2606 & _GEN_14;
  assign _T_2625 = _T_2623 != 56'h0;
  assign _T_2631 = _T_2606 & _GEN_15;
  assign _T_2633 = _T_2631 != 56'h0;
  assign _T_2635 = _T_2605 == 2'h1;
  assign _T_2636 = _T_2635 ? _T_2625 : _T_2615;
  assign _T_2638 = _T_2605 == 2'h2;
  assign _T_2639 = _T_2638 ? _T_2633 : _T_2636;
  assign _T_2641 = _T_2605 == 2'h3;
  assign _T_2642 = _T_2641 ? _T_2633 : _T_2639;
  assign _T_2645 = csr_io_counters_28_eventSel[1:0];
  assign _T_2646 = csr_io_counters_28_eventSel[63:8];
  assign _T_2653 = _T_2646 & _GEN_13;
  assign _T_2655 = _T_2653 != 56'h0;
  assign _T_2663 = _T_2646 & _GEN_14;
  assign _T_2665 = _T_2663 != 56'h0;
  assign _T_2671 = _T_2646 & _GEN_15;
  assign _T_2673 = _T_2671 != 56'h0;
  assign _T_2675 = _T_2645 == 2'h1;
  assign _T_2676 = _T_2675 ? _T_2665 : _T_2655;
  assign _T_2678 = _T_2645 == 2'h2;
  assign _T_2679 = _T_2678 ? _T_2673 : _T_2676;
  assign _T_2681 = _T_2645 == 2'h3;
  assign _T_2682 = _T_2681 ? _T_2673 : _T_2679;
  assign _T_2693 = debug_tsc_reg + 64'h1;
  assign _T_2694 = _T_2693[63:0];
  assign _T_2695 = {rob_io_commit_valids_1,rob_io_commit_valids_0};
  assign _T_2696 = _T_2695[0];
  assign _T_2697 = _T_2695[1];
  assign _T_2698 = _T_2696 + _T_2697;
  assign _GEN_100 = {{62'd0}, _T_2698};
  assign _T_2699 = debug_irt_reg + _GEN_100;
  assign _T_2700 = _T_2699[63:0];
  assign _T_2701 = br_unit_brinfo_mispredict | rob_io_flush_valid;
  assign _T_2702 = _T_2701 | fetch_unit_io_sfence_take_pc;
  assign _T_2705 = rob_io_flush_valid | _T_2704;
  assign _T_2706 = rob_io_commit_valids_0 & rob_io_commit_uops_0_is_fencei;
  assign _T_2707 = rob_io_commit_valids_1 & rob_io_commit_uops_1_is_fencei;
  assign _T_2708 = _T_2706 | _T_2707;
  assign _T_2710 = _T_1537 & csr_io_status_debug;
  assign _T_2711 = _T_2708 | _T_2710;
  assign _T_2731 = dec_serializer_io_deq_valid & dec_serializer_io_deq_bits_uops_0_valid;
  assign _T_2732 = dec_finished_mask[0];
  assign _T_2734 = _T_2732 == 1'h0;
  assign _T_2735 = _T_2731 & _T_2734;
  assign _T_2738 = rename_stage_io_inst_can_proceed_0 == 1'h0;
  assign _T_2739 = dec_valids_0 & dec_uops_0_is_unique;
  assign _T_2741 = rob_io_empty == 1'h0;
  assign _T_2743 = lsu_io_lsu_fencei_rdy == 1'h0;
  assign _T_2744 = _T_2741 | _T_2743;
  assign _T_2746 = _T_2739 & _T_2744;
  assign _T_2747 = _T_2738 | _T_2746;
  assign _T_2749 = rob_io_ready == 1'h0;
  assign _T_2750 = _T_2747 | _T_2749;
  assign _T_2751 = _T_2750 | lsu_io_laq_full;
  assign _T_2752 = _T_2751 | lsu_io_stq_full;
  assign _T_2753 = _T_2752 | branch_mask_full_0;
  assign _T_2754 = _T_2753 | br_unit_brinfo_mispredict;
  assign _T_2755 = _T_2754 | rob_io_flush_valid;
  assign _T_2758 = bpd_stage_io_brob_allocate_ready == 1'h0;
  assign _T_2759 = _T_2755 | _T_2758;
  assign _T_2760 = dec_valids_0 & dec_uops_0_is_fencei;
  assign _T_2763 = _T_2760 & _T_2743;
  assign _T_2764 = _T_2759 | _T_2763;
  assign _T_2765 = dec_valids_0 & _T_2764;
  assign _T_2768 = _T_2765 | _T_2739;
  assign _T_2770 = _T_2765 == 1'h0;
  assign _T_2771 = dec_valids_0 & _T_2770;
  assign _T_2773 = fetch_unit_io_clear_fetchbuffer == 1'h0;
  assign _T_2774 = _T_2771 & _T_2773;
  assign _T_2775 = dec_serializer_io_deq_valid & dec_serializer_io_deq_bits_uops_1_valid;
  assign _T_2776 = dec_finished_mask[1];
  assign _T_2778 = _T_2776 == 1'h0;
  assign _T_2779 = _T_2775 & _T_2778;
  assign _T_2783 = rename_stage_io_inst_can_proceed_1 == 1'h0;
  assign _T_2784 = dec_valids_1 & dec_uops_1_is_unique;
  assign _T_2790 = _T_2744 | dec_valids_0;
  assign _T_2791 = _T_2784 & _T_2790;
  assign _T_2792 = _T_2783 | _T_2791;
  assign _T_2795 = _T_2792 | _T_2749;
  assign _T_2796 = _T_2795 | lsu_io_laq_full;
  assign _T_2797 = _T_2796 | lsu_io_stq_full;
  assign _T_2798 = _T_2797 | branch_mask_full_1;
  assign _T_2799 = _T_2798 | br_unit_brinfo_mispredict;
  assign _T_2800 = _T_2799 | rob_io_flush_valid;
  assign _T_2801 = _T_2800 | _T_2768;
  assign _T_2804 = _T_2801 | _T_2758;
  assign _T_2805 = dec_valids_1 & dec_uops_1_is_fencei;
  assign _T_2808 = _T_2805 & _T_2743;
  assign _T_2809 = _T_2804 | _T_2808;
  assign _T_2810 = dec_valids_1 & _T_2809;
  assign dec_last_inst_was_stalled = _T_2810 | _T_2765;
  assign dec_stall_next_inst = dec_last_inst_was_stalled | _T_2784;
  assign _T_2813 = dec_last_inst_was_stalled == 1'h0;
  assign _T_2814 = dec_valids_1 & _T_2813;
  assign _T_2817 = _T_2814 & _T_2773;
  assign _T_2819 = dec_stall_next_inst == 1'h0;
  assign _T_2820 = dec_rdy | fetch_unit_io_clear_fetchbuffer;
  assign _T_2822 = {dec_will_fire_1,dec_will_fire_0};
  assign _T_2823 = _T_2822 | dec_finished_mask;
  assign _GEN_0 = _T_2820 ? 2'h0 : _T_2823;
  assign _T_2827 = _T_2734 & dec_uops_0_allocate_brtag;
  assign _T_2828 = dec_will_fire_0 & dec_uops_0_allocate_brtag;
  assign _T_2832 = _T_2778 & dec_uops_1_allocate_brtag;
  assign _T_2833 = dec_will_fire_1 & dec_uops_1_allocate_brtag;
  assign _T_2836 = dec_will_fire_0 & dec_uops_0_is_load;
  assign _T_2838 = new_ldq_idx + 4'h1;
  assign _T_2839 = _T_2838[3:0];
  assign _T_2841 = _T_2836 ? _T_2839 : new_ldq_idx;
  assign _T_2842 = dec_will_fire_0 & dec_uops_0_is_store;
  assign _T_2844 = new_stq_idx + 4'h1;
  assign _T_2845 = _T_2844[3:0];
  assign _T_2847 = _T_2842 ? _T_2845 : new_stq_idx;
  assign _T_2859 = {rob_io_curr_rob_tail,1'h0};
  assign _T_2861 = {rob_io_curr_rob_tail,1'h1};
  assign _T_2862 = dec_valids_0 & dec_uops_0_is_br_or_jmp;
  assign _T_2864 = dec_uops_0_is_jal == 1'h0;
  assign _T_2865 = _T_2862 & _T_2864;
  assign _T_2866 = dec_valids_1 & dec_uops_1_is_br_or_jmp;
  assign _T_2868 = dec_uops_1_is_jal == 1'h0;
  assign _T_2869 = _T_2866 & _T_2868;
  assign dec_has_br_or_jalr_in_packet = _T_2865 | _T_2869;
  assign _T_2870 = dec_will_fire_0 | dec_will_fire_1;
  assign _T_2872 = dec_finished_mask == 2'h0;
  assign _T_2873 = _T_2870 & _T_2872;
  assign _T_2874 = _T_2873 & dec_has_br_or_jalr_in_packet;
  assign _T_2882 = {issue_units_0_io_dis_readys_1,issue_units_0_io_dis_readys_0};
  assign _T_2883 = {issue_units_1_io_dis_readys_1,issue_units_1_io_dis_readys_0};
  assign _T_2884 = _T_2882 & _T_2883;
  assign _T_2885 = {fp_pipeline_io_dis_readys_1,fp_pipeline_io_dis_readys_0};
  assign dis_readys = _T_2884 & _T_2885;
  assign _T_2886 = dis_readys[0];
  assign _T_2887 = dis_readys[1];
  assign _T_2932 = ll_wbarb_io_out_ready & ll_wbarb_io_out_valid;
  assign _T_2933 = iss_valids_1 & iss_uops_1_bypassable;
  assign _T_2934 = iss_uops_1_dst_rtype == 2'h0;
  assign _T_2935 = _T_2933 & _T_2934;
  assign _T_2936 = _T_2935 & iss_uops_1_ldst_val;
  assign _T_2937 = iss_uops_1_dst_rtype == 2'h1;
  assign _T_2938 = _T_2937 & iss_uops_1_bypassable;
  assign _T_2940 = _T_2938 == 1'h0;
  assign _T_2942 = _T_2940 | reset;
  assign _T_2944 = _T_2942 == 1'h0;
  assign _T_2945 = csr_exe_unit_io_resp_0_valid & csr_exe_unit_io_resp_0_bits_uop_ctrl_rf_wen;
  assign _T_2947 = csr_exe_unit_io_resp_0_bits_uop_bypassable == 1'h0;
  assign _T_2948 = _T_2945 & _T_2947;
  assign _T_2949 = csr_exe_unit_io_resp_0_bits_uop_dst_rtype == 2'h0;
  assign _T_2950 = _T_2948 & _T_2949;
  assign _T_2951 = iss_valids_2 & iss_uops_2_bypassable;
  assign _T_2952 = iss_uops_2_dst_rtype == 2'h0;
  assign _T_2953 = _T_2951 & _T_2952;
  assign _T_2954 = _T_2953 & iss_uops_2_ldst_val;
  assign _T_2955 = iss_uops_2_dst_rtype == 2'h1;
  assign _T_2956 = _T_2955 & iss_uops_2_bypassable;
  assign _T_2958 = _T_2956 == 1'h0;
  assign _T_2960 = _T_2958 | reset;
  assign _T_2962 = _T_2960 == 1'h0;
  assign _T_2963 = ALUExeUnit_io_resp_0_valid & ALUExeUnit_io_resp_0_bits_uop_ctrl_rf_wen;
  assign _T_2965 = ALUExeUnit_io_resp_0_bits_uop_bypassable == 1'h0;
  assign _T_2966 = _T_2963 & _T_2965;
  assign _T_2967 = ALUExeUnit_io_resp_0_bits_uop_dst_rtype == 2'h0;
  assign _T_2968 = _T_2966 & _T_2967;
  assign _T_2979 = ~ br_unit_brinfo_mask;
  assign _T_2980 = rename_stage_io_ren2_uops_0_br_mask & _T_2979;
  assign _T_2981 = br_unit_brinfo_valid ? _T_2980 : rename_stage_io_ren2_uops_0_br_mask;
  assign _T_2993 = rename_stage_io_ren2_uops_1_br_mask & _T_2979;
  assign _T_2994 = br_unit_brinfo_valid ? _T_2993 : rename_stage_io_ren2_uops_1_br_mask;
  assign _T_2996 = dis_uops_0_iqtype == 2'h1;
  assign _T_2997 = dis_valids_0 & _T_2996;
  assign _T_2998 = dis_uops_0_uopc == 9'h2;
  assign _T_2999 = dis_uops_0_lrs2_rtype == 2'h1;
  assign _T_3000 = _T_2998 & _T_2999;
  assign _GEN_1 = _T_3000 ? 2'h2 : dis_uops_0_lrs2_rtype;
  assign _GEN_2 = _T_3000 ? 1'h0 : dis_uops_0_prs2_busy;
  assign _T_3003 = dis_uops_1_iqtype == 2'h1;
  assign _T_3004 = dis_valids_1 & _T_3003;
  assign _T_3005 = dis_uops_1_uopc == 9'h2;
  assign _T_3006 = dis_uops_1_lrs2_rtype == 2'h1;
  assign _T_3007 = _T_3005 & _T_3006;
  assign _GEN_3 = _T_3007 ? 2'h2 : dis_uops_1_lrs2_rtype;
  assign _GEN_4 = _T_3007 ? 1'h0 : dis_uops_1_prs2_busy;
  assign _T_3010 = dis_uops_0_iqtype == 2'h0;
  assign _T_3011 = dis_valids_0 & _T_3010;
  assign _T_3017 = dis_uops_1_iqtype == 2'h0;
  assign _T_3018 = dis_valids_1 & _T_3017;
  assign _T_3023 = iss_uops_1_fu_code == 10'h10;
  assign _T_3024 = iss_valids_1 & _T_3023;
  assign _T_3026 = _T_3024 ? 10'h10 : 10'h0;
  assign _T_3027 = ~ _T_3026;
  assign _T_3030 = csr_exe_unit_io_fu_types & _T_3029;
  assign _T_3033 = csr_exe_unit_io_resp_0_valid ? csr_exe_unit_io_resp_0_bits_uop_ctrl_csr_cmd : 3'h0;
  assign _T_3038 = iregister_read_io_exe_reqs_2_bits_uop_fu_code == 10'h100;
  assign _GEN_9 = _T_3038 ? 1'h0 : iregister_read_io_exe_reqs_2_valid;
  assign _T_3041 = iregister_read_io_exe_reqs_2_valid & _T_3038;
  assign _T_3042 = dec_will_fire_0 & rename_stage_io_inst_can_proceed_0;
  assign _T_3044 = rob_io_flush_valid == 1'h0;
  assign _T_3045 = _T_3042 & _T_3044;
  assign _T_3046 = _T_3045 & dec_uops_0_is_store;
  assign _T_3051 = _T_3045 & dec_uops_0_is_load;
  assign _T_3052 = dec_will_fire_1 & rename_stage_io_inst_can_proceed_1;
  assign _T_3055 = _T_3052 & _T_3044;
  assign _T_3056 = _T_3055 & dec_uops_1_is_store;
  assign _T_3061 = _T_3055 & dec_uops_1_is_load;
  assign _T_3064 = mem_unit_io_resp_0_valid & mem_unit_io_resp_0_bits_uop_ctrl_rf_wen;
  assign _T_3065 = mem_unit_io_resp_0_bits_uop_dst_rtype == 2'h0;
  assign _T_3066 = _T_3064 & _T_3065;
  assign _T_3067 = mem_unit_io_resp_0_bits_data[64];
  assign _T_3069 = _T_3066 & _T_3067;
  assign _T_3071 = _T_3069 == 1'h0;
  assign _T_3073 = _T_3071 | reset;
  assign _T_3075 = _T_3073 == 1'h0;
  assign _T_3077 = mem_unit_io_resp_0_bits_uop_dst_rtype == 2'h1;
  assign _T_3078 = _T_3064 & _T_3077;
  assign _T_3081 = mem_unit_io_resp_0_bits_uop_ctrl_rf_wen == 1'h0;
  assign _T_3082 = mem_unit_io_resp_0_valid & _T_3081;
  assign _T_3084 = _T_3082 & _T_3065;
  assign _T_3086 = _T_3084 == 1'h0;
  assign _T_3088 = _T_3086 | reset;
  assign _T_3090 = _T_3088 == 1'h0;
  assign _T_3092 = csr_exe_unit_io_resp_0_bits_uop_ctrl_csr_cmd != 3'h0;
  assign _T_3095 = _T_2945 & _T_2949;
  assign _T_3096 = _T_3092 ? csr_io_rw_rdata : csr_exe_unit_io_resp_0_bits_data;
  assign _T_3098 = csr_exe_unit_io_resp_0_bits_uop_dst_rtype == 2'h1;
  assign _T_3099 = _T_2945 & _T_3098;
  assign _T_3101 = _T_3099 == 1'h0;
  assign _T_3103 = _T_3101 | reset;
  assign _T_3105 = _T_3103 == 1'h0;
  assign _T_3107 = csr_exe_unit_io_resp_0_bits_uop_ctrl_rf_wen == 1'h0;
  assign _T_3108 = csr_exe_unit_io_resp_0_valid & _T_3107;
  assign _T_3110 = _T_3108 & _T_2949;
  assign _T_3112 = _T_3110 == 1'h0;
  assign _T_3114 = _T_3112 | reset;
  assign _T_3116 = _T_3114 == 1'h0;
  assign _T_3118 = csr_exe_unit_io_resp_0_bits_uop_dst_rtype != 2'h0;
  assign _T_3119 = _T_2945 & _T_3118;
  assign _T_3121 = _T_3119 == 1'h0;
  assign _T_3123 = _T_3121 | reset;
  assign _T_3125 = _T_3123 == 1'h0;
  assign _T_3130 = _T_2963 & _T_2967;
  assign _T_3132 = ALUExeUnit_io_resp_0_bits_uop_dst_rtype == 2'h1;
  assign _T_3133 = _T_2963 & _T_3132;
  assign _T_3135 = _T_3133 == 1'h0;
  assign _T_3137 = _T_3135 | reset;
  assign _T_3139 = _T_3137 == 1'h0;
  assign _T_3141 = ALUExeUnit_io_resp_0_bits_uop_ctrl_rf_wen == 1'h0;
  assign _T_3142 = ALUExeUnit_io_resp_0_valid & _T_3141;
  assign _T_3144 = _T_3142 & _T_2967;
  assign _T_3146 = _T_3144 == 1'h0;
  assign _T_3148 = _T_3146 | reset;
  assign _T_3150 = _T_3148 == 1'h0;
  assign _T_3152 = ALUExeUnit_io_resp_0_bits_uop_dst_rtype != 2'h0;
  assign _T_3153 = _T_2963 & _T_3152;
  assign _T_3155 = _T_3153 == 1'h0;
  assign _T_3157 = _T_3155 | reset;
  assign _T_3159 = _T_3157 == 1'h0;
  assign _T_3182 = dec_rdy == 1'h0;
  assign _T_3184 = dec_will_fire_1 == 1'h0;
  assign _T_3185 = _T_3182 & _T_3184;
  assign _T_3188 = dec_will_fire_0 == rename_stage_io_ren1_mask_0;
  assign _T_3189 = dec_will_fire_1 == rename_stage_io_ren1_mask_1;
  assign _T_3190 = _T_3188 | _T_3189;
  assign _T_3192 = _T_3190 | reset;
  assign _T_3194 = _T_3192 == 1'h0;
  assign _T_3196 = ll_wbarb_io_out_bits_uop_is_amo == 1'h0;
  assign _T_3197 = ll_wbarb_io_out_bits_uop_is_store & _T_3196;
  assign _T_3199 = _T_3197 == 1'h0;
  assign _T_3200 = ll_wbarb_io_out_valid & _T_3199;
  assign _T_3204 = mem_unit_io_resp_0_valid & mem_unit_io_resp_0_bits_uop_fp_val;
  assign _T_3206 = _T_3204 & _T_3077;
  assign _T_3207 = mem_unit_io_resp_0_bits_uop_uopc != 9'h1;
  assign _T_3208 = _T_3206 & _T_3207;
  assign _T_3210 = _T_3208 == 1'h0;
  assign _T_3212 = _T_3210 | reset;
  assign _T_3214 = _T_3212 == 1'h0;
  assign _T_3216 = csr_exe_unit_io_resp_0_bits_uop_is_amo == 1'h0;
  assign _T_3217 = csr_exe_unit_io_resp_0_bits_uop_is_store & _T_3216;
  assign _T_3219 = _T_3217 == 1'h0;
  assign _T_3220 = csr_exe_unit_io_resp_0_valid & _T_3219;
  assign _T_3228 = ALUExeUnit_io_resp_0_bits_uop_is_amo == 1'h0;
  assign _T_3229 = ALUExeUnit_io_resp_0_bits_uop_is_store & _T_3228;
  assign _T_3231 = _T_3229 == 1'h0;
  assign _T_3232 = ALUExeUnit_io_resp_0_valid & _T_3231;
  assign _T_3353 = fp_pipeline_io_wakeups_0_bits_uop_dst_rtype != 2'h1;
  assign _T_3354 = fp_pipeline_io_wakeups_0_valid & _T_3353;
  assign _T_3356 = _T_3354 == 1'h0;
  assign _T_3358 = _T_3356 | reset;
  assign _T_3360 = _T_3358 == 1'h0;
  assign _T_3362 = fp_pipeline_io_wakeups_0_bits_uop_fp_val == 1'h0;
  assign _T_3363 = fp_pipeline_io_wakeups_0_valid & _T_3362;
  assign _T_3365 = _T_3363 == 1'h0;
  assign _T_3367 = _T_3365 | reset;
  assign _T_3369 = _T_3367 == 1'h0;
  assign _T_3487 = fp_pipeline_io_wakeups_1_bits_uop_dst_rtype != 2'h1;
  assign _T_3488 = fp_pipeline_io_wakeups_1_valid & _T_3487;
  assign _T_3490 = _T_3488 == 1'h0;
  assign _T_3492 = _T_3490 | reset;
  assign _T_3494 = _T_3492 == 1'h0;
  assign _T_3496 = fp_pipeline_io_wakeups_1_bits_uop_fp_val == 1'h0;
  assign _T_3497 = fp_pipeline_io_wakeups_1_valid & _T_3496;
  assign _T_3499 = _T_3497 == 1'h0;
  assign _T_3501 = _T_3499 | reset;
  assign _T_3503 = _T_3501 == 1'h0;
  assign _T_3516 = csr_io_singleStep == 1'h0;
  assign _T_3518 = _T_3516 | reset;
  assign _T_3520 = _T_3518 == 1'h0;
  assign _T_3521 = rob_io_flush_valid | rob_io_clear_brob;
  assign _T_3526 = _T_3523 & _T_3044;
  assign _T_3528 = _T_3526 == 1'h0;
  assign _T_3530 = _T_3528 | reset;
  assign _T_3532 = _T_3530 == 1'h0;
  assign _T_3537 = _T_3536 + 5'h1;
  assign _T_3541 = _T_3537[5];
  assign _T_3543 = _T_3540 + 27'h1;
  assign _T_3544 = _T_3543[26:0];
  assign _GEN_10 = _T_3541 ? _T_3544 : _T_3540;
  assign _T_3545 = {_T_3540,_T_3536};
  assign _T_3548 = _T_2695 != 2'h0;
  assign _T_3549 = _T_3548 | csr_io_csr_stall;
  assign _T_3551 = _T_3549 | reset;
  assign _GEN_11 = _T_3551 ? 6'h0 : _T_3537;
  assign _GEN_12 = _T_3551 ? 27'h0 : _GEN_10;
  assign _T_3554 = _T_3545[13];
  assign _T_3556 = _T_3554 == 1'h0;
  assign _T_3558 = _T_3556 | reset;
  assign _T_3560 = _T_3558 == 1'h0;
  assign io_imem_req_valid = fetch_unit_io_imem_req_valid;
  assign io_imem_req_bits_pc = fetch_unit_io_imem_req_bits_pc;
  assign io_imem_req_bits_speculative = fetch_unit_io_imem_req_bits_speculative;
  assign io_imem_sfence_valid = _T_2715_valid;
  assign io_imem_sfence_bits_rs1 = _T_2715_bits_rs1;
  assign io_imem_sfence_bits_rs2 = _T_2715_bits_rs2;
  assign io_imem_sfence_bits_addr = _T_2715_bits_addr;
  assign io_imem_resp_ready = fetch_unit_io_imem_resp_ready;
  assign io_imem_flush_icache = _T_2711;
  assign io_dmem_req_valid = dc_shim_io_dmem_req_valid;
  assign io_dmem_req_bits_addr = dc_shim_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_tag = dc_shim_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_cmd = dc_shim_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_typ = dc_shim_io_dmem_req_bits_typ;
  assign io_dmem_s1_kill = dc_shim_io_dmem_s1_kill;
  assign io_dmem_s1_data_data = dc_shim_io_dmem_s1_data_data;
  assign io_dmem_invalidate_lr = dc_shim_io_dmem_invalidate_lr;
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_sfence_valid = io_imem_sfence_valid;
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1;
  assign io_ptw_status_dprv = csr_io_status_dprv;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_sum = csr_io_status_sum;
  assign io_ptw_tlb_req_valid = lsu_io_ptw_req_valid;
  assign io_ptw_tlb_req_bits_addr = lsu_io_ptw_req_bits_addr;
  assign mem_unit_io_req_valid = iregister_read_io_exe_reqs_0_valid;
  assign mem_unit_io_req_bits_uop_uopc = iregister_read_io_exe_reqs_0_bits_uop_uopc;
  assign mem_unit_io_req_bits_uop_ctrl_is_load = iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_load;
  assign mem_unit_io_req_bits_uop_ctrl_is_sta = iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_sta;
  assign mem_unit_io_req_bits_uop_ctrl_is_std = iregister_read_io_exe_reqs_0_bits_uop_ctrl_is_std;
  assign mem_unit_io_req_bits_uop_br_mask = iregister_read_io_exe_reqs_0_bits_uop_br_mask;
  assign mem_unit_io_req_bits_uop_imm_packed = iregister_read_io_exe_reqs_0_bits_uop_imm_packed;
  assign mem_unit_io_req_bits_uop_rob_idx = iregister_read_io_exe_reqs_0_bits_uop_rob_idx;
  assign mem_unit_io_req_bits_uop_ldq_idx = iregister_read_io_exe_reqs_0_bits_uop_ldq_idx;
  assign mem_unit_io_req_bits_uop_stq_idx = iregister_read_io_exe_reqs_0_bits_uop_stq_idx;
  assign mem_unit_io_req_bits_uop_pdst = iregister_read_io_exe_reqs_0_bits_uop_pdst;
  assign mem_unit_io_req_bits_uop_mem_cmd = iregister_read_io_exe_reqs_0_bits_uop_mem_cmd;
  assign mem_unit_io_req_bits_uop_mem_typ = iregister_read_io_exe_reqs_0_bits_uop_mem_typ;
  assign mem_unit_io_req_bits_uop_is_fence = iregister_read_io_exe_reqs_0_bits_uop_is_fence;
  assign mem_unit_io_req_bits_uop_is_store = iregister_read_io_exe_reqs_0_bits_uop_is_store;
  assign mem_unit_io_req_bits_uop_is_amo = iregister_read_io_exe_reqs_0_bits_uop_is_amo;
  assign mem_unit_io_req_bits_uop_is_load = iregister_read_io_exe_reqs_0_bits_uop_is_load;
  assign mem_unit_io_req_bits_uop_dst_rtype = iregister_read_io_exe_reqs_0_bits_uop_dst_rtype;
  assign mem_unit_io_req_bits_uop_fp_val = iregister_read_io_exe_reqs_0_bits_uop_fp_val;
  assign mem_unit_io_req_bits_rs1_data = {{1'd0}, iregister_read_io_exe_reqs_0_bits_rs1_data};
  assign mem_unit_io_req_bits_rs2_data = {{1'd0}, iregister_read_io_exe_reqs_0_bits_rs2_data};
  assign mem_unit_io_brinfo_valid = br_unit_brinfo_valid;
  assign mem_unit_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign mem_unit_io_brinfo_mask = br_unit_brinfo_mask;
  assign mem_unit_io_lsu_io_memreq_val = lsu_io_memreq_val;
  assign mem_unit_io_lsu_io_memreq_addr = lsu_io_memreq_addr;
  assign mem_unit_io_lsu_io_memreq_wdata = lsu_io_memreq_wdata;
  assign mem_unit_io_lsu_io_memreq_uop_uopc = lsu_io_memreq_uop_uopc;
  assign mem_unit_io_lsu_io_memreq_uop_br_mask = lsu_io_memreq_uop_br_mask;
  assign mem_unit_io_lsu_io_memreq_uop_rob_idx = lsu_io_memreq_uop_rob_idx;
  assign mem_unit_io_lsu_io_memreq_uop_ldq_idx = lsu_io_memreq_uop_ldq_idx;
  assign mem_unit_io_lsu_io_memreq_uop_stq_idx = lsu_io_memreq_uop_stq_idx;
  assign mem_unit_io_lsu_io_memreq_uop_pdst = lsu_io_memreq_uop_pdst;
  assign mem_unit_io_lsu_io_memreq_uop_mem_cmd = lsu_io_memreq_uop_mem_cmd;
  assign mem_unit_io_lsu_io_memreq_uop_mem_typ = lsu_io_memreq_uop_mem_typ;
  assign mem_unit_io_lsu_io_memreq_uop_is_store = lsu_io_memreq_uop_is_store;
  assign mem_unit_io_lsu_io_memreq_uop_is_amo = lsu_io_memreq_uop_is_amo;
  assign mem_unit_io_lsu_io_memreq_uop_is_load = lsu_io_memreq_uop_is_load;
  assign mem_unit_io_lsu_io_memreq_uop_dst_rtype = lsu_io_memreq_uop_dst_rtype;
  assign mem_unit_io_lsu_io_memreq_uop_fp_val = lsu_io_memreq_uop_fp_val;
  assign mem_unit_io_lsu_io_memreq_kill = lsu_io_memreq_kill;
  assign mem_unit_io_lsu_io_forward_val = lsu_io_forward_val;
  assign mem_unit_io_lsu_io_forward_data = lsu_io_forward_data;
  assign mem_unit_io_lsu_io_forward_uop_uopc = lsu_io_forward_uop_uopc;
  assign mem_unit_io_lsu_io_forward_uop_rob_idx = lsu_io_forward_uop_rob_idx;
  assign mem_unit_io_lsu_io_forward_uop_ldq_idx = lsu_io_forward_uop_ldq_idx;
  assign mem_unit_io_lsu_io_forward_uop_stq_idx = lsu_io_forward_uop_stq_idx;
  assign mem_unit_io_lsu_io_forward_uop_pdst = lsu_io_forward_uop_pdst;
  assign mem_unit_io_lsu_io_forward_uop_mem_typ = lsu_io_forward_uop_mem_typ;
  assign mem_unit_io_lsu_io_forward_uop_is_store = lsu_io_forward_uop_is_store;
  assign mem_unit_io_lsu_io_forward_uop_is_amo = lsu_io_forward_uop_is_amo;
  assign mem_unit_io_lsu_io_forward_uop_is_load = lsu_io_forward_uop_is_load;
  assign mem_unit_io_lsu_io_forward_uop_dst_rtype = lsu_io_forward_uop_dst_rtype;
  assign mem_unit_io_lsu_io_forward_uop_fp_val = lsu_io_forward_uop_fp_val;
  assign mem_unit_io_dmem_resp_valid = dc_shim_io_core_resp_valid;
  assign mem_unit_io_dmem_resp_bits_data_subword = dc_shim_io_core_resp_bits_data_subword;
  assign mem_unit_io_dmem_resp_bits_uop_uopc = dc_shim_io_core_resp_bits_uop_uopc;
  assign mem_unit_io_dmem_resp_bits_uop_rob_idx = dc_shim_io_core_resp_bits_uop_rob_idx;
  assign mem_unit_io_dmem_resp_bits_uop_ldq_idx = dc_shim_io_core_resp_bits_uop_ldq_idx;
  assign mem_unit_io_dmem_resp_bits_uop_stq_idx = dc_shim_io_core_resp_bits_uop_stq_idx;
  assign mem_unit_io_dmem_resp_bits_uop_pdst = dc_shim_io_core_resp_bits_uop_pdst;
  assign mem_unit_io_dmem_resp_bits_uop_mem_cmd = dc_shim_io_core_resp_bits_uop_mem_cmd;
  assign mem_unit_io_dmem_resp_bits_uop_mem_typ = dc_shim_io_core_resp_bits_uop_mem_typ;
  assign mem_unit_io_dmem_resp_bits_uop_is_store = dc_shim_io_core_resp_bits_uop_is_store;
  assign mem_unit_io_dmem_resp_bits_uop_is_amo = dc_shim_io_core_resp_bits_uop_is_amo;
  assign mem_unit_io_dmem_resp_bits_uop_is_load = dc_shim_io_core_resp_bits_uop_is_load;
  assign mem_unit_io_dmem_resp_bits_uop_dst_rtype = dc_shim_io_core_resp_bits_uop_dst_rtype;
  assign mem_unit_io_dmem_resp_bits_uop_fp_val = dc_shim_io_core_resp_bits_uop_fp_val;
  assign mem_unit_io_com_exception = rob_io_flush_valid;
  assign mem_unit_clock = clock;
  assign mem_unit_reset = reset;
  assign csr_exe_unit_io_req_valid = iregister_read_io_exe_reqs_1_valid;
  assign csr_exe_unit_io_req_bits_uop_valid = iregister_read_io_exe_reqs_1_bits_uop_valid;
  assign csr_exe_unit_io_req_bits_uop_iw_state = iregister_read_io_exe_reqs_1_bits_uop_iw_state;
  assign csr_exe_unit_io_req_bits_uop_uopc = iregister_read_io_exe_reqs_1_bits_uop_uopc;
  assign csr_exe_unit_io_req_bits_uop_inst = iregister_read_io_exe_reqs_1_bits_uop_inst;
  assign csr_exe_unit_io_req_bits_uop_pc = iregister_read_io_exe_reqs_1_bits_uop_pc;
  assign csr_exe_unit_io_req_bits_uop_iqtype = iregister_read_io_exe_reqs_1_bits_uop_iqtype;
  assign csr_exe_unit_io_req_bits_uop_fu_code = iregister_read_io_exe_reqs_1_bits_uop_fu_code;
  assign csr_exe_unit_io_req_bits_uop_ctrl_br_type = iregister_read_io_exe_reqs_1_bits_uop_ctrl_br_type;
  assign csr_exe_unit_io_req_bits_uop_ctrl_op1_sel = iregister_read_io_exe_reqs_1_bits_uop_ctrl_op1_sel;
  assign csr_exe_unit_io_req_bits_uop_ctrl_op2_sel = iregister_read_io_exe_reqs_1_bits_uop_ctrl_op2_sel;
  assign csr_exe_unit_io_req_bits_uop_ctrl_imm_sel = iregister_read_io_exe_reqs_1_bits_uop_ctrl_imm_sel;
  assign csr_exe_unit_io_req_bits_uop_ctrl_op_fcn = iregister_read_io_exe_reqs_1_bits_uop_ctrl_op_fcn;
  assign csr_exe_unit_io_req_bits_uop_ctrl_fcn_dw = iregister_read_io_exe_reqs_1_bits_uop_ctrl_fcn_dw;
  assign csr_exe_unit_io_req_bits_uop_ctrl_rf_wen = iregister_read_io_exe_reqs_1_bits_uop_ctrl_rf_wen;
  assign csr_exe_unit_io_req_bits_uop_ctrl_csr_cmd = iregister_read_io_exe_reqs_1_bits_uop_ctrl_csr_cmd;
  assign csr_exe_unit_io_req_bits_uop_ctrl_is_load = iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_load;
  assign csr_exe_unit_io_req_bits_uop_ctrl_is_sta = iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_sta;
  assign csr_exe_unit_io_req_bits_uop_ctrl_is_std = iregister_read_io_exe_reqs_1_bits_uop_ctrl_is_std;
  assign csr_exe_unit_io_req_bits_uop_allocate_brtag = iregister_read_io_exe_reqs_1_bits_uop_allocate_brtag;
  assign csr_exe_unit_io_req_bits_uop_is_br_or_jmp = iregister_read_io_exe_reqs_1_bits_uop_is_br_or_jmp;
  assign csr_exe_unit_io_req_bits_uop_is_jump = iregister_read_io_exe_reqs_1_bits_uop_is_jump;
  assign csr_exe_unit_io_req_bits_uop_is_jal = iregister_read_io_exe_reqs_1_bits_uop_is_jal;
  assign csr_exe_unit_io_req_bits_uop_is_ret = iregister_read_io_exe_reqs_1_bits_uop_is_ret;
  assign csr_exe_unit_io_req_bits_uop_is_call = iregister_read_io_exe_reqs_1_bits_uop_is_call;
  assign csr_exe_unit_io_req_bits_uop_br_mask = iregister_read_io_exe_reqs_1_bits_uop_br_mask;
  assign csr_exe_unit_io_req_bits_uop_br_tag = iregister_read_io_exe_reqs_1_bits_uop_br_tag;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_btb_blame = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_blame;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_btb_hit = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_hit;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_btb_taken = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_btb_taken;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_blame = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_blame;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_hit = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_hit;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_taken = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_taken;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_value = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_value;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_entry_idx = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_entry_idx;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bim_resp_way_idx = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bim_resp_way_idx;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_takens = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_takens;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_u = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_u;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_history_ptr;
  assign csr_exe_unit_io_req_bits_uop_br_prediction_bpd_resp_info = iregister_read_io_exe_reqs_1_bits_uop_br_prediction_bpd_resp_info;
  assign csr_exe_unit_io_req_bits_uop_stat_brjmp_mispredicted = iregister_read_io_exe_reqs_1_bits_uop_stat_brjmp_mispredicted;
  assign csr_exe_unit_io_req_bits_uop_stat_btb_made_pred = iregister_read_io_exe_reqs_1_bits_uop_stat_btb_made_pred;
  assign csr_exe_unit_io_req_bits_uop_stat_btb_mispredicted = iregister_read_io_exe_reqs_1_bits_uop_stat_btb_mispredicted;
  assign csr_exe_unit_io_req_bits_uop_stat_bpd_made_pred = iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_made_pred;
  assign csr_exe_unit_io_req_bits_uop_stat_bpd_mispredicted = iregister_read_io_exe_reqs_1_bits_uop_stat_bpd_mispredicted;
  assign csr_exe_unit_io_req_bits_uop_fetch_pc_lob = iregister_read_io_exe_reqs_1_bits_uop_fetch_pc_lob;
  assign csr_exe_unit_io_req_bits_uop_imm_packed = iregister_read_io_exe_reqs_1_bits_uop_imm_packed;
  assign csr_exe_unit_io_req_bits_uop_csr_addr = iregister_read_io_exe_reqs_1_bits_uop_csr_addr;
  assign csr_exe_unit_io_req_bits_uop_rob_idx = iregister_read_io_exe_reqs_1_bits_uop_rob_idx;
  assign csr_exe_unit_io_req_bits_uop_ldq_idx = iregister_read_io_exe_reqs_1_bits_uop_ldq_idx;
  assign csr_exe_unit_io_req_bits_uop_stq_idx = iregister_read_io_exe_reqs_1_bits_uop_stq_idx;
  assign csr_exe_unit_io_req_bits_uop_brob_idx = iregister_read_io_exe_reqs_1_bits_uop_brob_idx;
  assign csr_exe_unit_io_req_bits_uop_pdst = iregister_read_io_exe_reqs_1_bits_uop_pdst;
  assign csr_exe_unit_io_req_bits_uop_pop1 = iregister_read_io_exe_reqs_1_bits_uop_pop1;
  assign csr_exe_unit_io_req_bits_uop_pop2 = iregister_read_io_exe_reqs_1_bits_uop_pop2;
  assign csr_exe_unit_io_req_bits_uop_pop3 = iregister_read_io_exe_reqs_1_bits_uop_pop3;
  assign csr_exe_unit_io_req_bits_uop_prs1_busy = iregister_read_io_exe_reqs_1_bits_uop_prs1_busy;
  assign csr_exe_unit_io_req_bits_uop_prs2_busy = iregister_read_io_exe_reqs_1_bits_uop_prs2_busy;
  assign csr_exe_unit_io_req_bits_uop_prs3_busy = iregister_read_io_exe_reqs_1_bits_uop_prs3_busy;
  assign csr_exe_unit_io_req_bits_uop_stale_pdst = iregister_read_io_exe_reqs_1_bits_uop_stale_pdst;
  assign csr_exe_unit_io_req_bits_uop_exception = iregister_read_io_exe_reqs_1_bits_uop_exception;
  assign csr_exe_unit_io_req_bits_uop_exc_cause = iregister_read_io_exe_reqs_1_bits_uop_exc_cause;
  assign csr_exe_unit_io_req_bits_uop_bypassable = iregister_read_io_exe_reqs_1_bits_uop_bypassable;
  assign csr_exe_unit_io_req_bits_uop_mem_cmd = iregister_read_io_exe_reqs_1_bits_uop_mem_cmd;
  assign csr_exe_unit_io_req_bits_uop_mem_typ = iregister_read_io_exe_reqs_1_bits_uop_mem_typ;
  assign csr_exe_unit_io_req_bits_uop_is_fence = iregister_read_io_exe_reqs_1_bits_uop_is_fence;
  assign csr_exe_unit_io_req_bits_uop_is_fencei = iregister_read_io_exe_reqs_1_bits_uop_is_fencei;
  assign csr_exe_unit_io_req_bits_uop_is_store = iregister_read_io_exe_reqs_1_bits_uop_is_store;
  assign csr_exe_unit_io_req_bits_uop_is_amo = iregister_read_io_exe_reqs_1_bits_uop_is_amo;
  assign csr_exe_unit_io_req_bits_uop_is_load = iregister_read_io_exe_reqs_1_bits_uop_is_load;
  assign csr_exe_unit_io_req_bits_uop_is_sys_pc2epc = iregister_read_io_exe_reqs_1_bits_uop_is_sys_pc2epc;
  assign csr_exe_unit_io_req_bits_uop_is_unique = iregister_read_io_exe_reqs_1_bits_uop_is_unique;
  assign csr_exe_unit_io_req_bits_uop_flush_on_commit = iregister_read_io_exe_reqs_1_bits_uop_flush_on_commit;
  assign csr_exe_unit_io_req_bits_uop_ldst = iregister_read_io_exe_reqs_1_bits_uop_ldst;
  assign csr_exe_unit_io_req_bits_uop_lrs1 = iregister_read_io_exe_reqs_1_bits_uop_lrs1;
  assign csr_exe_unit_io_req_bits_uop_lrs2 = iregister_read_io_exe_reqs_1_bits_uop_lrs2;
  assign csr_exe_unit_io_req_bits_uop_lrs3 = iregister_read_io_exe_reqs_1_bits_uop_lrs3;
  assign csr_exe_unit_io_req_bits_uop_ldst_val = iregister_read_io_exe_reqs_1_bits_uop_ldst_val;
  assign csr_exe_unit_io_req_bits_uop_dst_rtype = iregister_read_io_exe_reqs_1_bits_uop_dst_rtype;
  assign csr_exe_unit_io_req_bits_uop_lrs1_rtype = iregister_read_io_exe_reqs_1_bits_uop_lrs1_rtype;
  assign csr_exe_unit_io_req_bits_uop_lrs2_rtype = iregister_read_io_exe_reqs_1_bits_uop_lrs2_rtype;
  assign csr_exe_unit_io_req_bits_uop_frs3_en = iregister_read_io_exe_reqs_1_bits_uop_frs3_en;
  assign csr_exe_unit_io_req_bits_uop_fp_val = iregister_read_io_exe_reqs_1_bits_uop_fp_val;
  assign csr_exe_unit_io_req_bits_uop_fp_single = iregister_read_io_exe_reqs_1_bits_uop_fp_single;
  assign csr_exe_unit_io_req_bits_uop_xcpt_pf_if = iregister_read_io_exe_reqs_1_bits_uop_xcpt_pf_if;
  assign csr_exe_unit_io_req_bits_uop_xcpt_ae_if = iregister_read_io_exe_reqs_1_bits_uop_xcpt_ae_if;
  assign csr_exe_unit_io_req_bits_uop_replay_if = iregister_read_io_exe_reqs_1_bits_uop_replay_if;
  assign csr_exe_unit_io_req_bits_uop_xcpt_ma_if = iregister_read_io_exe_reqs_1_bits_uop_xcpt_ma_if;
  assign csr_exe_unit_io_req_bits_uop_debug_wdata = iregister_read_io_exe_reqs_1_bits_uop_debug_wdata;
  assign csr_exe_unit_io_req_bits_uop_debug_events_fetch_seq = iregister_read_io_exe_reqs_1_bits_uop_debug_events_fetch_seq;
  assign csr_exe_unit_io_req_bits_rs1_data = iregister_read_io_exe_reqs_1_bits_rs1_data;
  assign csr_exe_unit_io_req_bits_rs2_data = iregister_read_io_exe_reqs_1_bits_rs2_data;
  assign csr_exe_unit_io_req_bits_kill = rob_io_flush_valid;
  assign csr_exe_unit_io_brinfo_valid = br_unit_brinfo_valid;
  assign csr_exe_unit_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign csr_exe_unit_io_brinfo_mask = br_unit_brinfo_mask;
  assign csr_exe_unit_io_get_rob_pc_curr_pc = _T_3507;
  assign csr_exe_unit_io_get_rob_pc_curr_brob_idx = _T_3509;
  assign csr_exe_unit_io_get_rob_pc_next_val = _T_3511;
  assign csr_exe_unit_io_get_rob_pc_next_pc = _T_3513;
  assign csr_exe_unit_io_get_pred_info_bim_resp_value = _T_2928_bim_resp_value;
  assign csr_exe_unit_io_get_pred_info_bim_resp_entry_idx = _T_2928_bim_resp_entry_idx;
  assign csr_exe_unit_io_get_pred_info_bim_resp_way_idx = _T_2928_bim_resp_way_idx;
  assign csr_exe_unit_io_get_pred_info_bpd_resp_history = _T_2928_bpd_resp_history;
  assign csr_exe_unit_io_get_pred_info_bpd_resp_history_ptr = _T_2928_bpd_resp_history_ptr;
  assign csr_exe_unit_io_status_debug = csr_io_status_debug;
  assign csr_exe_unit_clock = clock;
  assign csr_exe_unit_reset = reset;
  assign ALUExeUnit_io_req_valid = _GEN_9;
  assign ALUExeUnit_io_req_bits_uop_valid = iregister_read_io_exe_reqs_2_bits_uop_valid;
  assign ALUExeUnit_io_req_bits_uop_iw_state = iregister_read_io_exe_reqs_2_bits_uop_iw_state;
  assign ALUExeUnit_io_req_bits_uop_uopc = iregister_read_io_exe_reqs_2_bits_uop_uopc;
  assign ALUExeUnit_io_req_bits_uop_inst = iregister_read_io_exe_reqs_2_bits_uop_inst;
  assign ALUExeUnit_io_req_bits_uop_pc = iregister_read_io_exe_reqs_2_bits_uop_pc;
  assign ALUExeUnit_io_req_bits_uop_iqtype = iregister_read_io_exe_reqs_2_bits_uop_iqtype;
  assign ALUExeUnit_io_req_bits_uop_fu_code = iregister_read_io_exe_reqs_2_bits_uop_fu_code;
  assign ALUExeUnit_io_req_bits_uop_ctrl_op1_sel = iregister_read_io_exe_reqs_2_bits_uop_ctrl_op1_sel;
  assign ALUExeUnit_io_req_bits_uop_ctrl_op2_sel = iregister_read_io_exe_reqs_2_bits_uop_ctrl_op2_sel;
  assign ALUExeUnit_io_req_bits_uop_ctrl_imm_sel = iregister_read_io_exe_reqs_2_bits_uop_ctrl_imm_sel;
  assign ALUExeUnit_io_req_bits_uop_ctrl_op_fcn = iregister_read_io_exe_reqs_2_bits_uop_ctrl_op_fcn;
  assign ALUExeUnit_io_req_bits_uop_ctrl_fcn_dw = iregister_read_io_exe_reqs_2_bits_uop_ctrl_fcn_dw;
  assign ALUExeUnit_io_req_bits_uop_ctrl_rf_wen = iregister_read_io_exe_reqs_2_bits_uop_ctrl_rf_wen;
  assign ALUExeUnit_io_req_bits_uop_ctrl_is_load = iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_load;
  assign ALUExeUnit_io_req_bits_uop_ctrl_is_sta = iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_sta;
  assign ALUExeUnit_io_req_bits_uop_ctrl_is_std = iregister_read_io_exe_reqs_2_bits_uop_ctrl_is_std;
  assign ALUExeUnit_io_req_bits_uop_allocate_brtag = iregister_read_io_exe_reqs_2_bits_uop_allocate_brtag;
  assign ALUExeUnit_io_req_bits_uop_is_br_or_jmp = iregister_read_io_exe_reqs_2_bits_uop_is_br_or_jmp;
  assign ALUExeUnit_io_req_bits_uop_is_jump = iregister_read_io_exe_reqs_2_bits_uop_is_jump;
  assign ALUExeUnit_io_req_bits_uop_is_jal = iregister_read_io_exe_reqs_2_bits_uop_is_jal;
  assign ALUExeUnit_io_req_bits_uop_is_ret = iregister_read_io_exe_reqs_2_bits_uop_is_ret;
  assign ALUExeUnit_io_req_bits_uop_is_call = iregister_read_io_exe_reqs_2_bits_uop_is_call;
  assign ALUExeUnit_io_req_bits_uop_br_mask = iregister_read_io_exe_reqs_2_bits_uop_br_mask;
  assign ALUExeUnit_io_req_bits_uop_br_tag = iregister_read_io_exe_reqs_2_bits_uop_br_tag;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_btb_blame = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_blame;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_btb_hit = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_hit;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_btb_taken = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_btb_taken;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_blame = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_blame;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_hit = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_hit;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_taken = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_taken;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_value = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_value;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_entry_idx = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_entry_idx;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bim_resp_way_idx = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bim_resp_way_idx;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_takens = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_takens;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_u = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_u;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_history_ptr = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_history_ptr;
  assign ALUExeUnit_io_req_bits_uop_br_prediction_bpd_resp_info = iregister_read_io_exe_reqs_2_bits_uop_br_prediction_bpd_resp_info;
  assign ALUExeUnit_io_req_bits_uop_stat_brjmp_mispredicted = iregister_read_io_exe_reqs_2_bits_uop_stat_brjmp_mispredicted;
  assign ALUExeUnit_io_req_bits_uop_stat_btb_made_pred = iregister_read_io_exe_reqs_2_bits_uop_stat_btb_made_pred;
  assign ALUExeUnit_io_req_bits_uop_stat_btb_mispredicted = iregister_read_io_exe_reqs_2_bits_uop_stat_btb_mispredicted;
  assign ALUExeUnit_io_req_bits_uop_stat_bpd_made_pred = iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_made_pred;
  assign ALUExeUnit_io_req_bits_uop_stat_bpd_mispredicted = iregister_read_io_exe_reqs_2_bits_uop_stat_bpd_mispredicted;
  assign ALUExeUnit_io_req_bits_uop_fetch_pc_lob = iregister_read_io_exe_reqs_2_bits_uop_fetch_pc_lob;
  assign ALUExeUnit_io_req_bits_uop_imm_packed = iregister_read_io_exe_reqs_2_bits_uop_imm_packed;
  assign ALUExeUnit_io_req_bits_uop_csr_addr = iregister_read_io_exe_reqs_2_bits_uop_csr_addr;
  assign ALUExeUnit_io_req_bits_uop_rob_idx = iregister_read_io_exe_reqs_2_bits_uop_rob_idx;
  assign ALUExeUnit_io_req_bits_uop_ldq_idx = iregister_read_io_exe_reqs_2_bits_uop_ldq_idx;
  assign ALUExeUnit_io_req_bits_uop_stq_idx = iregister_read_io_exe_reqs_2_bits_uop_stq_idx;
  assign ALUExeUnit_io_req_bits_uop_brob_idx = iregister_read_io_exe_reqs_2_bits_uop_brob_idx;
  assign ALUExeUnit_io_req_bits_uop_pdst = iregister_read_io_exe_reqs_2_bits_uop_pdst;
  assign ALUExeUnit_io_req_bits_uop_pop1 = iregister_read_io_exe_reqs_2_bits_uop_pop1;
  assign ALUExeUnit_io_req_bits_uop_pop2 = iregister_read_io_exe_reqs_2_bits_uop_pop2;
  assign ALUExeUnit_io_req_bits_uop_pop3 = iregister_read_io_exe_reqs_2_bits_uop_pop3;
  assign ALUExeUnit_io_req_bits_uop_prs1_busy = iregister_read_io_exe_reqs_2_bits_uop_prs1_busy;
  assign ALUExeUnit_io_req_bits_uop_prs2_busy = iregister_read_io_exe_reqs_2_bits_uop_prs2_busy;
  assign ALUExeUnit_io_req_bits_uop_prs3_busy = iregister_read_io_exe_reqs_2_bits_uop_prs3_busy;
  assign ALUExeUnit_io_req_bits_uop_stale_pdst = iregister_read_io_exe_reqs_2_bits_uop_stale_pdst;
  assign ALUExeUnit_io_req_bits_uop_exception = iregister_read_io_exe_reqs_2_bits_uop_exception;
  assign ALUExeUnit_io_req_bits_uop_exc_cause = iregister_read_io_exe_reqs_2_bits_uop_exc_cause;
  assign ALUExeUnit_io_req_bits_uop_bypassable = iregister_read_io_exe_reqs_2_bits_uop_bypassable;
  assign ALUExeUnit_io_req_bits_uop_mem_cmd = iregister_read_io_exe_reqs_2_bits_uop_mem_cmd;
  assign ALUExeUnit_io_req_bits_uop_mem_typ = iregister_read_io_exe_reqs_2_bits_uop_mem_typ;
  assign ALUExeUnit_io_req_bits_uop_is_fence = iregister_read_io_exe_reqs_2_bits_uop_is_fence;
  assign ALUExeUnit_io_req_bits_uop_is_fencei = iregister_read_io_exe_reqs_2_bits_uop_is_fencei;
  assign ALUExeUnit_io_req_bits_uop_is_store = iregister_read_io_exe_reqs_2_bits_uop_is_store;
  assign ALUExeUnit_io_req_bits_uop_is_amo = iregister_read_io_exe_reqs_2_bits_uop_is_amo;
  assign ALUExeUnit_io_req_bits_uop_is_load = iregister_read_io_exe_reqs_2_bits_uop_is_load;
  assign ALUExeUnit_io_req_bits_uop_is_sys_pc2epc = iregister_read_io_exe_reqs_2_bits_uop_is_sys_pc2epc;
  assign ALUExeUnit_io_req_bits_uop_is_unique = iregister_read_io_exe_reqs_2_bits_uop_is_unique;
  assign ALUExeUnit_io_req_bits_uop_flush_on_commit = iregister_read_io_exe_reqs_2_bits_uop_flush_on_commit;
  assign ALUExeUnit_io_req_bits_uop_ldst = iregister_read_io_exe_reqs_2_bits_uop_ldst;
  assign ALUExeUnit_io_req_bits_uop_lrs1 = iregister_read_io_exe_reqs_2_bits_uop_lrs1;
  assign ALUExeUnit_io_req_bits_uop_lrs2 = iregister_read_io_exe_reqs_2_bits_uop_lrs2;
  assign ALUExeUnit_io_req_bits_uop_lrs3 = iregister_read_io_exe_reqs_2_bits_uop_lrs3;
  assign ALUExeUnit_io_req_bits_uop_ldst_val = iregister_read_io_exe_reqs_2_bits_uop_ldst_val;
  assign ALUExeUnit_io_req_bits_uop_dst_rtype = iregister_read_io_exe_reqs_2_bits_uop_dst_rtype;
  assign ALUExeUnit_io_req_bits_uop_lrs1_rtype = iregister_read_io_exe_reqs_2_bits_uop_lrs1_rtype;
  assign ALUExeUnit_io_req_bits_uop_lrs2_rtype = iregister_read_io_exe_reqs_2_bits_uop_lrs2_rtype;
  assign ALUExeUnit_io_req_bits_uop_frs3_en = iregister_read_io_exe_reqs_2_bits_uop_frs3_en;
  assign ALUExeUnit_io_req_bits_uop_fp_val = iregister_read_io_exe_reqs_2_bits_uop_fp_val;
  assign ALUExeUnit_io_req_bits_uop_fp_single = iregister_read_io_exe_reqs_2_bits_uop_fp_single;
  assign ALUExeUnit_io_req_bits_uop_xcpt_pf_if = iregister_read_io_exe_reqs_2_bits_uop_xcpt_pf_if;
  assign ALUExeUnit_io_req_bits_uop_xcpt_ae_if = iregister_read_io_exe_reqs_2_bits_uop_xcpt_ae_if;
  assign ALUExeUnit_io_req_bits_uop_replay_if = iregister_read_io_exe_reqs_2_bits_uop_replay_if;
  assign ALUExeUnit_io_req_bits_uop_xcpt_ma_if = iregister_read_io_exe_reqs_2_bits_uop_xcpt_ma_if;
  assign ALUExeUnit_io_req_bits_uop_debug_wdata = iregister_read_io_exe_reqs_2_bits_uop_debug_wdata;
  assign ALUExeUnit_io_req_bits_uop_debug_events_fetch_seq = iregister_read_io_exe_reqs_2_bits_uop_debug_events_fetch_seq;
  assign ALUExeUnit_io_req_bits_rs1_data = iregister_read_io_exe_reqs_2_bits_rs1_data;
  assign ALUExeUnit_io_req_bits_rs2_data = iregister_read_io_exe_reqs_2_bits_rs2_data;
  assign ALUExeUnit_io_req_bits_kill = rob_io_flush_valid;
  assign ALUExeUnit_io_brinfo_valid = br_unit_brinfo_valid;
  assign ALUExeUnit_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign ALUExeUnit_io_brinfo_mask = br_unit_brinfo_mask;
  assign ALUExeUnit_clock = clock;
  assign ALUExeUnit_reset = reset;
  assign fp_pipeline_io_brinfo_valid = br_unit_brinfo_valid;
  assign fp_pipeline_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign fp_pipeline_io_brinfo_mask = br_unit_brinfo_mask;
  assign fp_pipeline_io_flush_pipeline = rob_io_flush_valid;
  assign fp_pipeline_io_fcsr_rm = csr_io_fcsr_rm;
  assign fp_pipeline_io_dis_valids_0 = dis_valids_0;
  assign fp_pipeline_io_dis_valids_1 = dis_valids_1;
  assign fp_pipeline_io_dis_uops_0_valid = dis_uops_0_valid;
  assign fp_pipeline_io_dis_uops_0_uopc = dis_uops_0_uopc;
  assign fp_pipeline_io_dis_uops_0_inst = dis_uops_0_inst;
  assign fp_pipeline_io_dis_uops_0_pc = dis_uops_0_pc;
  assign fp_pipeline_io_dis_uops_0_iqtype = dis_uops_0_iqtype;
  assign fp_pipeline_io_dis_uops_0_fu_code = dis_uops_0_fu_code;
  assign fp_pipeline_io_dis_uops_0_allocate_brtag = dis_uops_0_allocate_brtag;
  assign fp_pipeline_io_dis_uops_0_is_br_or_jmp = dis_uops_0_is_br_or_jmp;
  assign fp_pipeline_io_dis_uops_0_is_jump = dis_uops_0_is_jump;
  assign fp_pipeline_io_dis_uops_0_is_jal = dis_uops_0_is_jal;
  assign fp_pipeline_io_dis_uops_0_is_ret = dis_uops_0_is_ret;
  assign fp_pipeline_io_dis_uops_0_is_call = dis_uops_0_is_call;
  assign fp_pipeline_io_dis_uops_0_br_mask = dis_uops_0_br_mask;
  assign fp_pipeline_io_dis_uops_0_br_tag = dis_uops_0_br_tag;
  assign fp_pipeline_io_dis_uops_0_br_prediction_btb_blame = dis_uops_0_br_prediction_btb_blame;
  assign fp_pipeline_io_dis_uops_0_br_prediction_btb_hit = dis_uops_0_br_prediction_btb_hit;
  assign fp_pipeline_io_dis_uops_0_br_prediction_btb_taken = dis_uops_0_br_prediction_btb_taken;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_blame = dis_uops_0_br_prediction_bpd_blame;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_hit = dis_uops_0_br_prediction_bpd_hit;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_taken = dis_uops_0_br_prediction_bpd_taken;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_value = dis_uops_0_br_prediction_bim_resp_value;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_entry_idx = dis_uops_0_br_prediction_bim_resp_entry_idx;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bim_resp_way_idx = dis_uops_0_br_prediction_bim_resp_way_idx;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_takens = dis_uops_0_br_prediction_bpd_resp_takens;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history = dis_uops_0_br_prediction_bpd_resp_history;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_u = dis_uops_0_br_prediction_bpd_resp_history_u;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_history_ptr = dis_uops_0_br_prediction_bpd_resp_history_ptr;
  assign fp_pipeline_io_dis_uops_0_br_prediction_bpd_resp_info = dis_uops_0_br_prediction_bpd_resp_info;
  assign fp_pipeline_io_dis_uops_0_stat_brjmp_mispredicted = dis_uops_0_stat_brjmp_mispredicted;
  assign fp_pipeline_io_dis_uops_0_stat_btb_made_pred = dis_uops_0_stat_btb_made_pred;
  assign fp_pipeline_io_dis_uops_0_stat_btb_mispredicted = dis_uops_0_stat_btb_mispredicted;
  assign fp_pipeline_io_dis_uops_0_stat_bpd_made_pred = dis_uops_0_stat_bpd_made_pred;
  assign fp_pipeline_io_dis_uops_0_stat_bpd_mispredicted = dis_uops_0_stat_bpd_mispredicted;
  assign fp_pipeline_io_dis_uops_0_fetch_pc_lob = dis_uops_0_fetch_pc_lob;
  assign fp_pipeline_io_dis_uops_0_imm_packed = dis_uops_0_imm_packed;
  assign fp_pipeline_io_dis_uops_0_csr_addr = dis_uops_0_csr_addr;
  assign fp_pipeline_io_dis_uops_0_rob_idx = dis_uops_0_rob_idx;
  assign fp_pipeline_io_dis_uops_0_ldq_idx = dis_uops_0_ldq_idx;
  assign fp_pipeline_io_dis_uops_0_stq_idx = dis_uops_0_stq_idx;
  assign fp_pipeline_io_dis_uops_0_brob_idx = dis_uops_0_brob_idx;
  assign fp_pipeline_io_dis_uops_0_pdst = dis_uops_0_pdst;
  assign fp_pipeline_io_dis_uops_0_pop1 = dis_uops_0_pop1;
  assign fp_pipeline_io_dis_uops_0_pop2 = dis_uops_0_pop2;
  assign fp_pipeline_io_dis_uops_0_pop3 = dis_uops_0_pop3;
  assign fp_pipeline_io_dis_uops_0_prs1_busy = dis_uops_0_prs1_busy;
  assign fp_pipeline_io_dis_uops_0_prs2_busy = dis_uops_0_prs2_busy;
  assign fp_pipeline_io_dis_uops_0_prs3_busy = dis_uops_0_prs3_busy;
  assign fp_pipeline_io_dis_uops_0_stale_pdst = dis_uops_0_stale_pdst;
  assign fp_pipeline_io_dis_uops_0_exception = dis_uops_0_exception;
  assign fp_pipeline_io_dis_uops_0_exc_cause = dis_uops_0_exc_cause;
  assign fp_pipeline_io_dis_uops_0_bypassable = dis_uops_0_bypassable;
  assign fp_pipeline_io_dis_uops_0_mem_cmd = dis_uops_0_mem_cmd;
  assign fp_pipeline_io_dis_uops_0_mem_typ = dis_uops_0_mem_typ;
  assign fp_pipeline_io_dis_uops_0_is_fence = dis_uops_0_is_fence;
  assign fp_pipeline_io_dis_uops_0_is_fencei = dis_uops_0_is_fencei;
  assign fp_pipeline_io_dis_uops_0_is_store = dis_uops_0_is_store;
  assign fp_pipeline_io_dis_uops_0_is_amo = dis_uops_0_is_amo;
  assign fp_pipeline_io_dis_uops_0_is_load = dis_uops_0_is_load;
  assign fp_pipeline_io_dis_uops_0_is_sys_pc2epc = dis_uops_0_is_sys_pc2epc;
  assign fp_pipeline_io_dis_uops_0_is_unique = dis_uops_0_is_unique;
  assign fp_pipeline_io_dis_uops_0_flush_on_commit = dis_uops_0_flush_on_commit;
  assign fp_pipeline_io_dis_uops_0_ldst = dis_uops_0_ldst;
  assign fp_pipeline_io_dis_uops_0_lrs1 = dis_uops_0_lrs1;
  assign fp_pipeline_io_dis_uops_0_lrs2 = dis_uops_0_lrs2;
  assign fp_pipeline_io_dis_uops_0_lrs3 = dis_uops_0_lrs3;
  assign fp_pipeline_io_dis_uops_0_ldst_val = dis_uops_0_ldst_val;
  assign fp_pipeline_io_dis_uops_0_dst_rtype = dis_uops_0_dst_rtype;
  assign fp_pipeline_io_dis_uops_0_lrs1_rtype = dis_uops_0_lrs1_rtype;
  assign fp_pipeline_io_dis_uops_0_lrs2_rtype = dis_uops_0_lrs2_rtype;
  assign fp_pipeline_io_dis_uops_0_frs3_en = dis_uops_0_frs3_en;
  assign fp_pipeline_io_dis_uops_0_fp_val = dis_uops_0_fp_val;
  assign fp_pipeline_io_dis_uops_0_fp_single = dis_uops_0_fp_single;
  assign fp_pipeline_io_dis_uops_0_xcpt_pf_if = dis_uops_0_xcpt_pf_if;
  assign fp_pipeline_io_dis_uops_0_xcpt_ae_if = dis_uops_0_xcpt_ae_if;
  assign fp_pipeline_io_dis_uops_0_replay_if = dis_uops_0_replay_if;
  assign fp_pipeline_io_dis_uops_0_xcpt_ma_if = dis_uops_0_xcpt_ma_if;
  assign fp_pipeline_io_dis_uops_0_debug_wdata = dis_uops_0_debug_wdata;
  assign fp_pipeline_io_dis_uops_0_debug_events_fetch_seq = dis_uops_0_debug_events_fetch_seq;
  assign fp_pipeline_io_dis_uops_1_valid = dis_uops_1_valid;
  assign fp_pipeline_io_dis_uops_1_uopc = dis_uops_1_uopc;
  assign fp_pipeline_io_dis_uops_1_inst = dis_uops_1_inst;
  assign fp_pipeline_io_dis_uops_1_pc = dis_uops_1_pc;
  assign fp_pipeline_io_dis_uops_1_iqtype = dis_uops_1_iqtype;
  assign fp_pipeline_io_dis_uops_1_fu_code = dis_uops_1_fu_code;
  assign fp_pipeline_io_dis_uops_1_allocate_brtag = dis_uops_1_allocate_brtag;
  assign fp_pipeline_io_dis_uops_1_is_br_or_jmp = dis_uops_1_is_br_or_jmp;
  assign fp_pipeline_io_dis_uops_1_is_jump = dis_uops_1_is_jump;
  assign fp_pipeline_io_dis_uops_1_is_jal = dis_uops_1_is_jal;
  assign fp_pipeline_io_dis_uops_1_is_ret = dis_uops_1_is_ret;
  assign fp_pipeline_io_dis_uops_1_is_call = dis_uops_1_is_call;
  assign fp_pipeline_io_dis_uops_1_br_mask = dis_uops_1_br_mask;
  assign fp_pipeline_io_dis_uops_1_br_tag = dis_uops_1_br_tag;
  assign fp_pipeline_io_dis_uops_1_br_prediction_btb_blame = dis_uops_1_br_prediction_btb_blame;
  assign fp_pipeline_io_dis_uops_1_br_prediction_btb_hit = dis_uops_1_br_prediction_btb_hit;
  assign fp_pipeline_io_dis_uops_1_br_prediction_btb_taken = dis_uops_1_br_prediction_btb_taken;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_blame = dis_uops_1_br_prediction_bpd_blame;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_hit = dis_uops_1_br_prediction_bpd_hit;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_taken = dis_uops_1_br_prediction_bpd_taken;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_value = dis_uops_1_br_prediction_bim_resp_value;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_entry_idx = dis_uops_1_br_prediction_bim_resp_entry_idx;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bim_resp_way_idx = dis_uops_1_br_prediction_bim_resp_way_idx;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_takens = dis_uops_1_br_prediction_bpd_resp_takens;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history = dis_uops_1_br_prediction_bpd_resp_history;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_u = dis_uops_1_br_prediction_bpd_resp_history_u;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_history_ptr = dis_uops_1_br_prediction_bpd_resp_history_ptr;
  assign fp_pipeline_io_dis_uops_1_br_prediction_bpd_resp_info = dis_uops_1_br_prediction_bpd_resp_info;
  assign fp_pipeline_io_dis_uops_1_stat_brjmp_mispredicted = dis_uops_1_stat_brjmp_mispredicted;
  assign fp_pipeline_io_dis_uops_1_stat_btb_made_pred = dis_uops_1_stat_btb_made_pred;
  assign fp_pipeline_io_dis_uops_1_stat_btb_mispredicted = dis_uops_1_stat_btb_mispredicted;
  assign fp_pipeline_io_dis_uops_1_stat_bpd_made_pred = dis_uops_1_stat_bpd_made_pred;
  assign fp_pipeline_io_dis_uops_1_stat_bpd_mispredicted = dis_uops_1_stat_bpd_mispredicted;
  assign fp_pipeline_io_dis_uops_1_fetch_pc_lob = dis_uops_1_fetch_pc_lob;
  assign fp_pipeline_io_dis_uops_1_imm_packed = dis_uops_1_imm_packed;
  assign fp_pipeline_io_dis_uops_1_csr_addr = dis_uops_1_csr_addr;
  assign fp_pipeline_io_dis_uops_1_rob_idx = dis_uops_1_rob_idx;
  assign fp_pipeline_io_dis_uops_1_ldq_idx = dis_uops_1_ldq_idx;
  assign fp_pipeline_io_dis_uops_1_stq_idx = dis_uops_1_stq_idx;
  assign fp_pipeline_io_dis_uops_1_brob_idx = dis_uops_1_brob_idx;
  assign fp_pipeline_io_dis_uops_1_pdst = dis_uops_1_pdst;
  assign fp_pipeline_io_dis_uops_1_pop1 = dis_uops_1_pop1;
  assign fp_pipeline_io_dis_uops_1_pop2 = dis_uops_1_pop2;
  assign fp_pipeline_io_dis_uops_1_pop3 = dis_uops_1_pop3;
  assign fp_pipeline_io_dis_uops_1_prs1_busy = dis_uops_1_prs1_busy;
  assign fp_pipeline_io_dis_uops_1_prs2_busy = dis_uops_1_prs2_busy;
  assign fp_pipeline_io_dis_uops_1_prs3_busy = dis_uops_1_prs3_busy;
  assign fp_pipeline_io_dis_uops_1_stale_pdst = dis_uops_1_stale_pdst;
  assign fp_pipeline_io_dis_uops_1_exception = dis_uops_1_exception;
  assign fp_pipeline_io_dis_uops_1_exc_cause = dis_uops_1_exc_cause;
  assign fp_pipeline_io_dis_uops_1_bypassable = dis_uops_1_bypassable;
  assign fp_pipeline_io_dis_uops_1_mem_cmd = dis_uops_1_mem_cmd;
  assign fp_pipeline_io_dis_uops_1_mem_typ = dis_uops_1_mem_typ;
  assign fp_pipeline_io_dis_uops_1_is_fence = dis_uops_1_is_fence;
  assign fp_pipeline_io_dis_uops_1_is_fencei = dis_uops_1_is_fencei;
  assign fp_pipeline_io_dis_uops_1_is_store = dis_uops_1_is_store;
  assign fp_pipeline_io_dis_uops_1_is_amo = dis_uops_1_is_amo;
  assign fp_pipeline_io_dis_uops_1_is_load = dis_uops_1_is_load;
  assign fp_pipeline_io_dis_uops_1_is_sys_pc2epc = dis_uops_1_is_sys_pc2epc;
  assign fp_pipeline_io_dis_uops_1_is_unique = dis_uops_1_is_unique;
  assign fp_pipeline_io_dis_uops_1_flush_on_commit = dis_uops_1_flush_on_commit;
  assign fp_pipeline_io_dis_uops_1_ldst = dis_uops_1_ldst;
  assign fp_pipeline_io_dis_uops_1_lrs1 = dis_uops_1_lrs1;
  assign fp_pipeline_io_dis_uops_1_lrs2 = dis_uops_1_lrs2;
  assign fp_pipeline_io_dis_uops_1_lrs3 = dis_uops_1_lrs3;
  assign fp_pipeline_io_dis_uops_1_ldst_val = dis_uops_1_ldst_val;
  assign fp_pipeline_io_dis_uops_1_dst_rtype = dis_uops_1_dst_rtype;
  assign fp_pipeline_io_dis_uops_1_lrs1_rtype = dis_uops_1_lrs1_rtype;
  assign fp_pipeline_io_dis_uops_1_lrs2_rtype = dis_uops_1_lrs2_rtype;
  assign fp_pipeline_io_dis_uops_1_frs3_en = dis_uops_1_frs3_en;
  assign fp_pipeline_io_dis_uops_1_fp_val = dis_uops_1_fp_val;
  assign fp_pipeline_io_dis_uops_1_fp_single = dis_uops_1_fp_single;
  assign fp_pipeline_io_dis_uops_1_xcpt_pf_if = dis_uops_1_xcpt_pf_if;
  assign fp_pipeline_io_dis_uops_1_xcpt_ae_if = dis_uops_1_xcpt_ae_if;
  assign fp_pipeline_io_dis_uops_1_replay_if = dis_uops_1_replay_if;
  assign fp_pipeline_io_dis_uops_1_xcpt_ma_if = dis_uops_1_xcpt_ma_if;
  assign fp_pipeline_io_dis_uops_1_debug_wdata = dis_uops_1_debug_wdata;
  assign fp_pipeline_io_dis_uops_1_debug_events_fetch_seq = dis_uops_1_debug_events_fetch_seq;
  assign fp_pipeline_io_ll_wport_valid = _T_3078;
  assign fp_pipeline_io_ll_wport_bits_uop_rob_idx = mem_unit_io_resp_0_bits_uop_rob_idx;
  assign fp_pipeline_io_ll_wport_bits_uop_pdst = mem_unit_io_resp_0_bits_uop_pdst;
  assign fp_pipeline_io_ll_wport_bits_uop_mem_typ = mem_unit_io_resp_0_bits_uop_mem_typ;
  assign fp_pipeline_io_ll_wport_bits_uop_dst_rtype = mem_unit_io_resp_0_bits_uop_dst_rtype;
  assign fp_pipeline_io_ll_wport_bits_uop_fp_val = mem_unit_io_resp_0_bits_uop_fp_val;
  assign fp_pipeline_io_ll_wport_bits_data = mem_unit_io_resp_0_bits_data;
  assign fp_pipeline_io_fromint_valid = _T_3041;
  assign fp_pipeline_io_fromint_bits_uop_uopc = iregister_read_io_exe_reqs_2_bits_uop_uopc;
  assign fp_pipeline_io_fromint_bits_uop_ctrl_rf_wen = iregister_read_io_exe_reqs_2_bits_uop_ctrl_rf_wen;
  assign fp_pipeline_io_fromint_bits_uop_br_mask = iregister_read_io_exe_reqs_2_bits_uop_br_mask;
  assign fp_pipeline_io_fromint_bits_uop_imm_packed = iregister_read_io_exe_reqs_2_bits_uop_imm_packed;
  assign fp_pipeline_io_fromint_bits_uop_rob_idx = iregister_read_io_exe_reqs_2_bits_uop_rob_idx;
  assign fp_pipeline_io_fromint_bits_uop_pdst = iregister_read_io_exe_reqs_2_bits_uop_pdst;
  assign fp_pipeline_io_fromint_bits_uop_dst_rtype = iregister_read_io_exe_reqs_2_bits_uop_dst_rtype;
  assign fp_pipeline_io_fromint_bits_uop_fp_val = iregister_read_io_exe_reqs_2_bits_uop_fp_val;
  assign fp_pipeline_io_fromint_bits_rs1_data = {{1'd0}, iregister_read_io_exe_reqs_2_bits_rs1_data};
  assign fp_pipeline_io_toint_ready = ll_wbarb_io_in_1_ready;
  assign fp_pipeline_clock = clock;
  assign fp_pipeline_reset = reset;
  assign fetch_unit_io_imem_resp_valid = io_imem_resp_valid;
  assign fetch_unit_io_imem_resp_bits_pc = io_imem_resp_bits_pc;
  assign fetch_unit_io_imem_resp_bits_data = io_imem_resp_bits_data;
  assign fetch_unit_io_imem_resp_bits_mask = io_imem_resp_bits_mask;
  assign fetch_unit_io_imem_resp_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst;
  assign fetch_unit_io_imem_resp_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
  assign fetch_unit_io_imem_resp_bits_replay = io_imem_resp_bits_replay;
  assign fetch_unit_io_f2_btb_resp_bits_bim_resp_value = bpd_stage_io_f2_btb_resp_bits_bim_resp_value;
  assign fetch_unit_io_f2_btb_resp_bits_bim_resp_entry_idx = bpd_stage_io_f2_btb_resp_bits_bim_resp_entry_idx;
  assign fetch_unit_io_f2_btb_resp_bits_bim_resp_way_idx = bpd_stage_io_f2_btb_resp_bits_bim_resp_way_idx;
  assign fetch_unit_io_f2_bpd_resp_bits_takens = bpd_stage_io_f2_bpd_resp_bits_takens;
  assign fetch_unit_io_f2_bpd_resp_bits_info = bpd_stage_io_f2_bpd_resp_bits_info;
  assign fetch_unit_io_f3_bpd_resp_bits_history = bpd_stage_io_f3_bpd_resp_bits_history;
  assign fetch_unit_io_f3_bpd_resp_bits_history_ptr = bpd_stage_io_f3_bpd_resp_bits_history_ptr;
  assign fetch_unit_io_br_unit_take_pc = br_unit_take_pc;
  assign fetch_unit_io_br_unit_target = br_unit_target;
  assign fetch_unit_io_clear_fetchbuffer = _T_2702;
  assign fetch_unit_io_flush_take_pc = _T_2705;
  assign fetch_unit_io_flush_pc = rob_io_flush_bits_pc[39:0];
  assign fetch_unit_io_sfence_take_pc = lsu_io_exe_resp_bits_sfence_valid;
  assign fetch_unit_io_sfence_addr = {{1'd0}, lsu_io_exe_resp_bits_sfence_bits_addr};
  assign fetch_unit_io_resp_ready = dec_serializer_io_enq_ready;
  assign fetch_unit_clock = clock;
  assign fetch_unit_reset = reset;
  assign bpd_stage_io_fetch_stalled = fetch_unit_io_stalled;
  assign bpd_stage_io_f3_btb_update_valid = fetch_unit_io_f3_btb_update_valid;
  assign bpd_stage_io_f3_btb_update_bits_pc = fetch_unit_io_f3_btb_update_bits_pc;
  assign bpd_stage_io_f3_btb_update_bits_target = fetch_unit_io_f3_btb_update_bits_target;
  assign bpd_stage_io_f3_btb_update_bits_cfi_pc = fetch_unit_io_f3_btb_update_bits_cfi_pc;
  assign bpd_stage_io_f3_btb_update_bits_bpd_type = fetch_unit_io_f3_btb_update_bits_bpd_type;
  assign bpd_stage_io_f3_btb_update_bits_cfi_type = fetch_unit_io_f3_btb_update_bits_cfi_type;
  assign bpd_stage_io_f3_hist_update_valid = fetch_unit_io_f3_hist_update_valid;
  assign bpd_stage_io_f3_hist_update_bits_taken = fetch_unit_io_f3_hist_update_bits_taken;
  assign bpd_stage_io_f3_bim_update_valid = fetch_unit_io_f3_bim_update_valid;
  assign bpd_stage_io_f3_bim_update_bits_taken = fetch_unit_io_f3_bim_update_bits_taken;
  assign bpd_stage_io_f3_bim_update_bits_bim_resp_value = fetch_unit_io_f3_bim_update_bits_bim_resp_value;
  assign bpd_stage_io_f3_bim_update_bits_bim_resp_entry_idx = fetch_unit_io_f3_bim_update_bits_bim_resp_entry_idx;
  assign bpd_stage_io_f3_bim_update_bits_bim_resp_way_idx = fetch_unit_io_f3_bim_update_bits_bim_resp_way_idx;
  assign bpd_stage_io_br_unit_btb_update_valid = br_unit_btb_update_valid;
  assign bpd_stage_io_br_unit_btb_update_bits_pc = br_unit_btb_update_bits_pc;
  assign bpd_stage_io_br_unit_btb_update_bits_target = br_unit_btb_update_bits_target;
  assign bpd_stage_io_br_unit_btb_update_bits_cfi_pc = br_unit_btb_update_bits_cfi_pc;
  assign bpd_stage_io_br_unit_btb_update_bits_bpd_type = br_unit_btb_update_bits_bpd_type;
  assign bpd_stage_io_br_unit_btb_update_bits_cfi_type = br_unit_btb_update_bits_cfi_type;
  assign bpd_stage_io_br_unit_bim_update_valid = br_unit_bim_update_valid;
  assign bpd_stage_io_br_unit_bim_update_bits_taken = br_unit_bim_update_bits_taken;
  assign bpd_stage_io_br_unit_bim_update_bits_bim_resp_value = br_unit_bim_update_bits_bim_resp_value;
  assign bpd_stage_io_br_unit_bim_update_bits_bim_resp_entry_idx = br_unit_bim_update_bits_bim_resp_entry_idx;
  assign bpd_stage_io_br_unit_bim_update_bits_bim_resp_way_idx = br_unit_bim_update_bits_bim_resp_way_idx;
  assign bpd_stage_io_br_unit_bpd_update_valid = br_unit_bpd_update_valid;
  assign bpd_stage_io_br_unit_bpd_update_bits_mispredict = br_unit_bpd_update_bits_mispredict;
  assign bpd_stage_io_br_unit_bpd_update_bits_history = br_unit_bpd_update_bits_history;
  assign bpd_stage_io_br_unit_bpd_update_bits_history_ptr = br_unit_bpd_update_bits_history_ptr;
  assign bpd_stage_io_br_unit_bpd_update_bits_bpd_mispredict = br_unit_bpd_update_bits_bpd_mispredict;
  assign bpd_stage_io_br_unit_bpd_update_bits_taken = br_unit_bpd_update_bits_taken;
  assign bpd_stage_io_br_unit_bpd_update_bits_new_pc_same_packet = br_unit_bpd_update_bits_new_pc_same_packet;
  assign bpd_stage_io_brob_allocate_valid = _T_2874;
  assign bpd_stage_io_brob_allocate_bits_ctrl_brob_idx = dec_uops_0_brob_idx;
  assign bpd_stage_io_brob_allocate_bits_info_info = dec_serializer_io_deq_bits_bpd_resp_info;
  assign bpd_stage_io_brob_deallocate_valid = rob_io_brob_deallocate_valid;
  assign bpd_stage_io_brob_deallocate_bits_brob_idx = rob_io_brob_deallocate_bits_brob_idx;
  assign bpd_stage_io_brob_bpd_update_valid = br_unit_bpd_update_valid;
  assign bpd_stage_io_brob_bpd_update_bits_br_pc = br_unit_bpd_update_bits_br_pc;
  assign bpd_stage_io_brob_bpd_update_bits_brob_idx = br_unit_bpd_update_bits_brob_idx;
  assign bpd_stage_io_brob_bpd_update_bits_mispredict = br_unit_bpd_update_bits_mispredict;
  assign bpd_stage_io_brob_bpd_update_bits_bpd_predict_val = br_unit_bpd_update_bits_bpd_predict_val;
  assign bpd_stage_io_brob_bpd_update_bits_bpd_mispredict = br_unit_bpd_update_bits_bpd_mispredict;
  assign bpd_stage_io_brob_bpd_update_bits_taken = br_unit_bpd_update_bits_taken;
  assign bpd_stage_io_brob_bpd_update_bits_is_br = br_unit_bpd_update_bits_is_br;
  assign bpd_stage_io_brob_flush = _T_3521;
  assign bpd_stage_io_flush = rob_io_flush_valid;
  assign bpd_stage_io_redirect = io_imem_req_valid;
  assign bpd_stage_io_status_debug = csr_io_status_debug;
  assign bpd_stage_clock = clock;
  assign bpd_stage_reset = reset;
  assign dec_serializer_io_enq_valid = fetch_unit_io_resp_valid;
  assign dec_serializer_io_enq_bits_pc = fetch_unit_io_resp_bits_pc;
  assign dec_serializer_io_enq_bits_insts_0 = fetch_unit_io_resp_bits_insts_0;
  assign dec_serializer_io_enq_bits_insts_1 = fetch_unit_io_resp_bits_insts_1;
  assign dec_serializer_io_enq_bits_mask = fetch_unit_io_resp_bits_mask;
  assign dec_serializer_io_enq_bits_xcpt_pf_if = fetch_unit_io_resp_bits_xcpt_pf_if;
  assign dec_serializer_io_enq_bits_xcpt_ae_if = fetch_unit_io_resp_bits_xcpt_ae_if;
  assign dec_serializer_io_enq_bits_replay_if = fetch_unit_io_resp_bits_replay_if;
  assign dec_serializer_io_enq_bits_xcpt_ma_if_oh = fetch_unit_io_resp_bits_xcpt_ma_if_oh;
  assign dec_serializer_io_enq_bits_bpu_info_0_btb_blame = fetch_unit_io_resp_bits_bpu_info_0_btb_blame;
  assign dec_serializer_io_enq_bits_bpu_info_0_btb_hit = fetch_unit_io_resp_bits_bpu_info_0_btb_hit;
  assign dec_serializer_io_enq_bits_bpu_info_0_btb_taken = fetch_unit_io_resp_bits_bpu_info_0_btb_taken;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_blame = fetch_unit_io_resp_bits_bpu_info_0_bpd_blame;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_hit = fetch_unit_io_resp_bits_bpu_info_0_bpd_hit;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_taken = fetch_unit_io_resp_bits_bpu_info_0_bpd_taken;
  assign dec_serializer_io_enq_bits_bpu_info_0_bim_resp_value = fetch_unit_io_resp_bits_bpu_info_0_bim_resp_value;
  assign dec_serializer_io_enq_bits_bpu_info_0_bim_resp_entry_idx = fetch_unit_io_resp_bits_bpu_info_0_bim_resp_entry_idx;
  assign dec_serializer_io_enq_bits_bpu_info_0_bim_resp_way_idx = fetch_unit_io_resp_bits_bpu_info_0_bim_resp_way_idx;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_takens = fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_takens;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history = fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_u = fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_u;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_history_ptr = fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_history_ptr;
  assign dec_serializer_io_enq_bits_bpu_info_0_bpd_resp_info = fetch_unit_io_resp_bits_bpu_info_0_bpd_resp_info;
  assign dec_serializer_io_enq_bits_bpu_info_1_btb_blame = fetch_unit_io_resp_bits_bpu_info_1_btb_blame;
  assign dec_serializer_io_enq_bits_bpu_info_1_btb_hit = fetch_unit_io_resp_bits_bpu_info_1_btb_hit;
  assign dec_serializer_io_enq_bits_bpu_info_1_btb_taken = fetch_unit_io_resp_bits_bpu_info_1_btb_taken;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_blame = fetch_unit_io_resp_bits_bpu_info_1_bpd_blame;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_hit = fetch_unit_io_resp_bits_bpu_info_1_bpd_hit;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_taken = fetch_unit_io_resp_bits_bpu_info_1_bpd_taken;
  assign dec_serializer_io_enq_bits_bpu_info_1_bim_resp_value = fetch_unit_io_resp_bits_bpu_info_1_bim_resp_value;
  assign dec_serializer_io_enq_bits_bpu_info_1_bim_resp_entry_idx = fetch_unit_io_resp_bits_bpu_info_1_bim_resp_entry_idx;
  assign dec_serializer_io_enq_bits_bpu_info_1_bim_resp_way_idx = fetch_unit_io_resp_bits_bpu_info_1_bim_resp_way_idx;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_takens = fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_takens;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history = fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_u = fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_u;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_history_ptr = fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_history_ptr;
  assign dec_serializer_io_enq_bits_bpu_info_1_bpd_resp_info = fetch_unit_io_resp_bits_bpu_info_1_bpd_resp_info;
  assign dec_serializer_io_enq_bits_debug_events_0_fetch_seq = fetch_unit_io_resp_bits_debug_events_0_fetch_seq;
  assign dec_serializer_io_enq_bits_debug_events_1_fetch_seq = fetch_unit_io_resp_bits_debug_events_1_fetch_seq;
  assign dec_serializer_io_deq_ready = dec_rdy;
  assign decode_units_0_io_enq_uop_valid = dec_serializer_io_deq_bits_uops_0_valid;
  assign decode_units_0_io_enq_uop_inst = dec_serializer_io_deq_bits_uops_0_inst;
  assign decode_units_0_io_enq_uop_pc = dec_serializer_io_deq_bits_uops_0_pc;
  assign decode_units_0_io_enq_uop_br_prediction_btb_blame = dec_serializer_io_deq_bits_uops_0_br_prediction_btb_blame;
  assign decode_units_0_io_enq_uop_br_prediction_btb_hit = dec_serializer_io_deq_bits_uops_0_br_prediction_btb_hit;
  assign decode_units_0_io_enq_uop_br_prediction_btb_taken = dec_serializer_io_deq_bits_uops_0_br_prediction_btb_taken;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_blame = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_blame;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_hit = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_hit;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_taken = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_taken;
  assign decode_units_0_io_enq_uop_br_prediction_bim_resp_value = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_value;
  assign decode_units_0_io_enq_uop_br_prediction_bim_resp_entry_idx = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_entry_idx;
  assign decode_units_0_io_enq_uop_br_prediction_bim_resp_way_idx = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_way_idx;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_resp_takens = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_takens;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_resp_history = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_u = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_u;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_resp_history_ptr = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_ptr;
  assign decode_units_0_io_enq_uop_br_prediction_bpd_resp_info = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_info;
  assign decode_units_0_io_enq_uop_fetch_pc_lob = dec_serializer_io_deq_bits_uops_0_fetch_pc_lob;
  assign decode_units_0_io_enq_uop_xcpt_pf_if = dec_serializer_io_deq_bits_uops_0_xcpt_pf_if;
  assign decode_units_0_io_enq_uop_xcpt_ae_if = dec_serializer_io_deq_bits_uops_0_xcpt_ae_if;
  assign decode_units_0_io_enq_uop_replay_if = dec_serializer_io_deq_bits_uops_0_replay_if;
  assign decode_units_0_io_enq_uop_xcpt_ma_if = dec_serializer_io_deq_bits_uops_0_xcpt_ma_if;
  assign decode_units_0_io_enq_uop_debug_events_fetch_seq = dec_serializer_io_deq_bits_uops_0_debug_events_fetch_seq;
  assign decode_units_0_io_status_isa = csr_io_status_isa;
  assign decode_units_0_io_csr_decode_fp_illegal = csr_io_decode_0_fp_illegal;
  assign decode_units_0_io_csr_decode_read_illegal = csr_io_decode_0_read_illegal;
  assign decode_units_0_io_csr_decode_write_illegal = csr_io_decode_0_write_illegal;
  assign decode_units_0_io_csr_decode_write_flush = csr_io_decode_0_write_flush;
  assign decode_units_0_io_csr_decode_system_illegal = csr_io_decode_0_system_illegal;
  assign decode_units_0_io_interrupt = csr_io_interrupt;
  assign decode_units_0_io_interrupt_cause = csr_io_interrupt_cause;
  assign decode_units_1_io_enq_uop_valid = dec_serializer_io_deq_bits_uops_1_valid;
  assign decode_units_1_io_enq_uop_inst = dec_serializer_io_deq_bits_uops_1_inst;
  assign decode_units_1_io_enq_uop_pc = dec_serializer_io_deq_bits_uops_1_pc;
  assign decode_units_1_io_enq_uop_br_prediction_btb_blame = dec_serializer_io_deq_bits_uops_1_br_prediction_btb_blame;
  assign decode_units_1_io_enq_uop_br_prediction_btb_hit = dec_serializer_io_deq_bits_uops_1_br_prediction_btb_hit;
  assign decode_units_1_io_enq_uop_br_prediction_btb_taken = dec_serializer_io_deq_bits_uops_1_br_prediction_btb_taken;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_blame = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_blame;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_hit = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_hit;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_taken = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_taken;
  assign decode_units_1_io_enq_uop_br_prediction_bim_resp_value = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_value;
  assign decode_units_1_io_enq_uop_br_prediction_bim_resp_entry_idx = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_entry_idx;
  assign decode_units_1_io_enq_uop_br_prediction_bim_resp_way_idx = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_way_idx;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_resp_takens = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_takens;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_resp_history = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_u = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_u;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_resp_history_ptr = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_ptr;
  assign decode_units_1_io_enq_uop_br_prediction_bpd_resp_info = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_info;
  assign decode_units_1_io_enq_uop_fetch_pc_lob = dec_serializer_io_deq_bits_uops_1_fetch_pc_lob;
  assign decode_units_1_io_enq_uop_xcpt_pf_if = dec_serializer_io_deq_bits_uops_1_xcpt_pf_if;
  assign decode_units_1_io_enq_uop_xcpt_ae_if = dec_serializer_io_deq_bits_uops_1_xcpt_ae_if;
  assign decode_units_1_io_enq_uop_replay_if = dec_serializer_io_deq_bits_uops_1_replay_if;
  assign decode_units_1_io_enq_uop_xcpt_ma_if = dec_serializer_io_deq_bits_uops_1_xcpt_ma_if;
  assign decode_units_1_io_enq_uop_debug_events_fetch_seq = dec_serializer_io_deq_bits_uops_1_debug_events_fetch_seq;
  assign decode_units_1_io_status_isa = csr_io_status_isa;
  assign decode_units_1_io_csr_decode_fp_illegal = csr_io_decode_1_fp_illegal;
  assign decode_units_1_io_csr_decode_read_illegal = csr_io_decode_1_read_illegal;
  assign decode_units_1_io_csr_decode_write_illegal = csr_io_decode_1_write_illegal;
  assign decode_units_1_io_csr_decode_write_flush = csr_io_decode_1_write_flush;
  assign decode_units_1_io_csr_decode_system_illegal = csr_io_decode_1_system_illegal;
  assign decode_units_1_io_interrupt = csr_io_interrupt;
  assign decode_units_1_io_interrupt_cause = csr_io_interrupt_cause;
  assign dec_brmask_logic_io_is_branch_0 = _T_2827;
  assign dec_brmask_logic_io_is_branch_1 = _T_2832;
  assign dec_brmask_logic_io_will_fire_0 = _T_2828;
  assign dec_brmask_logic_io_will_fire_1 = _T_2833;
  assign dec_brmask_logic_io_brinfo_valid = br_unit_brinfo_valid;
  assign dec_brmask_logic_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign dec_brmask_logic_io_brinfo_mask = br_unit_brinfo_mask;
  assign dec_brmask_logic_io_brinfo_exe_mask = br_unit_brinfo_exe_mask;
  assign dec_brmask_logic_io_flush_pipeline = rob_io_flush_valid;
  assign dec_brmask_logic_clock = clock;
  assign dec_brmask_logic_reset = reset;
  assign rename_stage_io_kill = fetch_unit_io_clear_fetchbuffer;
  assign rename_stage_io_dec_will_fire_0 = dec_will_fire_0;
  assign rename_stage_io_dec_will_fire_1 = dec_will_fire_1;
  assign rename_stage_io_dec_uops_0_valid = dec_uops_0_valid;
  assign rename_stage_io_dec_uops_0_uopc = dec_uops_0_uopc;
  assign rename_stage_io_dec_uops_0_inst = dec_uops_0_inst;
  assign rename_stage_io_dec_uops_0_pc = dec_uops_0_pc;
  assign rename_stage_io_dec_uops_0_iqtype = dec_uops_0_iqtype;
  assign rename_stage_io_dec_uops_0_fu_code = dec_uops_0_fu_code;
  assign rename_stage_io_dec_uops_0_allocate_brtag = dec_uops_0_allocate_brtag;
  assign rename_stage_io_dec_uops_0_is_br_or_jmp = dec_uops_0_is_br_or_jmp;
  assign rename_stage_io_dec_uops_0_is_jump = dec_uops_0_is_jump;
  assign rename_stage_io_dec_uops_0_is_jal = dec_uops_0_is_jal;
  assign rename_stage_io_dec_uops_0_is_ret = dec_uops_0_is_ret;
  assign rename_stage_io_dec_uops_0_is_call = dec_uops_0_is_call;
  assign rename_stage_io_dec_uops_0_br_mask = dec_uops_0_br_mask;
  assign rename_stage_io_dec_uops_0_br_tag = dec_uops_0_br_tag;
  assign rename_stage_io_dec_uops_0_br_prediction_btb_blame = dec_uops_0_br_prediction_btb_blame;
  assign rename_stage_io_dec_uops_0_br_prediction_btb_hit = dec_uops_0_br_prediction_btb_hit;
  assign rename_stage_io_dec_uops_0_br_prediction_btb_taken = dec_uops_0_br_prediction_btb_taken;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_blame = dec_uops_0_br_prediction_bpd_blame;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_hit = dec_uops_0_br_prediction_bpd_hit;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_taken = dec_uops_0_br_prediction_bpd_taken;
  assign rename_stage_io_dec_uops_0_br_prediction_bim_resp_value = dec_uops_0_br_prediction_bim_resp_value;
  assign rename_stage_io_dec_uops_0_br_prediction_bim_resp_entry_idx = dec_uops_0_br_prediction_bim_resp_entry_idx;
  assign rename_stage_io_dec_uops_0_br_prediction_bim_resp_way_idx = dec_uops_0_br_prediction_bim_resp_way_idx;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_resp_takens = dec_uops_0_br_prediction_bpd_resp_takens;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history = dec_uops_0_br_prediction_bpd_resp_history;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_u = dec_uops_0_br_prediction_bpd_resp_history_u;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_resp_history_ptr = dec_uops_0_br_prediction_bpd_resp_history_ptr;
  assign rename_stage_io_dec_uops_0_br_prediction_bpd_resp_info = dec_uops_0_br_prediction_bpd_resp_info;
  assign rename_stage_io_dec_uops_0_fetch_pc_lob = dec_uops_0_fetch_pc_lob;
  assign rename_stage_io_dec_uops_0_imm_packed = dec_uops_0_imm_packed;
  assign rename_stage_io_dec_uops_0_rob_idx = dec_uops_0_rob_idx;
  assign rename_stage_io_dec_uops_0_ldq_idx = dec_uops_0_ldq_idx;
  assign rename_stage_io_dec_uops_0_stq_idx = dec_uops_0_stq_idx;
  assign rename_stage_io_dec_uops_0_brob_idx = dec_uops_0_brob_idx;
  assign rename_stage_io_dec_uops_0_exception = dec_uops_0_exception;
  assign rename_stage_io_dec_uops_0_exc_cause = dec_uops_0_exc_cause;
  assign rename_stage_io_dec_uops_0_bypassable = dec_uops_0_bypassable;
  assign rename_stage_io_dec_uops_0_mem_cmd = dec_uops_0_mem_cmd;
  assign rename_stage_io_dec_uops_0_mem_typ = dec_uops_0_mem_typ;
  assign rename_stage_io_dec_uops_0_is_fence = dec_uops_0_is_fence;
  assign rename_stage_io_dec_uops_0_is_fencei = dec_uops_0_is_fencei;
  assign rename_stage_io_dec_uops_0_is_store = dec_uops_0_is_store;
  assign rename_stage_io_dec_uops_0_is_amo = dec_uops_0_is_amo;
  assign rename_stage_io_dec_uops_0_is_load = dec_uops_0_is_load;
  assign rename_stage_io_dec_uops_0_is_sys_pc2epc = dec_uops_0_is_sys_pc2epc;
  assign rename_stage_io_dec_uops_0_is_unique = dec_uops_0_is_unique;
  assign rename_stage_io_dec_uops_0_flush_on_commit = dec_uops_0_flush_on_commit;
  assign rename_stage_io_dec_uops_0_ldst = dec_uops_0_ldst;
  assign rename_stage_io_dec_uops_0_lrs1 = dec_uops_0_lrs1;
  assign rename_stage_io_dec_uops_0_lrs2 = dec_uops_0_lrs2;
  assign rename_stage_io_dec_uops_0_lrs3 = dec_uops_0_lrs3;
  assign rename_stage_io_dec_uops_0_ldst_val = dec_uops_0_ldst_val;
  assign rename_stage_io_dec_uops_0_dst_rtype = dec_uops_0_dst_rtype;
  assign rename_stage_io_dec_uops_0_lrs1_rtype = dec_uops_0_lrs1_rtype;
  assign rename_stage_io_dec_uops_0_lrs2_rtype = dec_uops_0_lrs2_rtype;
  assign rename_stage_io_dec_uops_0_frs3_en = dec_uops_0_frs3_en;
  assign rename_stage_io_dec_uops_0_fp_val = dec_uops_0_fp_val;
  assign rename_stage_io_dec_uops_0_fp_single = dec_uops_0_fp_single;
  assign rename_stage_io_dec_uops_0_xcpt_pf_if = dec_uops_0_xcpt_pf_if;
  assign rename_stage_io_dec_uops_0_xcpt_ae_if = dec_uops_0_xcpt_ae_if;
  assign rename_stage_io_dec_uops_0_replay_if = dec_uops_0_replay_if;
  assign rename_stage_io_dec_uops_0_xcpt_ma_if = dec_uops_0_xcpt_ma_if;
  assign rename_stage_io_dec_uops_0_debug_events_fetch_seq = dec_uops_0_debug_events_fetch_seq;
  assign rename_stage_io_dec_uops_1_valid = dec_uops_1_valid;
  assign rename_stage_io_dec_uops_1_uopc = dec_uops_1_uopc;
  assign rename_stage_io_dec_uops_1_inst = dec_uops_1_inst;
  assign rename_stage_io_dec_uops_1_pc = dec_uops_1_pc;
  assign rename_stage_io_dec_uops_1_iqtype = dec_uops_1_iqtype;
  assign rename_stage_io_dec_uops_1_fu_code = dec_uops_1_fu_code;
  assign rename_stage_io_dec_uops_1_allocate_brtag = dec_uops_1_allocate_brtag;
  assign rename_stage_io_dec_uops_1_is_br_or_jmp = dec_uops_1_is_br_or_jmp;
  assign rename_stage_io_dec_uops_1_is_jump = dec_uops_1_is_jump;
  assign rename_stage_io_dec_uops_1_is_jal = dec_uops_1_is_jal;
  assign rename_stage_io_dec_uops_1_is_ret = dec_uops_1_is_ret;
  assign rename_stage_io_dec_uops_1_is_call = dec_uops_1_is_call;
  assign rename_stage_io_dec_uops_1_br_mask = dec_uops_1_br_mask;
  assign rename_stage_io_dec_uops_1_br_tag = dec_uops_1_br_tag;
  assign rename_stage_io_dec_uops_1_br_prediction_btb_blame = dec_uops_1_br_prediction_btb_blame;
  assign rename_stage_io_dec_uops_1_br_prediction_btb_hit = dec_uops_1_br_prediction_btb_hit;
  assign rename_stage_io_dec_uops_1_br_prediction_btb_taken = dec_uops_1_br_prediction_btb_taken;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_blame = dec_uops_1_br_prediction_bpd_blame;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_hit = dec_uops_1_br_prediction_bpd_hit;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_taken = dec_uops_1_br_prediction_bpd_taken;
  assign rename_stage_io_dec_uops_1_br_prediction_bim_resp_value = dec_uops_1_br_prediction_bim_resp_value;
  assign rename_stage_io_dec_uops_1_br_prediction_bim_resp_entry_idx = dec_uops_1_br_prediction_bim_resp_entry_idx;
  assign rename_stage_io_dec_uops_1_br_prediction_bim_resp_way_idx = dec_uops_1_br_prediction_bim_resp_way_idx;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_resp_takens = dec_uops_1_br_prediction_bpd_resp_takens;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history = dec_uops_1_br_prediction_bpd_resp_history;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_u = dec_uops_1_br_prediction_bpd_resp_history_u;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_resp_history_ptr = dec_uops_1_br_prediction_bpd_resp_history_ptr;
  assign rename_stage_io_dec_uops_1_br_prediction_bpd_resp_info = dec_uops_1_br_prediction_bpd_resp_info;
  assign rename_stage_io_dec_uops_1_fetch_pc_lob = dec_uops_1_fetch_pc_lob;
  assign rename_stage_io_dec_uops_1_imm_packed = dec_uops_1_imm_packed;
  assign rename_stage_io_dec_uops_1_rob_idx = dec_uops_1_rob_idx;
  assign rename_stage_io_dec_uops_1_ldq_idx = dec_uops_1_ldq_idx;
  assign rename_stage_io_dec_uops_1_stq_idx = dec_uops_1_stq_idx;
  assign rename_stage_io_dec_uops_1_brob_idx = dec_uops_1_brob_idx;
  assign rename_stage_io_dec_uops_1_exception = dec_uops_1_exception;
  assign rename_stage_io_dec_uops_1_exc_cause = dec_uops_1_exc_cause;
  assign rename_stage_io_dec_uops_1_bypassable = dec_uops_1_bypassable;
  assign rename_stage_io_dec_uops_1_mem_cmd = dec_uops_1_mem_cmd;
  assign rename_stage_io_dec_uops_1_mem_typ = dec_uops_1_mem_typ;
  assign rename_stage_io_dec_uops_1_is_fence = dec_uops_1_is_fence;
  assign rename_stage_io_dec_uops_1_is_fencei = dec_uops_1_is_fencei;
  assign rename_stage_io_dec_uops_1_is_store = dec_uops_1_is_store;
  assign rename_stage_io_dec_uops_1_is_amo = dec_uops_1_is_amo;
  assign rename_stage_io_dec_uops_1_is_load = dec_uops_1_is_load;
  assign rename_stage_io_dec_uops_1_is_sys_pc2epc = dec_uops_1_is_sys_pc2epc;
  assign rename_stage_io_dec_uops_1_is_unique = dec_uops_1_is_unique;
  assign rename_stage_io_dec_uops_1_flush_on_commit = dec_uops_1_flush_on_commit;
  assign rename_stage_io_dec_uops_1_ldst = dec_uops_1_ldst;
  assign rename_stage_io_dec_uops_1_lrs1 = dec_uops_1_lrs1;
  assign rename_stage_io_dec_uops_1_lrs2 = dec_uops_1_lrs2;
  assign rename_stage_io_dec_uops_1_lrs3 = dec_uops_1_lrs3;
  assign rename_stage_io_dec_uops_1_ldst_val = dec_uops_1_ldst_val;
  assign rename_stage_io_dec_uops_1_dst_rtype = dec_uops_1_dst_rtype;
  assign rename_stage_io_dec_uops_1_lrs1_rtype = dec_uops_1_lrs1_rtype;
  assign rename_stage_io_dec_uops_1_lrs2_rtype = dec_uops_1_lrs2_rtype;
  assign rename_stage_io_dec_uops_1_frs3_en = dec_uops_1_frs3_en;
  assign rename_stage_io_dec_uops_1_fp_val = dec_uops_1_fp_val;
  assign rename_stage_io_dec_uops_1_fp_single = dec_uops_1_fp_single;
  assign rename_stage_io_dec_uops_1_xcpt_pf_if = dec_uops_1_xcpt_pf_if;
  assign rename_stage_io_dec_uops_1_xcpt_ae_if = dec_uops_1_xcpt_ae_if;
  assign rename_stage_io_dec_uops_1_replay_if = dec_uops_1_replay_if;
  assign rename_stage_io_dec_uops_1_xcpt_ma_if = dec_uops_1_xcpt_ma_if;
  assign rename_stage_io_dec_uops_1_debug_events_fetch_seq = dec_uops_1_debug_events_fetch_seq;
  assign rename_stage_io_ren_pred_info_0_bim_resp_value = _T_2899_0_bim_resp_value;
  assign rename_stage_io_ren_pred_info_0_bim_resp_entry_idx = _T_2899_0_bim_resp_entry_idx;
  assign rename_stage_io_ren_pred_info_0_bim_resp_way_idx = _T_2899_0_bim_resp_way_idx;
  assign rename_stage_io_ren_pred_info_0_bpd_resp_history = _T_2899_0_bpd_resp_history;
  assign rename_stage_io_ren_pred_info_0_bpd_resp_history_ptr = _T_2899_0_bpd_resp_history_ptr;
  assign rename_stage_io_ren_pred_info_1_bim_resp_value = _T_2899_1_bim_resp_value;
  assign rename_stage_io_ren_pred_info_1_bim_resp_entry_idx = _T_2899_1_bim_resp_entry_idx;
  assign rename_stage_io_ren_pred_info_1_bim_resp_way_idx = _T_2899_1_bim_resp_way_idx;
  assign rename_stage_io_ren_pred_info_1_bpd_resp_history = _T_2899_1_bpd_resp_history;
  assign rename_stage_io_ren_pred_info_1_bpd_resp_history_ptr = _T_2899_1_bpd_resp_history_ptr;
  assign rename_stage_io_brinfo_valid = br_unit_brinfo_valid;
  assign rename_stage_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign rename_stage_io_brinfo_mask = br_unit_brinfo_mask;
  assign rename_stage_io_brinfo_tag = br_unit_brinfo_tag;
  assign rename_stage_io_get_pred_br_tag = _T_2923;
  assign rename_stage_io_dis_inst_can_proceed_0 = _T_2886;
  assign rename_stage_io_dis_inst_can_proceed_1 = _T_2887;
  assign rename_stage_io_int_wakeups_0_valid = int_wakeups_0_valid;
  assign rename_stage_io_int_wakeups_0_bits_uop_pdst = int_wakeups_0_bits_uop_pdst;
  assign rename_stage_io_int_wakeups_0_bits_uop_dst_rtype = int_wakeups_0_bits_uop_dst_rtype;
  assign rename_stage_io_int_wakeups_1_valid = int_wakeups_1_valid;
  assign rename_stage_io_int_wakeups_1_bits_uop_pdst = int_wakeups_1_bits_uop_pdst;
  assign rename_stage_io_int_wakeups_1_bits_uop_dst_rtype = int_wakeups_1_bits_uop_dst_rtype;
  assign rename_stage_io_int_wakeups_2_valid = int_wakeups_2_valid;
  assign rename_stage_io_int_wakeups_2_bits_uop_pdst = int_wakeups_2_bits_uop_pdst;
  assign rename_stage_io_int_wakeups_2_bits_uop_dst_rtype = int_wakeups_2_bits_uop_dst_rtype;
  assign rename_stage_io_int_wakeups_3_valid = int_wakeups_3_valid;
  assign rename_stage_io_int_wakeups_3_bits_uop_pdst = int_wakeups_3_bits_uop_pdst;
  assign rename_stage_io_int_wakeups_3_bits_uop_dst_rtype = int_wakeups_3_bits_uop_dst_rtype;
  assign rename_stage_io_int_wakeups_4_valid = int_wakeups_4_valid;
  assign rename_stage_io_int_wakeups_4_bits_uop_pdst = int_wakeups_4_bits_uop_pdst;
  assign rename_stage_io_int_wakeups_4_bits_uop_dst_rtype = int_wakeups_4_bits_uop_dst_rtype;
  assign rename_stage_io_fp_wakeups_0_valid = fp_pipeline_io_wakeups_0_valid;
  assign rename_stage_io_fp_wakeups_0_bits_uop_pdst = fp_pipeline_io_wakeups_0_bits_uop_pdst;
  assign rename_stage_io_fp_wakeups_0_bits_uop_dst_rtype = fp_pipeline_io_wakeups_0_bits_uop_dst_rtype;
  assign rename_stage_io_fp_wakeups_1_valid = fp_pipeline_io_wakeups_1_valid;
  assign rename_stage_io_fp_wakeups_1_bits_uop_pdst = fp_pipeline_io_wakeups_1_bits_uop_pdst;
  assign rename_stage_io_fp_wakeups_1_bits_uop_dst_rtype = fp_pipeline_io_wakeups_1_bits_uop_dst_rtype;
  assign rename_stage_io_com_valids_0 = rob_io_commit_valids_0;
  assign rename_stage_io_com_valids_1 = rob_io_commit_valids_1;
  assign rename_stage_io_com_uops_0_pdst = rob_io_commit_uops_0_pdst;
  assign rename_stage_io_com_uops_0_stale_pdst = rob_io_commit_uops_0_stale_pdst;
  assign rename_stage_io_com_uops_0_ldst = rob_io_commit_uops_0_ldst;
  assign rename_stage_io_com_uops_0_dst_rtype = rob_io_commit_uops_0_dst_rtype;
  assign rename_stage_io_com_uops_1_pdst = rob_io_commit_uops_1_pdst;
  assign rename_stage_io_com_uops_1_stale_pdst = rob_io_commit_uops_1_stale_pdst;
  assign rename_stage_io_com_uops_1_ldst = rob_io_commit_uops_1_ldst;
  assign rename_stage_io_com_uops_1_dst_rtype = rob_io_commit_uops_1_dst_rtype;
  assign rename_stage_io_com_rbk_valids_0 = rob_io_commit_rbk_valids_0;
  assign rename_stage_io_com_rbk_valids_1 = rob_io_commit_rbk_valids_1;
  assign rename_stage_io_debug_rob_empty = rob_io_empty;
  assign rename_stage_clock = clock;
  assign rename_stage_reset = reset;
  assign issue_units_0_io_dis_valids_0 = _T_2997;
  assign issue_units_0_io_dis_valids_1 = _T_3004;
  assign issue_units_0_io_dis_uops_0_valid = dis_uops_0_valid;
  assign issue_units_0_io_dis_uops_0_uopc = dis_uops_0_uopc;
  assign issue_units_0_io_dis_uops_0_inst = dis_uops_0_inst;
  assign issue_units_0_io_dis_uops_0_pc = dis_uops_0_pc;
  assign issue_units_0_io_dis_uops_0_iqtype = dis_uops_0_iqtype;
  assign issue_units_0_io_dis_uops_0_fu_code = dis_uops_0_fu_code;
  assign issue_units_0_io_dis_uops_0_allocate_brtag = dis_uops_0_allocate_brtag;
  assign issue_units_0_io_dis_uops_0_is_br_or_jmp = dis_uops_0_is_br_or_jmp;
  assign issue_units_0_io_dis_uops_0_is_jump = dis_uops_0_is_jump;
  assign issue_units_0_io_dis_uops_0_is_jal = dis_uops_0_is_jal;
  assign issue_units_0_io_dis_uops_0_is_ret = dis_uops_0_is_ret;
  assign issue_units_0_io_dis_uops_0_is_call = dis_uops_0_is_call;
  assign issue_units_0_io_dis_uops_0_br_mask = dis_uops_0_br_mask;
  assign issue_units_0_io_dis_uops_0_br_tag = dis_uops_0_br_tag;
  assign issue_units_0_io_dis_uops_0_br_prediction_btb_blame = dis_uops_0_br_prediction_btb_blame;
  assign issue_units_0_io_dis_uops_0_br_prediction_btb_hit = dis_uops_0_br_prediction_btb_hit;
  assign issue_units_0_io_dis_uops_0_br_prediction_btb_taken = dis_uops_0_br_prediction_btb_taken;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_blame = dis_uops_0_br_prediction_bpd_blame;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_hit = dis_uops_0_br_prediction_bpd_hit;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_taken = dis_uops_0_br_prediction_bpd_taken;
  assign issue_units_0_io_dis_uops_0_br_prediction_bim_resp_value = dis_uops_0_br_prediction_bim_resp_value;
  assign issue_units_0_io_dis_uops_0_br_prediction_bim_resp_entry_idx = dis_uops_0_br_prediction_bim_resp_entry_idx;
  assign issue_units_0_io_dis_uops_0_br_prediction_bim_resp_way_idx = dis_uops_0_br_prediction_bim_resp_way_idx;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_takens = dis_uops_0_br_prediction_bpd_resp_takens;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history = dis_uops_0_br_prediction_bpd_resp_history;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_u = dis_uops_0_br_prediction_bpd_resp_history_u;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_history_ptr = dis_uops_0_br_prediction_bpd_resp_history_ptr;
  assign issue_units_0_io_dis_uops_0_br_prediction_bpd_resp_info = dis_uops_0_br_prediction_bpd_resp_info;
  assign issue_units_0_io_dis_uops_0_stat_brjmp_mispredicted = dis_uops_0_stat_brjmp_mispredicted;
  assign issue_units_0_io_dis_uops_0_stat_btb_made_pred = dis_uops_0_stat_btb_made_pred;
  assign issue_units_0_io_dis_uops_0_stat_btb_mispredicted = dis_uops_0_stat_btb_mispredicted;
  assign issue_units_0_io_dis_uops_0_stat_bpd_made_pred = dis_uops_0_stat_bpd_made_pred;
  assign issue_units_0_io_dis_uops_0_stat_bpd_mispredicted = dis_uops_0_stat_bpd_mispredicted;
  assign issue_units_0_io_dis_uops_0_fetch_pc_lob = dis_uops_0_fetch_pc_lob;
  assign issue_units_0_io_dis_uops_0_imm_packed = dis_uops_0_imm_packed;
  assign issue_units_0_io_dis_uops_0_csr_addr = dis_uops_0_csr_addr;
  assign issue_units_0_io_dis_uops_0_rob_idx = dis_uops_0_rob_idx;
  assign issue_units_0_io_dis_uops_0_ldq_idx = dis_uops_0_ldq_idx;
  assign issue_units_0_io_dis_uops_0_stq_idx = dis_uops_0_stq_idx;
  assign issue_units_0_io_dis_uops_0_brob_idx = dis_uops_0_brob_idx;
  assign issue_units_0_io_dis_uops_0_pdst = dis_uops_0_pdst;
  assign issue_units_0_io_dis_uops_0_pop1 = dis_uops_0_pop1;
  assign issue_units_0_io_dis_uops_0_pop2 = dis_uops_0_pop2;
  assign issue_units_0_io_dis_uops_0_pop3 = dis_uops_0_pop3;
  assign issue_units_0_io_dis_uops_0_prs1_busy = dis_uops_0_prs1_busy;
  assign issue_units_0_io_dis_uops_0_prs2_busy = _GEN_2;
  assign issue_units_0_io_dis_uops_0_prs3_busy = dis_uops_0_prs3_busy;
  assign issue_units_0_io_dis_uops_0_stale_pdst = dis_uops_0_stale_pdst;
  assign issue_units_0_io_dis_uops_0_exception = dis_uops_0_exception;
  assign issue_units_0_io_dis_uops_0_exc_cause = dis_uops_0_exc_cause;
  assign issue_units_0_io_dis_uops_0_bypassable = dis_uops_0_bypassable;
  assign issue_units_0_io_dis_uops_0_mem_cmd = dis_uops_0_mem_cmd;
  assign issue_units_0_io_dis_uops_0_mem_typ = dis_uops_0_mem_typ;
  assign issue_units_0_io_dis_uops_0_is_fence = dis_uops_0_is_fence;
  assign issue_units_0_io_dis_uops_0_is_fencei = dis_uops_0_is_fencei;
  assign issue_units_0_io_dis_uops_0_is_store = dis_uops_0_is_store;
  assign issue_units_0_io_dis_uops_0_is_amo = dis_uops_0_is_amo;
  assign issue_units_0_io_dis_uops_0_is_load = dis_uops_0_is_load;
  assign issue_units_0_io_dis_uops_0_is_sys_pc2epc = dis_uops_0_is_sys_pc2epc;
  assign issue_units_0_io_dis_uops_0_is_unique = dis_uops_0_is_unique;
  assign issue_units_0_io_dis_uops_0_flush_on_commit = dis_uops_0_flush_on_commit;
  assign issue_units_0_io_dis_uops_0_ldst = dis_uops_0_ldst;
  assign issue_units_0_io_dis_uops_0_lrs1 = dis_uops_0_lrs1;
  assign issue_units_0_io_dis_uops_0_lrs2 = dis_uops_0_lrs2;
  assign issue_units_0_io_dis_uops_0_lrs3 = dis_uops_0_lrs3;
  assign issue_units_0_io_dis_uops_0_ldst_val = dis_uops_0_ldst_val;
  assign issue_units_0_io_dis_uops_0_dst_rtype = dis_uops_0_dst_rtype;
  assign issue_units_0_io_dis_uops_0_lrs1_rtype = dis_uops_0_lrs1_rtype;
  assign issue_units_0_io_dis_uops_0_lrs2_rtype = _GEN_1;
  assign issue_units_0_io_dis_uops_0_frs3_en = dis_uops_0_frs3_en;
  assign issue_units_0_io_dis_uops_0_fp_val = dis_uops_0_fp_val;
  assign issue_units_0_io_dis_uops_0_fp_single = dis_uops_0_fp_single;
  assign issue_units_0_io_dis_uops_0_xcpt_pf_if = dis_uops_0_xcpt_pf_if;
  assign issue_units_0_io_dis_uops_0_xcpt_ae_if = dis_uops_0_xcpt_ae_if;
  assign issue_units_0_io_dis_uops_0_replay_if = dis_uops_0_replay_if;
  assign issue_units_0_io_dis_uops_0_xcpt_ma_if = dis_uops_0_xcpt_ma_if;
  assign issue_units_0_io_dis_uops_0_debug_wdata = dis_uops_0_debug_wdata;
  assign issue_units_0_io_dis_uops_0_debug_events_fetch_seq = dis_uops_0_debug_events_fetch_seq;
  assign issue_units_0_io_dis_uops_1_valid = dis_uops_1_valid;
  assign issue_units_0_io_dis_uops_1_uopc = dis_uops_1_uopc;
  assign issue_units_0_io_dis_uops_1_inst = dis_uops_1_inst;
  assign issue_units_0_io_dis_uops_1_pc = dis_uops_1_pc;
  assign issue_units_0_io_dis_uops_1_iqtype = dis_uops_1_iqtype;
  assign issue_units_0_io_dis_uops_1_fu_code = dis_uops_1_fu_code;
  assign issue_units_0_io_dis_uops_1_allocate_brtag = dis_uops_1_allocate_brtag;
  assign issue_units_0_io_dis_uops_1_is_br_or_jmp = dis_uops_1_is_br_or_jmp;
  assign issue_units_0_io_dis_uops_1_is_jump = dis_uops_1_is_jump;
  assign issue_units_0_io_dis_uops_1_is_jal = dis_uops_1_is_jal;
  assign issue_units_0_io_dis_uops_1_is_ret = dis_uops_1_is_ret;
  assign issue_units_0_io_dis_uops_1_is_call = dis_uops_1_is_call;
  assign issue_units_0_io_dis_uops_1_br_mask = dis_uops_1_br_mask;
  assign issue_units_0_io_dis_uops_1_br_tag = dis_uops_1_br_tag;
  assign issue_units_0_io_dis_uops_1_br_prediction_btb_blame = dis_uops_1_br_prediction_btb_blame;
  assign issue_units_0_io_dis_uops_1_br_prediction_btb_hit = dis_uops_1_br_prediction_btb_hit;
  assign issue_units_0_io_dis_uops_1_br_prediction_btb_taken = dis_uops_1_br_prediction_btb_taken;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_blame = dis_uops_1_br_prediction_bpd_blame;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_hit = dis_uops_1_br_prediction_bpd_hit;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_taken = dis_uops_1_br_prediction_bpd_taken;
  assign issue_units_0_io_dis_uops_1_br_prediction_bim_resp_value = dis_uops_1_br_prediction_bim_resp_value;
  assign issue_units_0_io_dis_uops_1_br_prediction_bim_resp_entry_idx = dis_uops_1_br_prediction_bim_resp_entry_idx;
  assign issue_units_0_io_dis_uops_1_br_prediction_bim_resp_way_idx = dis_uops_1_br_prediction_bim_resp_way_idx;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_takens = dis_uops_1_br_prediction_bpd_resp_takens;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history = dis_uops_1_br_prediction_bpd_resp_history;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_u = dis_uops_1_br_prediction_bpd_resp_history_u;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_history_ptr = dis_uops_1_br_prediction_bpd_resp_history_ptr;
  assign issue_units_0_io_dis_uops_1_br_prediction_bpd_resp_info = dis_uops_1_br_prediction_bpd_resp_info;
  assign issue_units_0_io_dis_uops_1_stat_brjmp_mispredicted = dis_uops_1_stat_brjmp_mispredicted;
  assign issue_units_0_io_dis_uops_1_stat_btb_made_pred = dis_uops_1_stat_btb_made_pred;
  assign issue_units_0_io_dis_uops_1_stat_btb_mispredicted = dis_uops_1_stat_btb_mispredicted;
  assign issue_units_0_io_dis_uops_1_stat_bpd_made_pred = dis_uops_1_stat_bpd_made_pred;
  assign issue_units_0_io_dis_uops_1_stat_bpd_mispredicted = dis_uops_1_stat_bpd_mispredicted;
  assign issue_units_0_io_dis_uops_1_fetch_pc_lob = dis_uops_1_fetch_pc_lob;
  assign issue_units_0_io_dis_uops_1_imm_packed = dis_uops_1_imm_packed;
  assign issue_units_0_io_dis_uops_1_csr_addr = dis_uops_1_csr_addr;
  assign issue_units_0_io_dis_uops_1_rob_idx = dis_uops_1_rob_idx;
  assign issue_units_0_io_dis_uops_1_ldq_idx = dis_uops_1_ldq_idx;
  assign issue_units_0_io_dis_uops_1_stq_idx = dis_uops_1_stq_idx;
  assign issue_units_0_io_dis_uops_1_brob_idx = dis_uops_1_brob_idx;
  assign issue_units_0_io_dis_uops_1_pdst = dis_uops_1_pdst;
  assign issue_units_0_io_dis_uops_1_pop1 = dis_uops_1_pop1;
  assign issue_units_0_io_dis_uops_1_pop2 = dis_uops_1_pop2;
  assign issue_units_0_io_dis_uops_1_pop3 = dis_uops_1_pop3;
  assign issue_units_0_io_dis_uops_1_prs1_busy = dis_uops_1_prs1_busy;
  assign issue_units_0_io_dis_uops_1_prs2_busy = _GEN_4;
  assign issue_units_0_io_dis_uops_1_prs3_busy = dis_uops_1_prs3_busy;
  assign issue_units_0_io_dis_uops_1_stale_pdst = dis_uops_1_stale_pdst;
  assign issue_units_0_io_dis_uops_1_exception = dis_uops_1_exception;
  assign issue_units_0_io_dis_uops_1_exc_cause = dis_uops_1_exc_cause;
  assign issue_units_0_io_dis_uops_1_bypassable = dis_uops_1_bypassable;
  assign issue_units_0_io_dis_uops_1_mem_cmd = dis_uops_1_mem_cmd;
  assign issue_units_0_io_dis_uops_1_mem_typ = dis_uops_1_mem_typ;
  assign issue_units_0_io_dis_uops_1_is_fence = dis_uops_1_is_fence;
  assign issue_units_0_io_dis_uops_1_is_fencei = dis_uops_1_is_fencei;
  assign issue_units_0_io_dis_uops_1_is_store = dis_uops_1_is_store;
  assign issue_units_0_io_dis_uops_1_is_amo = dis_uops_1_is_amo;
  assign issue_units_0_io_dis_uops_1_is_load = dis_uops_1_is_load;
  assign issue_units_0_io_dis_uops_1_is_sys_pc2epc = dis_uops_1_is_sys_pc2epc;
  assign issue_units_0_io_dis_uops_1_is_unique = dis_uops_1_is_unique;
  assign issue_units_0_io_dis_uops_1_flush_on_commit = dis_uops_1_flush_on_commit;
  assign issue_units_0_io_dis_uops_1_ldst = dis_uops_1_ldst;
  assign issue_units_0_io_dis_uops_1_lrs1 = dis_uops_1_lrs1;
  assign issue_units_0_io_dis_uops_1_lrs2 = dis_uops_1_lrs2;
  assign issue_units_0_io_dis_uops_1_lrs3 = dis_uops_1_lrs3;
  assign issue_units_0_io_dis_uops_1_ldst_val = dis_uops_1_ldst_val;
  assign issue_units_0_io_dis_uops_1_dst_rtype = dis_uops_1_dst_rtype;
  assign issue_units_0_io_dis_uops_1_lrs1_rtype = dis_uops_1_lrs1_rtype;
  assign issue_units_0_io_dis_uops_1_lrs2_rtype = _GEN_3;
  assign issue_units_0_io_dis_uops_1_frs3_en = dis_uops_1_frs3_en;
  assign issue_units_0_io_dis_uops_1_fp_val = dis_uops_1_fp_val;
  assign issue_units_0_io_dis_uops_1_fp_single = dis_uops_1_fp_single;
  assign issue_units_0_io_dis_uops_1_xcpt_pf_if = dis_uops_1_xcpt_pf_if;
  assign issue_units_0_io_dis_uops_1_xcpt_ae_if = dis_uops_1_xcpt_ae_if;
  assign issue_units_0_io_dis_uops_1_replay_if = dis_uops_1_replay_if;
  assign issue_units_0_io_dis_uops_1_xcpt_ma_if = dis_uops_1_xcpt_ma_if;
  assign issue_units_0_io_dis_uops_1_debug_wdata = dis_uops_1_debug_wdata;
  assign issue_units_0_io_dis_uops_1_debug_events_fetch_seq = dis_uops_1_debug_events_fetch_seq;
  assign issue_units_0_io_wakeup_pdsts_0_valid = int_wakeups_0_valid;
  assign issue_units_0_io_wakeup_pdsts_0_bits = int_wakeups_0_bits_uop_pdst;
  assign issue_units_0_io_wakeup_pdsts_1_valid = int_wakeups_1_valid;
  assign issue_units_0_io_wakeup_pdsts_1_bits = int_wakeups_1_bits_uop_pdst;
  assign issue_units_0_io_wakeup_pdsts_2_valid = int_wakeups_2_valid;
  assign issue_units_0_io_wakeup_pdsts_2_bits = int_wakeups_2_bits_uop_pdst;
  assign issue_units_0_io_wakeup_pdsts_3_valid = int_wakeups_3_valid;
  assign issue_units_0_io_wakeup_pdsts_3_bits = int_wakeups_3_bits_uop_pdst;
  assign issue_units_0_io_wakeup_pdsts_4_valid = int_wakeups_4_valid;
  assign issue_units_0_io_wakeup_pdsts_4_bits = int_wakeups_4_bits_uop_pdst;
  assign issue_units_0_io_brinfo_valid = br_unit_brinfo_valid;
  assign issue_units_0_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign issue_units_0_io_brinfo_mask = br_unit_brinfo_mask;
  assign issue_units_0_io_flush_pipeline = rob_io_flush_valid;
  assign issue_units_0_clock = clock;
  assign issue_units_0_reset = reset;
  assign issue_units_1_io_dis_valids_0 = _T_3011;
  assign issue_units_1_io_dis_valids_1 = _T_3018;
  assign issue_units_1_io_dis_uops_0_valid = dis_uops_0_valid;
  assign issue_units_1_io_dis_uops_0_uopc = dis_uops_0_uopc;
  assign issue_units_1_io_dis_uops_0_inst = dis_uops_0_inst;
  assign issue_units_1_io_dis_uops_0_pc = dis_uops_0_pc;
  assign issue_units_1_io_dis_uops_0_iqtype = dis_uops_0_iqtype;
  assign issue_units_1_io_dis_uops_0_fu_code = dis_uops_0_fu_code;
  assign issue_units_1_io_dis_uops_0_allocate_brtag = dis_uops_0_allocate_brtag;
  assign issue_units_1_io_dis_uops_0_is_br_or_jmp = dis_uops_0_is_br_or_jmp;
  assign issue_units_1_io_dis_uops_0_is_jump = dis_uops_0_is_jump;
  assign issue_units_1_io_dis_uops_0_is_jal = dis_uops_0_is_jal;
  assign issue_units_1_io_dis_uops_0_is_ret = dis_uops_0_is_ret;
  assign issue_units_1_io_dis_uops_0_is_call = dis_uops_0_is_call;
  assign issue_units_1_io_dis_uops_0_br_mask = dis_uops_0_br_mask;
  assign issue_units_1_io_dis_uops_0_br_tag = dis_uops_0_br_tag;
  assign issue_units_1_io_dis_uops_0_br_prediction_btb_blame = dis_uops_0_br_prediction_btb_blame;
  assign issue_units_1_io_dis_uops_0_br_prediction_btb_hit = dis_uops_0_br_prediction_btb_hit;
  assign issue_units_1_io_dis_uops_0_br_prediction_btb_taken = dis_uops_0_br_prediction_btb_taken;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_blame = dis_uops_0_br_prediction_bpd_blame;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_hit = dis_uops_0_br_prediction_bpd_hit;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_taken = dis_uops_0_br_prediction_bpd_taken;
  assign issue_units_1_io_dis_uops_0_br_prediction_bim_resp_value = dis_uops_0_br_prediction_bim_resp_value;
  assign issue_units_1_io_dis_uops_0_br_prediction_bim_resp_entry_idx = dis_uops_0_br_prediction_bim_resp_entry_idx;
  assign issue_units_1_io_dis_uops_0_br_prediction_bim_resp_way_idx = dis_uops_0_br_prediction_bim_resp_way_idx;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_takens = dis_uops_0_br_prediction_bpd_resp_takens;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history = dis_uops_0_br_prediction_bpd_resp_history;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_u = dis_uops_0_br_prediction_bpd_resp_history_u;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_history_ptr = dis_uops_0_br_prediction_bpd_resp_history_ptr;
  assign issue_units_1_io_dis_uops_0_br_prediction_bpd_resp_info = dis_uops_0_br_prediction_bpd_resp_info;
  assign issue_units_1_io_dis_uops_0_stat_brjmp_mispredicted = dis_uops_0_stat_brjmp_mispredicted;
  assign issue_units_1_io_dis_uops_0_stat_btb_made_pred = dis_uops_0_stat_btb_made_pred;
  assign issue_units_1_io_dis_uops_0_stat_btb_mispredicted = dis_uops_0_stat_btb_mispredicted;
  assign issue_units_1_io_dis_uops_0_stat_bpd_made_pred = dis_uops_0_stat_bpd_made_pred;
  assign issue_units_1_io_dis_uops_0_stat_bpd_mispredicted = dis_uops_0_stat_bpd_mispredicted;
  assign issue_units_1_io_dis_uops_0_fetch_pc_lob = dis_uops_0_fetch_pc_lob;
  assign issue_units_1_io_dis_uops_0_imm_packed = dis_uops_0_imm_packed;
  assign issue_units_1_io_dis_uops_0_csr_addr = dis_uops_0_csr_addr;
  assign issue_units_1_io_dis_uops_0_rob_idx = dis_uops_0_rob_idx;
  assign issue_units_1_io_dis_uops_0_ldq_idx = dis_uops_0_ldq_idx;
  assign issue_units_1_io_dis_uops_0_stq_idx = dis_uops_0_stq_idx;
  assign issue_units_1_io_dis_uops_0_brob_idx = dis_uops_0_brob_idx;
  assign issue_units_1_io_dis_uops_0_pdst = dis_uops_0_pdst;
  assign issue_units_1_io_dis_uops_0_pop1 = dis_uops_0_pop1;
  assign issue_units_1_io_dis_uops_0_pop2 = dis_uops_0_pop2;
  assign issue_units_1_io_dis_uops_0_pop3 = dis_uops_0_pop3;
  assign issue_units_1_io_dis_uops_0_prs1_busy = dis_uops_0_prs1_busy;
  assign issue_units_1_io_dis_uops_0_prs2_busy = _GEN_2;
  assign issue_units_1_io_dis_uops_0_prs3_busy = dis_uops_0_prs3_busy;
  assign issue_units_1_io_dis_uops_0_stale_pdst = dis_uops_0_stale_pdst;
  assign issue_units_1_io_dis_uops_0_exception = dis_uops_0_exception;
  assign issue_units_1_io_dis_uops_0_exc_cause = dis_uops_0_exc_cause;
  assign issue_units_1_io_dis_uops_0_bypassable = dis_uops_0_bypassable;
  assign issue_units_1_io_dis_uops_0_mem_cmd = dis_uops_0_mem_cmd;
  assign issue_units_1_io_dis_uops_0_mem_typ = dis_uops_0_mem_typ;
  assign issue_units_1_io_dis_uops_0_is_fence = dis_uops_0_is_fence;
  assign issue_units_1_io_dis_uops_0_is_fencei = dis_uops_0_is_fencei;
  assign issue_units_1_io_dis_uops_0_is_store = dis_uops_0_is_store;
  assign issue_units_1_io_dis_uops_0_is_amo = dis_uops_0_is_amo;
  assign issue_units_1_io_dis_uops_0_is_load = dis_uops_0_is_load;
  assign issue_units_1_io_dis_uops_0_is_sys_pc2epc = dis_uops_0_is_sys_pc2epc;
  assign issue_units_1_io_dis_uops_0_is_unique = dis_uops_0_is_unique;
  assign issue_units_1_io_dis_uops_0_flush_on_commit = dis_uops_0_flush_on_commit;
  assign issue_units_1_io_dis_uops_0_ldst = dis_uops_0_ldst;
  assign issue_units_1_io_dis_uops_0_lrs1 = dis_uops_0_lrs1;
  assign issue_units_1_io_dis_uops_0_lrs2 = dis_uops_0_lrs2;
  assign issue_units_1_io_dis_uops_0_lrs3 = dis_uops_0_lrs3;
  assign issue_units_1_io_dis_uops_0_ldst_val = dis_uops_0_ldst_val;
  assign issue_units_1_io_dis_uops_0_dst_rtype = dis_uops_0_dst_rtype;
  assign issue_units_1_io_dis_uops_0_lrs1_rtype = dis_uops_0_lrs1_rtype;
  assign issue_units_1_io_dis_uops_0_lrs2_rtype = _GEN_1;
  assign issue_units_1_io_dis_uops_0_frs3_en = dis_uops_0_frs3_en;
  assign issue_units_1_io_dis_uops_0_fp_val = dis_uops_0_fp_val;
  assign issue_units_1_io_dis_uops_0_fp_single = dis_uops_0_fp_single;
  assign issue_units_1_io_dis_uops_0_xcpt_pf_if = dis_uops_0_xcpt_pf_if;
  assign issue_units_1_io_dis_uops_0_xcpt_ae_if = dis_uops_0_xcpt_ae_if;
  assign issue_units_1_io_dis_uops_0_replay_if = dis_uops_0_replay_if;
  assign issue_units_1_io_dis_uops_0_xcpt_ma_if = dis_uops_0_xcpt_ma_if;
  assign issue_units_1_io_dis_uops_0_debug_wdata = dis_uops_0_debug_wdata;
  assign issue_units_1_io_dis_uops_0_debug_events_fetch_seq = dis_uops_0_debug_events_fetch_seq;
  assign issue_units_1_io_dis_uops_1_valid = dis_uops_1_valid;
  assign issue_units_1_io_dis_uops_1_uopc = dis_uops_1_uopc;
  assign issue_units_1_io_dis_uops_1_inst = dis_uops_1_inst;
  assign issue_units_1_io_dis_uops_1_pc = dis_uops_1_pc;
  assign issue_units_1_io_dis_uops_1_iqtype = dis_uops_1_iqtype;
  assign issue_units_1_io_dis_uops_1_fu_code = dis_uops_1_fu_code;
  assign issue_units_1_io_dis_uops_1_allocate_brtag = dis_uops_1_allocate_brtag;
  assign issue_units_1_io_dis_uops_1_is_br_or_jmp = dis_uops_1_is_br_or_jmp;
  assign issue_units_1_io_dis_uops_1_is_jump = dis_uops_1_is_jump;
  assign issue_units_1_io_dis_uops_1_is_jal = dis_uops_1_is_jal;
  assign issue_units_1_io_dis_uops_1_is_ret = dis_uops_1_is_ret;
  assign issue_units_1_io_dis_uops_1_is_call = dis_uops_1_is_call;
  assign issue_units_1_io_dis_uops_1_br_mask = dis_uops_1_br_mask;
  assign issue_units_1_io_dis_uops_1_br_tag = dis_uops_1_br_tag;
  assign issue_units_1_io_dis_uops_1_br_prediction_btb_blame = dis_uops_1_br_prediction_btb_blame;
  assign issue_units_1_io_dis_uops_1_br_prediction_btb_hit = dis_uops_1_br_prediction_btb_hit;
  assign issue_units_1_io_dis_uops_1_br_prediction_btb_taken = dis_uops_1_br_prediction_btb_taken;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_blame = dis_uops_1_br_prediction_bpd_blame;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_hit = dis_uops_1_br_prediction_bpd_hit;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_taken = dis_uops_1_br_prediction_bpd_taken;
  assign issue_units_1_io_dis_uops_1_br_prediction_bim_resp_value = dis_uops_1_br_prediction_bim_resp_value;
  assign issue_units_1_io_dis_uops_1_br_prediction_bim_resp_entry_idx = dis_uops_1_br_prediction_bim_resp_entry_idx;
  assign issue_units_1_io_dis_uops_1_br_prediction_bim_resp_way_idx = dis_uops_1_br_prediction_bim_resp_way_idx;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_takens = dis_uops_1_br_prediction_bpd_resp_takens;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history = dis_uops_1_br_prediction_bpd_resp_history;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_u = dis_uops_1_br_prediction_bpd_resp_history_u;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_history_ptr = dis_uops_1_br_prediction_bpd_resp_history_ptr;
  assign issue_units_1_io_dis_uops_1_br_prediction_bpd_resp_info = dis_uops_1_br_prediction_bpd_resp_info;
  assign issue_units_1_io_dis_uops_1_stat_brjmp_mispredicted = dis_uops_1_stat_brjmp_mispredicted;
  assign issue_units_1_io_dis_uops_1_stat_btb_made_pred = dis_uops_1_stat_btb_made_pred;
  assign issue_units_1_io_dis_uops_1_stat_btb_mispredicted = dis_uops_1_stat_btb_mispredicted;
  assign issue_units_1_io_dis_uops_1_stat_bpd_made_pred = dis_uops_1_stat_bpd_made_pred;
  assign issue_units_1_io_dis_uops_1_stat_bpd_mispredicted = dis_uops_1_stat_bpd_mispredicted;
  assign issue_units_1_io_dis_uops_1_fetch_pc_lob = dis_uops_1_fetch_pc_lob;
  assign issue_units_1_io_dis_uops_1_imm_packed = dis_uops_1_imm_packed;
  assign issue_units_1_io_dis_uops_1_csr_addr = dis_uops_1_csr_addr;
  assign issue_units_1_io_dis_uops_1_rob_idx = dis_uops_1_rob_idx;
  assign issue_units_1_io_dis_uops_1_ldq_idx = dis_uops_1_ldq_idx;
  assign issue_units_1_io_dis_uops_1_stq_idx = dis_uops_1_stq_idx;
  assign issue_units_1_io_dis_uops_1_brob_idx = dis_uops_1_brob_idx;
  assign issue_units_1_io_dis_uops_1_pdst = dis_uops_1_pdst;
  assign issue_units_1_io_dis_uops_1_pop1 = dis_uops_1_pop1;
  assign issue_units_1_io_dis_uops_1_pop2 = dis_uops_1_pop2;
  assign issue_units_1_io_dis_uops_1_pop3 = dis_uops_1_pop3;
  assign issue_units_1_io_dis_uops_1_prs1_busy = dis_uops_1_prs1_busy;
  assign issue_units_1_io_dis_uops_1_prs2_busy = _GEN_4;
  assign issue_units_1_io_dis_uops_1_prs3_busy = dis_uops_1_prs3_busy;
  assign issue_units_1_io_dis_uops_1_stale_pdst = dis_uops_1_stale_pdst;
  assign issue_units_1_io_dis_uops_1_exception = dis_uops_1_exception;
  assign issue_units_1_io_dis_uops_1_exc_cause = dis_uops_1_exc_cause;
  assign issue_units_1_io_dis_uops_1_bypassable = dis_uops_1_bypassable;
  assign issue_units_1_io_dis_uops_1_mem_cmd = dis_uops_1_mem_cmd;
  assign issue_units_1_io_dis_uops_1_mem_typ = dis_uops_1_mem_typ;
  assign issue_units_1_io_dis_uops_1_is_fence = dis_uops_1_is_fence;
  assign issue_units_1_io_dis_uops_1_is_fencei = dis_uops_1_is_fencei;
  assign issue_units_1_io_dis_uops_1_is_store = dis_uops_1_is_store;
  assign issue_units_1_io_dis_uops_1_is_amo = dis_uops_1_is_amo;
  assign issue_units_1_io_dis_uops_1_is_load = dis_uops_1_is_load;
  assign issue_units_1_io_dis_uops_1_is_sys_pc2epc = dis_uops_1_is_sys_pc2epc;
  assign issue_units_1_io_dis_uops_1_is_unique = dis_uops_1_is_unique;
  assign issue_units_1_io_dis_uops_1_flush_on_commit = dis_uops_1_flush_on_commit;
  assign issue_units_1_io_dis_uops_1_ldst = dis_uops_1_ldst;
  assign issue_units_1_io_dis_uops_1_lrs1 = dis_uops_1_lrs1;
  assign issue_units_1_io_dis_uops_1_lrs2 = dis_uops_1_lrs2;
  assign issue_units_1_io_dis_uops_1_lrs3 = dis_uops_1_lrs3;
  assign issue_units_1_io_dis_uops_1_ldst_val = dis_uops_1_ldst_val;
  assign issue_units_1_io_dis_uops_1_dst_rtype = dis_uops_1_dst_rtype;
  assign issue_units_1_io_dis_uops_1_lrs1_rtype = dis_uops_1_lrs1_rtype;
  assign issue_units_1_io_dis_uops_1_lrs2_rtype = _GEN_3;
  assign issue_units_1_io_dis_uops_1_frs3_en = dis_uops_1_frs3_en;
  assign issue_units_1_io_dis_uops_1_fp_val = dis_uops_1_fp_val;
  assign issue_units_1_io_dis_uops_1_fp_single = dis_uops_1_fp_single;
  assign issue_units_1_io_dis_uops_1_xcpt_pf_if = dis_uops_1_xcpt_pf_if;
  assign issue_units_1_io_dis_uops_1_xcpt_ae_if = dis_uops_1_xcpt_ae_if;
  assign issue_units_1_io_dis_uops_1_replay_if = dis_uops_1_replay_if;
  assign issue_units_1_io_dis_uops_1_xcpt_ma_if = dis_uops_1_xcpt_ma_if;
  assign issue_units_1_io_dis_uops_1_debug_wdata = dis_uops_1_debug_wdata;
  assign issue_units_1_io_dis_uops_1_debug_events_fetch_seq = dis_uops_1_debug_events_fetch_seq;
  assign issue_units_1_io_wakeup_pdsts_0_valid = int_wakeups_0_valid;
  assign issue_units_1_io_wakeup_pdsts_0_bits = int_wakeups_0_bits_uop_pdst;
  assign issue_units_1_io_wakeup_pdsts_1_valid = int_wakeups_1_valid;
  assign issue_units_1_io_wakeup_pdsts_1_bits = int_wakeups_1_bits_uop_pdst;
  assign issue_units_1_io_wakeup_pdsts_2_valid = int_wakeups_2_valid;
  assign issue_units_1_io_wakeup_pdsts_2_bits = int_wakeups_2_bits_uop_pdst;
  assign issue_units_1_io_wakeup_pdsts_3_valid = int_wakeups_3_valid;
  assign issue_units_1_io_wakeup_pdsts_3_bits = int_wakeups_3_bits_uop_pdst;
  assign issue_units_1_io_wakeup_pdsts_4_valid = int_wakeups_4_valid;
  assign issue_units_1_io_wakeup_pdsts_4_bits = int_wakeups_4_bits_uop_pdst;
  assign issue_units_1_io_fu_types_0 = _T_3030;
  assign issue_units_1_io_brinfo_valid = br_unit_brinfo_valid;
  assign issue_units_1_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign issue_units_1_io_brinfo_mask = br_unit_brinfo_mask;
  assign issue_units_1_io_flush_pipeline = rob_io_flush_valid;
  assign issue_units_1_clock = clock;
  assign issue_units_1_reset = reset;
  assign iregfile_io_read_ports_0_addr = iregister_read_io_rf_read_ports_0_addr;
  assign iregfile_io_read_ports_1_addr = iregister_read_io_rf_read_ports_1_addr;
  assign iregfile_io_read_ports_2_addr = iregister_read_io_rf_read_ports_2_addr;
  assign iregfile_io_read_ports_3_addr = iregister_read_io_rf_read_ports_3_addr;
  assign iregfile_io_read_ports_4_addr = iregister_read_io_rf_read_ports_4_addr;
  assign iregfile_io_read_ports_5_addr = iregister_read_io_rf_read_ports_5_addr;
  assign iregfile_io_write_ports_0_valid = _T_3175_valid;
  assign iregfile_io_write_ports_0_bits_addr = _T_3175_bits_addr;
  assign iregfile_io_write_ports_0_bits_data = _T_3175_bits_data;
  assign iregfile_io_write_ports_1_valid = _T_3095;
  assign iregfile_io_write_ports_1_bits_addr = csr_exe_unit_io_resp_0_bits_uop_pdst;
  assign iregfile_io_write_ports_1_bits_data = _T_3096;
  assign iregfile_io_write_ports_2_valid = _T_3130;
  assign iregfile_io_write_ports_2_bits_addr = ALUExeUnit_io_resp_0_bits_uop_pdst;
  assign iregfile_io_write_ports_2_bits_data = ALUExeUnit_io_resp_0_bits_data;
  assign iregfile_clock = clock;
  assign ll_wbarb_io_in_0_valid = _T_3066;
  assign ll_wbarb_io_in_0_bits_uop_rob_idx = mem_unit_io_resp_0_bits_uop_rob_idx;
  assign ll_wbarb_io_in_0_bits_uop_pdst = mem_unit_io_resp_0_bits_uop_pdst;
  assign ll_wbarb_io_in_0_bits_uop_is_store = mem_unit_io_resp_0_bits_uop_is_store;
  assign ll_wbarb_io_in_0_bits_uop_is_amo = mem_unit_io_resp_0_bits_uop_is_amo;
  assign ll_wbarb_io_in_0_bits_uop_dst_rtype = mem_unit_io_resp_0_bits_uop_dst_rtype;
  assign ll_wbarb_io_in_0_bits_data = mem_unit_io_resp_0_bits_data[63:0];
  assign ll_wbarb_io_in_1_valid = fp_pipeline_io_toint_valid;
  assign ll_wbarb_io_in_1_bits_uop_rob_idx = fp_pipeline_io_toint_bits_uop_rob_idx;
  assign ll_wbarb_io_in_1_bits_uop_pdst = fp_pipeline_io_toint_bits_uop_pdst;
  assign ll_wbarb_io_in_1_bits_uop_is_store = fp_pipeline_io_toint_bits_uop_is_store;
  assign ll_wbarb_io_in_1_bits_uop_is_amo = fp_pipeline_io_toint_bits_uop_is_amo;
  assign ll_wbarb_io_in_1_bits_uop_dst_rtype = fp_pipeline_io_toint_bits_uop_dst_rtype;
  assign ll_wbarb_io_in_1_bits_data = fp_pipeline_io_toint_bits_data;
  assign ll_wbarb_io_out_ready = 1'h1;
  assign iregister_read_io_iss_valids_0 = iss_valids_0;
  assign iregister_read_io_iss_valids_1 = iss_valids_1;
  assign iregister_read_io_iss_valids_2 = iss_valids_2;
  assign iregister_read_io_iss_uops_0_uopc = iss_uops_0_uopc;
  assign iregister_read_io_iss_uops_0_br_mask = iss_uops_0_br_mask;
  assign iregister_read_io_iss_uops_0_imm_packed = iss_uops_0_imm_packed;
  assign iregister_read_io_iss_uops_0_rob_idx = iss_uops_0_rob_idx;
  assign iregister_read_io_iss_uops_0_ldq_idx = iss_uops_0_ldq_idx;
  assign iregister_read_io_iss_uops_0_stq_idx = iss_uops_0_stq_idx;
  assign iregister_read_io_iss_uops_0_pdst = iss_uops_0_pdst;
  assign iregister_read_io_iss_uops_0_pop1 = iss_uops_0_pop1;
  assign iregister_read_io_iss_uops_0_pop2 = iss_uops_0_pop2;
  assign iregister_read_io_iss_uops_0_mem_cmd = iss_uops_0_mem_cmd;
  assign iregister_read_io_iss_uops_0_mem_typ = iss_uops_0_mem_typ;
  assign iregister_read_io_iss_uops_0_is_fence = iss_uops_0_is_fence;
  assign iregister_read_io_iss_uops_0_is_store = iss_uops_0_is_store;
  assign iregister_read_io_iss_uops_0_is_amo = iss_uops_0_is_amo;
  assign iregister_read_io_iss_uops_0_is_load = iss_uops_0_is_load;
  assign iregister_read_io_iss_uops_0_dst_rtype = iss_uops_0_dst_rtype;
  assign iregister_read_io_iss_uops_0_lrs1_rtype = iss_uops_0_lrs1_rtype;
  assign iregister_read_io_iss_uops_0_lrs2_rtype = iss_uops_0_lrs2_rtype;
  assign iregister_read_io_iss_uops_0_fp_val = iss_uops_0_fp_val;
  assign iregister_read_io_iss_uops_1_valid = iss_uops_1_valid;
  assign iregister_read_io_iss_uops_1_iw_state = iss_uops_1_iw_state;
  assign iregister_read_io_iss_uops_1_uopc = iss_uops_1_uopc;
  assign iregister_read_io_iss_uops_1_inst = iss_uops_1_inst;
  assign iregister_read_io_iss_uops_1_pc = iss_uops_1_pc;
  assign iregister_read_io_iss_uops_1_iqtype = iss_uops_1_iqtype;
  assign iregister_read_io_iss_uops_1_fu_code = iss_uops_1_fu_code;
  assign iregister_read_io_iss_uops_1_allocate_brtag = iss_uops_1_allocate_brtag;
  assign iregister_read_io_iss_uops_1_is_br_or_jmp = iss_uops_1_is_br_or_jmp;
  assign iregister_read_io_iss_uops_1_is_jump = iss_uops_1_is_jump;
  assign iregister_read_io_iss_uops_1_is_jal = iss_uops_1_is_jal;
  assign iregister_read_io_iss_uops_1_is_ret = iss_uops_1_is_ret;
  assign iregister_read_io_iss_uops_1_is_call = iss_uops_1_is_call;
  assign iregister_read_io_iss_uops_1_br_mask = iss_uops_1_br_mask;
  assign iregister_read_io_iss_uops_1_br_tag = iss_uops_1_br_tag;
  assign iregister_read_io_iss_uops_1_br_prediction_btb_blame = iss_uops_1_br_prediction_btb_blame;
  assign iregister_read_io_iss_uops_1_br_prediction_btb_hit = iss_uops_1_br_prediction_btb_hit;
  assign iregister_read_io_iss_uops_1_br_prediction_btb_taken = iss_uops_1_br_prediction_btb_taken;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_blame = iss_uops_1_br_prediction_bpd_blame;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_hit = iss_uops_1_br_prediction_bpd_hit;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_taken = iss_uops_1_br_prediction_bpd_taken;
  assign iregister_read_io_iss_uops_1_br_prediction_bim_resp_value = iss_uops_1_br_prediction_bim_resp_value;
  assign iregister_read_io_iss_uops_1_br_prediction_bim_resp_entry_idx = iss_uops_1_br_prediction_bim_resp_entry_idx;
  assign iregister_read_io_iss_uops_1_br_prediction_bim_resp_way_idx = iss_uops_1_br_prediction_bim_resp_way_idx;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_resp_takens = iss_uops_1_br_prediction_bpd_resp_takens;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history = iss_uops_1_br_prediction_bpd_resp_history;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_u = iss_uops_1_br_prediction_bpd_resp_history_u;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_resp_history_ptr = iss_uops_1_br_prediction_bpd_resp_history_ptr;
  assign iregister_read_io_iss_uops_1_br_prediction_bpd_resp_info = iss_uops_1_br_prediction_bpd_resp_info;
  assign iregister_read_io_iss_uops_1_stat_brjmp_mispredicted = iss_uops_1_stat_brjmp_mispredicted;
  assign iregister_read_io_iss_uops_1_stat_btb_made_pred = iss_uops_1_stat_btb_made_pred;
  assign iregister_read_io_iss_uops_1_stat_btb_mispredicted = iss_uops_1_stat_btb_mispredicted;
  assign iregister_read_io_iss_uops_1_stat_bpd_made_pred = iss_uops_1_stat_bpd_made_pred;
  assign iregister_read_io_iss_uops_1_stat_bpd_mispredicted = iss_uops_1_stat_bpd_mispredicted;
  assign iregister_read_io_iss_uops_1_fetch_pc_lob = iss_uops_1_fetch_pc_lob;
  assign iregister_read_io_iss_uops_1_imm_packed = iss_uops_1_imm_packed;
  assign iregister_read_io_iss_uops_1_csr_addr = iss_uops_1_csr_addr;
  assign iregister_read_io_iss_uops_1_rob_idx = iss_uops_1_rob_idx;
  assign iregister_read_io_iss_uops_1_ldq_idx = iss_uops_1_ldq_idx;
  assign iregister_read_io_iss_uops_1_stq_idx = iss_uops_1_stq_idx;
  assign iregister_read_io_iss_uops_1_brob_idx = iss_uops_1_brob_idx;
  assign iregister_read_io_iss_uops_1_pdst = iss_uops_1_pdst;
  assign iregister_read_io_iss_uops_1_pop1 = iss_uops_1_pop1;
  assign iregister_read_io_iss_uops_1_pop2 = iss_uops_1_pop2;
  assign iregister_read_io_iss_uops_1_pop3 = iss_uops_1_pop3;
  assign iregister_read_io_iss_uops_1_prs1_busy = iss_uops_1_prs1_busy;
  assign iregister_read_io_iss_uops_1_prs2_busy = iss_uops_1_prs2_busy;
  assign iregister_read_io_iss_uops_1_prs3_busy = iss_uops_1_prs3_busy;
  assign iregister_read_io_iss_uops_1_stale_pdst = iss_uops_1_stale_pdst;
  assign iregister_read_io_iss_uops_1_exception = iss_uops_1_exception;
  assign iregister_read_io_iss_uops_1_exc_cause = iss_uops_1_exc_cause;
  assign iregister_read_io_iss_uops_1_bypassable = iss_uops_1_bypassable;
  assign iregister_read_io_iss_uops_1_mem_cmd = iss_uops_1_mem_cmd;
  assign iregister_read_io_iss_uops_1_mem_typ = iss_uops_1_mem_typ;
  assign iregister_read_io_iss_uops_1_is_fence = iss_uops_1_is_fence;
  assign iregister_read_io_iss_uops_1_is_fencei = iss_uops_1_is_fencei;
  assign iregister_read_io_iss_uops_1_is_store = iss_uops_1_is_store;
  assign iregister_read_io_iss_uops_1_is_amo = iss_uops_1_is_amo;
  assign iregister_read_io_iss_uops_1_is_load = iss_uops_1_is_load;
  assign iregister_read_io_iss_uops_1_is_sys_pc2epc = iss_uops_1_is_sys_pc2epc;
  assign iregister_read_io_iss_uops_1_is_unique = iss_uops_1_is_unique;
  assign iregister_read_io_iss_uops_1_flush_on_commit = iss_uops_1_flush_on_commit;
  assign iregister_read_io_iss_uops_1_ldst = iss_uops_1_ldst;
  assign iregister_read_io_iss_uops_1_lrs1 = iss_uops_1_lrs1;
  assign iregister_read_io_iss_uops_1_lrs2 = iss_uops_1_lrs2;
  assign iregister_read_io_iss_uops_1_lrs3 = iss_uops_1_lrs3;
  assign iregister_read_io_iss_uops_1_ldst_val = iss_uops_1_ldst_val;
  assign iregister_read_io_iss_uops_1_dst_rtype = iss_uops_1_dst_rtype;
  assign iregister_read_io_iss_uops_1_lrs1_rtype = iss_uops_1_lrs1_rtype;
  assign iregister_read_io_iss_uops_1_lrs2_rtype = iss_uops_1_lrs2_rtype;
  assign iregister_read_io_iss_uops_1_frs3_en = iss_uops_1_frs3_en;
  assign iregister_read_io_iss_uops_1_fp_val = iss_uops_1_fp_val;
  assign iregister_read_io_iss_uops_1_fp_single = iss_uops_1_fp_single;
  assign iregister_read_io_iss_uops_1_xcpt_pf_if = iss_uops_1_xcpt_pf_if;
  assign iregister_read_io_iss_uops_1_xcpt_ae_if = iss_uops_1_xcpt_ae_if;
  assign iregister_read_io_iss_uops_1_replay_if = iss_uops_1_replay_if;
  assign iregister_read_io_iss_uops_1_xcpt_ma_if = iss_uops_1_xcpt_ma_if;
  assign iregister_read_io_iss_uops_1_debug_wdata = iss_uops_1_debug_wdata;
  assign iregister_read_io_iss_uops_1_debug_events_fetch_seq = iss_uops_1_debug_events_fetch_seq;
  assign iregister_read_io_iss_uops_2_valid = iss_uops_2_valid;
  assign iregister_read_io_iss_uops_2_iw_state = iss_uops_2_iw_state;
  assign iregister_read_io_iss_uops_2_uopc = iss_uops_2_uopc;
  assign iregister_read_io_iss_uops_2_inst = iss_uops_2_inst;
  assign iregister_read_io_iss_uops_2_pc = iss_uops_2_pc;
  assign iregister_read_io_iss_uops_2_iqtype = iss_uops_2_iqtype;
  assign iregister_read_io_iss_uops_2_fu_code = iss_uops_2_fu_code;
  assign iregister_read_io_iss_uops_2_allocate_brtag = iss_uops_2_allocate_brtag;
  assign iregister_read_io_iss_uops_2_is_br_or_jmp = iss_uops_2_is_br_or_jmp;
  assign iregister_read_io_iss_uops_2_is_jump = iss_uops_2_is_jump;
  assign iregister_read_io_iss_uops_2_is_jal = iss_uops_2_is_jal;
  assign iregister_read_io_iss_uops_2_is_ret = iss_uops_2_is_ret;
  assign iregister_read_io_iss_uops_2_is_call = iss_uops_2_is_call;
  assign iregister_read_io_iss_uops_2_br_mask = iss_uops_2_br_mask;
  assign iregister_read_io_iss_uops_2_br_tag = iss_uops_2_br_tag;
  assign iregister_read_io_iss_uops_2_br_prediction_btb_blame = iss_uops_2_br_prediction_btb_blame;
  assign iregister_read_io_iss_uops_2_br_prediction_btb_hit = iss_uops_2_br_prediction_btb_hit;
  assign iregister_read_io_iss_uops_2_br_prediction_btb_taken = iss_uops_2_br_prediction_btb_taken;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_blame = iss_uops_2_br_prediction_bpd_blame;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_hit = iss_uops_2_br_prediction_bpd_hit;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_taken = iss_uops_2_br_prediction_bpd_taken;
  assign iregister_read_io_iss_uops_2_br_prediction_bim_resp_value = iss_uops_2_br_prediction_bim_resp_value;
  assign iregister_read_io_iss_uops_2_br_prediction_bim_resp_entry_idx = iss_uops_2_br_prediction_bim_resp_entry_idx;
  assign iregister_read_io_iss_uops_2_br_prediction_bim_resp_way_idx = iss_uops_2_br_prediction_bim_resp_way_idx;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_resp_takens = iss_uops_2_br_prediction_bpd_resp_takens;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history = iss_uops_2_br_prediction_bpd_resp_history;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_u = iss_uops_2_br_prediction_bpd_resp_history_u;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_resp_history_ptr = iss_uops_2_br_prediction_bpd_resp_history_ptr;
  assign iregister_read_io_iss_uops_2_br_prediction_bpd_resp_info = iss_uops_2_br_prediction_bpd_resp_info;
  assign iregister_read_io_iss_uops_2_stat_brjmp_mispredicted = iss_uops_2_stat_brjmp_mispredicted;
  assign iregister_read_io_iss_uops_2_stat_btb_made_pred = iss_uops_2_stat_btb_made_pred;
  assign iregister_read_io_iss_uops_2_stat_btb_mispredicted = iss_uops_2_stat_btb_mispredicted;
  assign iregister_read_io_iss_uops_2_stat_bpd_made_pred = iss_uops_2_stat_bpd_made_pred;
  assign iregister_read_io_iss_uops_2_stat_bpd_mispredicted = iss_uops_2_stat_bpd_mispredicted;
  assign iregister_read_io_iss_uops_2_fetch_pc_lob = iss_uops_2_fetch_pc_lob;
  assign iregister_read_io_iss_uops_2_imm_packed = iss_uops_2_imm_packed;
  assign iregister_read_io_iss_uops_2_csr_addr = iss_uops_2_csr_addr;
  assign iregister_read_io_iss_uops_2_rob_idx = iss_uops_2_rob_idx;
  assign iregister_read_io_iss_uops_2_ldq_idx = iss_uops_2_ldq_idx;
  assign iregister_read_io_iss_uops_2_stq_idx = iss_uops_2_stq_idx;
  assign iregister_read_io_iss_uops_2_brob_idx = iss_uops_2_brob_idx;
  assign iregister_read_io_iss_uops_2_pdst = iss_uops_2_pdst;
  assign iregister_read_io_iss_uops_2_pop1 = iss_uops_2_pop1;
  assign iregister_read_io_iss_uops_2_pop2 = iss_uops_2_pop2;
  assign iregister_read_io_iss_uops_2_pop3 = iss_uops_2_pop3;
  assign iregister_read_io_iss_uops_2_prs1_busy = iss_uops_2_prs1_busy;
  assign iregister_read_io_iss_uops_2_prs2_busy = iss_uops_2_prs2_busy;
  assign iregister_read_io_iss_uops_2_prs3_busy = iss_uops_2_prs3_busy;
  assign iregister_read_io_iss_uops_2_stale_pdst = iss_uops_2_stale_pdst;
  assign iregister_read_io_iss_uops_2_exception = iss_uops_2_exception;
  assign iregister_read_io_iss_uops_2_exc_cause = iss_uops_2_exc_cause;
  assign iregister_read_io_iss_uops_2_bypassable = iss_uops_2_bypassable;
  assign iregister_read_io_iss_uops_2_mem_cmd = iss_uops_2_mem_cmd;
  assign iregister_read_io_iss_uops_2_mem_typ = iss_uops_2_mem_typ;
  assign iregister_read_io_iss_uops_2_is_fence = iss_uops_2_is_fence;
  assign iregister_read_io_iss_uops_2_is_fencei = iss_uops_2_is_fencei;
  assign iregister_read_io_iss_uops_2_is_store = iss_uops_2_is_store;
  assign iregister_read_io_iss_uops_2_is_amo = iss_uops_2_is_amo;
  assign iregister_read_io_iss_uops_2_is_load = iss_uops_2_is_load;
  assign iregister_read_io_iss_uops_2_is_sys_pc2epc = iss_uops_2_is_sys_pc2epc;
  assign iregister_read_io_iss_uops_2_is_unique = iss_uops_2_is_unique;
  assign iregister_read_io_iss_uops_2_flush_on_commit = iss_uops_2_flush_on_commit;
  assign iregister_read_io_iss_uops_2_ldst = iss_uops_2_ldst;
  assign iregister_read_io_iss_uops_2_lrs1 = iss_uops_2_lrs1;
  assign iregister_read_io_iss_uops_2_lrs2 = iss_uops_2_lrs2;
  assign iregister_read_io_iss_uops_2_lrs3 = iss_uops_2_lrs3;
  assign iregister_read_io_iss_uops_2_ldst_val = iss_uops_2_ldst_val;
  assign iregister_read_io_iss_uops_2_dst_rtype = iss_uops_2_dst_rtype;
  assign iregister_read_io_iss_uops_2_lrs1_rtype = iss_uops_2_lrs1_rtype;
  assign iregister_read_io_iss_uops_2_lrs2_rtype = iss_uops_2_lrs2_rtype;
  assign iregister_read_io_iss_uops_2_frs3_en = iss_uops_2_frs3_en;
  assign iregister_read_io_iss_uops_2_fp_val = iss_uops_2_fp_val;
  assign iregister_read_io_iss_uops_2_fp_single = iss_uops_2_fp_single;
  assign iregister_read_io_iss_uops_2_xcpt_pf_if = iss_uops_2_xcpt_pf_if;
  assign iregister_read_io_iss_uops_2_xcpt_ae_if = iss_uops_2_xcpt_ae_if;
  assign iregister_read_io_iss_uops_2_replay_if = iss_uops_2_replay_if;
  assign iregister_read_io_iss_uops_2_xcpt_ma_if = iss_uops_2_xcpt_ma_if;
  assign iregister_read_io_iss_uops_2_debug_wdata = iss_uops_2_debug_wdata;
  assign iregister_read_io_iss_uops_2_debug_events_fetch_seq = iss_uops_2_debug_events_fetch_seq;
  assign iregister_read_io_rf_read_ports_0_data = iregfile_io_read_ports_0_data;
  assign iregister_read_io_rf_read_ports_1_data = iregfile_io_read_ports_1_data;
  assign iregister_read_io_rf_read_ports_2_data = iregfile_io_read_ports_2_data;
  assign iregister_read_io_rf_read_ports_3_data = iregfile_io_read_ports_3_data;
  assign iregister_read_io_rf_read_ports_4_data = iregfile_io_read_ports_4_data;
  assign iregister_read_io_rf_read_ports_5_data = iregfile_io_read_ports_5_data;
  assign iregister_read_io_bypass_valid_0 = bypasses_valid_0;
  assign iregister_read_io_bypass_valid_1 = bypasses_valid_1;
  assign iregister_read_io_bypass_valid_2 = bypasses_valid_2;
  assign iregister_read_io_bypass_valid_3 = bypasses_valid_3;
  assign iregister_read_io_bypass_uop_0_ctrl_rf_wen = bypasses_uop_0_ctrl_rf_wen;
  assign iregister_read_io_bypass_uop_0_pdst = bypasses_uop_0_pdst;
  assign iregister_read_io_bypass_uop_0_dst_rtype = bypasses_uop_0_dst_rtype;
  assign iregister_read_io_bypass_uop_1_ctrl_rf_wen = bypasses_uop_1_ctrl_rf_wen;
  assign iregister_read_io_bypass_uop_1_pdst = bypasses_uop_1_pdst;
  assign iregister_read_io_bypass_uop_1_dst_rtype = bypasses_uop_1_dst_rtype;
  assign iregister_read_io_bypass_uop_2_ctrl_rf_wen = bypasses_uop_2_ctrl_rf_wen;
  assign iregister_read_io_bypass_uop_2_pdst = bypasses_uop_2_pdst;
  assign iregister_read_io_bypass_uop_2_dst_rtype = bypasses_uop_2_dst_rtype;
  assign iregister_read_io_bypass_uop_3_ctrl_rf_wen = bypasses_uop_3_ctrl_rf_wen;
  assign iregister_read_io_bypass_uop_3_pdst = bypasses_uop_3_pdst;
  assign iregister_read_io_bypass_uop_3_dst_rtype = bypasses_uop_3_dst_rtype;
  assign iregister_read_io_bypass_data_0 = bypasses_data_0;
  assign iregister_read_io_bypass_data_1 = bypasses_data_1;
  assign iregister_read_io_bypass_data_2 = bypasses_data_2;
  assign iregister_read_io_bypass_data_3 = bypasses_data_3;
  assign iregister_read_io_kill = rob_io_flush_valid;
  assign iregister_read_io_brinfo_valid = br_unit_brinfo_valid;
  assign iregister_read_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign iregister_read_io_brinfo_mask = br_unit_brinfo_mask;
  assign iregister_read_clock = clock;
  assign iregister_read_reset = reset;
  assign dc_shim_io_core_req_valid = mem_unit_io_dmem_req_valid;
  assign dc_shim_io_core_req_bits_addr = mem_unit_io_dmem_req_bits_addr;
  assign dc_shim_io_core_req_bits_uop_uopc = mem_unit_io_dmem_req_bits_uop_uopc;
  assign dc_shim_io_core_req_bits_uop_br_mask = mem_unit_io_dmem_req_bits_uop_br_mask;
  assign dc_shim_io_core_req_bits_uop_rob_idx = mem_unit_io_dmem_req_bits_uop_rob_idx;
  assign dc_shim_io_core_req_bits_uop_ldq_idx = mem_unit_io_dmem_req_bits_uop_ldq_idx;
  assign dc_shim_io_core_req_bits_uop_stq_idx = mem_unit_io_dmem_req_bits_uop_stq_idx;
  assign dc_shim_io_core_req_bits_uop_pdst = mem_unit_io_dmem_req_bits_uop_pdst;
  assign dc_shim_io_core_req_bits_uop_mem_cmd = mem_unit_io_dmem_req_bits_uop_mem_cmd;
  assign dc_shim_io_core_req_bits_uop_mem_typ = mem_unit_io_dmem_req_bits_uop_mem_typ;
  assign dc_shim_io_core_req_bits_uop_is_store = mem_unit_io_dmem_req_bits_uop_is_store;
  assign dc_shim_io_core_req_bits_uop_is_amo = mem_unit_io_dmem_req_bits_uop_is_amo;
  assign dc_shim_io_core_req_bits_uop_is_load = mem_unit_io_dmem_req_bits_uop_is_load;
  assign dc_shim_io_core_req_bits_uop_dst_rtype = mem_unit_io_dmem_req_bits_uop_dst_rtype;
  assign dc_shim_io_core_req_bits_uop_fp_val = mem_unit_io_dmem_req_bits_uop_fp_val;
  assign dc_shim_io_core_req_bits_data = mem_unit_io_dmem_req_bits_data;
  assign dc_shim_io_core_req_bits_kill = mem_unit_io_dmem_req_bits_kill;
  assign dc_shim_io_core_brinfo_valid = br_unit_brinfo_valid;
  assign dc_shim_io_core_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign dc_shim_io_core_brinfo_mask = br_unit_brinfo_mask;
  assign dc_shim_io_core_flush_pipe = rob_io_flush_valid;
  assign dc_shim_io_core_invalidate_lr = rob_io_com_xcpt_valid;
  assign dc_shim_io_dmem_req_ready = io_dmem_req_ready;
  assign dc_shim_io_dmem_s2_nack = io_dmem_s2_nack;
  assign dc_shim_io_dmem_resp_valid = io_dmem_resp_valid;
  assign dc_shim_io_dmem_resp_bits_tag = io_dmem_resp_bits_tag;
  assign dc_shim_io_dmem_resp_bits_data = io_dmem_resp_bits_data;
  assign dc_shim_io_dmem_resp_bits_has_data = io_dmem_resp_bits_has_data;
  assign dc_shim_io_dmem_s2_xcpt_ma_ld = io_dmem_s2_xcpt_ma_ld;
  assign dc_shim_io_dmem_s2_xcpt_ma_st = io_dmem_s2_xcpt_ma_st;
  assign dc_shim_io_dmem_s2_xcpt_pf_ld = io_dmem_s2_xcpt_pf_ld;
  assign dc_shim_io_dmem_s2_xcpt_pf_st = io_dmem_s2_xcpt_pf_st;
  assign dc_shim_io_dmem_ordered = io_dmem_ordered;
  assign dc_shim_clock = clock;
  assign dc_shim_reset = reset;
  assign lsu_io_dec_st_vals_0 = _T_3046;
  assign lsu_io_dec_st_vals_1 = _T_3056;
  assign lsu_io_dec_ld_vals_0 = _T_3051;
  assign lsu_io_dec_ld_vals_1 = _T_3061;
  assign lsu_io_dec_uops_0_uopc = dec_uops_0_uopc;
  assign lsu_io_dec_uops_0_br_mask = dec_uops_0_br_mask;
  assign lsu_io_dec_uops_0_rob_idx = dec_uops_0_rob_idx;
  assign lsu_io_dec_uops_0_ldq_idx = dec_uops_0_ldq_idx;
  assign lsu_io_dec_uops_0_stq_idx = dec_uops_0_stq_idx;
  assign lsu_io_dec_uops_0_mem_cmd = dec_uops_0_mem_cmd;
  assign lsu_io_dec_uops_0_mem_typ = dec_uops_0_mem_typ;
  assign lsu_io_dec_uops_0_is_fence = dec_uops_0_is_fence;
  assign lsu_io_dec_uops_0_is_store = dec_uops_0_is_store;
  assign lsu_io_dec_uops_0_is_amo = dec_uops_0_is_amo;
  assign lsu_io_dec_uops_0_is_load = dec_uops_0_is_load;
  assign lsu_io_dec_uops_0_dst_rtype = dec_uops_0_dst_rtype;
  assign lsu_io_dec_uops_0_fp_val = dec_uops_0_fp_val;
  assign lsu_io_dec_uops_1_uopc = dec_uops_1_uopc;
  assign lsu_io_dec_uops_1_br_mask = dec_uops_1_br_mask;
  assign lsu_io_dec_uops_1_rob_idx = dec_uops_1_rob_idx;
  assign lsu_io_dec_uops_1_ldq_idx = dec_uops_1_ldq_idx;
  assign lsu_io_dec_uops_1_stq_idx = dec_uops_1_stq_idx;
  assign lsu_io_dec_uops_1_mem_cmd = dec_uops_1_mem_cmd;
  assign lsu_io_dec_uops_1_mem_typ = dec_uops_1_mem_typ;
  assign lsu_io_dec_uops_1_is_fence = dec_uops_1_is_fence;
  assign lsu_io_dec_uops_1_is_store = dec_uops_1_is_store;
  assign lsu_io_dec_uops_1_is_amo = dec_uops_1_is_amo;
  assign lsu_io_dec_uops_1_is_load = dec_uops_1_is_load;
  assign lsu_io_dec_uops_1_dst_rtype = dec_uops_1_dst_rtype;
  assign lsu_io_dec_uops_1_fp_val = dec_uops_1_fp_val;
  assign lsu_io_exe_resp_valid = mem_unit_io_lsu_io_exe_resp_valid;
  assign lsu_io_exe_resp_bits_uop_uopc = mem_unit_io_lsu_io_exe_resp_bits_uop_uopc;
  assign lsu_io_exe_resp_bits_uop_ctrl_is_load = mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_load;
  assign lsu_io_exe_resp_bits_uop_ctrl_is_sta = mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_sta;
  assign lsu_io_exe_resp_bits_uop_ctrl_is_std = mem_unit_io_lsu_io_exe_resp_bits_uop_ctrl_is_std;
  assign lsu_io_exe_resp_bits_uop_br_mask = mem_unit_io_lsu_io_exe_resp_bits_uop_br_mask;
  assign lsu_io_exe_resp_bits_uop_rob_idx = mem_unit_io_lsu_io_exe_resp_bits_uop_rob_idx;
  assign lsu_io_exe_resp_bits_uop_ldq_idx = mem_unit_io_lsu_io_exe_resp_bits_uop_ldq_idx;
  assign lsu_io_exe_resp_bits_uop_stq_idx = mem_unit_io_lsu_io_exe_resp_bits_uop_stq_idx;
  assign lsu_io_exe_resp_bits_uop_pdst = mem_unit_io_lsu_io_exe_resp_bits_uop_pdst;
  assign lsu_io_exe_resp_bits_uop_mem_cmd = mem_unit_io_lsu_io_exe_resp_bits_uop_mem_cmd;
  assign lsu_io_exe_resp_bits_uop_mem_typ = mem_unit_io_lsu_io_exe_resp_bits_uop_mem_typ;
  assign lsu_io_exe_resp_bits_uop_is_fence = mem_unit_io_lsu_io_exe_resp_bits_uop_is_fence;
  assign lsu_io_exe_resp_bits_uop_is_store = mem_unit_io_lsu_io_exe_resp_bits_uop_is_store;
  assign lsu_io_exe_resp_bits_uop_is_amo = mem_unit_io_lsu_io_exe_resp_bits_uop_is_amo;
  assign lsu_io_exe_resp_bits_uop_is_load = mem_unit_io_lsu_io_exe_resp_bits_uop_is_load;
  assign lsu_io_exe_resp_bits_uop_dst_rtype = mem_unit_io_lsu_io_exe_resp_bits_uop_dst_rtype;
  assign lsu_io_exe_resp_bits_uop_fp_val = mem_unit_io_lsu_io_exe_resp_bits_uop_fp_val;
  assign lsu_io_exe_resp_bits_data = mem_unit_io_lsu_io_exe_resp_bits_data;
  assign lsu_io_exe_resp_bits_addr = mem_unit_io_lsu_io_exe_resp_bits_addr;
  assign lsu_io_exe_resp_bits_mxcpt_valid = mem_unit_io_lsu_io_exe_resp_bits_mxcpt_valid;
  assign lsu_io_exe_resp_bits_mxcpt_bits = mem_unit_io_lsu_io_exe_resp_bits_mxcpt_bits;
  assign lsu_io_exe_resp_bits_sfence_valid = mem_unit_io_lsu_io_exe_resp_bits_sfence_valid;
  assign lsu_io_exe_resp_bits_sfence_bits_rs1 = mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs1;
  assign lsu_io_exe_resp_bits_sfence_bits_rs2 = mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_rs2;
  assign lsu_io_exe_resp_bits_sfence_bits_addr = mem_unit_io_lsu_io_exe_resp_bits_sfence_bits_addr;
  assign lsu_io_fp_stdata_valid = fp_pipeline_io_tosdq_valid;
  assign lsu_io_fp_stdata_bits_uop_br_mask = fp_pipeline_io_tosdq_bits_uop_br_mask;
  assign lsu_io_fp_stdata_bits_uop_rob_idx = fp_pipeline_io_tosdq_bits_uop_rob_idx;
  assign lsu_io_fp_stdata_bits_uop_stq_idx = fp_pipeline_io_tosdq_bits_uop_stq_idx;
  assign lsu_io_fp_stdata_bits_uop_is_amo = fp_pipeline_io_tosdq_bits_uop_is_amo;
  assign lsu_io_fp_stdata_bits_data = fp_pipeline_io_tosdq_bits_data;
  assign lsu_io_commit_store_mask_0 = rob_io_commit_st_mask_0;
  assign lsu_io_commit_store_mask_1 = rob_io_commit_st_mask_1;
  assign lsu_io_commit_load_mask_0 = rob_io_commit_ld_mask_0;
  assign lsu_io_commit_load_mask_1 = rob_io_commit_ld_mask_1;
  assign lsu_io_commit_load_at_rob_head = rob_io_com_load_is_at_rob_head;
  assign lsu_io_memresp_valid = mem_unit_io_lsu_io_memresp_valid;
  assign lsu_io_memresp_bits_ldq_idx = mem_unit_io_lsu_io_memresp_bits_ldq_idx;
  assign lsu_io_memresp_bits_stq_idx = mem_unit_io_lsu_io_memresp_bits_stq_idx;
  assign lsu_io_memresp_bits_is_load = mem_unit_io_lsu_io_memresp_bits_is_load;
  assign lsu_io_brinfo_valid = br_unit_brinfo_valid;
  assign lsu_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign lsu_io_brinfo_mask = br_unit_brinfo_mask;
  assign lsu_io_brinfo_ldq_idx = br_unit_brinfo_ldq_idx;
  assign lsu_io_brinfo_stq_idx = br_unit_brinfo_stq_idx;
  assign lsu_io_exception = rob_io_flush_valid;
  assign lsu_io_nack_valid = dc_shim_io_core_nack_valid;
  assign lsu_io_nack_lsu_idx = dc_shim_io_core_nack_lsu_idx;
  assign lsu_io_nack_isload = dc_shim_io_core_nack_isload;
  assign lsu_io_nack_cache_nack = dc_shim_io_core_nack_cache_nack;
  assign lsu_io_dmem_is_ordered = dc_shim_io_core_ordered;
  assign lsu_io_ptw_req_ready = io_ptw_tlb_req_ready;
  assign lsu_io_ptw_resp_valid = io_ptw_tlb_resp_valid;
  assign lsu_io_ptw_resp_bits_ae = io_ptw_tlb_resp_bits_ae;
  assign lsu_io_ptw_resp_bits_pte_ppn = io_ptw_tlb_resp_bits_pte_ppn;
  assign lsu_io_ptw_resp_bits_pte_d = io_ptw_tlb_resp_bits_pte_d;
  assign lsu_io_ptw_resp_bits_pte_a = io_ptw_tlb_resp_bits_pte_a;
  assign lsu_io_ptw_resp_bits_pte_g = io_ptw_tlb_resp_bits_pte_g;
  assign lsu_io_ptw_resp_bits_pte_u = io_ptw_tlb_resp_bits_pte_u;
  assign lsu_io_ptw_resp_bits_pte_x = io_ptw_tlb_resp_bits_pte_x;
  assign lsu_io_ptw_resp_bits_pte_w = io_ptw_tlb_resp_bits_pte_w;
  assign lsu_io_ptw_resp_bits_pte_r = io_ptw_tlb_resp_bits_pte_r;
  assign lsu_io_ptw_resp_bits_pte_v = io_ptw_tlb_resp_bits_pte_v;
  assign lsu_io_ptw_resp_bits_level = io_ptw_tlb_resp_bits_level;
  assign lsu_io_ptw_resp_bits_homogeneous = io_ptw_tlb_resp_bits_homogeneous;
  assign lsu_io_ptw_ptbr_mode = io_ptw_tlb_ptbr_mode;
  assign lsu_io_ptw_status_dprv = io_ptw_tlb_status_dprv;
  assign lsu_io_ptw_status_mxr = io_ptw_tlb_status_mxr;
  assign lsu_io_ptw_status_sum = io_ptw_tlb_status_sum;
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign rob_io_enq_valids_0 = rename_stage_io_ren1_mask_0;
  assign rob_io_enq_valids_1 = rename_stage_io_ren1_mask_1;
  assign rob_io_enq_uops_0_pc = rename_stage_io_ren1_uops_0_pc;
  assign rob_io_enq_uops_0_br_mask = rename_stage_io_ren1_uops_0_br_mask;
  assign rob_io_enq_uops_0_rob_idx = rename_stage_io_ren1_uops_0_rob_idx;
  assign rob_io_enq_uops_0_brob_idx = rename_stage_io_ren1_uops_0_brob_idx;
  assign rob_io_enq_uops_0_pdst = rename_stage_io_ren1_uops_0_pdst;
  assign rob_io_enq_uops_0_stale_pdst = rename_stage_io_ren1_uops_0_stale_pdst;
  assign rob_io_enq_uops_0_exception = rename_stage_io_ren1_uops_0_exception;
  assign rob_io_enq_uops_0_exc_cause = rename_stage_io_ren1_uops_0_exc_cause;
  assign rob_io_enq_uops_0_is_fence = rename_stage_io_ren1_uops_0_is_fence;
  assign rob_io_enq_uops_0_is_fencei = rename_stage_io_ren1_uops_0_is_fencei;
  assign rob_io_enq_uops_0_is_store = rename_stage_io_ren1_uops_0_is_store;
  assign rob_io_enq_uops_0_is_load = rename_stage_io_ren1_uops_0_is_load;
  assign rob_io_enq_uops_0_is_sys_pc2epc = rename_stage_io_ren1_uops_0_is_sys_pc2epc;
  assign rob_io_enq_uops_0_is_unique = rename_stage_io_ren1_uops_0_is_unique;
  assign rob_io_enq_uops_0_flush_on_commit = rename_stage_io_ren1_uops_0_flush_on_commit;
  assign rob_io_enq_uops_0_ldst = rename_stage_io_ren1_uops_0_ldst;
  assign rob_io_enq_uops_0_ldst_val = rename_stage_io_ren1_uops_0_ldst_val;
  assign rob_io_enq_uops_0_dst_rtype = rename_stage_io_ren1_uops_0_dst_rtype;
  assign rob_io_enq_uops_0_fp_val = rename_stage_io_ren1_uops_0_fp_val;
  assign rob_io_enq_uops_1_br_mask = rename_stage_io_ren1_uops_1_br_mask;
  assign rob_io_enq_uops_1_rob_idx = rename_stage_io_ren1_uops_1_rob_idx;
  assign rob_io_enq_uops_1_pdst = rename_stage_io_ren1_uops_1_pdst;
  assign rob_io_enq_uops_1_stale_pdst = rename_stage_io_ren1_uops_1_stale_pdst;
  assign rob_io_enq_uops_1_exception = rename_stage_io_ren1_uops_1_exception;
  assign rob_io_enq_uops_1_exc_cause = rename_stage_io_ren1_uops_1_exc_cause;
  assign rob_io_enq_uops_1_is_fence = rename_stage_io_ren1_uops_1_is_fence;
  assign rob_io_enq_uops_1_is_fencei = rename_stage_io_ren1_uops_1_is_fencei;
  assign rob_io_enq_uops_1_is_store = rename_stage_io_ren1_uops_1_is_store;
  assign rob_io_enq_uops_1_is_load = rename_stage_io_ren1_uops_1_is_load;
  assign rob_io_enq_uops_1_is_sys_pc2epc = rename_stage_io_ren1_uops_1_is_sys_pc2epc;
  assign rob_io_enq_uops_1_is_unique = rename_stage_io_ren1_uops_1_is_unique;
  assign rob_io_enq_uops_1_flush_on_commit = rename_stage_io_ren1_uops_1_flush_on_commit;
  assign rob_io_enq_uops_1_ldst = rename_stage_io_ren1_uops_1_ldst;
  assign rob_io_enq_uops_1_ldst_val = rename_stage_io_ren1_uops_1_ldst_val;
  assign rob_io_enq_uops_1_dst_rtype = rename_stage_io_ren1_uops_1_dst_rtype;
  assign rob_io_enq_uops_1_fp_val = rename_stage_io_ren1_uops_1_fp_val;
  assign rob_io_enq_has_br_or_jalr_in_packet = dec_has_br_or_jalr_in_packet;
  assign rob_io_enq_partial_stall = _T_3185;
  assign rob_io_enq_new_packet = _T_2872;
  assign rob_io_brinfo_valid = br_unit_brinfo_valid;
  assign rob_io_brinfo_mispredict = br_unit_brinfo_mispredict;
  assign rob_io_brinfo_mask = br_unit_brinfo_mask;
  assign rob_io_brinfo_rob_idx = br_unit_brinfo_rob_idx;
  assign rob_io_get_pc_rob_idx = _T_3505;
  assign rob_io_wb_resps_0_valid = _T_3200;
  assign rob_io_wb_resps_0_bits_uop_rob_idx = ll_wbarb_io_out_bits_uop_rob_idx;
  assign rob_io_wb_resps_0_bits_uop_pdst = ll_wbarb_io_out_bits_uop_pdst;
  assign rob_io_wb_resps_1_valid = _T_3220;
  assign rob_io_wb_resps_1_bits_uop_rob_idx = csr_exe_unit_io_resp_0_bits_uop_rob_idx;
  assign rob_io_wb_resps_1_bits_uop_pdst = csr_exe_unit_io_resp_0_bits_uop_pdst;
  assign rob_io_wb_resps_2_valid = _T_3232;
  assign rob_io_wb_resps_2_bits_uop_rob_idx = ALUExeUnit_io_resp_0_bits_uop_rob_idx;
  assign rob_io_wb_resps_2_bits_uop_pdst = ALUExeUnit_io_resp_0_bits_uop_pdst;
  assign rob_io_wb_resps_3_valid = fp_pipeline_io_wakeups_0_valid;
  assign rob_io_wb_resps_3_bits_uop_rob_idx = fp_pipeline_io_wakeups_0_bits_uop_rob_idx;
  assign rob_io_wb_resps_3_bits_uop_pdst = fp_pipeline_io_wakeups_0_bits_uop_pdst;
  assign rob_io_wb_resps_4_valid = fp_pipeline_io_wakeups_1_valid;
  assign rob_io_wb_resps_4_bits_uop_rob_idx = fp_pipeline_io_wakeups_1_bits_uop_rob_idx;
  assign rob_io_wb_resps_4_bits_uop_pdst = fp_pipeline_io_wakeups_1_bits_uop_pdst;
  assign rob_io_lsu_clr_bsy_valid_0 = lsu_io_lsu_clr_bsy_valid_0;
  assign rob_io_lsu_clr_bsy_valid_1 = lsu_io_lsu_clr_bsy_valid_1;
  assign rob_io_lsu_clr_bsy_rob_idx_0 = lsu_io_lsu_clr_bsy_rob_idx_0;
  assign rob_io_lsu_clr_bsy_rob_idx_1 = lsu_io_lsu_clr_bsy_rob_idx_1;
  assign rob_io_fflags_0_valid = fp_pipeline_io_wakeups_0_bits_fflags_valid;
  assign rob_io_fflags_0_bits_uop_rob_idx = fp_pipeline_io_wakeups_0_bits_fflags_bits_uop_rob_idx;
  assign rob_io_fflags_0_bits_flags = fp_pipeline_io_wakeups_0_bits_fflags_bits_flags;
  assign rob_io_fflags_1_valid = fp_pipeline_io_wakeups_1_bits_fflags_valid;
  assign rob_io_fflags_1_bits_uop_rob_idx = fp_pipeline_io_wakeups_1_bits_fflags_bits_uop_rob_idx;
  assign rob_io_fflags_1_bits_flags = fp_pipeline_io_wakeups_1_bits_fflags_bits_flags;
  assign rob_io_lxcpt_valid = lsu_io_xcpt_valid;
  assign rob_io_lxcpt_bits_uop_br_mask = lsu_io_xcpt_bits_uop_br_mask;
  assign rob_io_lxcpt_bits_uop_rob_idx = lsu_io_xcpt_bits_uop_rob_idx;
  assign rob_io_lxcpt_bits_cause = lsu_io_xcpt_bits_cause;
  assign rob_io_lxcpt_bits_badvaddr = lsu_io_xcpt_bits_badvaddr;
  assign rob_io_bxcpt_valid = br_unit_xcpt_valid;
  assign rob_io_bxcpt_bits_uop_br_mask = br_unit_xcpt_bits_uop_br_mask;
  assign rob_io_bxcpt_bits_uop_rob_idx = br_unit_xcpt_bits_uop_rob_idx;
  assign rob_io_bxcpt_bits_badvaddr = br_unit_xcpt_bits_badvaddr;
  assign rob_io_csr_eret = csr_io_eret;
  assign rob_io_csr_evec = csr_io_evec;
  assign rob_io_csr_stall = csr_io_csr_stall;
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign int_wakeups_0_valid = _T_2932;
  assign int_wakeups_0_bits_uop_pdst = ll_wbarb_io_out_bits_uop_pdst;
  assign int_wakeups_0_bits_uop_dst_rtype = ll_wbarb_io_out_bits_uop_dst_rtype;
  assign int_wakeups_1_valid = _T_2936;
  assign int_wakeups_1_bits_uop_pdst = iss_uops_1_pdst;
  assign int_wakeups_1_bits_uop_dst_rtype = iss_uops_1_dst_rtype;
  assign int_wakeups_2_valid = _T_2950;
  assign int_wakeups_2_bits_uop_pdst = csr_exe_unit_io_resp_0_bits_uop_pdst;
  assign int_wakeups_2_bits_uop_dst_rtype = csr_exe_unit_io_resp_0_bits_uop_dst_rtype;
  assign int_wakeups_3_valid = _T_2954;
  assign int_wakeups_3_bits_uop_pdst = iss_uops_2_pdst;
  assign int_wakeups_3_bits_uop_dst_rtype = iss_uops_2_dst_rtype;
  assign int_wakeups_4_valid = _T_2968;
  assign int_wakeups_4_bits_uop_pdst = ALUExeUnit_io_resp_0_bits_uop_pdst;
  assign int_wakeups_4_bits_uop_dst_rtype = ALUExeUnit_io_resp_0_bits_uop_dst_rtype;
  assign dec_valids_0 = _T_2735;
  assign dec_valids_1 = _T_2779;
  assign dec_uops_0_valid = decode_units_0_io_deq_uop_valid;
  assign dec_uops_0_uopc = decode_units_0_io_deq_uop_uopc;
  assign dec_uops_0_inst = decode_units_0_io_deq_uop_inst;
  assign dec_uops_0_pc = decode_units_0_io_deq_uop_pc;
  assign dec_uops_0_iqtype = decode_units_0_io_deq_uop_iqtype;
  assign dec_uops_0_fu_code = decode_units_0_io_deq_uop_fu_code;
  assign dec_uops_0_allocate_brtag = decode_units_0_io_deq_uop_allocate_brtag;
  assign dec_uops_0_is_br_or_jmp = decode_units_0_io_deq_uop_is_br_or_jmp;
  assign dec_uops_0_is_jump = decode_units_0_io_deq_uop_is_jump;
  assign dec_uops_0_is_jal = decode_units_0_io_deq_uop_is_jal;
  assign dec_uops_0_is_ret = decode_units_0_io_deq_uop_is_ret;
  assign dec_uops_0_is_call = decode_units_0_io_deq_uop_is_call;
  assign dec_uops_0_br_mask = dec_brmask_logic_io_br_mask_0;
  assign dec_uops_0_br_tag = dec_brmask_logic_io_br_tag_0;
  assign dec_uops_0_br_prediction_btb_blame = decode_units_0_io_deq_uop_br_prediction_btb_blame;
  assign dec_uops_0_br_prediction_btb_hit = decode_units_0_io_deq_uop_br_prediction_btb_hit;
  assign dec_uops_0_br_prediction_btb_taken = decode_units_0_io_deq_uop_br_prediction_btb_taken;
  assign dec_uops_0_br_prediction_bpd_blame = decode_units_0_io_deq_uop_br_prediction_bpd_blame;
  assign dec_uops_0_br_prediction_bpd_hit = decode_units_0_io_deq_uop_br_prediction_bpd_hit;
  assign dec_uops_0_br_prediction_bpd_taken = decode_units_0_io_deq_uop_br_prediction_bpd_taken;
  assign dec_uops_0_br_prediction_bim_resp_value = decode_units_0_io_deq_uop_br_prediction_bim_resp_value;
  assign dec_uops_0_br_prediction_bim_resp_entry_idx = decode_units_0_io_deq_uop_br_prediction_bim_resp_entry_idx;
  assign dec_uops_0_br_prediction_bim_resp_way_idx = decode_units_0_io_deq_uop_br_prediction_bim_resp_way_idx;
  assign dec_uops_0_br_prediction_bpd_resp_takens = decode_units_0_io_deq_uop_br_prediction_bpd_resp_takens;
  assign dec_uops_0_br_prediction_bpd_resp_history = decode_units_0_io_deq_uop_br_prediction_bpd_resp_history;
  assign dec_uops_0_br_prediction_bpd_resp_history_u = decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_u;
  assign dec_uops_0_br_prediction_bpd_resp_history_ptr = decode_units_0_io_deq_uop_br_prediction_bpd_resp_history_ptr;
  assign dec_uops_0_br_prediction_bpd_resp_info = decode_units_0_io_deq_uop_br_prediction_bpd_resp_info;
  assign dec_uops_0_fetch_pc_lob = decode_units_0_io_deq_uop_fetch_pc_lob;
  assign dec_uops_0_imm_packed = decode_units_0_io_deq_uop_imm_packed;
  assign dec_uops_0_rob_idx = _T_2859[6:0];
  assign dec_uops_0_ldq_idx = new_ldq_idx;
  assign dec_uops_0_stq_idx = new_stq_idx;
  assign dec_uops_0_brob_idx = bpd_stage_io_brob_allocate_brob_tail;
  assign dec_uops_0_exception = decode_units_0_io_deq_uop_exception;
  assign dec_uops_0_exc_cause = decode_units_0_io_deq_uop_exc_cause;
  assign dec_uops_0_bypassable = decode_units_0_io_deq_uop_bypassable;
  assign dec_uops_0_mem_cmd = decode_units_0_io_deq_uop_mem_cmd;
  assign dec_uops_0_mem_typ = decode_units_0_io_deq_uop_mem_typ;
  assign dec_uops_0_is_fence = decode_units_0_io_deq_uop_is_fence;
  assign dec_uops_0_is_fencei = decode_units_0_io_deq_uop_is_fencei;
  assign dec_uops_0_is_store = decode_units_0_io_deq_uop_is_store;
  assign dec_uops_0_is_amo = decode_units_0_io_deq_uop_is_amo;
  assign dec_uops_0_is_load = decode_units_0_io_deq_uop_is_load;
  assign dec_uops_0_is_sys_pc2epc = decode_units_0_io_deq_uop_is_sys_pc2epc;
  assign dec_uops_0_is_unique = decode_units_0_io_deq_uop_is_unique;
  assign dec_uops_0_flush_on_commit = decode_units_0_io_deq_uop_flush_on_commit;
  assign dec_uops_0_ldst = decode_units_0_io_deq_uop_ldst;
  assign dec_uops_0_lrs1 = decode_units_0_io_deq_uop_lrs1;
  assign dec_uops_0_lrs2 = decode_units_0_io_deq_uop_lrs2;
  assign dec_uops_0_lrs3 = decode_units_0_io_deq_uop_lrs3;
  assign dec_uops_0_ldst_val = decode_units_0_io_deq_uop_ldst_val;
  assign dec_uops_0_dst_rtype = decode_units_0_io_deq_uop_dst_rtype;
  assign dec_uops_0_lrs1_rtype = decode_units_0_io_deq_uop_lrs1_rtype;
  assign dec_uops_0_lrs2_rtype = decode_units_0_io_deq_uop_lrs2_rtype;
  assign dec_uops_0_frs3_en = decode_units_0_io_deq_uop_frs3_en;
  assign dec_uops_0_fp_val = decode_units_0_io_deq_uop_fp_val;
  assign dec_uops_0_fp_single = decode_units_0_io_deq_uop_fp_single;
  assign dec_uops_0_xcpt_pf_if = decode_units_0_io_deq_uop_xcpt_pf_if;
  assign dec_uops_0_xcpt_ae_if = decode_units_0_io_deq_uop_xcpt_ae_if;
  assign dec_uops_0_replay_if = decode_units_0_io_deq_uop_replay_if;
  assign dec_uops_0_xcpt_ma_if = decode_units_0_io_deq_uop_xcpt_ma_if;
  assign dec_uops_0_debug_events_fetch_seq = decode_units_0_io_deq_uop_debug_events_fetch_seq;
  assign dec_uops_1_valid = decode_units_1_io_deq_uop_valid;
  assign dec_uops_1_uopc = decode_units_1_io_deq_uop_uopc;
  assign dec_uops_1_inst = decode_units_1_io_deq_uop_inst;
  assign dec_uops_1_pc = decode_units_1_io_deq_uop_pc;
  assign dec_uops_1_iqtype = decode_units_1_io_deq_uop_iqtype;
  assign dec_uops_1_fu_code = decode_units_1_io_deq_uop_fu_code;
  assign dec_uops_1_allocate_brtag = decode_units_1_io_deq_uop_allocate_brtag;
  assign dec_uops_1_is_br_or_jmp = decode_units_1_io_deq_uop_is_br_or_jmp;
  assign dec_uops_1_is_jump = decode_units_1_io_deq_uop_is_jump;
  assign dec_uops_1_is_jal = decode_units_1_io_deq_uop_is_jal;
  assign dec_uops_1_is_ret = decode_units_1_io_deq_uop_is_ret;
  assign dec_uops_1_is_call = decode_units_1_io_deq_uop_is_call;
  assign dec_uops_1_br_mask = dec_brmask_logic_io_br_mask_1;
  assign dec_uops_1_br_tag = dec_brmask_logic_io_br_tag_1;
  assign dec_uops_1_br_prediction_btb_blame = decode_units_1_io_deq_uop_br_prediction_btb_blame;
  assign dec_uops_1_br_prediction_btb_hit = decode_units_1_io_deq_uop_br_prediction_btb_hit;
  assign dec_uops_1_br_prediction_btb_taken = decode_units_1_io_deq_uop_br_prediction_btb_taken;
  assign dec_uops_1_br_prediction_bpd_blame = decode_units_1_io_deq_uop_br_prediction_bpd_blame;
  assign dec_uops_1_br_prediction_bpd_hit = decode_units_1_io_deq_uop_br_prediction_bpd_hit;
  assign dec_uops_1_br_prediction_bpd_taken = decode_units_1_io_deq_uop_br_prediction_bpd_taken;
  assign dec_uops_1_br_prediction_bim_resp_value = decode_units_1_io_deq_uop_br_prediction_bim_resp_value;
  assign dec_uops_1_br_prediction_bim_resp_entry_idx = decode_units_1_io_deq_uop_br_prediction_bim_resp_entry_idx;
  assign dec_uops_1_br_prediction_bim_resp_way_idx = decode_units_1_io_deq_uop_br_prediction_bim_resp_way_idx;
  assign dec_uops_1_br_prediction_bpd_resp_takens = decode_units_1_io_deq_uop_br_prediction_bpd_resp_takens;
  assign dec_uops_1_br_prediction_bpd_resp_history = decode_units_1_io_deq_uop_br_prediction_bpd_resp_history;
  assign dec_uops_1_br_prediction_bpd_resp_history_u = decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_u;
  assign dec_uops_1_br_prediction_bpd_resp_history_ptr = decode_units_1_io_deq_uop_br_prediction_bpd_resp_history_ptr;
  assign dec_uops_1_br_prediction_bpd_resp_info = decode_units_1_io_deq_uop_br_prediction_bpd_resp_info;
  assign dec_uops_1_fetch_pc_lob = decode_units_1_io_deq_uop_fetch_pc_lob;
  assign dec_uops_1_imm_packed = decode_units_1_io_deq_uop_imm_packed;
  assign dec_uops_1_rob_idx = _T_2861[6:0];
  assign dec_uops_1_ldq_idx = _T_2841;
  assign dec_uops_1_stq_idx = _T_2847;
  assign dec_uops_1_brob_idx = bpd_stage_io_brob_allocate_brob_tail;
  assign dec_uops_1_exception = decode_units_1_io_deq_uop_exception;
  assign dec_uops_1_exc_cause = decode_units_1_io_deq_uop_exc_cause;
  assign dec_uops_1_bypassable = decode_units_1_io_deq_uop_bypassable;
  assign dec_uops_1_mem_cmd = decode_units_1_io_deq_uop_mem_cmd;
  assign dec_uops_1_mem_typ = decode_units_1_io_deq_uop_mem_typ;
  assign dec_uops_1_is_fence = decode_units_1_io_deq_uop_is_fence;
  assign dec_uops_1_is_fencei = decode_units_1_io_deq_uop_is_fencei;
  assign dec_uops_1_is_store = decode_units_1_io_deq_uop_is_store;
  assign dec_uops_1_is_amo = decode_units_1_io_deq_uop_is_amo;
  assign dec_uops_1_is_load = decode_units_1_io_deq_uop_is_load;
  assign dec_uops_1_is_sys_pc2epc = decode_units_1_io_deq_uop_is_sys_pc2epc;
  assign dec_uops_1_is_unique = decode_units_1_io_deq_uop_is_unique;
  assign dec_uops_1_flush_on_commit = decode_units_1_io_deq_uop_flush_on_commit;
  assign dec_uops_1_ldst = decode_units_1_io_deq_uop_ldst;
  assign dec_uops_1_lrs1 = decode_units_1_io_deq_uop_lrs1;
  assign dec_uops_1_lrs2 = decode_units_1_io_deq_uop_lrs2;
  assign dec_uops_1_lrs3 = decode_units_1_io_deq_uop_lrs3;
  assign dec_uops_1_ldst_val = decode_units_1_io_deq_uop_ldst_val;
  assign dec_uops_1_dst_rtype = decode_units_1_io_deq_uop_dst_rtype;
  assign dec_uops_1_lrs1_rtype = decode_units_1_io_deq_uop_lrs1_rtype;
  assign dec_uops_1_lrs2_rtype = decode_units_1_io_deq_uop_lrs2_rtype;
  assign dec_uops_1_frs3_en = decode_units_1_io_deq_uop_frs3_en;
  assign dec_uops_1_fp_val = decode_units_1_io_deq_uop_fp_val;
  assign dec_uops_1_fp_single = decode_units_1_io_deq_uop_fp_single;
  assign dec_uops_1_xcpt_pf_if = decode_units_1_io_deq_uop_xcpt_pf_if;
  assign dec_uops_1_xcpt_ae_if = decode_units_1_io_deq_uop_xcpt_ae_if;
  assign dec_uops_1_replay_if = decode_units_1_io_deq_uop_replay_if;
  assign dec_uops_1_xcpt_ma_if = decode_units_1_io_deq_uop_xcpt_ma_if;
  assign dec_uops_1_debug_events_fetch_seq = decode_units_1_io_deq_uop_debug_events_fetch_seq;
  assign dec_will_fire_0 = _T_2774;
  assign dec_will_fire_1 = _T_2817;
  assign dec_rdy = _T_2819;
  assign dis_valids_0 = rename_stage_io_ren2_mask_0;
  assign dis_valids_1 = rename_stage_io_ren2_mask_1;
  assign dis_uops_0_valid = _T_2974_valid;
  assign dis_uops_0_uopc = _T_2974_uopc;
  assign dis_uops_0_inst = _T_2974_inst;
  assign dis_uops_0_pc = _T_2974_pc;
  assign dis_uops_0_iqtype = _T_2974_iqtype;
  assign dis_uops_0_fu_code = _T_2974_fu_code;
  assign dis_uops_0_allocate_brtag = _T_2974_allocate_brtag;
  assign dis_uops_0_is_br_or_jmp = _T_2974_is_br_or_jmp;
  assign dis_uops_0_is_jump = _T_2974_is_jump;
  assign dis_uops_0_is_jal = _T_2974_is_jal;
  assign dis_uops_0_is_ret = _T_2974_is_ret;
  assign dis_uops_0_is_call = _T_2974_is_call;
  assign dis_uops_0_br_mask = _T_2974_br_mask;
  assign dis_uops_0_br_tag = _T_2974_br_tag;
  assign dis_uops_0_br_prediction_btb_blame = _T_2974_br_prediction_btb_blame;
  assign dis_uops_0_br_prediction_btb_hit = _T_2974_br_prediction_btb_hit;
  assign dis_uops_0_br_prediction_btb_taken = _T_2974_br_prediction_btb_taken;
  assign dis_uops_0_br_prediction_bpd_blame = _T_2974_br_prediction_bpd_blame;
  assign dis_uops_0_br_prediction_bpd_hit = _T_2974_br_prediction_bpd_hit;
  assign dis_uops_0_br_prediction_bpd_taken = _T_2974_br_prediction_bpd_taken;
  assign dis_uops_0_br_prediction_bim_resp_value = _T_2974_br_prediction_bim_resp_value;
  assign dis_uops_0_br_prediction_bim_resp_entry_idx = _T_2974_br_prediction_bim_resp_entry_idx;
  assign dis_uops_0_br_prediction_bim_resp_way_idx = _T_2974_br_prediction_bim_resp_way_idx;
  assign dis_uops_0_br_prediction_bpd_resp_takens = _T_2974_br_prediction_bpd_resp_takens;
  assign dis_uops_0_br_prediction_bpd_resp_history = _T_2974_br_prediction_bpd_resp_history;
  assign dis_uops_0_br_prediction_bpd_resp_history_u = _T_2974_br_prediction_bpd_resp_history_u;
  assign dis_uops_0_br_prediction_bpd_resp_history_ptr = _T_2974_br_prediction_bpd_resp_history_ptr;
  assign dis_uops_0_br_prediction_bpd_resp_info = _T_2974_br_prediction_bpd_resp_info;
  assign dis_uops_0_stat_brjmp_mispredicted = _T_2974_stat_brjmp_mispredicted;
  assign dis_uops_0_stat_btb_made_pred = _T_2974_stat_btb_made_pred;
  assign dis_uops_0_stat_btb_mispredicted = _T_2974_stat_btb_mispredicted;
  assign dis_uops_0_stat_bpd_made_pred = _T_2974_stat_bpd_made_pred;
  assign dis_uops_0_stat_bpd_mispredicted = _T_2974_stat_bpd_mispredicted;
  assign dis_uops_0_fetch_pc_lob = _T_2974_fetch_pc_lob;
  assign dis_uops_0_imm_packed = _T_2974_imm_packed;
  assign dis_uops_0_csr_addr = _T_2974_csr_addr;
  assign dis_uops_0_rob_idx = _T_2974_rob_idx;
  assign dis_uops_0_ldq_idx = _T_2974_ldq_idx;
  assign dis_uops_0_stq_idx = _T_2974_stq_idx;
  assign dis_uops_0_brob_idx = _T_2974_brob_idx;
  assign dis_uops_0_pdst = _T_2974_pdst;
  assign dis_uops_0_pop1 = _T_2974_pop1;
  assign dis_uops_0_pop2 = _T_2974_pop2;
  assign dis_uops_0_pop3 = _T_2974_pop3;
  assign dis_uops_0_prs1_busy = _T_2974_prs1_busy;
  assign dis_uops_0_prs2_busy = _T_2974_prs2_busy;
  assign dis_uops_0_prs3_busy = _T_2974_prs3_busy;
  assign dis_uops_0_stale_pdst = _T_2974_stale_pdst;
  assign dis_uops_0_exception = _T_2974_exception;
  assign dis_uops_0_exc_cause = _T_2974_exc_cause;
  assign dis_uops_0_bypassable = _T_2974_bypassable;
  assign dis_uops_0_mem_cmd = _T_2974_mem_cmd;
  assign dis_uops_0_mem_typ = _T_2974_mem_typ;
  assign dis_uops_0_is_fence = _T_2974_is_fence;
  assign dis_uops_0_is_fencei = _T_2974_is_fencei;
  assign dis_uops_0_is_store = _T_2974_is_store;
  assign dis_uops_0_is_amo = _T_2974_is_amo;
  assign dis_uops_0_is_load = _T_2974_is_load;
  assign dis_uops_0_is_sys_pc2epc = _T_2974_is_sys_pc2epc;
  assign dis_uops_0_is_unique = _T_2974_is_unique;
  assign dis_uops_0_flush_on_commit = _T_2974_flush_on_commit;
  assign dis_uops_0_ldst = _T_2974_ldst;
  assign dis_uops_0_lrs1 = _T_2974_lrs1;
  assign dis_uops_0_lrs2 = _T_2974_lrs2;
  assign dis_uops_0_lrs3 = _T_2974_lrs3;
  assign dis_uops_0_ldst_val = _T_2974_ldst_val;
  assign dis_uops_0_dst_rtype = _T_2974_dst_rtype;
  assign dis_uops_0_lrs1_rtype = _T_2974_lrs1_rtype;
  assign dis_uops_0_lrs2_rtype = _T_2974_lrs2_rtype;
  assign dis_uops_0_frs3_en = _T_2974_frs3_en;
  assign dis_uops_0_fp_val = _T_2974_fp_val;
  assign dis_uops_0_fp_single = _T_2974_fp_single;
  assign dis_uops_0_xcpt_pf_if = _T_2974_xcpt_pf_if;
  assign dis_uops_0_xcpt_ae_if = _T_2974_xcpt_ae_if;
  assign dis_uops_0_replay_if = _T_2974_replay_if;
  assign dis_uops_0_xcpt_ma_if = _T_2974_xcpt_ma_if;
  assign dis_uops_0_debug_wdata = _T_2974_debug_wdata;
  assign dis_uops_0_debug_events_fetch_seq = _T_2974_debug_events_fetch_seq;
  assign dis_uops_1_valid = _T_2987_valid;
  assign dis_uops_1_uopc = _T_2987_uopc;
  assign dis_uops_1_inst = _T_2987_inst;
  assign dis_uops_1_pc = _T_2987_pc;
  assign dis_uops_1_iqtype = _T_2987_iqtype;
  assign dis_uops_1_fu_code = _T_2987_fu_code;
  assign dis_uops_1_allocate_brtag = _T_2987_allocate_brtag;
  assign dis_uops_1_is_br_or_jmp = _T_2987_is_br_or_jmp;
  assign dis_uops_1_is_jump = _T_2987_is_jump;
  assign dis_uops_1_is_jal = _T_2987_is_jal;
  assign dis_uops_1_is_ret = _T_2987_is_ret;
  assign dis_uops_1_is_call = _T_2987_is_call;
  assign dis_uops_1_br_mask = _T_2987_br_mask;
  assign dis_uops_1_br_tag = _T_2987_br_tag;
  assign dis_uops_1_br_prediction_btb_blame = _T_2987_br_prediction_btb_blame;
  assign dis_uops_1_br_prediction_btb_hit = _T_2987_br_prediction_btb_hit;
  assign dis_uops_1_br_prediction_btb_taken = _T_2987_br_prediction_btb_taken;
  assign dis_uops_1_br_prediction_bpd_blame = _T_2987_br_prediction_bpd_blame;
  assign dis_uops_1_br_prediction_bpd_hit = _T_2987_br_prediction_bpd_hit;
  assign dis_uops_1_br_prediction_bpd_taken = _T_2987_br_prediction_bpd_taken;
  assign dis_uops_1_br_prediction_bim_resp_value = _T_2987_br_prediction_bim_resp_value;
  assign dis_uops_1_br_prediction_bim_resp_entry_idx = _T_2987_br_prediction_bim_resp_entry_idx;
  assign dis_uops_1_br_prediction_bim_resp_way_idx = _T_2987_br_prediction_bim_resp_way_idx;
  assign dis_uops_1_br_prediction_bpd_resp_takens = _T_2987_br_prediction_bpd_resp_takens;
  assign dis_uops_1_br_prediction_bpd_resp_history = _T_2987_br_prediction_bpd_resp_history;
  assign dis_uops_1_br_prediction_bpd_resp_history_u = _T_2987_br_prediction_bpd_resp_history_u;
  assign dis_uops_1_br_prediction_bpd_resp_history_ptr = _T_2987_br_prediction_bpd_resp_history_ptr;
  assign dis_uops_1_br_prediction_bpd_resp_info = _T_2987_br_prediction_bpd_resp_info;
  assign dis_uops_1_stat_brjmp_mispredicted = _T_2987_stat_brjmp_mispredicted;
  assign dis_uops_1_stat_btb_made_pred = _T_2987_stat_btb_made_pred;
  assign dis_uops_1_stat_btb_mispredicted = _T_2987_stat_btb_mispredicted;
  assign dis_uops_1_stat_bpd_made_pred = _T_2987_stat_bpd_made_pred;
  assign dis_uops_1_stat_bpd_mispredicted = _T_2987_stat_bpd_mispredicted;
  assign dis_uops_1_fetch_pc_lob = _T_2987_fetch_pc_lob;
  assign dis_uops_1_imm_packed = _T_2987_imm_packed;
  assign dis_uops_1_csr_addr = _T_2987_csr_addr;
  assign dis_uops_1_rob_idx = _T_2987_rob_idx;
  assign dis_uops_1_ldq_idx = _T_2987_ldq_idx;
  assign dis_uops_1_stq_idx = _T_2987_stq_idx;
  assign dis_uops_1_brob_idx = _T_2987_brob_idx;
  assign dis_uops_1_pdst = _T_2987_pdst;
  assign dis_uops_1_pop1 = _T_2987_pop1;
  assign dis_uops_1_pop2 = _T_2987_pop2;
  assign dis_uops_1_pop3 = _T_2987_pop3;
  assign dis_uops_1_prs1_busy = _T_2987_prs1_busy;
  assign dis_uops_1_prs2_busy = _T_2987_prs2_busy;
  assign dis_uops_1_prs3_busy = _T_2987_prs3_busy;
  assign dis_uops_1_stale_pdst = _T_2987_stale_pdst;
  assign dis_uops_1_exception = _T_2987_exception;
  assign dis_uops_1_exc_cause = _T_2987_exc_cause;
  assign dis_uops_1_bypassable = _T_2987_bypassable;
  assign dis_uops_1_mem_cmd = _T_2987_mem_cmd;
  assign dis_uops_1_mem_typ = _T_2987_mem_typ;
  assign dis_uops_1_is_fence = _T_2987_is_fence;
  assign dis_uops_1_is_fencei = _T_2987_is_fencei;
  assign dis_uops_1_is_store = _T_2987_is_store;
  assign dis_uops_1_is_amo = _T_2987_is_amo;
  assign dis_uops_1_is_load = _T_2987_is_load;
  assign dis_uops_1_is_sys_pc2epc = _T_2987_is_sys_pc2epc;
  assign dis_uops_1_is_unique = _T_2987_is_unique;
  assign dis_uops_1_flush_on_commit = _T_2987_flush_on_commit;
  assign dis_uops_1_ldst = _T_2987_ldst;
  assign dis_uops_1_lrs1 = _T_2987_lrs1;
  assign dis_uops_1_lrs2 = _T_2987_lrs2;
  assign dis_uops_1_lrs3 = _T_2987_lrs3;
  assign dis_uops_1_ldst_val = _T_2987_ldst_val;
  assign dis_uops_1_dst_rtype = _T_2987_dst_rtype;
  assign dis_uops_1_lrs1_rtype = _T_2987_lrs1_rtype;
  assign dis_uops_1_lrs2_rtype = _T_2987_lrs2_rtype;
  assign dis_uops_1_frs3_en = _T_2987_frs3_en;
  assign dis_uops_1_fp_val = _T_2987_fp_val;
  assign dis_uops_1_fp_single = _T_2987_fp_single;
  assign dis_uops_1_xcpt_pf_if = _T_2987_xcpt_pf_if;
  assign dis_uops_1_xcpt_ae_if = _T_2987_xcpt_ae_if;
  assign dis_uops_1_replay_if = _T_2987_replay_if;
  assign dis_uops_1_xcpt_ma_if = _T_2987_xcpt_ma_if;
  assign dis_uops_1_debug_wdata = _T_2987_debug_wdata;
  assign dis_uops_1_debug_events_fetch_seq = _T_2987_debug_events_fetch_seq;
  assign iss_valids_0 = issue_units_0_io_iss_valids_0;
  assign iss_valids_1 = issue_units_1_io_iss_valids_0;
  assign iss_valids_2 = issue_units_1_io_iss_valids_1;
  assign iss_uops_0_uopc = issue_units_0_io_iss_uops_0_uopc;
  assign iss_uops_0_br_mask = issue_units_0_io_iss_uops_0_br_mask;
  assign iss_uops_0_imm_packed = issue_units_0_io_iss_uops_0_imm_packed;
  assign iss_uops_0_rob_idx = issue_units_0_io_iss_uops_0_rob_idx;
  assign iss_uops_0_ldq_idx = issue_units_0_io_iss_uops_0_ldq_idx;
  assign iss_uops_0_stq_idx = issue_units_0_io_iss_uops_0_stq_idx;
  assign iss_uops_0_pdst = issue_units_0_io_iss_uops_0_pdst;
  assign iss_uops_0_pop1 = issue_units_0_io_iss_uops_0_pop1;
  assign iss_uops_0_pop2 = issue_units_0_io_iss_uops_0_pop2;
  assign iss_uops_0_mem_cmd = issue_units_0_io_iss_uops_0_mem_cmd;
  assign iss_uops_0_mem_typ = issue_units_0_io_iss_uops_0_mem_typ;
  assign iss_uops_0_is_fence = issue_units_0_io_iss_uops_0_is_fence;
  assign iss_uops_0_is_store = issue_units_0_io_iss_uops_0_is_store;
  assign iss_uops_0_is_amo = issue_units_0_io_iss_uops_0_is_amo;
  assign iss_uops_0_is_load = issue_units_0_io_iss_uops_0_is_load;
  assign iss_uops_0_dst_rtype = issue_units_0_io_iss_uops_0_dst_rtype;
  assign iss_uops_0_lrs1_rtype = issue_units_0_io_iss_uops_0_lrs1_rtype;
  assign iss_uops_0_lrs2_rtype = issue_units_0_io_iss_uops_0_lrs2_rtype;
  assign iss_uops_0_fp_val = issue_units_0_io_iss_uops_0_fp_val;
  assign iss_uops_1_valid = issue_units_1_io_iss_uops_0_valid;
  assign iss_uops_1_iw_state = issue_units_1_io_iss_uops_0_iw_state;
  assign iss_uops_1_uopc = issue_units_1_io_iss_uops_0_uopc;
  assign iss_uops_1_inst = issue_units_1_io_iss_uops_0_inst;
  assign iss_uops_1_pc = issue_units_1_io_iss_uops_0_pc;
  assign iss_uops_1_iqtype = issue_units_1_io_iss_uops_0_iqtype;
  assign iss_uops_1_fu_code = issue_units_1_io_iss_uops_0_fu_code;
  assign iss_uops_1_allocate_brtag = issue_units_1_io_iss_uops_0_allocate_brtag;
  assign iss_uops_1_is_br_or_jmp = issue_units_1_io_iss_uops_0_is_br_or_jmp;
  assign iss_uops_1_is_jump = issue_units_1_io_iss_uops_0_is_jump;
  assign iss_uops_1_is_jal = issue_units_1_io_iss_uops_0_is_jal;
  assign iss_uops_1_is_ret = issue_units_1_io_iss_uops_0_is_ret;
  assign iss_uops_1_is_call = issue_units_1_io_iss_uops_0_is_call;
  assign iss_uops_1_br_mask = issue_units_1_io_iss_uops_0_br_mask;
  assign iss_uops_1_br_tag = issue_units_1_io_iss_uops_0_br_tag;
  assign iss_uops_1_br_prediction_btb_blame = issue_units_1_io_iss_uops_0_br_prediction_btb_blame;
  assign iss_uops_1_br_prediction_btb_hit = issue_units_1_io_iss_uops_0_br_prediction_btb_hit;
  assign iss_uops_1_br_prediction_btb_taken = issue_units_1_io_iss_uops_0_br_prediction_btb_taken;
  assign iss_uops_1_br_prediction_bpd_blame = issue_units_1_io_iss_uops_0_br_prediction_bpd_blame;
  assign iss_uops_1_br_prediction_bpd_hit = issue_units_1_io_iss_uops_0_br_prediction_bpd_hit;
  assign iss_uops_1_br_prediction_bpd_taken = issue_units_1_io_iss_uops_0_br_prediction_bpd_taken;
  assign iss_uops_1_br_prediction_bim_resp_value = issue_units_1_io_iss_uops_0_br_prediction_bim_resp_value;
  assign iss_uops_1_br_prediction_bim_resp_entry_idx = issue_units_1_io_iss_uops_0_br_prediction_bim_resp_entry_idx;
  assign iss_uops_1_br_prediction_bim_resp_way_idx = issue_units_1_io_iss_uops_0_br_prediction_bim_resp_way_idx;
  assign iss_uops_1_br_prediction_bpd_resp_takens = issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_takens;
  assign iss_uops_1_br_prediction_bpd_resp_history = issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history;
  assign iss_uops_1_br_prediction_bpd_resp_history_u = issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_u;
  assign iss_uops_1_br_prediction_bpd_resp_history_ptr = issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_history_ptr;
  assign iss_uops_1_br_prediction_bpd_resp_info = issue_units_1_io_iss_uops_0_br_prediction_bpd_resp_info;
  assign iss_uops_1_stat_brjmp_mispredicted = issue_units_1_io_iss_uops_0_stat_brjmp_mispredicted;
  assign iss_uops_1_stat_btb_made_pred = issue_units_1_io_iss_uops_0_stat_btb_made_pred;
  assign iss_uops_1_stat_btb_mispredicted = issue_units_1_io_iss_uops_0_stat_btb_mispredicted;
  assign iss_uops_1_stat_bpd_made_pred = issue_units_1_io_iss_uops_0_stat_bpd_made_pred;
  assign iss_uops_1_stat_bpd_mispredicted = issue_units_1_io_iss_uops_0_stat_bpd_mispredicted;
  assign iss_uops_1_fetch_pc_lob = issue_units_1_io_iss_uops_0_fetch_pc_lob;
  assign iss_uops_1_imm_packed = issue_units_1_io_iss_uops_0_imm_packed;
  assign iss_uops_1_csr_addr = issue_units_1_io_iss_uops_0_csr_addr;
  assign iss_uops_1_rob_idx = issue_units_1_io_iss_uops_0_rob_idx;
  assign iss_uops_1_ldq_idx = issue_units_1_io_iss_uops_0_ldq_idx;
  assign iss_uops_1_stq_idx = issue_units_1_io_iss_uops_0_stq_idx;
  assign iss_uops_1_brob_idx = issue_units_1_io_iss_uops_0_brob_idx;
  assign iss_uops_1_pdst = issue_units_1_io_iss_uops_0_pdst;
  assign iss_uops_1_pop1 = issue_units_1_io_iss_uops_0_pop1;
  assign iss_uops_1_pop2 = issue_units_1_io_iss_uops_0_pop2;
  assign iss_uops_1_pop3 = issue_units_1_io_iss_uops_0_pop3;
  assign iss_uops_1_prs1_busy = issue_units_1_io_iss_uops_0_prs1_busy;
  assign iss_uops_1_prs2_busy = issue_units_1_io_iss_uops_0_prs2_busy;
  assign iss_uops_1_prs3_busy = issue_units_1_io_iss_uops_0_prs3_busy;
  assign iss_uops_1_stale_pdst = issue_units_1_io_iss_uops_0_stale_pdst;
  assign iss_uops_1_exception = issue_units_1_io_iss_uops_0_exception;
  assign iss_uops_1_exc_cause = issue_units_1_io_iss_uops_0_exc_cause;
  assign iss_uops_1_bypassable = issue_units_1_io_iss_uops_0_bypassable;
  assign iss_uops_1_mem_cmd = issue_units_1_io_iss_uops_0_mem_cmd;
  assign iss_uops_1_mem_typ = issue_units_1_io_iss_uops_0_mem_typ;
  assign iss_uops_1_is_fence = issue_units_1_io_iss_uops_0_is_fence;
  assign iss_uops_1_is_fencei = issue_units_1_io_iss_uops_0_is_fencei;
  assign iss_uops_1_is_store = issue_units_1_io_iss_uops_0_is_store;
  assign iss_uops_1_is_amo = issue_units_1_io_iss_uops_0_is_amo;
  assign iss_uops_1_is_load = issue_units_1_io_iss_uops_0_is_load;
  assign iss_uops_1_is_sys_pc2epc = issue_units_1_io_iss_uops_0_is_sys_pc2epc;
  assign iss_uops_1_is_unique = issue_units_1_io_iss_uops_0_is_unique;
  assign iss_uops_1_flush_on_commit = issue_units_1_io_iss_uops_0_flush_on_commit;
  assign iss_uops_1_ldst = issue_units_1_io_iss_uops_0_ldst;
  assign iss_uops_1_lrs1 = issue_units_1_io_iss_uops_0_lrs1;
  assign iss_uops_1_lrs2 = issue_units_1_io_iss_uops_0_lrs2;
  assign iss_uops_1_lrs3 = issue_units_1_io_iss_uops_0_lrs3;
  assign iss_uops_1_ldst_val = issue_units_1_io_iss_uops_0_ldst_val;
  assign iss_uops_1_dst_rtype = issue_units_1_io_iss_uops_0_dst_rtype;
  assign iss_uops_1_lrs1_rtype = issue_units_1_io_iss_uops_0_lrs1_rtype;
  assign iss_uops_1_lrs2_rtype = issue_units_1_io_iss_uops_0_lrs2_rtype;
  assign iss_uops_1_frs3_en = issue_units_1_io_iss_uops_0_frs3_en;
  assign iss_uops_1_fp_val = issue_units_1_io_iss_uops_0_fp_val;
  assign iss_uops_1_fp_single = issue_units_1_io_iss_uops_0_fp_single;
  assign iss_uops_1_xcpt_pf_if = issue_units_1_io_iss_uops_0_xcpt_pf_if;
  assign iss_uops_1_xcpt_ae_if = issue_units_1_io_iss_uops_0_xcpt_ae_if;
  assign iss_uops_1_replay_if = issue_units_1_io_iss_uops_0_replay_if;
  assign iss_uops_1_xcpt_ma_if = issue_units_1_io_iss_uops_0_xcpt_ma_if;
  assign iss_uops_1_debug_wdata = issue_units_1_io_iss_uops_0_debug_wdata;
  assign iss_uops_1_debug_events_fetch_seq = issue_units_1_io_iss_uops_0_debug_events_fetch_seq;
  assign iss_uops_2_valid = issue_units_1_io_iss_uops_1_valid;
  assign iss_uops_2_iw_state = issue_units_1_io_iss_uops_1_iw_state;
  assign iss_uops_2_uopc = issue_units_1_io_iss_uops_1_uopc;
  assign iss_uops_2_inst = issue_units_1_io_iss_uops_1_inst;
  assign iss_uops_2_pc = issue_units_1_io_iss_uops_1_pc;
  assign iss_uops_2_iqtype = issue_units_1_io_iss_uops_1_iqtype;
  assign iss_uops_2_fu_code = issue_units_1_io_iss_uops_1_fu_code;
  assign iss_uops_2_allocate_brtag = issue_units_1_io_iss_uops_1_allocate_brtag;
  assign iss_uops_2_is_br_or_jmp = issue_units_1_io_iss_uops_1_is_br_or_jmp;
  assign iss_uops_2_is_jump = issue_units_1_io_iss_uops_1_is_jump;
  assign iss_uops_2_is_jal = issue_units_1_io_iss_uops_1_is_jal;
  assign iss_uops_2_is_ret = issue_units_1_io_iss_uops_1_is_ret;
  assign iss_uops_2_is_call = issue_units_1_io_iss_uops_1_is_call;
  assign iss_uops_2_br_mask = issue_units_1_io_iss_uops_1_br_mask;
  assign iss_uops_2_br_tag = issue_units_1_io_iss_uops_1_br_tag;
  assign iss_uops_2_br_prediction_btb_blame = issue_units_1_io_iss_uops_1_br_prediction_btb_blame;
  assign iss_uops_2_br_prediction_btb_hit = issue_units_1_io_iss_uops_1_br_prediction_btb_hit;
  assign iss_uops_2_br_prediction_btb_taken = issue_units_1_io_iss_uops_1_br_prediction_btb_taken;
  assign iss_uops_2_br_prediction_bpd_blame = issue_units_1_io_iss_uops_1_br_prediction_bpd_blame;
  assign iss_uops_2_br_prediction_bpd_hit = issue_units_1_io_iss_uops_1_br_prediction_bpd_hit;
  assign iss_uops_2_br_prediction_bpd_taken = issue_units_1_io_iss_uops_1_br_prediction_bpd_taken;
  assign iss_uops_2_br_prediction_bim_resp_value = issue_units_1_io_iss_uops_1_br_prediction_bim_resp_value;
  assign iss_uops_2_br_prediction_bim_resp_entry_idx = issue_units_1_io_iss_uops_1_br_prediction_bim_resp_entry_idx;
  assign iss_uops_2_br_prediction_bim_resp_way_idx = issue_units_1_io_iss_uops_1_br_prediction_bim_resp_way_idx;
  assign iss_uops_2_br_prediction_bpd_resp_takens = issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_takens;
  assign iss_uops_2_br_prediction_bpd_resp_history = issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history;
  assign iss_uops_2_br_prediction_bpd_resp_history_u = issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_u;
  assign iss_uops_2_br_prediction_bpd_resp_history_ptr = issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_history_ptr;
  assign iss_uops_2_br_prediction_bpd_resp_info = issue_units_1_io_iss_uops_1_br_prediction_bpd_resp_info;
  assign iss_uops_2_stat_brjmp_mispredicted = issue_units_1_io_iss_uops_1_stat_brjmp_mispredicted;
  assign iss_uops_2_stat_btb_made_pred = issue_units_1_io_iss_uops_1_stat_btb_made_pred;
  assign iss_uops_2_stat_btb_mispredicted = issue_units_1_io_iss_uops_1_stat_btb_mispredicted;
  assign iss_uops_2_stat_bpd_made_pred = issue_units_1_io_iss_uops_1_stat_bpd_made_pred;
  assign iss_uops_2_stat_bpd_mispredicted = issue_units_1_io_iss_uops_1_stat_bpd_mispredicted;
  assign iss_uops_2_fetch_pc_lob = issue_units_1_io_iss_uops_1_fetch_pc_lob;
  assign iss_uops_2_imm_packed = issue_units_1_io_iss_uops_1_imm_packed;
  assign iss_uops_2_csr_addr = issue_units_1_io_iss_uops_1_csr_addr;
  assign iss_uops_2_rob_idx = issue_units_1_io_iss_uops_1_rob_idx;
  assign iss_uops_2_ldq_idx = issue_units_1_io_iss_uops_1_ldq_idx;
  assign iss_uops_2_stq_idx = issue_units_1_io_iss_uops_1_stq_idx;
  assign iss_uops_2_brob_idx = issue_units_1_io_iss_uops_1_brob_idx;
  assign iss_uops_2_pdst = issue_units_1_io_iss_uops_1_pdst;
  assign iss_uops_2_pop1 = issue_units_1_io_iss_uops_1_pop1;
  assign iss_uops_2_pop2 = issue_units_1_io_iss_uops_1_pop2;
  assign iss_uops_2_pop3 = issue_units_1_io_iss_uops_1_pop3;
  assign iss_uops_2_prs1_busy = issue_units_1_io_iss_uops_1_prs1_busy;
  assign iss_uops_2_prs2_busy = issue_units_1_io_iss_uops_1_prs2_busy;
  assign iss_uops_2_prs3_busy = issue_units_1_io_iss_uops_1_prs3_busy;
  assign iss_uops_2_stale_pdst = issue_units_1_io_iss_uops_1_stale_pdst;
  assign iss_uops_2_exception = issue_units_1_io_iss_uops_1_exception;
  assign iss_uops_2_exc_cause = issue_units_1_io_iss_uops_1_exc_cause;
  assign iss_uops_2_bypassable = issue_units_1_io_iss_uops_1_bypassable;
  assign iss_uops_2_mem_cmd = issue_units_1_io_iss_uops_1_mem_cmd;
  assign iss_uops_2_mem_typ = issue_units_1_io_iss_uops_1_mem_typ;
  assign iss_uops_2_is_fence = issue_units_1_io_iss_uops_1_is_fence;
  assign iss_uops_2_is_fencei = issue_units_1_io_iss_uops_1_is_fencei;
  assign iss_uops_2_is_store = issue_units_1_io_iss_uops_1_is_store;
  assign iss_uops_2_is_amo = issue_units_1_io_iss_uops_1_is_amo;
  assign iss_uops_2_is_load = issue_units_1_io_iss_uops_1_is_load;
  assign iss_uops_2_is_sys_pc2epc = issue_units_1_io_iss_uops_1_is_sys_pc2epc;
  assign iss_uops_2_is_unique = issue_units_1_io_iss_uops_1_is_unique;
  assign iss_uops_2_flush_on_commit = issue_units_1_io_iss_uops_1_flush_on_commit;
  assign iss_uops_2_ldst = issue_units_1_io_iss_uops_1_ldst;
  assign iss_uops_2_lrs1 = issue_units_1_io_iss_uops_1_lrs1;
  assign iss_uops_2_lrs2 = issue_units_1_io_iss_uops_1_lrs2;
  assign iss_uops_2_lrs3 = issue_units_1_io_iss_uops_1_lrs3;
  assign iss_uops_2_ldst_val = issue_units_1_io_iss_uops_1_ldst_val;
  assign iss_uops_2_dst_rtype = issue_units_1_io_iss_uops_1_dst_rtype;
  assign iss_uops_2_lrs1_rtype = issue_units_1_io_iss_uops_1_lrs1_rtype;
  assign iss_uops_2_lrs2_rtype = issue_units_1_io_iss_uops_1_lrs2_rtype;
  assign iss_uops_2_frs3_en = issue_units_1_io_iss_uops_1_frs3_en;
  assign iss_uops_2_fp_val = issue_units_1_io_iss_uops_1_fp_val;
  assign iss_uops_2_fp_single = issue_units_1_io_iss_uops_1_fp_single;
  assign iss_uops_2_xcpt_pf_if = issue_units_1_io_iss_uops_1_xcpt_pf_if;
  assign iss_uops_2_xcpt_ae_if = issue_units_1_io_iss_uops_1_xcpt_ae_if;
  assign iss_uops_2_replay_if = issue_units_1_io_iss_uops_1_replay_if;
  assign iss_uops_2_xcpt_ma_if = issue_units_1_io_iss_uops_1_xcpt_ma_if;
  assign iss_uops_2_debug_wdata = issue_units_1_io_iss_uops_1_debug_wdata;
  assign iss_uops_2_debug_events_fetch_seq = issue_units_1_io_iss_uops_1_debug_events_fetch_seq;
  assign bypasses_valid_0 = csr_exe_unit_io_bypass_valid_0;
  assign bypasses_valid_1 = csr_exe_unit_io_bypass_valid_1;
  assign bypasses_valid_2 = csr_exe_unit_io_bypass_valid_2;
  assign bypasses_valid_3 = ALUExeUnit_io_bypass_valid_0;
  assign bypasses_uop_0_ctrl_rf_wen = csr_exe_unit_io_bypass_uop_0_ctrl_rf_wen;
  assign bypasses_uop_0_pdst = csr_exe_unit_io_bypass_uop_0_pdst;
  assign bypasses_uop_0_dst_rtype = csr_exe_unit_io_bypass_uop_0_dst_rtype;
  assign bypasses_uop_1_ctrl_rf_wen = csr_exe_unit_io_bypass_uop_1_ctrl_rf_wen;
  assign bypasses_uop_1_pdst = csr_exe_unit_io_bypass_uop_1_pdst;
  assign bypasses_uop_1_dst_rtype = csr_exe_unit_io_bypass_uop_1_dst_rtype;
  assign bypasses_uop_2_ctrl_rf_wen = csr_exe_unit_io_bypass_uop_2_ctrl_rf_wen;
  assign bypasses_uop_2_pdst = csr_exe_unit_io_bypass_uop_2_pdst;
  assign bypasses_uop_2_dst_rtype = csr_exe_unit_io_bypass_uop_2_dst_rtype;
  assign bypasses_uop_3_ctrl_rf_wen = ALUExeUnit_io_bypass_uop_0_ctrl_rf_wen;
  assign bypasses_uop_3_pdst = ALUExeUnit_io_bypass_uop_0_pdst;
  assign bypasses_uop_3_dst_rtype = ALUExeUnit_io_bypass_uop_0_dst_rtype;
  assign bypasses_data_0 = csr_exe_unit_io_bypass_data_0;
  assign bypasses_data_1 = csr_exe_unit_io_bypass_data_1;
  assign bypasses_data_2 = csr_exe_unit_io_bypass_data_2;
  assign bypasses_data_3 = ALUExeUnit_io_bypass_data_0;
  assign br_unit_take_pc = csr_exe_unit_io_br_unit_take_pc;
  assign br_unit_target = csr_exe_unit_io_br_unit_target;
  assign br_unit_brinfo_valid = csr_exe_unit_io_br_unit_brinfo_valid;
  assign br_unit_brinfo_mispredict = csr_exe_unit_io_br_unit_brinfo_mispredict;
  assign br_unit_brinfo_mask = csr_exe_unit_io_br_unit_brinfo_mask;
  assign br_unit_brinfo_tag = csr_exe_unit_io_br_unit_brinfo_tag;
  assign br_unit_brinfo_exe_mask = csr_exe_unit_io_br_unit_brinfo_exe_mask;
  assign br_unit_brinfo_rob_idx = csr_exe_unit_io_br_unit_brinfo_rob_idx;
  assign br_unit_brinfo_ldq_idx = csr_exe_unit_io_br_unit_brinfo_ldq_idx;
  assign br_unit_brinfo_stq_idx = csr_exe_unit_io_br_unit_brinfo_stq_idx;
  assign br_unit_brinfo_is_jr = csr_exe_unit_io_br_unit_brinfo_is_jr;
  assign br_unit_btb_update_valid = csr_exe_unit_io_br_unit_btb_update_valid;
  assign br_unit_btb_update_bits_pc = csr_exe_unit_io_br_unit_btb_update_bits_pc;
  assign br_unit_btb_update_bits_target = csr_exe_unit_io_br_unit_btb_update_bits_target;
  assign br_unit_btb_update_bits_cfi_pc = csr_exe_unit_io_br_unit_btb_update_bits_cfi_pc;
  assign br_unit_btb_update_bits_bpd_type = csr_exe_unit_io_br_unit_btb_update_bits_bpd_type;
  assign br_unit_btb_update_bits_cfi_type = csr_exe_unit_io_br_unit_btb_update_bits_cfi_type;
  assign br_unit_bim_update_valid = csr_exe_unit_io_br_unit_bim_update_valid;
  assign br_unit_bim_update_bits_taken = csr_exe_unit_io_br_unit_bim_update_bits_taken;
  assign br_unit_bim_update_bits_bim_resp_value = csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_value;
  assign br_unit_bim_update_bits_bim_resp_entry_idx = csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_entry_idx;
  assign br_unit_bim_update_bits_bim_resp_way_idx = csr_exe_unit_io_br_unit_bim_update_bits_bim_resp_way_idx;
  assign br_unit_bpd_update_valid = csr_exe_unit_io_br_unit_bpd_update_valid;
  assign br_unit_bpd_update_bits_br_pc = csr_exe_unit_io_br_unit_bpd_update_bits_br_pc;
  assign br_unit_bpd_update_bits_brob_idx = csr_exe_unit_io_br_unit_bpd_update_bits_brob_idx;
  assign br_unit_bpd_update_bits_mispredict = csr_exe_unit_io_br_unit_bpd_update_bits_mispredict;
  assign br_unit_bpd_update_bits_history = csr_exe_unit_io_br_unit_bpd_update_bits_history;
  assign br_unit_bpd_update_bits_history_ptr = csr_exe_unit_io_br_unit_bpd_update_bits_history_ptr;
  assign br_unit_bpd_update_bits_bpd_predict_val = csr_exe_unit_io_br_unit_bpd_update_bits_bpd_predict_val;
  assign br_unit_bpd_update_bits_bpd_mispredict = csr_exe_unit_io_br_unit_bpd_update_bits_bpd_mispredict;
  assign br_unit_bpd_update_bits_taken = csr_exe_unit_io_br_unit_bpd_update_bits_taken;
  assign br_unit_bpd_update_bits_is_br = csr_exe_unit_io_br_unit_bpd_update_bits_is_br;
  assign br_unit_bpd_update_bits_new_pc_same_packet = csr_exe_unit_io_br_unit_bpd_update_bits_new_pc_same_packet;
  assign br_unit_xcpt_valid = csr_exe_unit_io_br_unit_xcpt_valid;
  assign br_unit_xcpt_bits_uop_br_mask = csr_exe_unit_io_br_unit_xcpt_bits_uop_br_mask;
  assign br_unit_xcpt_bits_uop_rob_idx = csr_exe_unit_io_br_unit_xcpt_bits_uop_rob_idx;
  assign br_unit_xcpt_bits_badvaddr = csr_exe_unit_io_br_unit_xcpt_bits_badvaddr;
  assign csr_io_interrupts_debug = io_interrupts_debug;
  assign csr_io_interrupts_mtip = io_interrupts_mtip;
  assign csr_io_interrupts_msip = io_interrupts_msip;
  assign csr_io_interrupts_meip = io_interrupts_meip;
  assign csr_io_interrupts_seip = io_interrupts_seip;
  assign csr_io_rw_addr = csr_exe_unit_io_resp_0_bits_uop_csr_addr;
  assign csr_io_rw_cmd = _T_3033;
  assign csr_io_rw_wdata = csr_exe_unit_io_resp_0_bits_data;
  assign csr_io_decode_0_csr = decode_units_0_io_csr_decode_csr;
  assign csr_io_decode_1_csr = decode_units_1_io_csr_decode_csr;
  assign csr_io_exception = rob_io_com_xcpt_valid;
  assign csr_io_retire = _T_2698;
  assign csr_io_cause = rob_io_com_xcpt_bits_cause;
  assign csr_io_pc = rob_io_com_xcpt_bits_pc[39:0];
  assign csr_io_badaddr = rob_io_com_xcpt_bits_badvaddr[39:0];
  assign csr_io_fcsr_flags_valid = rob_io_commit_fflags_valid;
  assign csr_io_fcsr_flags_bits = rob_io_commit_fflags_bits;
  assign csr_io_counters_0_inc = {{1'd0}, _T_1564};
  assign csr_io_counters_1_inc = {{1'd0}, _T_1604};
  assign csr_io_counters_2_inc = {{1'd0}, _T_1644};
  assign csr_io_counters_3_inc = {{1'd0}, _T_1684};
  assign csr_io_counters_4_inc = {{1'd0}, _T_1724};
  assign csr_io_counters_5_inc = {{1'd0}, _T_1764};
  assign csr_io_counters_6_inc = {{1'd0}, _T_1804};
  assign csr_io_counters_7_inc = {{1'd0}, _T_1844};
  assign csr_io_counters_8_inc = {{1'd0}, _T_1884};
  assign csr_io_counters_9_inc = {{1'd0}, _T_1924};
  assign csr_io_counters_10_inc = {{1'd0}, _T_1964};
  assign csr_io_counters_11_inc = {{1'd0}, _T_2004};
  assign csr_io_counters_12_inc = {{1'd0}, _T_2044};
  assign csr_io_counters_13_inc = {{1'd0}, _T_2084};
  assign csr_io_counters_14_inc = {{1'd0}, _T_2124};
  assign csr_io_counters_15_inc = {{1'd0}, _T_2164};
  assign csr_io_counters_16_inc = {{1'd0}, _T_2204};
  assign csr_io_counters_17_inc = {{1'd0}, _T_2244};
  assign csr_io_counters_18_inc = {{1'd0}, _T_2284};
  assign csr_io_counters_19_inc = {{1'd0}, _T_2324};
  assign csr_io_counters_20_inc = {{1'd0}, _T_2364};
  assign csr_io_counters_21_inc = {{1'd0}, _T_2404};
  assign csr_io_counters_22_inc = {{1'd0}, _T_2444};
  assign csr_io_counters_23_inc = {{1'd0}, _T_2484};
  assign csr_io_counters_24_inc = {{1'd0}, _T_2524};
  assign csr_io_counters_25_inc = {{1'd0}, _T_2564};
  assign csr_io_counters_26_inc = {{1'd0}, _T_2604};
  assign csr_io_counters_27_inc = {{1'd0}, _T_2644};
  assign csr_io_counters_28_inc = {{1'd0}, _T_2684};
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign branch_mask_full_0 = dec_brmask_logic_io_is_full_0;
  assign branch_mask_full_1 = dec_brmask_logic_io_is_full_1;
  assign new_ldq_idx = lsu_io_new_ldq_idx;
  assign new_stq_idx = lsu_io_new_stq_idx;
  assign _T_2899_0_bim_resp_value = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_value;
  assign _T_2899_0_bim_resp_entry_idx = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_entry_idx;
  assign _T_2899_0_bim_resp_way_idx = dec_serializer_io_deq_bits_uops_0_br_prediction_bim_resp_way_idx;
  assign _T_2899_0_bpd_resp_history = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history;
  assign _T_2899_0_bpd_resp_history_ptr = dec_serializer_io_deq_bits_uops_0_br_prediction_bpd_resp_history_ptr;
  assign _T_2899_1_bim_resp_value = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_value;
  assign _T_2899_1_bim_resp_entry_idx = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_entry_idx;
  assign _T_2899_1_bim_resp_way_idx = dec_serializer_io_deq_bits_uops_1_br_prediction_bim_resp_way_idx;
  assign _T_2899_1_bpd_resp_history = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history;
  assign _T_2899_1_bpd_resp_history_ptr = dec_serializer_io_deq_bits_uops_1_br_prediction_bpd_resp_history_ptr;
  assign _T_2974_valid = rename_stage_io_ren2_uops_0_valid;
  assign _T_2974_uopc = rename_stage_io_ren2_uops_0_uopc;
  assign _T_2974_inst = rename_stage_io_ren2_uops_0_inst;
  assign _T_2974_pc = rename_stage_io_ren2_uops_0_pc;
  assign _T_2974_iqtype = rename_stage_io_ren2_uops_0_iqtype;
  assign _T_2974_fu_code = rename_stage_io_ren2_uops_0_fu_code;
  assign _T_2974_allocate_brtag = rename_stage_io_ren2_uops_0_allocate_brtag;
  assign _T_2974_is_br_or_jmp = rename_stage_io_ren2_uops_0_is_br_or_jmp;
  assign _T_2974_is_jump = rename_stage_io_ren2_uops_0_is_jump;
  assign _T_2974_is_jal = rename_stage_io_ren2_uops_0_is_jal;
  assign _T_2974_is_ret = rename_stage_io_ren2_uops_0_is_ret;
  assign _T_2974_is_call = rename_stage_io_ren2_uops_0_is_call;
  assign _T_2974_br_mask = _T_2981;
  assign _T_2974_br_tag = rename_stage_io_ren2_uops_0_br_tag;
  assign _T_2974_br_prediction_btb_blame = rename_stage_io_ren2_uops_0_br_prediction_btb_blame;
  assign _T_2974_br_prediction_btb_hit = rename_stage_io_ren2_uops_0_br_prediction_btb_hit;
  assign _T_2974_br_prediction_btb_taken = rename_stage_io_ren2_uops_0_br_prediction_btb_taken;
  assign _T_2974_br_prediction_bpd_blame = rename_stage_io_ren2_uops_0_br_prediction_bpd_blame;
  assign _T_2974_br_prediction_bpd_hit = rename_stage_io_ren2_uops_0_br_prediction_bpd_hit;
  assign _T_2974_br_prediction_bpd_taken = rename_stage_io_ren2_uops_0_br_prediction_bpd_taken;
  assign _T_2974_br_prediction_bim_resp_value = rename_stage_io_ren2_uops_0_br_prediction_bim_resp_value;
  assign _T_2974_br_prediction_bim_resp_entry_idx = rename_stage_io_ren2_uops_0_br_prediction_bim_resp_entry_idx;
  assign _T_2974_br_prediction_bim_resp_way_idx = rename_stage_io_ren2_uops_0_br_prediction_bim_resp_way_idx;
  assign _T_2974_br_prediction_bpd_resp_takens = rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_takens;
  assign _T_2974_br_prediction_bpd_resp_history = rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history;
  assign _T_2974_br_prediction_bpd_resp_history_u = rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_u;
  assign _T_2974_br_prediction_bpd_resp_history_ptr = rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_history_ptr;
  assign _T_2974_br_prediction_bpd_resp_info = rename_stage_io_ren2_uops_0_br_prediction_bpd_resp_info;
  assign _T_2974_stat_brjmp_mispredicted = rename_stage_io_ren2_uops_0_stat_brjmp_mispredicted;
  assign _T_2974_stat_btb_made_pred = rename_stage_io_ren2_uops_0_stat_btb_made_pred;
  assign _T_2974_stat_btb_mispredicted = rename_stage_io_ren2_uops_0_stat_btb_mispredicted;
  assign _T_2974_stat_bpd_made_pred = rename_stage_io_ren2_uops_0_stat_bpd_made_pred;
  assign _T_2974_stat_bpd_mispredicted = rename_stage_io_ren2_uops_0_stat_bpd_mispredicted;
  assign _T_2974_fetch_pc_lob = rename_stage_io_ren2_uops_0_fetch_pc_lob;
  assign _T_2974_imm_packed = rename_stage_io_ren2_uops_0_imm_packed;
  assign _T_2974_csr_addr = rename_stage_io_ren2_uops_0_csr_addr;
  assign _T_2974_rob_idx = rename_stage_io_ren2_uops_0_rob_idx;
  assign _T_2974_ldq_idx = rename_stage_io_ren2_uops_0_ldq_idx;
  assign _T_2974_stq_idx = rename_stage_io_ren2_uops_0_stq_idx;
  assign _T_2974_brob_idx = rename_stage_io_ren2_uops_0_brob_idx;
  assign _T_2974_pdst = rename_stage_io_ren2_uops_0_pdst;
  assign _T_2974_pop1 = rename_stage_io_ren2_uops_0_pop1;
  assign _T_2974_pop2 = rename_stage_io_ren2_uops_0_pop2;
  assign _T_2974_pop3 = rename_stage_io_ren2_uops_0_pop3;
  assign _T_2974_prs1_busy = rename_stage_io_ren2_uops_0_prs1_busy;
  assign _T_2974_prs2_busy = rename_stage_io_ren2_uops_0_prs2_busy;
  assign _T_2974_prs3_busy = rename_stage_io_ren2_uops_0_prs3_busy;
  assign _T_2974_stale_pdst = rename_stage_io_ren2_uops_0_stale_pdst;
  assign _T_2974_exception = rename_stage_io_ren2_uops_0_exception;
  assign _T_2974_exc_cause = rename_stage_io_ren2_uops_0_exc_cause;
  assign _T_2974_bypassable = rename_stage_io_ren2_uops_0_bypassable;
  assign _T_2974_mem_cmd = rename_stage_io_ren2_uops_0_mem_cmd;
  assign _T_2974_mem_typ = rename_stage_io_ren2_uops_0_mem_typ;
  assign _T_2974_is_fence = rename_stage_io_ren2_uops_0_is_fence;
  assign _T_2974_is_fencei = rename_stage_io_ren2_uops_0_is_fencei;
  assign _T_2974_is_store = rename_stage_io_ren2_uops_0_is_store;
  assign _T_2974_is_amo = rename_stage_io_ren2_uops_0_is_amo;
  assign _T_2974_is_load = rename_stage_io_ren2_uops_0_is_load;
  assign _T_2974_is_sys_pc2epc = rename_stage_io_ren2_uops_0_is_sys_pc2epc;
  assign _T_2974_is_unique = rename_stage_io_ren2_uops_0_is_unique;
  assign _T_2974_flush_on_commit = rename_stage_io_ren2_uops_0_flush_on_commit;
  assign _T_2974_ldst = rename_stage_io_ren2_uops_0_ldst;
  assign _T_2974_lrs1 = rename_stage_io_ren2_uops_0_lrs1;
  assign _T_2974_lrs2 = rename_stage_io_ren2_uops_0_lrs2;
  assign _T_2974_lrs3 = rename_stage_io_ren2_uops_0_lrs3;
  assign _T_2974_ldst_val = rename_stage_io_ren2_uops_0_ldst_val;
  assign _T_2974_dst_rtype = rename_stage_io_ren2_uops_0_dst_rtype;
  assign _T_2974_lrs1_rtype = rename_stage_io_ren2_uops_0_lrs1_rtype;
  assign _T_2974_lrs2_rtype = rename_stage_io_ren2_uops_0_lrs2_rtype;
  assign _T_2974_frs3_en = rename_stage_io_ren2_uops_0_frs3_en;
  assign _T_2974_fp_val = rename_stage_io_ren2_uops_0_fp_val;
  assign _T_2974_fp_single = rename_stage_io_ren2_uops_0_fp_single;
  assign _T_2974_xcpt_pf_if = rename_stage_io_ren2_uops_0_xcpt_pf_if;
  assign _T_2974_xcpt_ae_if = rename_stage_io_ren2_uops_0_xcpt_ae_if;
  assign _T_2974_replay_if = rename_stage_io_ren2_uops_0_replay_if;
  assign _T_2974_xcpt_ma_if = rename_stage_io_ren2_uops_0_xcpt_ma_if;
  assign _T_2974_debug_wdata = rename_stage_io_ren2_uops_0_debug_wdata;
  assign _T_2974_debug_events_fetch_seq = rename_stage_io_ren2_uops_0_debug_events_fetch_seq;
  assign _T_2987_valid = rename_stage_io_ren2_uops_1_valid;
  assign _T_2987_uopc = rename_stage_io_ren2_uops_1_uopc;
  assign _T_2987_inst = rename_stage_io_ren2_uops_1_inst;
  assign _T_2987_pc = rename_stage_io_ren2_uops_1_pc;
  assign _T_2987_iqtype = rename_stage_io_ren2_uops_1_iqtype;
  assign _T_2987_fu_code = rename_stage_io_ren2_uops_1_fu_code;
  assign _T_2987_allocate_brtag = rename_stage_io_ren2_uops_1_allocate_brtag;
  assign _T_2987_is_br_or_jmp = rename_stage_io_ren2_uops_1_is_br_or_jmp;
  assign _T_2987_is_jump = rename_stage_io_ren2_uops_1_is_jump;
  assign _T_2987_is_jal = rename_stage_io_ren2_uops_1_is_jal;
  assign _T_2987_is_ret = rename_stage_io_ren2_uops_1_is_ret;
  assign _T_2987_is_call = rename_stage_io_ren2_uops_1_is_call;
  assign _T_2987_br_mask = _T_2994;
  assign _T_2987_br_tag = rename_stage_io_ren2_uops_1_br_tag;
  assign _T_2987_br_prediction_btb_blame = rename_stage_io_ren2_uops_1_br_prediction_btb_blame;
  assign _T_2987_br_prediction_btb_hit = rename_stage_io_ren2_uops_1_br_prediction_btb_hit;
  assign _T_2987_br_prediction_btb_taken = rename_stage_io_ren2_uops_1_br_prediction_btb_taken;
  assign _T_2987_br_prediction_bpd_blame = rename_stage_io_ren2_uops_1_br_prediction_bpd_blame;
  assign _T_2987_br_prediction_bpd_hit = rename_stage_io_ren2_uops_1_br_prediction_bpd_hit;
  assign _T_2987_br_prediction_bpd_taken = rename_stage_io_ren2_uops_1_br_prediction_bpd_taken;
  assign _T_2987_br_prediction_bim_resp_value = rename_stage_io_ren2_uops_1_br_prediction_bim_resp_value;
  assign _T_2987_br_prediction_bim_resp_entry_idx = rename_stage_io_ren2_uops_1_br_prediction_bim_resp_entry_idx;
  assign _T_2987_br_prediction_bim_resp_way_idx = rename_stage_io_ren2_uops_1_br_prediction_bim_resp_way_idx;
  assign _T_2987_br_prediction_bpd_resp_takens = rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_takens;
  assign _T_2987_br_prediction_bpd_resp_history = rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history;
  assign _T_2987_br_prediction_bpd_resp_history_u = rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_u;
  assign _T_2987_br_prediction_bpd_resp_history_ptr = rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_history_ptr;
  assign _T_2987_br_prediction_bpd_resp_info = rename_stage_io_ren2_uops_1_br_prediction_bpd_resp_info;
  assign _T_2987_stat_brjmp_mispredicted = rename_stage_io_ren2_uops_1_stat_brjmp_mispredicted;
  assign _T_2987_stat_btb_made_pred = rename_stage_io_ren2_uops_1_stat_btb_made_pred;
  assign _T_2987_stat_btb_mispredicted = rename_stage_io_ren2_uops_1_stat_btb_mispredicted;
  assign _T_2987_stat_bpd_made_pred = rename_stage_io_ren2_uops_1_stat_bpd_made_pred;
  assign _T_2987_stat_bpd_mispredicted = rename_stage_io_ren2_uops_1_stat_bpd_mispredicted;
  assign _T_2987_fetch_pc_lob = rename_stage_io_ren2_uops_1_fetch_pc_lob;
  assign _T_2987_imm_packed = rename_stage_io_ren2_uops_1_imm_packed;
  assign _T_2987_csr_addr = rename_stage_io_ren2_uops_1_csr_addr;
  assign _T_2987_rob_idx = rename_stage_io_ren2_uops_1_rob_idx;
  assign _T_2987_ldq_idx = rename_stage_io_ren2_uops_1_ldq_idx;
  assign _T_2987_stq_idx = rename_stage_io_ren2_uops_1_stq_idx;
  assign _T_2987_brob_idx = rename_stage_io_ren2_uops_1_brob_idx;
  assign _T_2987_pdst = rename_stage_io_ren2_uops_1_pdst;
  assign _T_2987_pop1 = rename_stage_io_ren2_uops_1_pop1;
  assign _T_2987_pop2 = rename_stage_io_ren2_uops_1_pop2;
  assign _T_2987_pop3 = rename_stage_io_ren2_uops_1_pop3;
  assign _T_2987_prs1_busy = rename_stage_io_ren2_uops_1_prs1_busy;
  assign _T_2987_prs2_busy = rename_stage_io_ren2_uops_1_prs2_busy;
  assign _T_2987_prs3_busy = rename_stage_io_ren2_uops_1_prs3_busy;
  assign _T_2987_stale_pdst = rename_stage_io_ren2_uops_1_stale_pdst;
  assign _T_2987_exception = rename_stage_io_ren2_uops_1_exception;
  assign _T_2987_exc_cause = rename_stage_io_ren2_uops_1_exc_cause;
  assign _T_2987_bypassable = rename_stage_io_ren2_uops_1_bypassable;
  assign _T_2987_mem_cmd = rename_stage_io_ren2_uops_1_mem_cmd;
  assign _T_2987_mem_typ = rename_stage_io_ren2_uops_1_mem_typ;
  assign _T_2987_is_fence = rename_stage_io_ren2_uops_1_is_fence;
  assign _T_2987_is_fencei = rename_stage_io_ren2_uops_1_is_fencei;
  assign _T_2987_is_store = rename_stage_io_ren2_uops_1_is_store;
  assign _T_2987_is_amo = rename_stage_io_ren2_uops_1_is_amo;
  assign _T_2987_is_load = rename_stage_io_ren2_uops_1_is_load;
  assign _T_2987_is_sys_pc2epc = rename_stage_io_ren2_uops_1_is_sys_pc2epc;
  assign _T_2987_is_unique = rename_stage_io_ren2_uops_1_is_unique;
  assign _T_2987_flush_on_commit = rename_stage_io_ren2_uops_1_flush_on_commit;
  assign _T_2987_ldst = rename_stage_io_ren2_uops_1_ldst;
  assign _T_2987_lrs1 = rename_stage_io_ren2_uops_1_lrs1;
  assign _T_2987_lrs2 = rename_stage_io_ren2_uops_1_lrs2;
  assign _T_2987_lrs3 = rename_stage_io_ren2_uops_1_lrs3;
  assign _T_2987_ldst_val = rename_stage_io_ren2_uops_1_ldst_val;
  assign _T_2987_dst_rtype = rename_stage_io_ren2_uops_1_dst_rtype;
  assign _T_2987_lrs1_rtype = rename_stage_io_ren2_uops_1_lrs1_rtype;
  assign _T_2987_lrs2_rtype = rename_stage_io_ren2_uops_1_lrs2_rtype;
  assign _T_2987_frs3_en = rename_stage_io_ren2_uops_1_frs3_en;
  assign _T_2987_fp_val = rename_stage_io_ren2_uops_1_fp_val;
  assign _T_2987_fp_single = rename_stage_io_ren2_uops_1_fp_single;
  assign _T_2987_xcpt_pf_if = rename_stage_io_ren2_uops_1_xcpt_pf_if;
  assign _T_2987_xcpt_ae_if = rename_stage_io_ren2_uops_1_xcpt_ae_if;
  assign _T_2987_replay_if = rename_stage_io_ren2_uops_1_replay_if;
  assign _T_2987_xcpt_ma_if = rename_stage_io_ren2_uops_1_xcpt_ma_if;
  assign _T_2987_debug_wdata = rename_stage_io_ren2_uops_1_debug_wdata;
  assign _T_2987_debug_events_fetch_seq = rename_stage_io_ren2_uops_1_debug_events_fetch_seq;
  assign _T_3175_valid = ll_wbarb_io_out_valid;
  assign _T_3175_bits_addr = ll_wbarb_io_out_bits_uop_pdst;
  assign _T_3175_bits_data = ll_wbarb_io_out_bits_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1522 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1564 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_1604 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_1644 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_1684 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_1724 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_1764 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_1804 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_1844 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_1884 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_1924 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_1964 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_2004 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_2044 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_2084 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_2124 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_2164 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_2204 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_2244 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_2284 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_2324 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_2364 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_2404 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_2444 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_2484 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_2524 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_2564 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_2604 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_2644 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_2684 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{$random}};
  debug_tsc_reg = _RAND_30[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{$random}};
  debug_irt_reg = _RAND_31[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_2704 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_2715_valid = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_2715_bits_rs1 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_2715_bits_rs2 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{$random}};
  _T_2715_bits_addr = _RAND_36[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  dec_finished_mask = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_2923 = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_2928_bim_resp_value = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_2928_bim_resp_entry_idx = _RAND_40[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_2928_bim_resp_way_idx = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_2928_bpd_resp_history = _RAND_42[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_2928_bpd_resp_history_ptr = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_3029 = _RAND_44[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_3505 = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{$random}};
  _T_3507 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_3509 = _RAND_47[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_3511 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{$random}};
  _T_3513 = _RAND_49[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_3523 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_3536 = _RAND_51[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_3540 = _RAND_52[26:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_1522 <= io_imem_resp_valid;
    if (_T_1561) begin
      _T_1564 <= _T_1553;
    end else begin
      if (_T_1558) begin
        _T_1564 <= _T_1553;
      end else begin
        if (_T_1555) begin
          _T_1564 <= _T_1545;
        end else begin
          _T_1564 <= _T_1535;
        end
      end
    end
    if (_T_1601) begin
      _T_1604 <= _T_1593;
    end else begin
      if (_T_1598) begin
        _T_1604 <= _T_1593;
      end else begin
        if (_T_1595) begin
          _T_1604 <= _T_1585;
        end else begin
          _T_1604 <= _T_1575;
        end
      end
    end
    if (_T_1641) begin
      _T_1644 <= _T_1633;
    end else begin
      if (_T_1638) begin
        _T_1644 <= _T_1633;
      end else begin
        if (_T_1635) begin
          _T_1644 <= _T_1625;
        end else begin
          _T_1644 <= _T_1615;
        end
      end
    end
    if (_T_1681) begin
      _T_1684 <= _T_1673;
    end else begin
      if (_T_1678) begin
        _T_1684 <= _T_1673;
      end else begin
        if (_T_1675) begin
          _T_1684 <= _T_1665;
        end else begin
          _T_1684 <= _T_1655;
        end
      end
    end
    if (_T_1721) begin
      _T_1724 <= _T_1713;
    end else begin
      if (_T_1718) begin
        _T_1724 <= _T_1713;
      end else begin
        if (_T_1715) begin
          _T_1724 <= _T_1705;
        end else begin
          _T_1724 <= _T_1695;
        end
      end
    end
    if (_T_1761) begin
      _T_1764 <= _T_1753;
    end else begin
      if (_T_1758) begin
        _T_1764 <= _T_1753;
      end else begin
        if (_T_1755) begin
          _T_1764 <= _T_1745;
        end else begin
          _T_1764 <= _T_1735;
        end
      end
    end
    if (_T_1801) begin
      _T_1804 <= _T_1793;
    end else begin
      if (_T_1798) begin
        _T_1804 <= _T_1793;
      end else begin
        if (_T_1795) begin
          _T_1804 <= _T_1785;
        end else begin
          _T_1804 <= _T_1775;
        end
      end
    end
    if (_T_1841) begin
      _T_1844 <= _T_1833;
    end else begin
      if (_T_1838) begin
        _T_1844 <= _T_1833;
      end else begin
        if (_T_1835) begin
          _T_1844 <= _T_1825;
        end else begin
          _T_1844 <= _T_1815;
        end
      end
    end
    if (_T_1881) begin
      _T_1884 <= _T_1873;
    end else begin
      if (_T_1878) begin
        _T_1884 <= _T_1873;
      end else begin
        if (_T_1875) begin
          _T_1884 <= _T_1865;
        end else begin
          _T_1884 <= _T_1855;
        end
      end
    end
    if (_T_1921) begin
      _T_1924 <= _T_1913;
    end else begin
      if (_T_1918) begin
        _T_1924 <= _T_1913;
      end else begin
        if (_T_1915) begin
          _T_1924 <= _T_1905;
        end else begin
          _T_1924 <= _T_1895;
        end
      end
    end
    if (_T_1961) begin
      _T_1964 <= _T_1953;
    end else begin
      if (_T_1958) begin
        _T_1964 <= _T_1953;
      end else begin
        if (_T_1955) begin
          _T_1964 <= _T_1945;
        end else begin
          _T_1964 <= _T_1935;
        end
      end
    end
    if (_T_2001) begin
      _T_2004 <= _T_1993;
    end else begin
      if (_T_1998) begin
        _T_2004 <= _T_1993;
      end else begin
        if (_T_1995) begin
          _T_2004 <= _T_1985;
        end else begin
          _T_2004 <= _T_1975;
        end
      end
    end
    if (_T_2041) begin
      _T_2044 <= _T_2033;
    end else begin
      if (_T_2038) begin
        _T_2044 <= _T_2033;
      end else begin
        if (_T_2035) begin
          _T_2044 <= _T_2025;
        end else begin
          _T_2044 <= _T_2015;
        end
      end
    end
    if (_T_2081) begin
      _T_2084 <= _T_2073;
    end else begin
      if (_T_2078) begin
        _T_2084 <= _T_2073;
      end else begin
        if (_T_2075) begin
          _T_2084 <= _T_2065;
        end else begin
          _T_2084 <= _T_2055;
        end
      end
    end
    if (_T_2121) begin
      _T_2124 <= _T_2113;
    end else begin
      if (_T_2118) begin
        _T_2124 <= _T_2113;
      end else begin
        if (_T_2115) begin
          _T_2124 <= _T_2105;
        end else begin
          _T_2124 <= _T_2095;
        end
      end
    end
    if (_T_2161) begin
      _T_2164 <= _T_2153;
    end else begin
      if (_T_2158) begin
        _T_2164 <= _T_2153;
      end else begin
        if (_T_2155) begin
          _T_2164 <= _T_2145;
        end else begin
          _T_2164 <= _T_2135;
        end
      end
    end
    if (_T_2201) begin
      _T_2204 <= _T_2193;
    end else begin
      if (_T_2198) begin
        _T_2204 <= _T_2193;
      end else begin
        if (_T_2195) begin
          _T_2204 <= _T_2185;
        end else begin
          _T_2204 <= _T_2175;
        end
      end
    end
    if (_T_2241) begin
      _T_2244 <= _T_2233;
    end else begin
      if (_T_2238) begin
        _T_2244 <= _T_2233;
      end else begin
        if (_T_2235) begin
          _T_2244 <= _T_2225;
        end else begin
          _T_2244 <= _T_2215;
        end
      end
    end
    if (_T_2281) begin
      _T_2284 <= _T_2273;
    end else begin
      if (_T_2278) begin
        _T_2284 <= _T_2273;
      end else begin
        if (_T_2275) begin
          _T_2284 <= _T_2265;
        end else begin
          _T_2284 <= _T_2255;
        end
      end
    end
    if (_T_2321) begin
      _T_2324 <= _T_2313;
    end else begin
      if (_T_2318) begin
        _T_2324 <= _T_2313;
      end else begin
        if (_T_2315) begin
          _T_2324 <= _T_2305;
        end else begin
          _T_2324 <= _T_2295;
        end
      end
    end
    if (_T_2361) begin
      _T_2364 <= _T_2353;
    end else begin
      if (_T_2358) begin
        _T_2364 <= _T_2353;
      end else begin
        if (_T_2355) begin
          _T_2364 <= _T_2345;
        end else begin
          _T_2364 <= _T_2335;
        end
      end
    end
    if (_T_2401) begin
      _T_2404 <= _T_2393;
    end else begin
      if (_T_2398) begin
        _T_2404 <= _T_2393;
      end else begin
        if (_T_2395) begin
          _T_2404 <= _T_2385;
        end else begin
          _T_2404 <= _T_2375;
        end
      end
    end
    if (_T_2441) begin
      _T_2444 <= _T_2433;
    end else begin
      if (_T_2438) begin
        _T_2444 <= _T_2433;
      end else begin
        if (_T_2435) begin
          _T_2444 <= _T_2425;
        end else begin
          _T_2444 <= _T_2415;
        end
      end
    end
    if (_T_2481) begin
      _T_2484 <= _T_2473;
    end else begin
      if (_T_2478) begin
        _T_2484 <= _T_2473;
      end else begin
        if (_T_2475) begin
          _T_2484 <= _T_2465;
        end else begin
          _T_2484 <= _T_2455;
        end
      end
    end
    if (_T_2521) begin
      _T_2524 <= _T_2513;
    end else begin
      if (_T_2518) begin
        _T_2524 <= _T_2513;
      end else begin
        if (_T_2515) begin
          _T_2524 <= _T_2505;
        end else begin
          _T_2524 <= _T_2495;
        end
      end
    end
    if (_T_2561) begin
      _T_2564 <= _T_2553;
    end else begin
      if (_T_2558) begin
        _T_2564 <= _T_2553;
      end else begin
        if (_T_2555) begin
          _T_2564 <= _T_2545;
        end else begin
          _T_2564 <= _T_2535;
        end
      end
    end
    if (_T_2601) begin
      _T_2604 <= _T_2593;
    end else begin
      if (_T_2598) begin
        _T_2604 <= _T_2593;
      end else begin
        if (_T_2595) begin
          _T_2604 <= _T_2585;
        end else begin
          _T_2604 <= _T_2575;
        end
      end
    end
    if (_T_2641) begin
      _T_2644 <= _T_2633;
    end else begin
      if (_T_2638) begin
        _T_2644 <= _T_2633;
      end else begin
        if (_T_2635) begin
          _T_2644 <= _T_2625;
        end else begin
          _T_2644 <= _T_2615;
        end
      end
    end
    if (_T_2681) begin
      _T_2684 <= _T_2673;
    end else begin
      if (_T_2678) begin
        _T_2684 <= _T_2673;
      end else begin
        if (_T_2675) begin
          _T_2684 <= _T_2665;
        end else begin
          _T_2684 <= _T_2655;
        end
      end
    end
    if (reset) begin
      debug_tsc_reg <= 64'h0;
    end else begin
      debug_tsc_reg <= _T_2694;
    end
    if (reset) begin
      debug_irt_reg <= 64'h0;
    end else begin
      debug_irt_reg <= _T_2700;
    end
    _T_2704 <= lsu_io_exe_resp_bits_sfence_valid;
    _T_2715_valid <= lsu_io_exe_resp_bits_sfence_valid;
    _T_2715_bits_rs1 <= lsu_io_exe_resp_bits_sfence_bits_rs1;
    _T_2715_bits_rs2 <= lsu_io_exe_resp_bits_sfence_bits_rs2;
    _T_2715_bits_addr <= lsu_io_exe_resp_bits_sfence_bits_addr;
    if (reset) begin
      dec_finished_mask <= 2'h0;
    end else begin
      if (_T_2820) begin
        dec_finished_mask <= 2'h0;
      end else begin
        dec_finished_mask <= _T_2823;
      end
    end
    _T_2923 <= iss_uops_1_br_tag;
    _T_2928_bim_resp_value <= rename_stage_io_get_pred_info_bim_resp_value;
    _T_2928_bim_resp_entry_idx <= rename_stage_io_get_pred_info_bim_resp_entry_idx;
    _T_2928_bim_resp_way_idx <= rename_stage_io_get_pred_info_bim_resp_way_idx;
    _T_2928_bpd_resp_history <= rename_stage_io_get_pred_info_bpd_resp_history;
    _T_2928_bpd_resp_history_ptr <= rename_stage_io_get_pred_info_bpd_resp_history_ptr;
    _T_3029 <= _T_3027;
    _T_3505 <= iss_uops_1_rob_idx;
    _T_3507 <= rob_io_get_pc_curr_pc;
    _T_3509 <= rob_io_get_pc_curr_brob_idx;
    _T_3511 <= rob_io_get_pc_next_val;
    _T_3513 <= rob_io_get_pc_next_pc;
    _T_3523 <= rob_io_com_xcpt_valid;
    if (reset) begin
      _T_3536 <= 5'h0;
    end else begin
      _T_3536 <= _GEN_11[4:0];
    end
    if (reset) begin
      _T_3540 <= 27'h0;
    end else begin
      if (_T_3551) begin
        _T_3540 <= 27'h0;
      end else begin
        if (_T_3541) begin
          _T_3540 <= _T_3544;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2944) begin
          $fwrite(32'h80000002,"Assertion failed: Bypassing FP is not supported.\n    at core.scala:545 assert (!(iss_uops(i).dst_rtype === RT_FLT && iss_uops(i).bypassable), \"Bypassing FP is not supported.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2944) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2962) begin
          $fwrite(32'h80000002,"Assertion failed: Bypassing FP is not supported.\n    at core.scala:545 assert (!(iss_uops(i).dst_rtype === RT_FLT && iss_uops(i).bypassable), \"Bypassing FP is not supported.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2962) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3075) begin
          $fwrite(32'h80000002,"Assertion failed: the 65th bit was set on a fixed point write-back to the regfile.\n    at core.scala:842 assert (!(wbIsValid(RT_FIX) && exe_units(i).io.resp(j).bits.data(64).toBool),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3075) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3090) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] An Int writeback is being attempted with rf_wen disabled.\n    at core.scala:878 assert (!(exe_units(i).io.resp(j).valid &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3090) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3105) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] An FP writeback is being attempted to the Int Regfile.\n    at core.scala:875 assert (!wbIsValid(RT_FLT), \"[fppipeline] An FP writeback is being attempted to the Int Regfile.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3116) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] An Int writeback is being attempted with rf_wen disabled.\n    at core.scala:878 assert (!(exe_units(i).io.resp(j).valid &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3125) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] writeback being attempted to Int RF with dst != Int type exe_units(1).resp(0)\n    at core.scala:884 assert (!(exe_units(i).io.resp(j).valid &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3139) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] An FP writeback is being attempted to the Int Regfile.\n    at core.scala:875 assert (!wbIsValid(RT_FLT), \"[fppipeline] An FP writeback is being attempted to the Int Regfile.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3150) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] An Int writeback is being attempted with rf_wen disabled.\n    at core.scala:878 assert (!(exe_units(i).io.resp(j).valid &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3159) begin
          $fwrite(32'h80000002,"Assertion failed: [fppipeline] writeback being attempted to Int RF with dst != Int type exe_units(2).resp(0)\n    at core.scala:884 assert (!(exe_units(i).io.resp(j).valid &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at core.scala:902 assert (ll_wbarb.io.in(0).ready) // never backpressure the memory unit.\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3194) begin
          $fwrite(32'h80000002,"Assertion failed: [core] Assumption that dec_will_fire and ren1_mask are equal is being violated.\n    at core.scala:923 assert ((dec_will_fire zip rename_stage.io.ren1_mask map {case(d,r) => d === r}).reduce(_|_),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3214) begin
          $fwrite(32'h80000002,"Assertion failed: [core] I think we never use FP now.\n    at core.scala:964 assert (!(resp.valid && resp.bits.uop.fp_val && wb_uop.dst_rtype === RT_FLT && wb_uop.uopc =/= uopLD),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3360) begin
          $fwrite(32'h80000002,"Assertion failed: [core] FP wakeup does not write back to a FP register.\n    at core.scala:999 assert (!(wakeup.valid && wakeup.bits.uop.dst_rtype =/= RT_FLT),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3369) begin
          $fwrite(32'h80000002,"Assertion failed: [core] FP wakeup does not involve an FP instruction.\n    at core.scala:1002 assert (!(wakeup.valid && !wakeup.bits.uop.fp_val),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3369) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3494) begin
          $fwrite(32'h80000002,"Assertion failed: [core] FP wakeup does not write back to a FP register.\n    at core.scala:999 assert (!(wakeup.valid && wakeup.bits.uop.dst_rtype =/= RT_FLT),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3494) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3503) begin
          $fwrite(32'h80000002,"Assertion failed: [core] FP wakeup does not involve an FP instruction.\n    at core.scala:1002 assert (!(wakeup.valid && !wakeup.bits.uop.fp_val),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3503) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3520) begin
          $fwrite(32'h80000002,"Assertion failed: [core] single-step is unsupported.\n    at core.scala:1030 assert (!(csr.io.singleStep), \"[core] single-step is unsupported.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3520) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3532) begin
          $fwrite(32'h80000002,"Assertion failed: [core] exception occurred, but pipeline flush signal not set!\n    at core.scala:1049 assert (!(RegNext(rob.io.com_xcpt.valid) && !rob.io.flush.valid),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3532) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3560) begin
          $fwrite(32'h80000002,"Assertion failed: Pipeline has hung.\n    at core.scala:1061 assert (!(idle_cycles.value(13)), \"Pipeline has hung.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3560) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BoomTile_boom(
  input         clock,
  input         reset,
  input         auto_master_out_a_ready,
  output        auto_master_out_a_valid,
  output [2:0]  auto_master_out_a_bits_opcode,
  output [2:0]  auto_master_out_a_bits_param,
  output [3:0]  auto_master_out_a_bits_size,
  output [3:0]  auto_master_out_a_bits_source,
  output [31:0] auto_master_out_a_bits_address,
  output [7:0]  auto_master_out_a_bits_mask,
  output [63:0] auto_master_out_a_bits_data,
  output        auto_master_out_b_ready,
  input         auto_master_out_b_valid,
  input  [1:0]  auto_master_out_b_bits_param,
  input  [3:0]  auto_master_out_b_bits_size,
  input  [3:0]  auto_master_out_b_bits_source,
  input  [31:0] auto_master_out_b_bits_address,
  input         auto_master_out_c_ready,
  output        auto_master_out_c_valid,
  output [2:0]  auto_master_out_c_bits_opcode,
  output [2:0]  auto_master_out_c_bits_param,
  output [3:0]  auto_master_out_c_bits_size,
  output [3:0]  auto_master_out_c_bits_source,
  output [31:0] auto_master_out_c_bits_address,
  output [63:0] auto_master_out_c_bits_data,
  output        auto_master_out_d_ready,
  input         auto_master_out_d_valid,
  input  [2:0]  auto_master_out_d_bits_opcode,
  input  [1:0]  auto_master_out_d_bits_param,
  input  [3:0]  auto_master_out_d_bits_size,
  input  [3:0]  auto_master_out_d_bits_source,
  input  [2:0]  auto_master_out_d_bits_sink,
  input  [63:0] auto_master_out_d_bits_data,
  input         auto_master_out_d_bits_error,
  input         auto_master_out_e_ready,
  output        auto_master_out_e_valid,
  output [2:0]  auto_master_out_e_bits_sink,
  input         auto_int_in_0,
  input         auto_int_in_1,
  input         auto_int_in_2,
  input         auto_int_in_3,
  input         auto_int_in_4
);
  wire  tileBus_clock;
  wire  tileBus_reset;
  wire  tileBus_auto_in_1_a_ready;
  wire  tileBus_auto_in_1_a_valid;
  wire [31:0] tileBus_auto_in_1_a_bits_address;
  wire  tileBus_auto_in_1_d_valid;
  wire [2:0] tileBus_auto_in_1_d_bits_opcode;
  wire [3:0] tileBus_auto_in_1_d_bits_size;
  wire [63:0] tileBus_auto_in_1_d_bits_data;
  wire  tileBus_auto_in_1_d_bits_error;
  wire  tileBus_auto_in_0_a_ready;
  wire  tileBus_auto_in_0_a_valid;
  wire [2:0] tileBus_auto_in_0_a_bits_opcode;
  wire [2:0] tileBus_auto_in_0_a_bits_param;
  wire [3:0] tileBus_auto_in_0_a_bits_size;
  wire [2:0] tileBus_auto_in_0_a_bits_source;
  wire [31:0] tileBus_auto_in_0_a_bits_address;
  wire [7:0] tileBus_auto_in_0_a_bits_mask;
  wire [63:0] tileBus_auto_in_0_a_bits_data;
  wire  tileBus_auto_in_0_b_ready;
  wire  tileBus_auto_in_0_b_valid;
  wire [1:0] tileBus_auto_in_0_b_bits_param;
  wire [3:0] tileBus_auto_in_0_b_bits_size;
  wire [2:0] tileBus_auto_in_0_b_bits_source;
  wire [31:0] tileBus_auto_in_0_b_bits_address;
  wire  tileBus_auto_in_0_c_ready;
  wire  tileBus_auto_in_0_c_valid;
  wire [2:0] tileBus_auto_in_0_c_bits_opcode;
  wire [2:0] tileBus_auto_in_0_c_bits_param;
  wire [3:0] tileBus_auto_in_0_c_bits_size;
  wire [2:0] tileBus_auto_in_0_c_bits_source;
  wire [31:0] tileBus_auto_in_0_c_bits_address;
  wire [63:0] tileBus_auto_in_0_c_bits_data;
  wire  tileBus_auto_in_0_d_ready;
  wire  tileBus_auto_in_0_d_valid;
  wire [2:0] tileBus_auto_in_0_d_bits_opcode;
  wire [1:0] tileBus_auto_in_0_d_bits_param;
  wire [3:0] tileBus_auto_in_0_d_bits_size;
  wire [2:0] tileBus_auto_in_0_d_bits_source;
  wire [2:0] tileBus_auto_in_0_d_bits_sink;
  wire [63:0] tileBus_auto_in_0_d_bits_data;
  wire  tileBus_auto_in_0_e_ready;
  wire  tileBus_auto_in_0_e_valid;
  wire [2:0] tileBus_auto_in_0_e_bits_sink;
  wire  tileBus_auto_out_a_ready;
  wire  tileBus_auto_out_a_valid;
  wire [2:0] tileBus_auto_out_a_bits_opcode;
  wire [2:0] tileBus_auto_out_a_bits_param;
  wire [3:0] tileBus_auto_out_a_bits_size;
  wire [3:0] tileBus_auto_out_a_bits_source;
  wire [31:0] tileBus_auto_out_a_bits_address;
  wire [7:0] tileBus_auto_out_a_bits_mask;
  wire [63:0] tileBus_auto_out_a_bits_data;
  wire  tileBus_auto_out_b_ready;
  wire  tileBus_auto_out_b_valid;
  wire [1:0] tileBus_auto_out_b_bits_param;
  wire [3:0] tileBus_auto_out_b_bits_size;
  wire [3:0] tileBus_auto_out_b_bits_source;
  wire [31:0] tileBus_auto_out_b_bits_address;
  wire  tileBus_auto_out_c_ready;
  wire  tileBus_auto_out_c_valid;
  wire [2:0] tileBus_auto_out_c_bits_opcode;
  wire [2:0] tileBus_auto_out_c_bits_param;
  wire [3:0] tileBus_auto_out_c_bits_size;
  wire [3:0] tileBus_auto_out_c_bits_source;
  wire [31:0] tileBus_auto_out_c_bits_address;
  wire [63:0] tileBus_auto_out_c_bits_data;
  wire  tileBus_auto_out_d_ready;
  wire  tileBus_auto_out_d_valid;
  wire [2:0] tileBus_auto_out_d_bits_opcode;
  wire [1:0] tileBus_auto_out_d_bits_param;
  wire [3:0] tileBus_auto_out_d_bits_size;
  wire [3:0] tileBus_auto_out_d_bits_source;
  wire [2:0] tileBus_auto_out_d_bits_sink;
  wire [63:0] tileBus_auto_out_d_bits_data;
  wire  tileBus_auto_out_d_bits_error;
  wire  tileBus_auto_out_e_ready;
  wire  tileBus_auto_out_e_valid;
  wire [2:0] tileBus_auto_out_e_bits_sink;
  wire  dcache_clock;
  wire  dcache_reset;
  wire  dcache_auto_out_a_ready;
  wire  dcache_auto_out_a_valid;
  wire [2:0] dcache_auto_out_a_bits_opcode;
  wire [2:0] dcache_auto_out_a_bits_param;
  wire [3:0] dcache_auto_out_a_bits_size;
  wire [2:0] dcache_auto_out_a_bits_source;
  wire [31:0] dcache_auto_out_a_bits_address;
  wire [7:0] dcache_auto_out_a_bits_mask;
  wire [63:0] dcache_auto_out_a_bits_data;
  wire  dcache_auto_out_b_ready;
  wire  dcache_auto_out_b_valid;
  wire [1:0] dcache_auto_out_b_bits_param;
  wire [3:0] dcache_auto_out_b_bits_size;
  wire [2:0] dcache_auto_out_b_bits_source;
  wire [31:0] dcache_auto_out_b_bits_address;
  wire  dcache_auto_out_c_ready;
  wire  dcache_auto_out_c_valid;
  wire [2:0] dcache_auto_out_c_bits_opcode;
  wire [2:0] dcache_auto_out_c_bits_param;
  wire [3:0] dcache_auto_out_c_bits_size;
  wire [2:0] dcache_auto_out_c_bits_source;
  wire [31:0] dcache_auto_out_c_bits_address;
  wire [63:0] dcache_auto_out_c_bits_data;
  wire  dcache_auto_out_d_ready;
  wire  dcache_auto_out_d_valid;
  wire [2:0] dcache_auto_out_d_bits_opcode;
  wire [1:0] dcache_auto_out_d_bits_param;
  wire [3:0] dcache_auto_out_d_bits_size;
  wire [2:0] dcache_auto_out_d_bits_source;
  wire [2:0] dcache_auto_out_d_bits_sink;
  wire [63:0] dcache_auto_out_d_bits_data;
  wire  dcache_auto_out_e_ready;
  wire  dcache_auto_out_e_valid;
  wire [2:0] dcache_auto_out_e_bits_sink;
  wire  dcache_io_cpu_req_ready;
  wire  dcache_io_cpu_req_valid;
  wire [39:0] dcache_io_cpu_req_bits_addr;
  wire [6:0] dcache_io_cpu_req_bits_tag;
  wire [4:0] dcache_io_cpu_req_bits_cmd;
  wire [2:0] dcache_io_cpu_req_bits_typ;
  wire  dcache_io_cpu_s1_kill;
  wire [63:0] dcache_io_cpu_s1_data_data;
  wire  dcache_io_cpu_s2_nack;
  wire  dcache_io_cpu_resp_valid;
  wire [6:0] dcache_io_cpu_resp_bits_tag;
  wire [63:0] dcache_io_cpu_resp_bits_data;
  wire  dcache_io_cpu_resp_bits_has_data;
  wire  dcache_io_cpu_s2_xcpt_ma_ld;
  wire  dcache_io_cpu_s2_xcpt_ma_st;
  wire  dcache_io_cpu_s2_xcpt_pf_ld;
  wire  dcache_io_cpu_s2_xcpt_pf_st;
  wire  dcache_io_cpu_s2_xcpt_ae_ld;
  wire  dcache_io_cpu_s2_xcpt_ae_st;
  wire  dcache_io_cpu_invalidate_lr;
  wire  dcache_io_cpu_ordered;
  wire  dcache_io_cpu_perf_acquire;
  wire  dcache_io_cpu_perf_release;
  wire  dcache_io_cpu_perf_tlbMiss;
  wire  dcache_io_ptw_req_ready;
  wire  dcache_io_ptw_req_valid;
  wire [26:0] dcache_io_ptw_req_bits_addr;
  wire  dcache_io_ptw_resp_valid;
  wire  dcache_io_ptw_resp_bits_ae;
  wire [53:0] dcache_io_ptw_resp_bits_pte_ppn;
  wire  dcache_io_ptw_resp_bits_pte_d;
  wire  dcache_io_ptw_resp_bits_pte_a;
  wire  dcache_io_ptw_resp_bits_pte_g;
  wire  dcache_io_ptw_resp_bits_pte_u;
  wire  dcache_io_ptw_resp_bits_pte_x;
  wire  dcache_io_ptw_resp_bits_pte_w;
  wire  dcache_io_ptw_resp_bits_pte_r;
  wire  dcache_io_ptw_resp_bits_pte_v;
  wire [1:0] dcache_io_ptw_resp_bits_level;
  wire  dcache_io_ptw_resp_bits_homogeneous;
  wire [3:0] dcache_io_ptw_ptbr_mode;
  wire [1:0] dcache_io_ptw_status_dprv;
  wire  dcache_io_ptw_status_mxr;
  wire  dcache_io_ptw_status_sum;
  wire  frontend_clock;
  wire  frontend_reset;
  wire  frontend_auto_icache_master_out_a_ready;
  wire  frontend_auto_icache_master_out_a_valid;
  wire [31:0] frontend_auto_icache_master_out_a_bits_address;
  wire  frontend_auto_icache_master_out_d_valid;
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode;
  wire [3:0] frontend_auto_icache_master_out_d_bits_size;
  wire [63:0] frontend_auto_icache_master_out_d_bits_data;
  wire  frontend_auto_icache_master_out_d_bits_error;
  wire  frontend_io_cpu_req_valid;
  wire [39:0] frontend_io_cpu_req_bits_pc;
  wire  frontend_io_cpu_req_bits_speculative;
  wire  frontend_io_cpu_sfence_valid;
  wire  frontend_io_cpu_sfence_bits_rs1;
  wire  frontend_io_cpu_sfence_bits_rs2;
  wire [38:0] frontend_io_cpu_sfence_bits_addr;
  wire  frontend_io_cpu_resp_ready;
  wire  frontend_io_cpu_resp_valid;
  wire [39:0] frontend_io_cpu_resp_bits_pc;
  wire [63:0] frontend_io_cpu_resp_bits_data;
  wire [1:0] frontend_io_cpu_resp_bits_mask;
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst;
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst;
  wire  frontend_io_cpu_resp_bits_replay;
  wire  frontend_io_cpu_flush_icache;
  wire [39:0] frontend_io_cpu_npc;
  wire  frontend_io_cpu_perf_acquire;
  wire  frontend_io_cpu_perf_tlbMiss;
  wire  frontend_io_ptw_req_ready;
  wire  frontend_io_ptw_req_valid;
  wire [26:0] frontend_io_ptw_req_bits_addr;
  wire  frontend_io_ptw_resp_valid;
  wire  frontend_io_ptw_resp_bits_ae;
  wire [53:0] frontend_io_ptw_resp_bits_pte_ppn;
  wire  frontend_io_ptw_resp_bits_pte_d;
  wire  frontend_io_ptw_resp_bits_pte_a;
  wire  frontend_io_ptw_resp_bits_pte_g;
  wire  frontend_io_ptw_resp_bits_pte_u;
  wire  frontend_io_ptw_resp_bits_pte_x;
  wire  frontend_io_ptw_resp_bits_pte_w;
  wire  frontend_io_ptw_resp_bits_pte_r;
  wire  frontend_io_ptw_resp_bits_pte_v;
  wire [1:0] frontend_io_ptw_resp_bits_level;
  wire  frontend_io_ptw_resp_bits_homogeneous;
  wire [3:0] frontend_io_ptw_ptbr_mode;
  wire [1:0] frontend_io_ptw_status_prv;
  wire  _T_5_0;
  wire  _T_5_1;
  wire  _T_5_2;
  wire  _T_5_3;
  wire  _T_5_4;
  wire  _T_42_a_ready;
  wire  _T_42_a_valid;
  wire [2:0] _T_42_a_bits_opcode;
  wire [2:0] _T_42_a_bits_param;
  wire [3:0] _T_42_a_bits_size;
  wire [3:0] _T_42_a_bits_source;
  wire [31:0] _T_42_a_bits_address;
  wire [7:0] _T_42_a_bits_mask;
  wire [63:0] _T_42_a_bits_data;
  wire  _T_42_b_ready;
  wire  _T_42_b_valid;
  wire [1:0] _T_42_b_bits_param;
  wire [3:0] _T_42_b_bits_size;
  wire [3:0] _T_42_b_bits_source;
  wire [31:0] _T_42_b_bits_address;
  wire  _T_42_c_ready;
  wire  _T_42_c_valid;
  wire [2:0] _T_42_c_bits_opcode;
  wire [2:0] _T_42_c_bits_param;
  wire [3:0] _T_42_c_bits_size;
  wire [3:0] _T_42_c_bits_source;
  wire [31:0] _T_42_c_bits_address;
  wire [63:0] _T_42_c_bits_data;
  wire  _T_42_d_ready;
  wire  _T_42_d_valid;
  wire [2:0] _T_42_d_bits_opcode;
  wire [1:0] _T_42_d_bits_param;
  wire [3:0] _T_42_d_bits_size;
  wire [3:0] _T_42_d_bits_source;
  wire [2:0] _T_42_d_bits_sink;
  wire [63:0] _T_42_d_bits_data;
  wire  _T_42_d_bits_error;
  wire  _T_42_e_ready;
  wire  _T_42_e_valid;
  wire [2:0] _T_42_e_bits_sink;
  wire  _T_100_a_ready;
  wire  _T_100_a_valid;
  wire [2:0] _T_100_a_bits_opcode;
  wire [2:0] _T_100_a_bits_param;
  wire [3:0] _T_100_a_bits_size;
  wire [3:0] _T_100_a_bits_source;
  wire [31:0] _T_100_a_bits_address;
  wire [7:0] _T_100_a_bits_mask;
  wire [63:0] _T_100_a_bits_data;
  wire  _T_100_b_ready;
  wire  _T_100_b_valid;
  wire [1:0] _T_100_b_bits_param;
  wire [3:0] _T_100_b_bits_size;
  wire [3:0] _T_100_b_bits_source;
  wire [31:0] _T_100_b_bits_address;
  wire  _T_100_c_ready;
  wire  _T_100_c_valid;
  wire [2:0] _T_100_c_bits_opcode;
  wire [2:0] _T_100_c_bits_param;
  wire [3:0] _T_100_c_bits_size;
  wire [3:0] _T_100_c_bits_source;
  wire [31:0] _T_100_c_bits_address;
  wire [63:0] _T_100_c_bits_data;
  wire  _T_100_d_ready;
  wire  _T_100_d_valid;
  wire [2:0] _T_100_d_bits_opcode;
  wire [1:0] _T_100_d_bits_param;
  wire [3:0] _T_100_d_bits_size;
  wire [3:0] _T_100_d_bits_source;
  wire [2:0] _T_100_d_bits_sink;
  wire [63:0] _T_100_d_bits_data;
  wire  _T_100_d_bits_error;
  wire  _T_100_e_ready;
  wire  _T_100_e_valid;
  wire [2:0] _T_100_e_bits_sink;
  wire  fpuOpt_clock;
  wire  fpuOpt_reset;
  wire  fpuOpt_io_nack_mem;
  wire  dcacheArb_clock;
  wire  dcacheArb_io_requestor_0_req_ready;
  wire  dcacheArb_io_requestor_0_req_valid;
  wire [39:0] dcacheArb_io_requestor_0_req_bits_addr;
  wire  dcacheArb_io_requestor_0_s1_kill;
  wire  dcacheArb_io_requestor_0_s2_nack;
  wire  dcacheArb_io_requestor_0_resp_valid;
  wire [63:0] dcacheArb_io_requestor_0_resp_bits_data;
  wire  dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
  wire  dcacheArb_io_requestor_1_req_ready;
  wire  dcacheArb_io_requestor_1_req_valid;
  wire [39:0] dcacheArb_io_requestor_1_req_bits_addr;
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag;
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd;
  wire [2:0] dcacheArb_io_requestor_1_req_bits_typ;
  wire  dcacheArb_io_requestor_1_s1_kill;
  wire [63:0] dcacheArb_io_requestor_1_s1_data_data;
  wire  dcacheArb_io_requestor_1_s2_nack;
  wire  dcacheArb_io_requestor_1_resp_valid;
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag;
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data;
  wire  dcacheArb_io_requestor_1_resp_bits_has_data;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  wire  dcacheArb_io_requestor_1_invalidate_lr;
  wire  dcacheArb_io_requestor_1_ordered;
  wire  dcacheArb_io_requestor_1_perf_acquire;
  wire  dcacheArb_io_requestor_1_perf_release;
  wire  dcacheArb_io_requestor_1_perf_tlbMiss;
  wire  dcacheArb_io_mem_req_ready;
  wire  dcacheArb_io_mem_req_valid;
  wire [39:0] dcacheArb_io_mem_req_bits_addr;
  wire [6:0] dcacheArb_io_mem_req_bits_tag;
  wire [4:0] dcacheArb_io_mem_req_bits_cmd;
  wire [2:0] dcacheArb_io_mem_req_bits_typ;
  wire  dcacheArb_io_mem_s1_kill;
  wire [63:0] dcacheArb_io_mem_s1_data_data;
  wire  dcacheArb_io_mem_s2_nack;
  wire  dcacheArb_io_mem_resp_valid;
  wire [6:0] dcacheArb_io_mem_resp_bits_tag;
  wire [63:0] dcacheArb_io_mem_resp_bits_data;
  wire  dcacheArb_io_mem_resp_bits_has_data;
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld;
  wire  dcacheArb_io_mem_s2_xcpt_ma_st;
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld;
  wire  dcacheArb_io_mem_s2_xcpt_pf_st;
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld;
  wire  dcacheArb_io_mem_invalidate_lr;
  wire  dcacheArb_io_mem_ordered;
  wire  dcacheArb_io_mem_perf_acquire;
  wire  dcacheArb_io_mem_perf_release;
  wire  dcacheArb_io_mem_perf_tlbMiss;
  wire  ptw_clock;
  wire  ptw_reset;
  wire  ptw_io_requestor_0_req_ready;
  wire  ptw_io_requestor_0_req_valid;
  wire [26:0] ptw_io_requestor_0_req_bits_addr;
  wire  ptw_io_requestor_0_resp_valid;
  wire  ptw_io_requestor_0_resp_bits_ae;
  wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn;
  wire  ptw_io_requestor_0_resp_bits_pte_d;
  wire  ptw_io_requestor_0_resp_bits_pte_a;
  wire  ptw_io_requestor_0_resp_bits_pte_g;
  wire  ptw_io_requestor_0_resp_bits_pte_u;
  wire  ptw_io_requestor_0_resp_bits_pte_x;
  wire  ptw_io_requestor_0_resp_bits_pte_w;
  wire  ptw_io_requestor_0_resp_bits_pte_r;
  wire  ptw_io_requestor_0_resp_bits_pte_v;
  wire [1:0] ptw_io_requestor_0_resp_bits_level;
  wire  ptw_io_requestor_0_resp_bits_homogeneous;
  wire [3:0] ptw_io_requestor_0_ptbr_mode;
  wire [1:0] ptw_io_requestor_0_status_dprv;
  wire  ptw_io_requestor_0_status_mxr;
  wire  ptw_io_requestor_0_status_sum;
  wire  ptw_io_requestor_1_req_ready;
  wire  ptw_io_requestor_1_req_valid;
  wire [26:0] ptw_io_requestor_1_req_bits_addr;
  wire  ptw_io_requestor_1_resp_valid;
  wire  ptw_io_requestor_1_resp_bits_ae;
  wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn;
  wire  ptw_io_requestor_1_resp_bits_pte_d;
  wire  ptw_io_requestor_1_resp_bits_pte_a;
  wire  ptw_io_requestor_1_resp_bits_pte_g;
  wire  ptw_io_requestor_1_resp_bits_pte_u;
  wire  ptw_io_requestor_1_resp_bits_pte_x;
  wire  ptw_io_requestor_1_resp_bits_pte_w;
  wire  ptw_io_requestor_1_resp_bits_pte_r;
  wire  ptw_io_requestor_1_resp_bits_pte_v;
  wire [1:0] ptw_io_requestor_1_resp_bits_level;
  wire  ptw_io_requestor_1_resp_bits_homogeneous;
  wire [3:0] ptw_io_requestor_1_ptbr_mode;
  wire [1:0] ptw_io_requestor_1_status_prv;
  wire  ptw_io_requestor_2_req_ready;
  wire  ptw_io_requestor_2_req_valid;
  wire [26:0] ptw_io_requestor_2_req_bits_addr;
  wire  ptw_io_requestor_2_resp_valid;
  wire  ptw_io_requestor_2_resp_bits_ae;
  wire [53:0] ptw_io_requestor_2_resp_bits_pte_ppn;
  wire  ptw_io_requestor_2_resp_bits_pte_d;
  wire  ptw_io_requestor_2_resp_bits_pte_a;
  wire  ptw_io_requestor_2_resp_bits_pte_g;
  wire  ptw_io_requestor_2_resp_bits_pte_u;
  wire  ptw_io_requestor_2_resp_bits_pte_x;
  wire  ptw_io_requestor_2_resp_bits_pte_w;
  wire  ptw_io_requestor_2_resp_bits_pte_r;
  wire  ptw_io_requestor_2_resp_bits_pte_v;
  wire [1:0] ptw_io_requestor_2_resp_bits_level;
  wire  ptw_io_requestor_2_resp_bits_homogeneous;
  wire [3:0] ptw_io_requestor_2_ptbr_mode;
  wire [1:0] ptw_io_requestor_2_status_dprv;
  wire  ptw_io_requestor_2_status_mxr;
  wire  ptw_io_requestor_2_status_sum;
  wire  ptw_io_mem_req_ready;
  wire  ptw_io_mem_req_valid;
  wire [39:0] ptw_io_mem_req_bits_addr;
  wire  ptw_io_mem_s1_kill;
  wire  ptw_io_mem_s2_nack;
  wire  ptw_io_mem_resp_valid;
  wire [63:0] ptw_io_mem_resp_bits_data;
  wire  ptw_io_mem_s2_xcpt_ae_ld;
  wire [3:0] ptw_io_dpath_ptbr_mode;
  wire [43:0] ptw_io_dpath_ptbr_ppn;
  wire  ptw_io_dpath_sfence_valid;
  wire  ptw_io_dpath_sfence_bits_rs1;
  wire [1:0] ptw_io_dpath_status_dprv;
  wire [1:0] ptw_io_dpath_status_prv;
  wire  ptw_io_dpath_status_mxr;
  wire  ptw_io_dpath_status_sum;
  wire  core_clock;
  wire  core_reset;
  wire  core_io_interrupts_debug;
  wire  core_io_interrupts_mtip;
  wire  core_io_interrupts_msip;
  wire  core_io_interrupts_meip;
  wire  core_io_interrupts_seip;
  wire  core_io_imem_req_valid;
  wire [39:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_sfence_valid;
  wire  core_io_imem_sfence_bits_rs1;
  wire  core_io_imem_sfence_bits_rs2;
  wire [38:0] core_io_imem_sfence_bits_addr;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire [39:0] core_io_imem_resp_bits_pc;
  wire [63:0] core_io_imem_resp_bits_data;
  wire [1:0] core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_pf_inst;
  wire  core_io_imem_resp_bits_xcpt_ae_inst;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_perf_acquire;
  wire  core_io_imem_perf_tlbMiss;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [39:0] core_io_dmem_req_bits_addr;
  wire [6:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_s1_kill;
  wire [63:0] core_io_dmem_s1_data_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [6:0] core_io_dmem_resp_bits_tag;
  wire [63:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_has_data;
  wire  core_io_dmem_s2_xcpt_ma_ld;
  wire  core_io_dmem_s2_xcpt_ma_st;
  wire  core_io_dmem_s2_xcpt_pf_ld;
  wire  core_io_dmem_s2_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire  core_io_dmem_perf_acquire;
  wire  core_io_dmem_perf_release;
  wire  core_io_dmem_perf_tlbMiss;
  wire [3:0] core_io_ptw_ptbr_mode;
  wire [43:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_sfence_valid;
  wire  core_io_ptw_sfence_bits_rs1;
  wire [1:0] core_io_ptw_status_dprv;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_sum;
  wire  core_io_ptw_tlb_req_ready;
  wire  core_io_ptw_tlb_req_valid;
  wire [26:0] core_io_ptw_tlb_req_bits_addr;
  wire  core_io_ptw_tlb_resp_valid;
  wire  core_io_ptw_tlb_resp_bits_ae;
  wire [53:0] core_io_ptw_tlb_resp_bits_pte_ppn;
  wire  core_io_ptw_tlb_resp_bits_pte_d;
  wire  core_io_ptw_tlb_resp_bits_pte_a;
  wire  core_io_ptw_tlb_resp_bits_pte_g;
  wire  core_io_ptw_tlb_resp_bits_pte_u;
  wire  core_io_ptw_tlb_resp_bits_pte_x;
  wire  core_io_ptw_tlb_resp_bits_pte_w;
  wire  core_io_ptw_tlb_resp_bits_pte_r;
  wire  core_io_ptw_tlb_resp_bits_pte_v;
  wire [1:0] core_io_ptw_tlb_resp_bits_level;
  wire  core_io_ptw_tlb_resp_bits_homogeneous;
  wire [3:0] core_io_ptw_tlb_ptbr_mode;
  wire [1:0] core_io_ptw_tlb_status_dprv;
  wire  core_io_ptw_tlb_status_mxr;
  wire  core_io_ptw_tlb_status_sum;
  TLXbar_tileBus tileBus (
    .clock(tileBus_clock),
    .reset(tileBus_reset),
    .auto_in_1_a_ready(tileBus_auto_in_1_a_ready),
    .auto_in_1_a_valid(tileBus_auto_in_1_a_valid),
    .auto_in_1_a_bits_address(tileBus_auto_in_1_a_bits_address),
    .auto_in_1_d_valid(tileBus_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tileBus_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(tileBus_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_data(tileBus_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_error(tileBus_auto_in_1_d_bits_error),
    .auto_in_0_a_ready(tileBus_auto_in_0_a_ready),
    .auto_in_0_a_valid(tileBus_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tileBus_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tileBus_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tileBus_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tileBus_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tileBus_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tileBus_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tileBus_auto_in_0_a_bits_data),
    .auto_in_0_b_ready(tileBus_auto_in_0_b_ready),
    .auto_in_0_b_valid(tileBus_auto_in_0_b_valid),
    .auto_in_0_b_bits_param(tileBus_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tileBus_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tileBus_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tileBus_auto_in_0_b_bits_address),
    .auto_in_0_c_ready(tileBus_auto_in_0_c_ready),
    .auto_in_0_c_valid(tileBus_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tileBus_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tileBus_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tileBus_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tileBus_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tileBus_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tileBus_auto_in_0_c_bits_data),
    .auto_in_0_d_ready(tileBus_auto_in_0_d_ready),
    .auto_in_0_d_valid(tileBus_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tileBus_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tileBus_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tileBus_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tileBus_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tileBus_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_data(tileBus_auto_in_0_d_bits_data),
    .auto_in_0_e_ready(tileBus_auto_in_0_e_ready),
    .auto_in_0_e_valid(tileBus_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tileBus_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tileBus_auto_out_a_ready),
    .auto_out_a_valid(tileBus_auto_out_a_valid),
    .auto_out_a_bits_opcode(tileBus_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tileBus_auto_out_a_bits_param),
    .auto_out_a_bits_size(tileBus_auto_out_a_bits_size),
    .auto_out_a_bits_source(tileBus_auto_out_a_bits_source),
    .auto_out_a_bits_address(tileBus_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tileBus_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tileBus_auto_out_a_bits_data),
    .auto_out_b_ready(tileBus_auto_out_b_ready),
    .auto_out_b_valid(tileBus_auto_out_b_valid),
    .auto_out_b_bits_param(tileBus_auto_out_b_bits_param),
    .auto_out_b_bits_size(tileBus_auto_out_b_bits_size),
    .auto_out_b_bits_source(tileBus_auto_out_b_bits_source),
    .auto_out_b_bits_address(tileBus_auto_out_b_bits_address),
    .auto_out_c_ready(tileBus_auto_out_c_ready),
    .auto_out_c_valid(tileBus_auto_out_c_valid),
    .auto_out_c_bits_opcode(tileBus_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tileBus_auto_out_c_bits_param),
    .auto_out_c_bits_size(tileBus_auto_out_c_bits_size),
    .auto_out_c_bits_source(tileBus_auto_out_c_bits_source),
    .auto_out_c_bits_address(tileBus_auto_out_c_bits_address),
    .auto_out_c_bits_data(tileBus_auto_out_c_bits_data),
    .auto_out_d_ready(tileBus_auto_out_d_ready),
    .auto_out_d_valid(tileBus_auto_out_d_valid),
    .auto_out_d_bits_opcode(tileBus_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tileBus_auto_out_d_bits_param),
    .auto_out_d_bits_size(tileBus_auto_out_d_bits_size),
    .auto_out_d_bits_source(tileBus_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tileBus_auto_out_d_bits_sink),
    .auto_out_d_bits_data(tileBus_auto_out_d_bits_data),
    .auto_out_d_bits_error(tileBus_auto_out_d_bits_error),
    .auto_out_e_ready(tileBus_auto_out_e_ready),
    .auto_out_e_valid(tileBus_auto_out_e_valid),
    .auto_out_e_bits_sink(tileBus_auto_out_e_bits_sink)
  );
  NonBlockingDCache_dcache dcache (
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(dcache_io_cpu_req_bits_typ),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_invalidate_lr(dcache_io_cpu_invalidate_lr),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_cpu_perf_acquire(dcache_io_cpu_perf_acquire),
    .io_cpu_perf_release(dcache_io_cpu_perf_release),
    .io_cpu_perf_tlbMiss(dcache_io_cpu_perf_tlbMiss),
    .io_ptw_req_ready(dcache_io_ptw_req_ready),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dcache_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),
    .io_ptw_status_dprv(dcache_io_ptw_status_dprv),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum)
  );
  Frontend_frontend frontend (
    .clock(frontend_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_error(frontend_auto_icache_master_out_d_bits_error),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_mask(frontend_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_cpu_perf_acquire(frontend_io_cpu_perf_acquire),
    .io_cpu_perf_tlbMiss(frontend_io_cpu_perf_tlbMiss),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_addr(frontend_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_status_prv(frontend_io_ptw_status_prv)
  );
  FPU fpuOpt (
    .clock(fpuOpt_clock),
    .reset(fpuOpt_reset),
    .io_nack_mem(fpuOpt_io_nack_mem)
  );
  HellaCacheArbiter dcacheArb (
    .clock(dcacheArb_clock),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_invalidate_lr(dcacheArb_io_requestor_1_invalidate_lr),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_requestor_1_perf_acquire(dcacheArb_io_requestor_1_perf_acquire),
    .io_requestor_1_perf_release(dcacheArb_io_requestor_1_perf_release),
    .io_requestor_1_perf_tlbMiss(dcacheArb_io_requestor_1_perf_tlbMiss),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcacheArb_io_mem_req_bits_typ),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_invalidate_lr(dcacheArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcacheArb_io_mem_ordered),
    .io_mem_perf_acquire(dcacheArb_io_mem_perf_acquire),
    .io_mem_perf_release(dcacheArb_io_mem_perf_release),
    .io_mem_perf_tlbMiss(dcacheArb_io_mem_perf_tlbMiss)
  );
  PTW ptw (
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(ptw_io_requestor_0_req_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(ptw_io_requestor_1_req_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_2_req_ready(ptw_io_requestor_2_req_ready),
    .io_requestor_2_req_valid(ptw_io_requestor_2_req_valid),
    .io_requestor_2_req_bits_addr(ptw_io_requestor_2_req_bits_addr),
    .io_requestor_2_resp_valid(ptw_io_requestor_2_resp_valid),
    .io_requestor_2_resp_bits_ae(ptw_io_requestor_2_resp_bits_ae),
    .io_requestor_2_resp_bits_pte_ppn(ptw_io_requestor_2_resp_bits_pte_ppn),
    .io_requestor_2_resp_bits_pte_d(ptw_io_requestor_2_resp_bits_pte_d),
    .io_requestor_2_resp_bits_pte_a(ptw_io_requestor_2_resp_bits_pte_a),
    .io_requestor_2_resp_bits_pte_g(ptw_io_requestor_2_resp_bits_pte_g),
    .io_requestor_2_resp_bits_pte_u(ptw_io_requestor_2_resp_bits_pte_u),
    .io_requestor_2_resp_bits_pte_x(ptw_io_requestor_2_resp_bits_pte_x),
    .io_requestor_2_resp_bits_pte_w(ptw_io_requestor_2_resp_bits_pte_w),
    .io_requestor_2_resp_bits_pte_r(ptw_io_requestor_2_resp_bits_pte_r),
    .io_requestor_2_resp_bits_pte_v(ptw_io_requestor_2_resp_bits_pte_v),
    .io_requestor_2_resp_bits_level(ptw_io_requestor_2_resp_bits_level),
    .io_requestor_2_resp_bits_homogeneous(ptw_io_requestor_2_resp_bits_homogeneous),
    .io_requestor_2_ptbr_mode(ptw_io_requestor_2_ptbr_mode),
    .io_requestor_2_status_dprv(ptw_io_requestor_2_status_dprv),
    .io_requestor_2_status_mxr(ptw_io_requestor_2_status_mxr),
    .io_requestor_2_status_sum(ptw_io_requestor_2_status_sum),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum)
  );
  BoomCore core (
    .clock(core_clock),
    .reset(core_reset),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_interrupts_seip(core_io_interrupts_seip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),
    .io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_perf_acquire(core_io_imem_perf_acquire),
    .io_imem_perf_tlbMiss(core_io_imem_perf_tlbMiss),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_dmem_perf_acquire(core_io_dmem_perf_acquire),
    .io_dmem_perf_release(core_io_dmem_perf_release),
    .io_dmem_perf_tlbMiss(core_io_dmem_perf_tlbMiss),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_tlb_req_ready(core_io_ptw_tlb_req_ready),
    .io_ptw_tlb_req_valid(core_io_ptw_tlb_req_valid),
    .io_ptw_tlb_req_bits_addr(core_io_ptw_tlb_req_bits_addr),
    .io_ptw_tlb_resp_valid(core_io_ptw_tlb_resp_valid),
    .io_ptw_tlb_resp_bits_ae(core_io_ptw_tlb_resp_bits_ae),
    .io_ptw_tlb_resp_bits_pte_ppn(core_io_ptw_tlb_resp_bits_pte_ppn),
    .io_ptw_tlb_resp_bits_pte_d(core_io_ptw_tlb_resp_bits_pte_d),
    .io_ptw_tlb_resp_bits_pte_a(core_io_ptw_tlb_resp_bits_pte_a),
    .io_ptw_tlb_resp_bits_pte_g(core_io_ptw_tlb_resp_bits_pte_g),
    .io_ptw_tlb_resp_bits_pte_u(core_io_ptw_tlb_resp_bits_pte_u),
    .io_ptw_tlb_resp_bits_pte_x(core_io_ptw_tlb_resp_bits_pte_x),
    .io_ptw_tlb_resp_bits_pte_w(core_io_ptw_tlb_resp_bits_pte_w),
    .io_ptw_tlb_resp_bits_pte_r(core_io_ptw_tlb_resp_bits_pte_r),
    .io_ptw_tlb_resp_bits_pte_v(core_io_ptw_tlb_resp_bits_pte_v),
    .io_ptw_tlb_resp_bits_level(core_io_ptw_tlb_resp_bits_level),
    .io_ptw_tlb_resp_bits_homogeneous(core_io_ptw_tlb_resp_bits_homogeneous),
    .io_ptw_tlb_ptbr_mode(core_io_ptw_tlb_ptbr_mode),
    .io_ptw_tlb_status_dprv(core_io_ptw_tlb_status_dprv),
    .io_ptw_tlb_status_mxr(core_io_ptw_tlb_status_mxr),
    .io_ptw_tlb_status_sum(core_io_ptw_tlb_status_sum)
  );
  assign auto_master_out_a_valid = _T_42_a_valid;
  assign auto_master_out_a_bits_opcode = _T_42_a_bits_opcode;
  assign auto_master_out_a_bits_param = _T_42_a_bits_param;
  assign auto_master_out_a_bits_size = _T_42_a_bits_size;
  assign auto_master_out_a_bits_source = _T_42_a_bits_source;
  assign auto_master_out_a_bits_address = _T_42_a_bits_address;
  assign auto_master_out_a_bits_mask = _T_42_a_bits_mask;
  assign auto_master_out_a_bits_data = _T_42_a_bits_data;
  assign auto_master_out_b_ready = _T_42_b_ready;
  assign auto_master_out_c_valid = _T_42_c_valid;
  assign auto_master_out_c_bits_opcode = _T_42_c_bits_opcode;
  assign auto_master_out_c_bits_param = _T_42_c_bits_param;
  assign auto_master_out_c_bits_size = _T_42_c_bits_size;
  assign auto_master_out_c_bits_source = _T_42_c_bits_source;
  assign auto_master_out_c_bits_address = _T_42_c_bits_address;
  assign auto_master_out_c_bits_data = _T_42_c_bits_data;
  assign auto_master_out_d_ready = _T_42_d_ready;
  assign auto_master_out_e_valid = _T_42_e_valid;
  assign auto_master_out_e_bits_sink = _T_42_e_bits_sink;
  assign tileBus_clock = clock;
  assign tileBus_reset = reset;
  assign tileBus_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid;
  assign tileBus_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address;
  assign tileBus_auto_in_0_a_valid = dcache_auto_out_a_valid;
  assign tileBus_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode;
  assign tileBus_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param;
  assign tileBus_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size;
  assign tileBus_auto_in_0_a_bits_source = dcache_auto_out_a_bits_source;
  assign tileBus_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address;
  assign tileBus_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask;
  assign tileBus_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data;
  assign tileBus_auto_in_0_b_ready = dcache_auto_out_b_ready;
  assign tileBus_auto_in_0_c_valid = dcache_auto_out_c_valid;
  assign tileBus_auto_in_0_c_bits_opcode = dcache_auto_out_c_bits_opcode;
  assign tileBus_auto_in_0_c_bits_param = dcache_auto_out_c_bits_param;
  assign tileBus_auto_in_0_c_bits_size = dcache_auto_out_c_bits_size;
  assign tileBus_auto_in_0_c_bits_source = dcache_auto_out_c_bits_source;
  assign tileBus_auto_in_0_c_bits_address = dcache_auto_out_c_bits_address;
  assign tileBus_auto_in_0_c_bits_data = dcache_auto_out_c_bits_data;
  assign tileBus_auto_in_0_d_ready = dcache_auto_out_d_ready;
  assign tileBus_auto_in_0_e_valid = dcache_auto_out_e_valid;
  assign tileBus_auto_in_0_e_bits_sink = dcache_auto_out_e_bits_sink;
  assign tileBus_auto_out_a_ready = _T_100_a_ready;
  assign tileBus_auto_out_b_valid = _T_100_b_valid;
  assign tileBus_auto_out_b_bits_param = _T_100_b_bits_param;
  assign tileBus_auto_out_b_bits_size = _T_100_b_bits_size;
  assign tileBus_auto_out_b_bits_source = _T_100_b_bits_source;
  assign tileBus_auto_out_b_bits_address = _T_100_b_bits_address;
  assign tileBus_auto_out_c_ready = _T_100_c_ready;
  assign tileBus_auto_out_d_valid = _T_100_d_valid;
  assign tileBus_auto_out_d_bits_opcode = _T_100_d_bits_opcode;
  assign tileBus_auto_out_d_bits_param = _T_100_d_bits_param;
  assign tileBus_auto_out_d_bits_size = _T_100_d_bits_size;
  assign tileBus_auto_out_d_bits_source = _T_100_d_bits_source;
  assign tileBus_auto_out_d_bits_sink = _T_100_d_bits_sink;
  assign tileBus_auto_out_d_bits_data = _T_100_d_bits_data;
  assign tileBus_auto_out_d_bits_error = _T_100_d_bits_error;
  assign tileBus_auto_out_e_ready = _T_100_e_ready;
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = tileBus_auto_in_0_a_ready;
  assign dcache_auto_out_b_valid = tileBus_auto_in_0_b_valid;
  assign dcache_auto_out_b_bits_param = tileBus_auto_in_0_b_bits_param;
  assign dcache_auto_out_b_bits_size = tileBus_auto_in_0_b_bits_size;
  assign dcache_auto_out_b_bits_source = tileBus_auto_in_0_b_bits_source;
  assign dcache_auto_out_b_bits_address = tileBus_auto_in_0_b_bits_address;
  assign dcache_auto_out_c_ready = tileBus_auto_in_0_c_ready;
  assign dcache_auto_out_d_valid = tileBus_auto_in_0_d_valid;
  assign dcache_auto_out_d_bits_opcode = tileBus_auto_in_0_d_bits_opcode;
  assign dcache_auto_out_d_bits_param = tileBus_auto_in_0_d_bits_param;
  assign dcache_auto_out_d_bits_size = tileBus_auto_in_0_d_bits_size;
  assign dcache_auto_out_d_bits_source = tileBus_auto_in_0_d_bits_source;
  assign dcache_auto_out_d_bits_sink = tileBus_auto_in_0_d_bits_sink;
  assign dcache_auto_out_d_bits_data = tileBus_auto_in_0_d_bits_data;
  assign dcache_auto_out_e_ready = tileBus_auto_in_0_e_ready;
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid;
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr;
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag;
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd;
  assign dcache_io_cpu_req_bits_typ = dcacheArb_io_mem_req_bits_typ;
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill;
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data;
  assign dcache_io_cpu_invalidate_lr = dcacheArb_io_mem_invalidate_lr;
  assign dcache_io_ptw_req_ready = ptw_io_requestor_0_req_ready;
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid;
  assign dcache_io_ptw_resp_bits_ae = ptw_io_requestor_0_resp_bits_ae;
  assign dcache_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn;
  assign dcache_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d;
  assign dcache_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a;
  assign dcache_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g;
  assign dcache_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u;
  assign dcache_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x;
  assign dcache_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w;
  assign dcache_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r;
  assign dcache_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v;
  assign dcache_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level;
  assign dcache_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous;
  assign dcache_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode;
  assign dcache_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv;
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr;
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = tileBus_auto_in_1_a_ready;
  assign frontend_auto_icache_master_out_d_valid = tileBus_auto_in_1_d_valid;
  assign frontend_auto_icache_master_out_d_bits_opcode = tileBus_auto_in_1_d_bits_opcode;
  assign frontend_auto_icache_master_out_d_bits_size = tileBus_auto_in_1_d_bits_size;
  assign frontend_auto_icache_master_out_d_bits_data = tileBus_auto_in_1_d_bits_data;
  assign frontend_auto_icache_master_out_d_bits_error = tileBus_auto_in_1_d_bits_error;
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid;
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign frontend_io_cpu_sfence_valid = core_io_imem_sfence_valid;
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1;
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2;
  assign frontend_io_cpu_sfence_bits_addr = core_io_imem_sfence_bits_addr;
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready;
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid;
  assign frontend_io_ptw_resp_bits_ae = ptw_io_requestor_1_resp_bits_ae;
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn;
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d;
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a;
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g;
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u;
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x;
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w;
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r;
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v;
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level;
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous;
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode;
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv;
  assign _T_5_0 = auto_int_in_0;
  assign _T_5_1 = auto_int_in_1;
  assign _T_5_2 = auto_int_in_2;
  assign _T_5_3 = auto_int_in_3;
  assign _T_5_4 = auto_int_in_4;
  assign _T_42_a_ready = auto_master_out_a_ready;
  assign _T_42_a_valid = _T_100_a_valid;
  assign _T_42_a_bits_opcode = _T_100_a_bits_opcode;
  assign _T_42_a_bits_param = _T_100_a_bits_param;
  assign _T_42_a_bits_size = _T_100_a_bits_size;
  assign _T_42_a_bits_source = _T_100_a_bits_source;
  assign _T_42_a_bits_address = _T_100_a_bits_address;
  assign _T_42_a_bits_mask = _T_100_a_bits_mask;
  assign _T_42_a_bits_data = _T_100_a_bits_data;
  assign _T_42_b_ready = _T_100_b_ready;
  assign _T_42_b_valid = auto_master_out_b_valid;
  assign _T_42_b_bits_param = auto_master_out_b_bits_param;
  assign _T_42_b_bits_size = auto_master_out_b_bits_size;
  assign _T_42_b_bits_source = auto_master_out_b_bits_source;
  assign _T_42_b_bits_address = auto_master_out_b_bits_address;
  assign _T_42_c_ready = auto_master_out_c_ready;
  assign _T_42_c_valid = _T_100_c_valid;
  assign _T_42_c_bits_opcode = _T_100_c_bits_opcode;
  assign _T_42_c_bits_param = _T_100_c_bits_param;
  assign _T_42_c_bits_size = _T_100_c_bits_size;
  assign _T_42_c_bits_source = _T_100_c_bits_source;
  assign _T_42_c_bits_address = _T_100_c_bits_address;
  assign _T_42_c_bits_data = _T_100_c_bits_data;
  assign _T_42_d_ready = _T_100_d_ready;
  assign _T_42_d_valid = auto_master_out_d_valid;
  assign _T_42_d_bits_opcode = auto_master_out_d_bits_opcode;
  assign _T_42_d_bits_param = auto_master_out_d_bits_param;
  assign _T_42_d_bits_size = auto_master_out_d_bits_size;
  assign _T_42_d_bits_source = auto_master_out_d_bits_source;
  assign _T_42_d_bits_sink = auto_master_out_d_bits_sink;
  assign _T_42_d_bits_data = auto_master_out_d_bits_data;
  assign _T_42_d_bits_error = auto_master_out_d_bits_error;
  assign _T_42_e_ready = auto_master_out_e_ready;
  assign _T_42_e_valid = _T_100_e_valid;
  assign _T_42_e_bits_sink = _T_100_e_bits_sink;
  assign _T_100_a_ready = _T_42_a_ready;
  assign _T_100_a_valid = tileBus_auto_out_a_valid;
  assign _T_100_a_bits_opcode = tileBus_auto_out_a_bits_opcode;
  assign _T_100_a_bits_param = tileBus_auto_out_a_bits_param;
  assign _T_100_a_bits_size = tileBus_auto_out_a_bits_size;
  assign _T_100_a_bits_source = tileBus_auto_out_a_bits_source;
  assign _T_100_a_bits_address = tileBus_auto_out_a_bits_address;
  assign _T_100_a_bits_mask = tileBus_auto_out_a_bits_mask;
  assign _T_100_a_bits_data = tileBus_auto_out_a_bits_data;
  assign _T_100_b_ready = tileBus_auto_out_b_ready;
  assign _T_100_b_valid = _T_42_b_valid;
  assign _T_100_b_bits_param = _T_42_b_bits_param;
  assign _T_100_b_bits_size = _T_42_b_bits_size;
  assign _T_100_b_bits_source = _T_42_b_bits_source;
  assign _T_100_b_bits_address = _T_42_b_bits_address;
  assign _T_100_c_ready = _T_42_c_ready;
  assign _T_100_c_valid = tileBus_auto_out_c_valid;
  assign _T_100_c_bits_opcode = tileBus_auto_out_c_bits_opcode;
  assign _T_100_c_bits_param = tileBus_auto_out_c_bits_param;
  assign _T_100_c_bits_size = tileBus_auto_out_c_bits_size;
  assign _T_100_c_bits_source = tileBus_auto_out_c_bits_source;
  assign _T_100_c_bits_address = tileBus_auto_out_c_bits_address;
  assign _T_100_c_bits_data = tileBus_auto_out_c_bits_data;
  assign _T_100_d_ready = tileBus_auto_out_d_ready;
  assign _T_100_d_valid = _T_42_d_valid;
  assign _T_100_d_bits_opcode = _T_42_d_bits_opcode;
  assign _T_100_d_bits_param = _T_42_d_bits_param;
  assign _T_100_d_bits_size = _T_42_d_bits_size;
  assign _T_100_d_bits_source = _T_42_d_bits_source;
  assign _T_100_d_bits_sink = _T_42_d_bits_sink;
  assign _T_100_d_bits_data = _T_42_d_bits_data;
  assign _T_100_d_bits_error = _T_42_d_bits_error;
  assign _T_100_e_ready = _T_42_e_ready;
  assign _T_100_e_valid = tileBus_auto_out_e_valid;
  assign _T_100_e_bits_sink = tileBus_auto_out_e_bits_sink;
  assign fpuOpt_clock = clock;
  assign fpuOpt_reset = reset;
  assign dcacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid;
  assign dcacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr;
  assign dcacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill;
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid;
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcacheArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill;
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data;
  assign dcacheArb_io_requestor_1_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready;
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack;
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid;
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag;
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data;
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data;
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld;
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st;
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld;
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st;
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld;
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered;
  assign dcacheArb_io_mem_perf_acquire = dcache_io_cpu_perf_acquire;
  assign dcacheArb_io_mem_perf_release = dcache_io_cpu_perf_release;
  assign dcacheArb_io_mem_perf_tlbMiss = dcache_io_cpu_perf_tlbMiss;
  assign dcacheArb_clock = clock;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid;
  assign ptw_io_requestor_0_req_bits_addr = dcache_io_ptw_req_bits_addr;
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid;
  assign ptw_io_requestor_1_req_bits_addr = frontend_io_ptw_req_bits_addr;
  assign ptw_io_requestor_2_req_valid = core_io_ptw_tlb_req_valid;
  assign ptw_io_requestor_2_req_bits_addr = core_io_ptw_tlb_req_bits_addr;
  assign ptw_io_mem_req_ready = dcacheArb_io_requestor_0_req_ready;
  assign ptw_io_mem_s2_nack = dcacheArb_io_requestor_0_s2_nack;
  assign ptw_io_mem_resp_valid = dcacheArb_io_requestor_0_resp_valid;
  assign ptw_io_mem_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data;
  assign ptw_io_mem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode;
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn;
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid;
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1;
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv;
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv;
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr;
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum;
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign core_io_interrupts_debug = _T_5_0;
  assign core_io_interrupts_mtip = _T_5_2;
  assign core_io_interrupts_msip = _T_5_1;
  assign core_io_interrupts_meip = _T_5_3;
  assign core_io_interrupts_seip = _T_5_4;
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data;
  assign core_io_imem_resp_bits_mask = frontend_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst;
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst;
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay;
  assign core_io_imem_perf_acquire = frontend_io_cpu_perf_acquire;
  assign core_io_imem_perf_tlbMiss = frontend_io_cpu_perf_tlbMiss;
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready;
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack;
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid;
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag;
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data;
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data;
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered;
  assign core_io_dmem_perf_acquire = dcacheArb_io_requestor_1_perf_acquire;
  assign core_io_dmem_perf_release = dcacheArb_io_requestor_1_perf_release;
  assign core_io_dmem_perf_tlbMiss = dcacheArb_io_requestor_1_perf_tlbMiss;
  assign core_io_ptw_tlb_req_ready = ptw_io_requestor_2_req_ready;
  assign core_io_ptw_tlb_resp_valid = ptw_io_requestor_2_resp_valid;
  assign core_io_ptw_tlb_resp_bits_ae = ptw_io_requestor_2_resp_bits_ae;
  assign core_io_ptw_tlb_resp_bits_pte_ppn = ptw_io_requestor_2_resp_bits_pte_ppn;
  assign core_io_ptw_tlb_resp_bits_pte_d = ptw_io_requestor_2_resp_bits_pte_d;
  assign core_io_ptw_tlb_resp_bits_pte_a = ptw_io_requestor_2_resp_bits_pte_a;
  assign core_io_ptw_tlb_resp_bits_pte_g = ptw_io_requestor_2_resp_bits_pte_g;
  assign core_io_ptw_tlb_resp_bits_pte_u = ptw_io_requestor_2_resp_bits_pte_u;
  assign core_io_ptw_tlb_resp_bits_pte_x = ptw_io_requestor_2_resp_bits_pte_x;
  assign core_io_ptw_tlb_resp_bits_pte_w = ptw_io_requestor_2_resp_bits_pte_w;
  assign core_io_ptw_tlb_resp_bits_pte_r = ptw_io_requestor_2_resp_bits_pte_r;
  assign core_io_ptw_tlb_resp_bits_pte_v = ptw_io_requestor_2_resp_bits_pte_v;
  assign core_io_ptw_tlb_resp_bits_level = ptw_io_requestor_2_resp_bits_level;
  assign core_io_ptw_tlb_resp_bits_homogeneous = ptw_io_requestor_2_resp_bits_homogeneous;
  assign core_io_ptw_tlb_ptbr_mode = ptw_io_requestor_2_ptbr_mode;
  assign core_io_ptw_tlb_status_dprv = ptw_io_requestor_2_status_dprv;
  assign core_io_ptw_tlb_status_mxr = ptw_io_requestor_2_status_mxr;
  assign core_io_ptw_tlb_status_sum = ptw_io_requestor_2_status_sum;
  assign core_clock = clock;
  assign core_reset = reset;
endmodule
module IntXbar_intXbar(
  input   auto_int_in_3_0,
  input   auto_int_in_2_0,
  input   auto_int_in_1_0,
  input   auto_int_in_1_1,
  input   auto_int_in_0_0,
  output  auto_int_out_0,
  output  auto_int_out_1,
  output  auto_int_out_2,
  output  auto_int_out_3,
  output  auto_int_out_4
);
  wire  _T_5_0;
  wire  _T_12_0;
  wire  _T_12_1;
  wire  _T_20_0;
  wire  _T_27_0;
  wire  _T_34_0;
  wire  _T_34_1;
  wire  _T_34_2;
  wire  _T_34_3;
  wire  _T_34_4;
  assign auto_int_out_0 = _T_34_0;
  assign auto_int_out_1 = _T_34_1;
  assign auto_int_out_2 = _T_34_2;
  assign auto_int_out_3 = _T_34_3;
  assign auto_int_out_4 = _T_34_4;
  assign _T_5_0 = auto_int_in_0_0;
  assign _T_12_0 = auto_int_in_1_0;
  assign _T_12_1 = auto_int_in_1_1;
  assign _T_20_0 = auto_int_in_2_0;
  assign _T_27_0 = auto_int_in_3_0;
  assign _T_34_0 = _T_5_0;
  assign _T_34_1 = _T_12_0;
  assign _T_34_2 = _T_12_1;
  assign _T_34_3 = _T_20_0;
  assign _T_34_4 = _T_27_0;
endmodule
module Queue_27(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_50_data;
  wire  ram_opcode__T_50_addr;
  wire [2:0] ram_opcode__T_36_data;
  wire  ram_opcode__T_36_addr;
  wire  ram_opcode__T_36_mask;
  wire  ram_opcode__T_36_en;
  reg [2:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_50_data;
  wire  ram_param__T_50_addr;
  wire [2:0] ram_param__T_36_data;
  wire  ram_param__T_36_addr;
  wire  ram_param__T_36_mask;
  wire  ram_param__T_36_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [3:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] ram_source__T_50_data;
  wire  ram_source__T_50_addr;
  wire [3:0] ram_source__T_36_data;
  wire  ram_source__T_36_addr;
  wire  ram_source__T_36_mask;
  wire  ram_source__T_36_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_50_data;
  wire  ram_address__T_50_addr;
  wire [31:0] ram_address__T_36_data;
  wire  ram_address__T_36_addr;
  wire  ram_address__T_36_mask;
  wire  ram_address__T_36_en;
  reg [7:0] ram_mask [0:1];
  reg [31:0] _RAND_5;
  wire [7:0] ram_mask__T_50_data;
  wire  ram_mask__T_50_addr;
  wire [7:0] ram_mask__T_36_data;
  wire  ram_mask__T_36_addr;
  wire  ram_mask__T_36_mask;
  wire  ram_mask__T_36_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_6;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_10;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_11;
  wire  _T_45;
  wire  _GEN_12;
  wire  _T_47;
  wire  _T_49;
  assign ram_opcode__T_50_addr = value_1;
  assign ram_opcode__T_50_data = ram_opcode[ram_opcode__T_50_addr];
  assign ram_opcode__T_36_data = io_enq_bits_opcode;
  assign ram_opcode__T_36_addr = value;
  assign ram_opcode__T_36_mask = do_enq;
  assign ram_opcode__T_36_en = do_enq;
  assign ram_param__T_50_addr = value_1;
  assign ram_param__T_50_data = ram_param[ram_param__T_50_addr];
  assign ram_param__T_36_data = io_enq_bits_param;
  assign ram_param__T_36_addr = value;
  assign ram_param__T_36_mask = do_enq;
  assign ram_param__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_source__T_50_addr = value_1;
  assign ram_source__T_50_data = ram_source[ram_source__T_50_addr];
  assign ram_source__T_36_data = io_enq_bits_source;
  assign ram_source__T_36_addr = value;
  assign ram_source__T_36_mask = do_enq;
  assign ram_source__T_36_en = do_enq;
  assign ram_address__T_50_addr = value_1;
  assign ram_address__T_50_data = ram_address[ram_address__T_50_addr];
  assign ram_address__T_36_data = io_enq_bits_address;
  assign ram_address__T_36_addr = value;
  assign ram_address__T_36_mask = do_enq;
  assign ram_address__T_36_en = do_enq;
  assign ram_mask__T_50_addr = value_1;
  assign ram_mask__T_50_data = ram_mask[ram_mask__T_50_addr];
  assign ram_mask__T_36_data = io_enq_bits_mask;
  assign ram_mask__T_36_addr = value;
  assign ram_mask__T_36_mask = do_enq;
  assign ram_mask__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_10 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_11 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_12 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_opcode = ram_opcode__T_50_data;
  assign io_deq_bits_param = ram_param__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_source = ram_source__T_50_data;
  assign io_deq_bits_address = ram_address__T_50_data;
  assign io_deq_bits_mask = ram_mask__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_36_en & ram_opcode__T_36_mask) begin
      ram_opcode[ram_opcode__T_36_addr] <= ram_opcode__T_36_data;
    end
    if(ram_param__T_36_en & ram_param__T_36_mask) begin
      ram_param[ram_param__T_36_addr] <= ram_param__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_source__T_36_en & ram_source__T_36_mask) begin
      ram_source[ram_source__T_36_addr] <= ram_source__T_36_data;
    end
    if(ram_address__T_36_en & ram_address__T_36_mask) begin
      ram_address[ram_address__T_36_addr] <= ram_address__T_36_data;
    end
    if(ram_mask__T_36_en & ram_mask__T_36_mask) begin
      ram_mask[ram_mask__T_36_addr] <= ram_mask__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_28(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [2:0]  io_enq_bits_sink,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [2:0]  io_deq_bits_sink,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_50_data;
  wire  ram_opcode__T_50_addr;
  wire [2:0] ram_opcode__T_36_data;
  wire  ram_opcode__T_36_addr;
  wire  ram_opcode__T_36_mask;
  wire  ram_opcode__T_36_en;
  reg [1:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_50_data;
  wire  ram_param__T_50_addr;
  wire [1:0] ram_param__T_36_data;
  wire  ram_param__T_36_addr;
  wire  ram_param__T_36_mask;
  wire  ram_param__T_36_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [3:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] ram_source__T_50_data;
  wire  ram_source__T_50_addr;
  wire [3:0] ram_source__T_36_data;
  wire  ram_source__T_36_addr;
  wire  ram_source__T_36_mask;
  wire  ram_source__T_36_en;
  reg [2:0] ram_sink [0:1];
  reg [31:0] _RAND_4;
  wire [2:0] ram_sink__T_50_data;
  wire  ram_sink__T_50_addr;
  wire [2:0] ram_sink__T_36_data;
  wire  ram_sink__T_36_addr;
  wire  ram_sink__T_36_mask;
  wire  ram_sink__T_36_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_5;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg  ram_error [0:1];
  reg [31:0] _RAND_6;
  wire  ram_error__T_50_data;
  wire  ram_error__T_50_addr;
  wire  ram_error__T_36_data;
  wire  ram_error__T_36_addr;
  wire  ram_error__T_36_mask;
  wire  ram_error__T_36_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_10;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_11;
  wire  _T_45;
  wire  _GEN_12;
  wire  _T_47;
  wire  _T_49;
  assign ram_opcode__T_50_addr = value_1;
  assign ram_opcode__T_50_data = ram_opcode[ram_opcode__T_50_addr];
  assign ram_opcode__T_36_data = io_enq_bits_opcode;
  assign ram_opcode__T_36_addr = value;
  assign ram_opcode__T_36_mask = do_enq;
  assign ram_opcode__T_36_en = do_enq;
  assign ram_param__T_50_addr = value_1;
  assign ram_param__T_50_data = ram_param[ram_param__T_50_addr];
  assign ram_param__T_36_data = io_enq_bits_param;
  assign ram_param__T_36_addr = value;
  assign ram_param__T_36_mask = do_enq;
  assign ram_param__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_source__T_50_addr = value_1;
  assign ram_source__T_50_data = ram_source[ram_source__T_50_addr];
  assign ram_source__T_36_data = io_enq_bits_source;
  assign ram_source__T_36_addr = value;
  assign ram_source__T_36_mask = do_enq;
  assign ram_source__T_36_en = do_enq;
  assign ram_sink__T_50_addr = value_1;
  assign ram_sink__T_50_data = ram_sink[ram_sink__T_50_addr];
  assign ram_sink__T_36_data = io_enq_bits_sink;
  assign ram_sink__T_36_addr = value;
  assign ram_sink__T_36_mask = do_enq;
  assign ram_sink__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign ram_error__T_50_addr = value_1;
  assign ram_error__T_50_data = ram_error[ram_error__T_50_addr];
  assign ram_error__T_36_data = io_enq_bits_error;
  assign ram_error__T_36_addr = value;
  assign ram_error__T_36_mask = do_enq;
  assign ram_error__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_10 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_11 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_12 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_opcode = ram_opcode__T_50_data;
  assign io_deq_bits_param = ram_param__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_source = ram_source__T_50_data;
  assign io_deq_bits_sink = ram_sink__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign io_deq_bits_error = ram_error__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_error[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_36_en & ram_opcode__T_36_mask) begin
      ram_opcode[ram_opcode__T_36_addr] <= ram_opcode__T_36_data;
    end
    if(ram_param__T_36_en & ram_param__T_36_mask) begin
      ram_param[ram_param__T_36_addr] <= ram_param__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_source__T_36_en & ram_source__T_36_mask) begin
      ram_source[ram_source__T_36_addr] <= ram_source__T_36_data;
    end
    if(ram_sink__T_36_en & ram_sink__T_36_mask) begin
      ram_sink[ram_sink__T_36_addr] <= ram_sink__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if(ram_error__T_36_en & ram_error__T_36_mask) begin
      ram_error[ram_error__T_36_addr] <= ram_error__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_29(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address
);
  reg [1:0] ram_param [0:1];
  reg [31:0] _RAND_0;
  wire [1:0] ram_param__T_50_data;
  wire  ram_param__T_50_addr;
  wire [1:0] ram_param__T_36_data;
  wire  ram_param__T_36_addr;
  wire  ram_param__T_36_mask;
  wire  ram_param__T_36_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [3:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_source__T_50_data;
  wire  ram_source__T_50_addr;
  wire [3:0] ram_source__T_36_data;
  wire  ram_source__T_36_addr;
  wire  ram_source__T_36_mask;
  wire  ram_source__T_36_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_3;
  wire [31:0] ram_address__T_50_data;
  wire  ram_address__T_50_addr;
  wire [31:0] ram_address__T_36_data;
  wire  ram_address__T_36_addr;
  wire  ram_address__T_36_mask;
  wire  ram_address__T_36_en;
  reg  value;
  reg [31:0] _RAND_4;
  reg  value_1;
  reg [31:0] _RAND_5;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_10;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_11;
  wire  _T_45;
  wire  _GEN_12;
  wire  _T_47;
  wire  _T_49;
  assign ram_param__T_50_addr = value_1;
  assign ram_param__T_50_data = ram_param[ram_param__T_50_addr];
  assign ram_param__T_36_data = io_enq_bits_param;
  assign ram_param__T_36_addr = value;
  assign ram_param__T_36_mask = do_enq;
  assign ram_param__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_source__T_50_addr = value_1;
  assign ram_source__T_50_data = ram_source[ram_source__T_50_addr];
  assign ram_source__T_36_data = io_enq_bits_source;
  assign ram_source__T_36_addr = value;
  assign ram_source__T_36_mask = do_enq;
  assign ram_source__T_36_en = do_enq;
  assign ram_address__T_50_addr = value_1;
  assign ram_address__T_50_data = ram_address[ram_address__T_50_addr];
  assign ram_address__T_36_data = io_enq_bits_address;
  assign ram_address__T_36_addr = value;
  assign ram_address__T_36_mask = do_enq;
  assign ram_address__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_10 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_11 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_12 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_param = ram_param__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_source = ram_source__T_50_data;
  assign io_deq_bits_address = ram_address__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_param__T_36_en & ram_param__T_36_mask) begin
      ram_param[ram_param__T_36_addr] <= ram_param__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_source__T_36_en & ram_source__T_36_mask) begin
      ram_source[ram_source__T_36_addr] <= ram_source__T_36_data;
    end
    if(ram_address__T_36_en & ram_address__T_36_mask) begin
      ram_address[ram_address__T_36_addr] <= ram_address__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_30(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [63:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_50_data;
  wire  ram_opcode__T_50_addr;
  wire [2:0] ram_opcode__T_36_data;
  wire  ram_opcode__T_36_addr;
  wire  ram_opcode__T_36_mask;
  wire  ram_opcode__T_36_en;
  reg [2:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_50_data;
  wire  ram_param__T_50_addr;
  wire [2:0] ram_param__T_36_data;
  wire  ram_param__T_36_addr;
  wire  ram_param__T_36_mask;
  wire  ram_param__T_36_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [3:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] ram_source__T_50_data;
  wire  ram_source__T_50_addr;
  wire [3:0] ram_source__T_36_data;
  wire  ram_source__T_36_addr;
  wire  ram_source__T_36_mask;
  wire  ram_source__T_36_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_50_data;
  wire  ram_address__T_50_addr;
  wire [31:0] ram_address__T_36_data;
  wire  ram_address__T_36_addr;
  wire  ram_address__T_36_mask;
  wire  ram_address__T_36_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_5;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg  value;
  reg [31:0] _RAND_6;
  reg  value_1;
  reg [31:0] _RAND_7;
  reg  maybe_full;
  reg [31:0] _RAND_8;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_10;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_11;
  wire  _T_45;
  wire  _GEN_12;
  wire  _T_47;
  wire  _T_49;
  assign ram_opcode__T_50_addr = value_1;
  assign ram_opcode__T_50_data = ram_opcode[ram_opcode__T_50_addr];
  assign ram_opcode__T_36_data = io_enq_bits_opcode;
  assign ram_opcode__T_36_addr = value;
  assign ram_opcode__T_36_mask = do_enq;
  assign ram_opcode__T_36_en = do_enq;
  assign ram_param__T_50_addr = value_1;
  assign ram_param__T_50_data = ram_param[ram_param__T_50_addr];
  assign ram_param__T_36_data = io_enq_bits_param;
  assign ram_param__T_36_addr = value;
  assign ram_param__T_36_mask = do_enq;
  assign ram_param__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_source__T_50_addr = value_1;
  assign ram_source__T_50_data = ram_source[ram_source__T_50_addr];
  assign ram_source__T_36_data = io_enq_bits_source;
  assign ram_source__T_36_addr = value;
  assign ram_source__T_36_mask = do_enq;
  assign ram_source__T_36_en = do_enq;
  assign ram_address__T_50_addr = value_1;
  assign ram_address__T_50_data = ram_address[ram_address__T_50_addr];
  assign ram_address__T_36_data = io_enq_bits_address;
  assign ram_address__T_36_addr = value;
  assign ram_address__T_36_mask = do_enq;
  assign ram_address__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_10 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_11 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_12 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_opcode = ram_opcode__T_50_data;
  assign io_deq_bits_param = ram_param__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_source = ram_source__T_50_data;
  assign io_deq_bits_address = ram_address__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  maybe_full = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_36_en & ram_opcode__T_36_mask) begin
      ram_opcode[ram_opcode__T_36_addr] <= ram_opcode__T_36_data;
    end
    if(ram_param__T_36_en & ram_param__T_36_mask) begin
      ram_param[ram_param__T_36_addr] <= ram_param__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_source__T_36_en & ram_source__T_36_mask) begin
      ram_source[ram_source__T_36_addr] <= ram_source__T_36_data;
    end
    if(ram_address__T_36_en & ram_address__T_36_mask) begin
      ram_address[ram_address__T_36_addr] <= ram_address__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_31(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_sink,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_sink
);
  reg [2:0] ram_sink [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_sink__T_50_data;
  wire  ram_sink__T_50_addr;
  wire [2:0] ram_sink__T_36_data;
  wire  ram_sink__T_36_addr;
  wire  ram_sink__T_36_mask;
  wire  ram_sink__T_36_en;
  reg  value;
  reg [31:0] _RAND_1;
  reg  value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_4;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_5;
  wire  _T_45;
  wire  _GEN_6;
  wire  _T_47;
  wire  _T_49;
  assign ram_sink__T_50_addr = value_1;
  assign ram_sink__T_50_data = ram_sink[ram_sink__T_50_addr];
  assign ram_sink__T_36_data = io_enq_bits_sink;
  assign ram_sink__T_36_addr = value;
  assign ram_sink__T_36_mask = do_enq;
  assign ram_sink__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_4 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_5 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_6 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_sink = ram_sink__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_sink__T_36_en & ram_sink__T_36_mask) begin
      ram_sink[ram_sink__T_36_addr] <= ram_sink__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TLBuffer_SystemBus(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_param,
  output [3:0]  auto_in_b_bits_size,
  output [3:0]  auto_in_b_bits_source,
  output [31:0] auto_in_b_bits_address,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [3:0]  auto_in_c_bits_size,
  input  [3:0]  auto_in_c_bits_source,
  input  [31:0] auto_in_c_bits_address,
  input  [63:0] auto_in_c_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [3:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output [2:0]  auto_in_d_bits_sink,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error,
  output        auto_in_e_ready,
  input         auto_in_e_valid,
  input  [2:0]  auto_in_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [3:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [3:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [2:0]  auto_out_d_bits_sink,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_error,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [2:0]  auto_out_e_bits_sink
);
  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [2:0] _T_31_a_bits_param;
  wire [3:0] _T_31_a_bits_size;
  wire [3:0] _T_31_a_bits_source;
  wire [31:0] _T_31_a_bits_address;
  wire [7:0] _T_31_a_bits_mask;
  wire [63:0] _T_31_a_bits_data;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [1:0] _T_31_b_bits_param;
  wire [3:0] _T_31_b_bits_size;
  wire [3:0] _T_31_b_bits_source;
  wire [31:0] _T_31_b_bits_address;
  wire  _T_31_c_ready;
  wire  _T_31_c_valid;
  wire [2:0] _T_31_c_bits_opcode;
  wire [2:0] _T_31_c_bits_param;
  wire [3:0] _T_31_c_bits_size;
  wire [3:0] _T_31_c_bits_source;
  wire [31:0] _T_31_c_bits_address;
  wire [63:0] _T_31_c_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [1:0] _T_31_d_bits_param;
  wire [3:0] _T_31_d_bits_size;
  wire [3:0] _T_31_d_bits_source;
  wire [2:0] _T_31_d_bits_sink;
  wire [63:0] _T_31_d_bits_data;
  wire  _T_31_d_bits_error;
  wire  _T_31_e_ready;
  wire  _T_31_e_valid;
  wire [2:0] _T_31_e_bits_sink;
  wire  _T_89_a_ready;
  wire  _T_89_a_valid;
  wire [2:0] _T_89_a_bits_opcode;
  wire [2:0] _T_89_a_bits_param;
  wire [3:0] _T_89_a_bits_size;
  wire [3:0] _T_89_a_bits_source;
  wire [31:0] _T_89_a_bits_address;
  wire [7:0] _T_89_a_bits_mask;
  wire [63:0] _T_89_a_bits_data;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [1:0] _T_89_b_bits_param;
  wire [3:0] _T_89_b_bits_size;
  wire [3:0] _T_89_b_bits_source;
  wire [31:0] _T_89_b_bits_address;
  wire  _T_89_c_ready;
  wire  _T_89_c_valid;
  wire [2:0] _T_89_c_bits_opcode;
  wire [2:0] _T_89_c_bits_param;
  wire [3:0] _T_89_c_bits_size;
  wire [3:0] _T_89_c_bits_source;
  wire [31:0] _T_89_c_bits_address;
  wire [63:0] _T_89_c_bits_data;
  wire  _T_89_d_ready;
  wire  _T_89_d_valid;
  wire [2:0] _T_89_d_bits_opcode;
  wire [1:0] _T_89_d_bits_param;
  wire [3:0] _T_89_d_bits_size;
  wire [3:0] _T_89_d_bits_source;
  wire [2:0] _T_89_d_bits_sink;
  wire [63:0] _T_89_d_bits_data;
  wire  _T_89_d_bits_error;
  wire  _T_89_e_ready;
  wire  _T_89_e_valid;
  wire [2:0] _T_89_e_bits_sink;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [3:0] Queue_io_enq_bits_size;
  wire [3:0] Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [7:0] Queue_io_enq_bits_mask;
  wire [63:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [3:0] Queue_io_deq_bits_size;
  wire [3:0] Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [7:0] Queue_io_deq_bits_mask;
  wire [63:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [1:0] Queue_1_io_enq_bits_param;
  wire [3:0] Queue_1_io_enq_bits_size;
  wire [3:0] Queue_1_io_enq_bits_source;
  wire [2:0] Queue_1_io_enq_bits_sink;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [1:0] Queue_1_io_deq_bits_param;
  wire [3:0] Queue_1_io_deq_bits_size;
  wire [3:0] Queue_1_io_deq_bits_source;
  wire [2:0] Queue_1_io_deq_bits_sink;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [1:0] Queue_2_io_enq_bits_param;
  wire [3:0] Queue_2_io_enq_bits_size;
  wire [3:0] Queue_2_io_enq_bits_source;
  wire [31:0] Queue_2_io_enq_bits_address;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [1:0] Queue_2_io_deq_bits_param;
  wire [3:0] Queue_2_io_deq_bits_size;
  wire [3:0] Queue_2_io_deq_bits_source;
  wire [31:0] Queue_2_io_deq_bits_address;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [2:0] Queue_3_io_enq_bits_opcode;
  wire [2:0] Queue_3_io_enq_bits_param;
  wire [3:0] Queue_3_io_enq_bits_size;
  wire [3:0] Queue_3_io_enq_bits_source;
  wire [31:0] Queue_3_io_enq_bits_address;
  wire [63:0] Queue_3_io_enq_bits_data;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [2:0] Queue_3_io_deq_bits_opcode;
  wire [2:0] Queue_3_io_deq_bits_param;
  wire [3:0] Queue_3_io_deq_bits_size;
  wire [3:0] Queue_3_io_deq_bits_source;
  wire [31:0] Queue_3_io_deq_bits_address;
  wire [63:0] Queue_3_io_deq_bits_data;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [2:0] Queue_4_io_enq_bits_sink;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [2:0] Queue_4_io_deq_bits_sink;
  Queue_27 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_28 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  Queue_29 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_param(Queue_2_io_enq_bits_param),
    .io_enq_bits_size(Queue_2_io_enq_bits_size),
    .io_enq_bits_source(Queue_2_io_enq_bits_source),
    .io_enq_bits_address(Queue_2_io_enq_bits_address),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_param(Queue_2_io_deq_bits_param),
    .io_deq_bits_size(Queue_2_io_deq_bits_size),
    .io_deq_bits_source(Queue_2_io_deq_bits_source),
    .io_deq_bits_address(Queue_2_io_deq_bits_address)
  );
  Queue_30 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_opcode(Queue_3_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_3_io_enq_bits_param),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_source(Queue_3_io_enq_bits_source),
    .io_enq_bits_address(Queue_3_io_enq_bits_address),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_opcode(Queue_3_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_3_io_deq_bits_param),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_source(Queue_3_io_deq_bits_source),
    .io_deq_bits_address(Queue_3_io_deq_bits_address),
    .io_deq_bits_data(Queue_3_io_deq_bits_data)
  );
  Queue_31 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_sink(Queue_4_io_enq_bits_sink),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_sink(Queue_4_io_deq_bits_sink)
  );
  assign auto_in_a_ready = _T_31_a_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_param = _T_31_b_bits_param;
  assign auto_in_b_bits_size = _T_31_b_bits_size;
  assign auto_in_b_bits_source = _T_31_b_bits_source;
  assign auto_in_b_bits_address = _T_31_b_bits_address;
  assign auto_in_c_ready = _T_31_c_ready;
  assign auto_in_d_valid = _T_31_d_valid;
  assign auto_in_d_bits_opcode = _T_31_d_bits_opcode;
  assign auto_in_d_bits_param = _T_31_d_bits_param;
  assign auto_in_d_bits_size = _T_31_d_bits_size;
  assign auto_in_d_bits_source = _T_31_d_bits_source;
  assign auto_in_d_bits_sink = _T_31_d_bits_sink;
  assign auto_in_d_bits_data = _T_31_d_bits_data;
  assign auto_in_d_bits_error = _T_31_d_bits_error;
  assign auto_in_e_ready = _T_31_e_ready;
  assign auto_out_a_valid = _T_89_a_valid;
  assign auto_out_a_bits_opcode = _T_89_a_bits_opcode;
  assign auto_out_a_bits_param = _T_89_a_bits_param;
  assign auto_out_a_bits_size = _T_89_a_bits_size;
  assign auto_out_a_bits_source = _T_89_a_bits_source;
  assign auto_out_a_bits_address = _T_89_a_bits_address;
  assign auto_out_a_bits_mask = _T_89_a_bits_mask;
  assign auto_out_a_bits_data = _T_89_a_bits_data;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_c_valid = _T_89_c_valid;
  assign auto_out_c_bits_opcode = _T_89_c_bits_opcode;
  assign auto_out_c_bits_param = _T_89_c_bits_param;
  assign auto_out_c_bits_size = _T_89_c_bits_size;
  assign auto_out_c_bits_source = _T_89_c_bits_source;
  assign auto_out_c_bits_address = _T_89_c_bits_address;
  assign auto_out_c_bits_data = _T_89_c_bits_data;
  assign auto_out_d_ready = _T_89_d_ready;
  assign auto_out_e_valid = _T_89_e_valid;
  assign auto_out_e_bits_sink = _T_89_e_bits_sink;
  assign _T_31_a_ready = Queue_io_enq_ready;
  assign _T_31_a_valid = auto_in_a_valid;
  assign _T_31_a_bits_opcode = auto_in_a_bits_opcode;
  assign _T_31_a_bits_param = auto_in_a_bits_param;
  assign _T_31_a_bits_size = auto_in_a_bits_size;
  assign _T_31_a_bits_source = auto_in_a_bits_source;
  assign _T_31_a_bits_address = auto_in_a_bits_address;
  assign _T_31_a_bits_mask = auto_in_a_bits_mask;
  assign _T_31_a_bits_data = auto_in_a_bits_data;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = Queue_2_io_deq_valid;
  assign _T_31_b_bits_param = Queue_2_io_deq_bits_param;
  assign _T_31_b_bits_size = Queue_2_io_deq_bits_size;
  assign _T_31_b_bits_source = Queue_2_io_deq_bits_source;
  assign _T_31_b_bits_address = Queue_2_io_deq_bits_address;
  assign _T_31_c_ready = Queue_3_io_enq_ready;
  assign _T_31_c_valid = auto_in_c_valid;
  assign _T_31_c_bits_opcode = auto_in_c_bits_opcode;
  assign _T_31_c_bits_param = auto_in_c_bits_param;
  assign _T_31_c_bits_size = auto_in_c_bits_size;
  assign _T_31_c_bits_source = auto_in_c_bits_source;
  assign _T_31_c_bits_address = auto_in_c_bits_address;
  assign _T_31_c_bits_data = auto_in_c_bits_data;
  assign _T_31_d_ready = auto_in_d_ready;
  assign _T_31_d_valid = Queue_1_io_deq_valid;
  assign _T_31_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign _T_31_d_bits_param = Queue_1_io_deq_bits_param;
  assign _T_31_d_bits_size = Queue_1_io_deq_bits_size;
  assign _T_31_d_bits_source = Queue_1_io_deq_bits_source;
  assign _T_31_d_bits_sink = Queue_1_io_deq_bits_sink;
  assign _T_31_d_bits_data = Queue_1_io_deq_bits_data;
  assign _T_31_d_bits_error = Queue_1_io_deq_bits_error;
  assign _T_31_e_ready = Queue_4_io_enq_ready;
  assign _T_31_e_valid = auto_in_e_valid;
  assign _T_31_e_bits_sink = auto_in_e_bits_sink;
  assign _T_89_a_ready = auto_out_a_ready;
  assign _T_89_a_valid = Queue_io_deq_valid;
  assign _T_89_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign _T_89_a_bits_param = Queue_io_deq_bits_param;
  assign _T_89_a_bits_size = Queue_io_deq_bits_size;
  assign _T_89_a_bits_source = Queue_io_deq_bits_source;
  assign _T_89_a_bits_address = Queue_io_deq_bits_address;
  assign _T_89_a_bits_mask = Queue_io_deq_bits_mask;
  assign _T_89_a_bits_data = Queue_io_deq_bits_data;
  assign _T_89_b_ready = Queue_2_io_enq_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_param = auto_out_b_bits_param;
  assign _T_89_b_bits_size = auto_out_b_bits_size;
  assign _T_89_b_bits_source = auto_out_b_bits_source;
  assign _T_89_b_bits_address = auto_out_b_bits_address;
  assign _T_89_c_ready = auto_out_c_ready;
  assign _T_89_c_valid = Queue_3_io_deq_valid;
  assign _T_89_c_bits_opcode = Queue_3_io_deq_bits_opcode;
  assign _T_89_c_bits_param = Queue_3_io_deq_bits_param;
  assign _T_89_c_bits_size = Queue_3_io_deq_bits_size;
  assign _T_89_c_bits_source = Queue_3_io_deq_bits_source;
  assign _T_89_c_bits_address = Queue_3_io_deq_bits_address;
  assign _T_89_c_bits_data = Queue_3_io_deq_bits_data;
  assign _T_89_d_ready = Queue_1_io_enq_ready;
  assign _T_89_d_valid = auto_out_d_valid;
  assign _T_89_d_bits_opcode = auto_out_d_bits_opcode;
  assign _T_89_d_bits_param = auto_out_d_bits_param;
  assign _T_89_d_bits_size = auto_out_d_bits_size;
  assign _T_89_d_bits_source = auto_out_d_bits_source;
  assign _T_89_d_bits_sink = auto_out_d_bits_sink;
  assign _T_89_d_bits_data = auto_out_d_bits_data;
  assign _T_89_d_bits_error = auto_out_d_bits_error;
  assign _T_89_e_ready = auto_out_e_ready;
  assign _T_89_e_valid = Queue_4_io_deq_valid;
  assign _T_89_e_bits_sink = Queue_4_io_deq_bits_sink;
  assign Queue_io_enq_valid = _T_31_a_valid;
  assign Queue_io_enq_bits_opcode = _T_31_a_bits_opcode;
  assign Queue_io_enq_bits_param = _T_31_a_bits_param;
  assign Queue_io_enq_bits_size = _T_31_a_bits_size;
  assign Queue_io_enq_bits_source = _T_31_a_bits_source;
  assign Queue_io_enq_bits_address = _T_31_a_bits_address;
  assign Queue_io_enq_bits_mask = _T_31_a_bits_mask;
  assign Queue_io_enq_bits_data = _T_31_a_bits_data;
  assign Queue_io_deq_ready = _T_89_a_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_89_d_valid;
  assign Queue_1_io_enq_bits_opcode = _T_89_d_bits_opcode;
  assign Queue_1_io_enq_bits_param = _T_89_d_bits_param;
  assign Queue_1_io_enq_bits_size = _T_89_d_bits_size;
  assign Queue_1_io_enq_bits_source = _T_89_d_bits_source;
  assign Queue_1_io_enq_bits_sink = _T_89_d_bits_sink;
  assign Queue_1_io_enq_bits_data = _T_89_d_bits_data;
  assign Queue_1_io_enq_bits_error = _T_89_d_bits_error;
  assign Queue_1_io_deq_ready = _T_31_d_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_2_io_enq_valid = _T_89_b_valid;
  assign Queue_2_io_enq_bits_param = _T_89_b_bits_param;
  assign Queue_2_io_enq_bits_size = _T_89_b_bits_size;
  assign Queue_2_io_enq_bits_source = _T_89_b_bits_source;
  assign Queue_2_io_enq_bits_address = _T_89_b_bits_address;
  assign Queue_2_io_deq_ready = _T_31_b_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_3_io_enq_valid = _T_31_c_valid;
  assign Queue_3_io_enq_bits_opcode = _T_31_c_bits_opcode;
  assign Queue_3_io_enq_bits_param = _T_31_c_bits_param;
  assign Queue_3_io_enq_bits_size = _T_31_c_bits_size;
  assign Queue_3_io_enq_bits_source = _T_31_c_bits_source;
  assign Queue_3_io_enq_bits_address = _T_31_c_bits_address;
  assign Queue_3_io_enq_bits_data = _T_31_c_bits_data;
  assign Queue_3_io_deq_ready = _T_89_c_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_4_io_enq_valid = _T_31_e_valid;
  assign Queue_4_io_enq_bits_sink = _T_31_e_bits_sink;
  assign Queue_4_io_deq_ready = _T_89_e_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
endmodule
module SynchronizerShiftReg_w1_d3(
  input   clock,
  input   io_d,
  output  io_q
);
  reg  sync_0;
  reg [31:0] _RAND_0;
  reg  sync_1;
  reg [31:0] _RAND_1;
  reg  sync_2;
  reg [31:0] _RAND_2;
  assign io_q = sync_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  sync_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  sync_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  sync_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= sync_1;
    sync_1 <= sync_2;
    sync_2 <= io_d;
  end
endmodule
module IntSyncCrossingSink(
  input   clock,
  input   auto_in_sync_0,
  output  auto_out_0
);
  wire  _T_5_sync_0;
  wire  _T_11_0;
  wire  SynchronizerShiftReg_w1_d3_clock;
  wire  SynchronizerShiftReg_w1_d3_io_d;
  wire  SynchronizerShiftReg_w1_d3_io_q;
  wire  _T_29_0;
  wire  _T_36;
  SynchronizerShiftReg_w1_d3 SynchronizerShiftReg_w1_d3 (
    .clock(SynchronizerShiftReg_w1_d3_clock),
    .io_d(SynchronizerShiftReg_w1_d3_io_d),
    .io_q(SynchronizerShiftReg_w1_d3_io_q)
  );
  assign auto_out_0 = _T_11_0;
  assign _T_5_sync_0 = auto_in_sync_0;
  assign _T_11_0 = _T_29_0;
  assign SynchronizerShiftReg_w1_d3_io_d = _T_5_sync_0;
  assign SynchronizerShiftReg_w1_d3_clock = clock;
  assign _T_29_0 = _T_36;
  assign _T_36 = SynchronizerShiftReg_w1_d3_io_q;
endmodule
module IntSyncCrossingSink_1(
  input   auto_in_2_sync_0,
  input   auto_in_1_sync_0,
  input   auto_in_0_sync_0,
  input   auto_in_0_sync_1,
  output  auto_out_2_0,
  output  auto_out_1_0,
  output  auto_out_0_0,
  output  auto_out_0_1
);
  wire  _T_5_sync_0;
  wire  _T_5_sync_1;
  wire  _T_11_sync_0;
  wire  _T_17_sync_0;
  wire  _T_23_0;
  wire  _T_23_1;
  wire  _T_31_0;
  wire  _T_38_0;
  assign auto_out_2_0 = _T_38_0;
  assign auto_out_1_0 = _T_31_0;
  assign auto_out_0_0 = _T_23_0;
  assign auto_out_0_1 = _T_23_1;
  assign _T_5_sync_0 = auto_in_0_sync_0;
  assign _T_5_sync_1 = auto_in_0_sync_1;
  assign _T_11_sync_0 = auto_in_1_sync_0;
  assign _T_17_sync_0 = auto_in_2_sync_0;
  assign _T_23_0 = _T_5_sync_0;
  assign _T_23_1 = _T_5_sync_1;
  assign _T_31_0 = _T_11_sync_0;
  assign _T_38_0 = _T_17_sync_0;
endmodule
module BoomTileWrapper_tile(
  input         clock,
  input         reset,
  input         auto_anon_in_3_sync_0,
  input         auto_anon_in_2_sync_0,
  input         auto_anon_in_1_sync_0,
  input         auto_anon_in_1_sync_1,
  input         auto_anon_in_0_sync_0,
  input         auto_anon_out_a_ready,
  output        auto_anon_out_a_valid,
  output [2:0]  auto_anon_out_a_bits_opcode,
  output [2:0]  auto_anon_out_a_bits_param,
  output [3:0]  auto_anon_out_a_bits_size,
  output [3:0]  auto_anon_out_a_bits_source,
  output [31:0] auto_anon_out_a_bits_address,
  output [7:0]  auto_anon_out_a_bits_mask,
  output [63:0] auto_anon_out_a_bits_data,
  output        auto_anon_out_b_ready,
  input         auto_anon_out_b_valid,
  input  [1:0]  auto_anon_out_b_bits_param,
  input  [3:0]  auto_anon_out_b_bits_size,
  input  [3:0]  auto_anon_out_b_bits_source,
  input  [31:0] auto_anon_out_b_bits_address,
  input         auto_anon_out_c_ready,
  output        auto_anon_out_c_valid,
  output [2:0]  auto_anon_out_c_bits_opcode,
  output [2:0]  auto_anon_out_c_bits_param,
  output [3:0]  auto_anon_out_c_bits_size,
  output [3:0]  auto_anon_out_c_bits_source,
  output [31:0] auto_anon_out_c_bits_address,
  output [63:0] auto_anon_out_c_bits_data,
  output        auto_anon_out_d_ready,
  input         auto_anon_out_d_valid,
  input  [2:0]  auto_anon_out_d_bits_opcode,
  input  [1:0]  auto_anon_out_d_bits_param,
  input  [3:0]  auto_anon_out_d_bits_size,
  input  [3:0]  auto_anon_out_d_bits_source,
  input  [2:0]  auto_anon_out_d_bits_sink,
  input  [63:0] auto_anon_out_d_bits_data,
  input         auto_anon_out_d_bits_error,
  input         auto_anon_out_e_ready,
  output        auto_anon_out_e_valid,
  output [2:0]  auto_anon_out_e_bits_sink
);
  wire  boom_clock;
  wire  boom_reset;
  wire  boom_auto_master_out_a_ready;
  wire  boom_auto_master_out_a_valid;
  wire [2:0] boom_auto_master_out_a_bits_opcode;
  wire [2:0] boom_auto_master_out_a_bits_param;
  wire [3:0] boom_auto_master_out_a_bits_size;
  wire [3:0] boom_auto_master_out_a_bits_source;
  wire [31:0] boom_auto_master_out_a_bits_address;
  wire [7:0] boom_auto_master_out_a_bits_mask;
  wire [63:0] boom_auto_master_out_a_bits_data;
  wire  boom_auto_master_out_b_ready;
  wire  boom_auto_master_out_b_valid;
  wire [1:0] boom_auto_master_out_b_bits_param;
  wire [3:0] boom_auto_master_out_b_bits_size;
  wire [3:0] boom_auto_master_out_b_bits_source;
  wire [31:0] boom_auto_master_out_b_bits_address;
  wire  boom_auto_master_out_c_ready;
  wire  boom_auto_master_out_c_valid;
  wire [2:0] boom_auto_master_out_c_bits_opcode;
  wire [2:0] boom_auto_master_out_c_bits_param;
  wire [3:0] boom_auto_master_out_c_bits_size;
  wire [3:0] boom_auto_master_out_c_bits_source;
  wire [31:0] boom_auto_master_out_c_bits_address;
  wire [63:0] boom_auto_master_out_c_bits_data;
  wire  boom_auto_master_out_d_ready;
  wire  boom_auto_master_out_d_valid;
  wire [2:0] boom_auto_master_out_d_bits_opcode;
  wire [1:0] boom_auto_master_out_d_bits_param;
  wire [3:0] boom_auto_master_out_d_bits_size;
  wire [3:0] boom_auto_master_out_d_bits_source;
  wire [2:0] boom_auto_master_out_d_bits_sink;
  wire [63:0] boom_auto_master_out_d_bits_data;
  wire  boom_auto_master_out_d_bits_error;
  wire  boom_auto_master_out_e_ready;
  wire  boom_auto_master_out_e_valid;
  wire [2:0] boom_auto_master_out_e_bits_sink;
  wire  boom_auto_int_in_0;
  wire  boom_auto_int_in_1;
  wire  boom_auto_int_in_2;
  wire  boom_auto_int_in_3;
  wire  boom_auto_int_in_4;
  wire  intXbar_auto_int_in_3_0;
  wire  intXbar_auto_int_in_2_0;
  wire  intXbar_auto_int_in_1_0;
  wire  intXbar_auto_int_in_1_1;
  wire  intXbar_auto_int_in_0_0;
  wire  intXbar_auto_int_out_0;
  wire  intXbar_auto_int_out_1;
  wire  intXbar_auto_int_out_2;
  wire  intXbar_auto_int_out_3;
  wire  intXbar_auto_int_out_4;
  wire  SystemBus_TLBuffer_clock;
  wire  SystemBus_TLBuffer_reset;
  wire  SystemBus_TLBuffer_auto_in_a_ready;
  wire  SystemBus_TLBuffer_auto_in_a_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_a_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_in_a_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_in_a_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_a_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_in_a_bits_address;
  wire [7:0] SystemBus_TLBuffer_auto_in_a_bits_mask;
  wire [63:0] SystemBus_TLBuffer_auto_in_a_bits_data;
  wire  SystemBus_TLBuffer_auto_in_b_ready;
  wire  SystemBus_TLBuffer_auto_in_b_valid;
  wire [1:0] SystemBus_TLBuffer_auto_in_b_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_in_b_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_b_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_in_b_bits_address;
  wire  SystemBus_TLBuffer_auto_in_c_ready;
  wire  SystemBus_TLBuffer_auto_in_c_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_c_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_in_c_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_in_c_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_c_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_in_c_bits_address;
  wire [63:0] SystemBus_TLBuffer_auto_in_c_bits_data;
  wire  SystemBus_TLBuffer_auto_in_d_ready;
  wire  SystemBus_TLBuffer_auto_in_d_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_d_bits_opcode;
  wire [1:0] SystemBus_TLBuffer_auto_in_d_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_in_d_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_d_bits_source;
  wire [2:0] SystemBus_TLBuffer_auto_in_d_bits_sink;
  wire [63:0] SystemBus_TLBuffer_auto_in_d_bits_data;
  wire  SystemBus_TLBuffer_auto_in_d_bits_error;
  wire  SystemBus_TLBuffer_auto_in_e_ready;
  wire  SystemBus_TLBuffer_auto_in_e_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_e_bits_sink;
  wire  SystemBus_TLBuffer_auto_out_a_ready;
  wire  SystemBus_TLBuffer_auto_out_a_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_a_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_out_a_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_a_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_a_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_out_a_bits_address;
  wire [7:0] SystemBus_TLBuffer_auto_out_a_bits_mask;
  wire [63:0] SystemBus_TLBuffer_auto_out_a_bits_data;
  wire  SystemBus_TLBuffer_auto_out_b_ready;
  wire  SystemBus_TLBuffer_auto_out_b_valid;
  wire [1:0] SystemBus_TLBuffer_auto_out_b_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_b_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_b_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_out_b_bits_address;
  wire  SystemBus_TLBuffer_auto_out_c_ready;
  wire  SystemBus_TLBuffer_auto_out_c_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_c_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_out_c_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_c_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_c_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_out_c_bits_address;
  wire [63:0] SystemBus_TLBuffer_auto_out_c_bits_data;
  wire  SystemBus_TLBuffer_auto_out_d_ready;
  wire  SystemBus_TLBuffer_auto_out_d_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_d_bits_opcode;
  wire [1:0] SystemBus_TLBuffer_auto_out_d_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_d_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_d_bits_source;
  wire [2:0] SystemBus_TLBuffer_auto_out_d_bits_sink;
  wire [63:0] SystemBus_TLBuffer_auto_out_d_bits_data;
  wire  SystemBus_TLBuffer_auto_out_d_bits_error;
  wire  SystemBus_TLBuffer_auto_out_e_ready;
  wire  SystemBus_TLBuffer_auto_out_e_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_e_bits_sink;
  wire  IntSyncCrossingSink_clock;
  wire  IntSyncCrossingSink_auto_in_sync_0;
  wire  IntSyncCrossingSink_auto_out_0;
  wire  IntSyncCrossingSink_1_auto_in_2_sync_0;
  wire  IntSyncCrossingSink_1_auto_in_1_sync_0;
  wire  IntSyncCrossingSink_1_auto_in_0_sync_0;
  wire  IntSyncCrossingSink_1_auto_in_0_sync_1;
  wire  IntSyncCrossingSink_1_auto_out_2_0;
  wire  IntSyncCrossingSink_1_auto_out_1_0;
  wire  IntSyncCrossingSink_1_auto_out_0_0;
  wire  IntSyncCrossingSink_1_auto_out_0_1;
  BoomTile_boom boom (
    .clock(boom_clock),
    .reset(boom_reset),
    .auto_master_out_a_ready(boom_auto_master_out_a_ready),
    .auto_master_out_a_valid(boom_auto_master_out_a_valid),
    .auto_master_out_a_bits_opcode(boom_auto_master_out_a_bits_opcode),
    .auto_master_out_a_bits_param(boom_auto_master_out_a_bits_param),
    .auto_master_out_a_bits_size(boom_auto_master_out_a_bits_size),
    .auto_master_out_a_bits_source(boom_auto_master_out_a_bits_source),
    .auto_master_out_a_bits_address(boom_auto_master_out_a_bits_address),
    .auto_master_out_a_bits_mask(boom_auto_master_out_a_bits_mask),
    .auto_master_out_a_bits_data(boom_auto_master_out_a_bits_data),
    .auto_master_out_b_ready(boom_auto_master_out_b_ready),
    .auto_master_out_b_valid(boom_auto_master_out_b_valid),
    .auto_master_out_b_bits_param(boom_auto_master_out_b_bits_param),
    .auto_master_out_b_bits_size(boom_auto_master_out_b_bits_size),
    .auto_master_out_b_bits_source(boom_auto_master_out_b_bits_source),
    .auto_master_out_b_bits_address(boom_auto_master_out_b_bits_address),
    .auto_master_out_c_ready(boom_auto_master_out_c_ready),
    .auto_master_out_c_valid(boom_auto_master_out_c_valid),
    .auto_master_out_c_bits_opcode(boom_auto_master_out_c_bits_opcode),
    .auto_master_out_c_bits_param(boom_auto_master_out_c_bits_param),
    .auto_master_out_c_bits_size(boom_auto_master_out_c_bits_size),
    .auto_master_out_c_bits_source(boom_auto_master_out_c_bits_source),
    .auto_master_out_c_bits_address(boom_auto_master_out_c_bits_address),
    .auto_master_out_c_bits_data(boom_auto_master_out_c_bits_data),
    .auto_master_out_d_ready(boom_auto_master_out_d_ready),
    .auto_master_out_d_valid(boom_auto_master_out_d_valid),
    .auto_master_out_d_bits_opcode(boom_auto_master_out_d_bits_opcode),
    .auto_master_out_d_bits_param(boom_auto_master_out_d_bits_param),
    .auto_master_out_d_bits_size(boom_auto_master_out_d_bits_size),
    .auto_master_out_d_bits_source(boom_auto_master_out_d_bits_source),
    .auto_master_out_d_bits_sink(boom_auto_master_out_d_bits_sink),
    .auto_master_out_d_bits_data(boom_auto_master_out_d_bits_data),
    .auto_master_out_d_bits_error(boom_auto_master_out_d_bits_error),
    .auto_master_out_e_ready(boom_auto_master_out_e_ready),
    .auto_master_out_e_valid(boom_auto_master_out_e_valid),
    .auto_master_out_e_bits_sink(boom_auto_master_out_e_bits_sink),
    .auto_int_in_0(boom_auto_int_in_0),
    .auto_int_in_1(boom_auto_int_in_1),
    .auto_int_in_2(boom_auto_int_in_2),
    .auto_int_in_3(boom_auto_int_in_3),
    .auto_int_in_4(boom_auto_int_in_4)
  );
  IntXbar_intXbar intXbar (
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_in_0_0(intXbar_auto_int_in_0_0),
    .auto_int_out_0(intXbar_auto_int_out_0),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4)
  );
  TLBuffer_SystemBus SystemBus_TLBuffer (
    .clock(SystemBus_TLBuffer_clock),
    .reset(SystemBus_TLBuffer_reset),
    .auto_in_a_ready(SystemBus_TLBuffer_auto_in_a_ready),
    .auto_in_a_valid(SystemBus_TLBuffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(SystemBus_TLBuffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(SystemBus_TLBuffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(SystemBus_TLBuffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(SystemBus_TLBuffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(SystemBus_TLBuffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(SystemBus_TLBuffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(SystemBus_TLBuffer_auto_in_a_bits_data),
    .auto_in_b_ready(SystemBus_TLBuffer_auto_in_b_ready),
    .auto_in_b_valid(SystemBus_TLBuffer_auto_in_b_valid),
    .auto_in_b_bits_param(SystemBus_TLBuffer_auto_in_b_bits_param),
    .auto_in_b_bits_size(SystemBus_TLBuffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(SystemBus_TLBuffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(SystemBus_TLBuffer_auto_in_b_bits_address),
    .auto_in_c_ready(SystemBus_TLBuffer_auto_in_c_ready),
    .auto_in_c_valid(SystemBus_TLBuffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(SystemBus_TLBuffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(SystemBus_TLBuffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(SystemBus_TLBuffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(SystemBus_TLBuffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(SystemBus_TLBuffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(SystemBus_TLBuffer_auto_in_c_bits_data),
    .auto_in_d_ready(SystemBus_TLBuffer_auto_in_d_ready),
    .auto_in_d_valid(SystemBus_TLBuffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(SystemBus_TLBuffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(SystemBus_TLBuffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(SystemBus_TLBuffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(SystemBus_TLBuffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(SystemBus_TLBuffer_auto_in_d_bits_sink),
    .auto_in_d_bits_data(SystemBus_TLBuffer_auto_in_d_bits_data),
    .auto_in_d_bits_error(SystemBus_TLBuffer_auto_in_d_bits_error),
    .auto_in_e_ready(SystemBus_TLBuffer_auto_in_e_ready),
    .auto_in_e_valid(SystemBus_TLBuffer_auto_in_e_valid),
    .auto_in_e_bits_sink(SystemBus_TLBuffer_auto_in_e_bits_sink),
    .auto_out_a_ready(SystemBus_TLBuffer_auto_out_a_ready),
    .auto_out_a_valid(SystemBus_TLBuffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(SystemBus_TLBuffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(SystemBus_TLBuffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(SystemBus_TLBuffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(SystemBus_TLBuffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(SystemBus_TLBuffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(SystemBus_TLBuffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(SystemBus_TLBuffer_auto_out_a_bits_data),
    .auto_out_b_ready(SystemBus_TLBuffer_auto_out_b_ready),
    .auto_out_b_valid(SystemBus_TLBuffer_auto_out_b_valid),
    .auto_out_b_bits_param(SystemBus_TLBuffer_auto_out_b_bits_param),
    .auto_out_b_bits_size(SystemBus_TLBuffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(SystemBus_TLBuffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(SystemBus_TLBuffer_auto_out_b_bits_address),
    .auto_out_c_ready(SystemBus_TLBuffer_auto_out_c_ready),
    .auto_out_c_valid(SystemBus_TLBuffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(SystemBus_TLBuffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(SystemBus_TLBuffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(SystemBus_TLBuffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(SystemBus_TLBuffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(SystemBus_TLBuffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(SystemBus_TLBuffer_auto_out_c_bits_data),
    .auto_out_d_ready(SystemBus_TLBuffer_auto_out_d_ready),
    .auto_out_d_valid(SystemBus_TLBuffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(SystemBus_TLBuffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(SystemBus_TLBuffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(SystemBus_TLBuffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(SystemBus_TLBuffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(SystemBus_TLBuffer_auto_out_d_bits_sink),
    .auto_out_d_bits_data(SystemBus_TLBuffer_auto_out_d_bits_data),
    .auto_out_d_bits_error(SystemBus_TLBuffer_auto_out_d_bits_error),
    .auto_out_e_ready(SystemBus_TLBuffer_auto_out_e_ready),
    .auto_out_e_valid(SystemBus_TLBuffer_auto_out_e_valid),
    .auto_out_e_bits_sink(SystemBus_TLBuffer_auto_out_e_bits_sink)
  );
  IntSyncCrossingSink IntSyncCrossingSink (
    .clock(IntSyncCrossingSink_clock),
    .auto_in_sync_0(IntSyncCrossingSink_auto_in_sync_0),
    .auto_out_0(IntSyncCrossingSink_auto_out_0)
  );
  IntSyncCrossingSink_1 IntSyncCrossingSink_1 (
    .auto_in_2_sync_0(IntSyncCrossingSink_1_auto_in_2_sync_0),
    .auto_in_1_sync_0(IntSyncCrossingSink_1_auto_in_1_sync_0),
    .auto_in_0_sync_0(IntSyncCrossingSink_1_auto_in_0_sync_0),
    .auto_in_0_sync_1(IntSyncCrossingSink_1_auto_in_0_sync_1),
    .auto_out_2_0(IntSyncCrossingSink_1_auto_out_2_0),
    .auto_out_1_0(IntSyncCrossingSink_1_auto_out_1_0),
    .auto_out_0_0(IntSyncCrossingSink_1_auto_out_0_0),
    .auto_out_0_1(IntSyncCrossingSink_1_auto_out_0_1)
  );
  assign auto_anon_out_a_valid = SystemBus_TLBuffer_auto_out_a_valid;
  assign auto_anon_out_a_bits_opcode = SystemBus_TLBuffer_auto_out_a_bits_opcode;
  assign auto_anon_out_a_bits_param = SystemBus_TLBuffer_auto_out_a_bits_param;
  assign auto_anon_out_a_bits_size = SystemBus_TLBuffer_auto_out_a_bits_size;
  assign auto_anon_out_a_bits_source = SystemBus_TLBuffer_auto_out_a_bits_source;
  assign auto_anon_out_a_bits_address = SystemBus_TLBuffer_auto_out_a_bits_address;
  assign auto_anon_out_a_bits_mask = SystemBus_TLBuffer_auto_out_a_bits_mask;
  assign auto_anon_out_a_bits_data = SystemBus_TLBuffer_auto_out_a_bits_data;
  assign auto_anon_out_b_ready = SystemBus_TLBuffer_auto_out_b_ready;
  assign auto_anon_out_c_valid = SystemBus_TLBuffer_auto_out_c_valid;
  assign auto_anon_out_c_bits_opcode = SystemBus_TLBuffer_auto_out_c_bits_opcode;
  assign auto_anon_out_c_bits_param = SystemBus_TLBuffer_auto_out_c_bits_param;
  assign auto_anon_out_c_bits_size = SystemBus_TLBuffer_auto_out_c_bits_size;
  assign auto_anon_out_c_bits_source = SystemBus_TLBuffer_auto_out_c_bits_source;
  assign auto_anon_out_c_bits_address = SystemBus_TLBuffer_auto_out_c_bits_address;
  assign auto_anon_out_c_bits_data = SystemBus_TLBuffer_auto_out_c_bits_data;
  assign auto_anon_out_d_ready = SystemBus_TLBuffer_auto_out_d_ready;
  assign auto_anon_out_e_valid = SystemBus_TLBuffer_auto_out_e_valid;
  assign auto_anon_out_e_bits_sink = SystemBus_TLBuffer_auto_out_e_bits_sink;
  assign boom_clock = clock;
  assign boom_reset = reset;
  assign boom_auto_master_out_a_ready = SystemBus_TLBuffer_auto_in_a_ready;
  assign boom_auto_master_out_b_valid = SystemBus_TLBuffer_auto_in_b_valid;
  assign boom_auto_master_out_b_bits_param = SystemBus_TLBuffer_auto_in_b_bits_param;
  assign boom_auto_master_out_b_bits_size = SystemBus_TLBuffer_auto_in_b_bits_size;
  assign boom_auto_master_out_b_bits_source = SystemBus_TLBuffer_auto_in_b_bits_source;
  assign boom_auto_master_out_b_bits_address = SystemBus_TLBuffer_auto_in_b_bits_address;
  assign boom_auto_master_out_c_ready = SystemBus_TLBuffer_auto_in_c_ready;
  assign boom_auto_master_out_d_valid = SystemBus_TLBuffer_auto_in_d_valid;
  assign boom_auto_master_out_d_bits_opcode = SystemBus_TLBuffer_auto_in_d_bits_opcode;
  assign boom_auto_master_out_d_bits_param = SystemBus_TLBuffer_auto_in_d_bits_param;
  assign boom_auto_master_out_d_bits_size = SystemBus_TLBuffer_auto_in_d_bits_size;
  assign boom_auto_master_out_d_bits_source = SystemBus_TLBuffer_auto_in_d_bits_source;
  assign boom_auto_master_out_d_bits_sink = SystemBus_TLBuffer_auto_in_d_bits_sink;
  assign boom_auto_master_out_d_bits_data = SystemBus_TLBuffer_auto_in_d_bits_data;
  assign boom_auto_master_out_d_bits_error = SystemBus_TLBuffer_auto_in_d_bits_error;
  assign boom_auto_master_out_e_ready = SystemBus_TLBuffer_auto_in_e_ready;
  assign boom_auto_int_in_0 = intXbar_auto_int_out_0;
  assign boom_auto_int_in_1 = intXbar_auto_int_out_1;
  assign boom_auto_int_in_2 = intXbar_auto_int_out_2;
  assign boom_auto_int_in_3 = intXbar_auto_int_out_3;
  assign boom_auto_int_in_4 = intXbar_auto_int_out_4;
  assign intXbar_auto_int_in_3_0 = IntSyncCrossingSink_1_auto_out_2_0;
  assign intXbar_auto_int_in_2_0 = IntSyncCrossingSink_1_auto_out_1_0;
  assign intXbar_auto_int_in_1_0 = IntSyncCrossingSink_1_auto_out_0_0;
  assign intXbar_auto_int_in_1_1 = IntSyncCrossingSink_1_auto_out_0_1;
  assign intXbar_auto_int_in_0_0 = IntSyncCrossingSink_auto_out_0;
  assign SystemBus_TLBuffer_clock = clock;
  assign SystemBus_TLBuffer_reset = reset;
  assign SystemBus_TLBuffer_auto_in_a_valid = boom_auto_master_out_a_valid;
  assign SystemBus_TLBuffer_auto_in_a_bits_opcode = boom_auto_master_out_a_bits_opcode;
  assign SystemBus_TLBuffer_auto_in_a_bits_param = boom_auto_master_out_a_bits_param;
  assign SystemBus_TLBuffer_auto_in_a_bits_size = boom_auto_master_out_a_bits_size;
  assign SystemBus_TLBuffer_auto_in_a_bits_source = boom_auto_master_out_a_bits_source;
  assign SystemBus_TLBuffer_auto_in_a_bits_address = boom_auto_master_out_a_bits_address;
  assign SystemBus_TLBuffer_auto_in_a_bits_mask = boom_auto_master_out_a_bits_mask;
  assign SystemBus_TLBuffer_auto_in_a_bits_data = boom_auto_master_out_a_bits_data;
  assign SystemBus_TLBuffer_auto_in_b_ready = boom_auto_master_out_b_ready;
  assign SystemBus_TLBuffer_auto_in_c_valid = boom_auto_master_out_c_valid;
  assign SystemBus_TLBuffer_auto_in_c_bits_opcode = boom_auto_master_out_c_bits_opcode;
  assign SystemBus_TLBuffer_auto_in_c_bits_param = boom_auto_master_out_c_bits_param;
  assign SystemBus_TLBuffer_auto_in_c_bits_size = boom_auto_master_out_c_bits_size;
  assign SystemBus_TLBuffer_auto_in_c_bits_source = boom_auto_master_out_c_bits_source;
  assign SystemBus_TLBuffer_auto_in_c_bits_address = boom_auto_master_out_c_bits_address;
  assign SystemBus_TLBuffer_auto_in_c_bits_data = boom_auto_master_out_c_bits_data;
  assign SystemBus_TLBuffer_auto_in_d_ready = boom_auto_master_out_d_ready;
  assign SystemBus_TLBuffer_auto_in_e_valid = boom_auto_master_out_e_valid;
  assign SystemBus_TLBuffer_auto_in_e_bits_sink = boom_auto_master_out_e_bits_sink;
  assign SystemBus_TLBuffer_auto_out_a_ready = auto_anon_out_a_ready;
  assign SystemBus_TLBuffer_auto_out_b_valid = auto_anon_out_b_valid;
  assign SystemBus_TLBuffer_auto_out_b_bits_param = auto_anon_out_b_bits_param;
  assign SystemBus_TLBuffer_auto_out_b_bits_size = auto_anon_out_b_bits_size;
  assign SystemBus_TLBuffer_auto_out_b_bits_source = auto_anon_out_b_bits_source;
  assign SystemBus_TLBuffer_auto_out_b_bits_address = auto_anon_out_b_bits_address;
  assign SystemBus_TLBuffer_auto_out_c_ready = auto_anon_out_c_ready;
  assign SystemBus_TLBuffer_auto_out_d_valid = auto_anon_out_d_valid;
  assign SystemBus_TLBuffer_auto_out_d_bits_opcode = auto_anon_out_d_bits_opcode;
  assign SystemBus_TLBuffer_auto_out_d_bits_param = auto_anon_out_d_bits_param;
  assign SystemBus_TLBuffer_auto_out_d_bits_size = auto_anon_out_d_bits_size;
  assign SystemBus_TLBuffer_auto_out_d_bits_source = auto_anon_out_d_bits_source;
  assign SystemBus_TLBuffer_auto_out_d_bits_sink = auto_anon_out_d_bits_sink;
  assign SystemBus_TLBuffer_auto_out_d_bits_data = auto_anon_out_d_bits_data;
  assign SystemBus_TLBuffer_auto_out_d_bits_error = auto_anon_out_d_bits_error;
  assign SystemBus_TLBuffer_auto_out_e_ready = auto_anon_out_e_ready;
  assign IntSyncCrossingSink_clock = clock;
  assign IntSyncCrossingSink_auto_in_sync_0 = auto_anon_in_0_sync_0;
  assign IntSyncCrossingSink_1_auto_in_2_sync_0 = auto_anon_in_3_sync_0;
  assign IntSyncCrossingSink_1_auto_in_1_sync_0 = auto_anon_in_2_sync_0;
  assign IntSyncCrossingSink_1_auto_in_0_sync_0 = auto_anon_in_1_sync_0;
  assign IntSyncCrossingSink_1_auto_in_0_sync_1 = auto_anon_in_1_sync_1;
endmodule
module AsyncResetRegVec_w2_i0(
  input        clock,
  input        reset,
  input  [1:0] io_d,
  output [1:0] io_q
);
  wire  reg_0_rst;
  wire  reg_0_clk;
  wire  reg_0_en;
  wire  reg_0_q;
  wire  reg_0_d;
  wire  reg_1_rst;
  wire  reg_1_clk;
  wire  reg_1_en;
  wire  reg_1_q;
  wire  reg_1_d;
  wire  _T_5;
  wire  _T_6;
  wire [1:0] _T_7;
  AsyncResetReg reg_0 (
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  AsyncResetReg reg_1 (
    .rst(reg_1_rst),
    .clk(reg_1_clk),
    .en(reg_1_en),
    .q(reg_1_q),
    .d(reg_1_d)
  );
  assign _T_5 = io_d[0];
  assign _T_6 = io_d[1];
  assign _T_7 = {reg_1_q,reg_0_q};
  assign io_q = _T_7;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = 1'h1;
  assign reg_0_d = _T_5;
  assign reg_1_rst = reset;
  assign reg_1_clk = clock;
  assign reg_1_en = 1'h1;
  assign reg_1_d = _T_6;
endmodule
module IntSyncCrossingSource_1(
  input   clock,
  input   reset,
  input   auto_in_2_0,
  input   auto_in_1_0,
  input   auto_in_0_0,
  input   auto_in_0_1,
  output  auto_out_2_sync_0,
  output  auto_out_1_sync_0,
  output  auto_out_0_sync_0,
  output  auto_out_0_sync_1
);
  wire  _T_5_0;
  wire  _T_5_1;
  wire  _T_13_0;
  wire  _T_20_0;
  wire  _T_27_sync_0;
  wire  _T_27_sync_1;
  wire  _T_33_sync_0;
  wire  _T_39_sync_0;
  wire [1:0] _T_92;
  wire  AsyncResetRegVec_w2_i0_clock;
  wire  AsyncResetRegVec_w2_i0_reset;
  wire [1:0] AsyncResetRegVec_w2_i0_io_d;
  wire [1:0] AsyncResetRegVec_w2_i0_io_q;
  wire  _T_94;
  wire  _T_95;
  wire  AsyncResetRegVec_w1_i0_clock;
  wire  AsyncResetRegVec_w1_i0_reset;
  wire  AsyncResetRegVec_w1_i0_io_d;
  wire  AsyncResetRegVec_w1_i0_io_q;
  wire  _T_97;
  wire  AsyncResetRegVec_w1_i0_1_clock;
  wire  AsyncResetRegVec_w1_i0_1_reset;
  wire  AsyncResetRegVec_w1_i0_1_io_d;
  wire  AsyncResetRegVec_w1_i0_1_io_q;
  wire  _T_99;
  AsyncResetRegVec_w2_i0 AsyncResetRegVec_w2_i0 (
    .clock(AsyncResetRegVec_w2_i0_clock),
    .reset(AsyncResetRegVec_w2_i0_reset),
    .io_d(AsyncResetRegVec_w2_i0_io_d),
    .io_q(AsyncResetRegVec_w2_i0_io_q)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 (
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0_1 (
    .clock(AsyncResetRegVec_w1_i0_1_clock),
    .reset(AsyncResetRegVec_w1_i0_1_reset),
    .io_d(AsyncResetRegVec_w1_i0_1_io_d),
    .io_q(AsyncResetRegVec_w1_i0_1_io_q)
  );
  assign _T_92 = {_T_5_1,_T_5_0};
  assign _T_94 = AsyncResetRegVec_w2_i0_io_q[0];
  assign _T_95 = AsyncResetRegVec_w2_i0_io_q[1];
  assign _T_97 = AsyncResetRegVec_w1_i0_io_q;
  assign _T_99 = AsyncResetRegVec_w1_i0_1_io_q;
  assign auto_out_2_sync_0 = _T_39_sync_0;
  assign auto_out_1_sync_0 = _T_33_sync_0;
  assign auto_out_0_sync_0 = _T_27_sync_0;
  assign auto_out_0_sync_1 = _T_27_sync_1;
  assign _T_5_0 = auto_in_0_0;
  assign _T_5_1 = auto_in_0_1;
  assign _T_13_0 = auto_in_1_0;
  assign _T_20_0 = auto_in_2_0;
  assign _T_27_sync_0 = _T_94;
  assign _T_27_sync_1 = _T_95;
  assign _T_33_sync_0 = _T_97;
  assign _T_39_sync_0 = _T_99;
  assign AsyncResetRegVec_w2_i0_io_d = _T_92;
  assign AsyncResetRegVec_w2_i0_clock = clock;
  assign AsyncResetRegVec_w2_i0_reset = reset;
  assign AsyncResetRegVec_w1_i0_io_d = _T_13_0;
  assign AsyncResetRegVec_w1_i0_clock = clock;
  assign AsyncResetRegVec_w1_i0_reset = reset;
  assign AsyncResetRegVec_w1_i0_1_io_d = _T_20_0;
  assign AsyncResetRegVec_w1_i0_1_clock = clock;
  assign AsyncResetRegVec_w1_i0_1_reset = reset;
endmodule
module SynchronizerShiftReg_w2_d3(
  input        clock,
  input  [1:0] io_d,
  output [1:0] io_q
);
  reg [1:0] sync_0;
  reg [31:0] _RAND_0;
  reg [1:0] sync_1;
  reg [31:0] _RAND_1;
  reg [1:0] sync_2;
  reg [31:0] _RAND_2;
  assign io_q = sync_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  sync_0 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  sync_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  sync_2 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= sync_1;
    sync_1 <= sync_2;
    sync_2 <= io_d;
  end
endmodule
module IntXing(
  input   clock,
  input   auto_int_in_0,
  input   auto_int_in_1,
  output  auto_int_out_0,
  output  auto_int_out_1
);
  wire  _T_5_0;
  wire  _T_5_1;
  wire  _T_13_0;
  wire  _T_13_1;
  wire  SynchronizerShiftReg_w2_d3_clock;
  wire [1:0] SynchronizerShiftReg_w2_d3_io_d;
  wire [1:0] SynchronizerShiftReg_w2_d3_io_q;
  wire [1:0] _T_43;
  wire  _T_52_0;
  wire  _T_52_1;
  wire [1:0] _T_64;
  wire  _T_65;
  wire  _T_66;
  SynchronizerShiftReg_w2_d3 SynchronizerShiftReg_w2_d3 (
    .clock(SynchronizerShiftReg_w2_d3_clock),
    .io_d(SynchronizerShiftReg_w2_d3_io_d),
    .io_q(SynchronizerShiftReg_w2_d3_io_q)
  );
  assign _T_43 = {_T_5_1,_T_5_0};
  assign _T_65 = _T_64[0];
  assign _T_66 = _T_64[1];
  assign auto_int_out_0 = _T_13_0;
  assign auto_int_out_1 = _T_13_1;
  assign _T_5_0 = auto_int_in_0;
  assign _T_5_1 = auto_int_in_1;
  assign _T_13_0 = _T_52_0;
  assign _T_13_1 = _T_52_1;
  assign SynchronizerShiftReg_w2_d3_io_d = _T_43;
  assign SynchronizerShiftReg_w2_d3_clock = clock;
  assign _T_52_0 = _T_65;
  assign _T_52_1 = _T_66;
  assign _T_64 = SynchronizerShiftReg_w2_d3_io_q;
endmodule
module Queue_32(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [63:0] ram_data [0:0];
  reg [63:0] _RAND_0;
  wire [63:0] ram_data__T_42_data;
  wire  ram_data__T_42_addr;
  wire [63:0] ram_data__T_33_data;
  wire  ram_data__T_33_addr;
  wire  ram_data__T_33_mask;
  wire  ram_data__T_33_en;
  reg [7:0] ram_strb [0:0];
  reg [31:0] _RAND_1;
  wire [7:0] ram_strb__T_42_data;
  wire  ram_strb__T_42_addr;
  wire [7:0] ram_strb__T_33_data;
  wire  ram_strb__T_33_addr;
  wire  ram_strb__T_33_mask;
  wire  ram_strb__T_33_en;
  reg  ram_last [0:0];
  reg [31:0] _RAND_2;
  wire  ram_last__T_42_data;
  wire  ram_last__T_42_addr;
  wire  ram_last__T_33_data;
  wire  ram_last__T_33_addr;
  wire  ram_last__T_33_mask;
  wire  ram_last__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_6;
  wire  _T_38;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire [7:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  assign ram_data__T_42_addr = 1'h0;
  assign ram_data__T_42_data = ram_data[ram_data__T_42_addr];
  assign ram_data__T_33_data = io_enq_bits_data;
  assign ram_data__T_33_addr = 1'h0;
  assign ram_data__T_33_mask = do_enq;
  assign ram_data__T_33_en = do_enq;
  assign ram_strb__T_42_addr = 1'h0;
  assign ram_strb__T_42_data = ram_strb[ram_strb__T_42_addr];
  assign ram_strb__T_33_data = io_enq_bits_strb;
  assign ram_strb__T_33_addr = 1'h0;
  assign ram_strb__T_33_mask = do_enq;
  assign ram_strb__T_33_en = do_enq;
  assign ram_last__T_42_addr = 1'h0;
  assign ram_last__T_42_data = ram_last[ram_last__T_42_addr];
  assign ram_last__T_33_data = io_enq_bits_last;
  assign ram_last__T_33_addr = 1'h0;
  assign ram_last__T_33_mask = do_enq;
  assign ram_last__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_6 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_7 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_8 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_9 = empty ? io_enq_bits_last : ram_last__T_42_data;
  assign _GEN_10 = empty ? io_enq_bits_strb : ram_strb__T_42_data;
  assign _GEN_11 = empty ? io_enq_bits_data : ram_data__T_42_data;
  assign _GEN_12 = empty ? 1'h0 : _T_30;
  assign _GEN_13 = empty ? _GEN_8 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_7;
  assign io_deq_bits_data = _GEN_11;
  assign io_deq_bits_strb = _GEN_10;
  assign io_deq_bits_last = _GEN_9;
  assign do_enq = _GEN_13;
  assign do_deq = _GEN_12;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_data__T_33_en & ram_data__T_33_mask) begin
      ram_data[ram_data__T_33_addr] <= ram_data__T_33_data;
    end
    if(ram_strb__T_33_en & ram_strb__T_33_mask) begin
      ram_strb[ram_strb__T_33_addr] <= ram_strb__T_33_data;
    end
    if(ram_last__T_33_en & ram_last__T_33_mask) begin
      ram_last[ram_last__T_33_addr] <= ram_last__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_33(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [6:0]  io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [10:0] io_enq_bits_user,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [6:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [10:0] io_deq_bits_user,
  output        io_deq_bits_wen
);
  reg [6:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [6:0] ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire [6:0] ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [31:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [31:0] ram_addr__T_42_data;
  wire  ram_addr__T_42_addr;
  wire [31:0] ram_addr__T_33_data;
  wire  ram_addr__T_33_addr;
  wire  ram_addr__T_33_mask;
  wire  ram_addr__T_33_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_42_data;
  wire  ram_len__T_42_addr;
  wire [7:0] ram_len__T_33_data;
  wire  ram_len__T_33_addr;
  wire  ram_len__T_33_mask;
  wire  ram_len__T_33_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [2:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_42_data;
  wire  ram_burst__T_42_addr;
  wire [1:0] ram_burst__T_33_data;
  wire  ram_burst__T_33_addr;
  wire  ram_burst__T_33_mask;
  wire  ram_burst__T_33_en;
  reg  ram_lock [0:0];
  reg [31:0] _RAND_5;
  wire  ram_lock__T_42_data;
  wire  ram_lock__T_42_addr;
  wire  ram_lock__T_33_data;
  wire  ram_lock__T_33_addr;
  wire  ram_lock__T_33_mask;
  wire  ram_lock__T_33_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] _RAND_6;
  wire [3:0] ram_cache__T_42_data;
  wire  ram_cache__T_42_addr;
  wire [3:0] ram_cache__T_33_data;
  wire  ram_cache__T_33_addr;
  wire  ram_cache__T_33_mask;
  wire  ram_cache__T_33_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] _RAND_7;
  wire [2:0] ram_prot__T_42_data;
  wire  ram_prot__T_42_addr;
  wire [2:0] ram_prot__T_33_data;
  wire  ram_prot__T_33_addr;
  wire  ram_prot__T_33_mask;
  wire  ram_prot__T_33_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] _RAND_8;
  wire [3:0] ram_qos__T_42_data;
  wire  ram_qos__T_42_addr;
  wire [3:0] ram_qos__T_33_data;
  wire  ram_qos__T_33_addr;
  wire  ram_qos__T_33_mask;
  wire  ram_qos__T_33_en;
  reg [10:0] ram_user [0:0];
  reg [31:0] _RAND_9;
  wire [10:0] ram_user__T_42_data;
  wire  ram_user__T_42_addr;
  wire [10:0] ram_user__T_33_data;
  wire  ram_user__T_33_addr;
  wire  ram_user__T_33_mask;
  wire  ram_user__T_33_en;
  reg  ram_wen [0:0];
  reg [31:0] _RAND_10;
  wire  ram_wen__T_42_data;
  wire  ram_wen__T_42_addr;
  wire  ram_wen__T_33_data;
  wire  ram_wen__T_33_addr;
  wire  ram_wen__T_33_mask;
  wire  ram_wen__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_11;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_14;
  wire  _T_38;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire [10:0] _GEN_18;
  wire [3:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [3:0] _GEN_21;
  wire  _GEN_22;
  wire [1:0] _GEN_23;
  wire [2:0] _GEN_24;
  wire [7:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [6:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_addr__T_42_addr = 1'h0;
  assign ram_addr__T_42_data = ram_addr[ram_addr__T_42_addr];
  assign ram_addr__T_33_data = io_enq_bits_addr;
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_mask = do_enq;
  assign ram_addr__T_33_en = do_enq;
  assign ram_len__T_42_addr = 1'h0;
  assign ram_len__T_42_data = ram_len[ram_len__T_42_addr];
  assign ram_len__T_33_data = io_enq_bits_len;
  assign ram_len__T_33_addr = 1'h0;
  assign ram_len__T_33_mask = do_enq;
  assign ram_len__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_burst__T_42_addr = 1'h0;
  assign ram_burst__T_42_data = ram_burst[ram_burst__T_42_addr];
  assign ram_burst__T_33_data = 2'h1;
  assign ram_burst__T_33_addr = 1'h0;
  assign ram_burst__T_33_mask = do_enq;
  assign ram_burst__T_33_en = do_enq;
  assign ram_lock__T_42_addr = 1'h0;
  assign ram_lock__T_42_data = ram_lock[ram_lock__T_42_addr];
  assign ram_lock__T_33_data = 1'h0;
  assign ram_lock__T_33_addr = 1'h0;
  assign ram_lock__T_33_mask = do_enq;
  assign ram_lock__T_33_en = do_enq;
  assign ram_cache__T_42_addr = 1'h0;
  assign ram_cache__T_42_data = ram_cache[ram_cache__T_42_addr];
  assign ram_cache__T_33_data = 4'h0;
  assign ram_cache__T_33_addr = 1'h0;
  assign ram_cache__T_33_mask = do_enq;
  assign ram_cache__T_33_en = do_enq;
  assign ram_prot__T_42_addr = 1'h0;
  assign ram_prot__T_42_data = ram_prot[ram_prot__T_42_addr];
  assign ram_prot__T_33_data = 3'h1;
  assign ram_prot__T_33_addr = 1'h0;
  assign ram_prot__T_33_mask = do_enq;
  assign ram_prot__T_33_en = do_enq;
  assign ram_qos__T_42_addr = 1'h0;
  assign ram_qos__T_42_data = ram_qos[ram_qos__T_42_addr];
  assign ram_qos__T_33_data = 4'h0;
  assign ram_qos__T_33_addr = 1'h0;
  assign ram_qos__T_33_mask = do_enq;
  assign ram_qos__T_33_en = do_enq;
  assign ram_user__T_42_addr = 1'h0;
  assign ram_user__T_42_data = ram_user[ram_user__T_42_addr];
  assign ram_user__T_33_data = io_enq_bits_user;
  assign ram_user__T_33_addr = 1'h0;
  assign ram_user__T_33_mask = do_enq;
  assign ram_user__T_33_en = do_enq;
  assign ram_wen__T_42_addr = 1'h0;
  assign ram_wen__T_42_data = ram_wen[ram_wen__T_42_addr];
  assign ram_wen__T_33_data = io_enq_bits_wen;
  assign ram_wen__T_33_addr = 1'h0;
  assign ram_wen__T_33_mask = do_enq;
  assign ram_wen__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_14 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_15 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_16 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_17 = empty ? io_enq_bits_wen : ram_wen__T_42_data;
  assign _GEN_18 = empty ? io_enq_bits_user : ram_user__T_42_data;
  assign _GEN_19 = empty ? 4'h0 : ram_qos__T_42_data;
  assign _GEN_20 = empty ? 3'h1 : ram_prot__T_42_data;
  assign _GEN_21 = empty ? 4'h0 : ram_cache__T_42_data;
  assign _GEN_22 = empty ? 1'h0 : ram_lock__T_42_data;
  assign _GEN_23 = empty ? 2'h1 : ram_burst__T_42_data;
  assign _GEN_24 = empty ? io_enq_bits_size : ram_size__T_42_data;
  assign _GEN_25 = empty ? io_enq_bits_len : ram_len__T_42_data;
  assign _GEN_26 = empty ? io_enq_bits_addr : ram_addr__T_42_data;
  assign _GEN_27 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_28 = empty ? 1'h0 : _T_30;
  assign _GEN_29 = empty ? _GEN_16 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_15;
  assign io_deq_bits_id = _GEN_27;
  assign io_deq_bits_addr = _GEN_26;
  assign io_deq_bits_len = _GEN_25;
  assign io_deq_bits_size = _GEN_24;
  assign io_deq_bits_burst = _GEN_23;
  assign io_deq_bits_lock = _GEN_22;
  assign io_deq_bits_cache = _GEN_21;
  assign io_deq_bits_prot = _GEN_20;
  assign io_deq_bits_qos = _GEN_19;
  assign io_deq_bits_user = _GEN_18;
  assign io_deq_bits_wen = _GEN_17;
  assign do_enq = _GEN_29;
  assign do_deq = _GEN_28;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[6:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = _RAND_9[10:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  maybe_full = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_addr__T_33_en & ram_addr__T_33_mask) begin
      ram_addr[ram_addr__T_33_addr] <= ram_addr__T_33_data;
    end
    if(ram_len__T_33_en & ram_len__T_33_mask) begin
      ram_len[ram_len__T_33_addr] <= ram_len__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_burst__T_33_en & ram_burst__T_33_mask) begin
      ram_burst[ram_burst__T_33_addr] <= ram_burst__T_33_data;
    end
    if(ram_lock__T_33_en & ram_lock__T_33_mask) begin
      ram_lock[ram_lock__T_33_addr] <= ram_lock__T_33_data;
    end
    if(ram_cache__T_33_en & ram_cache__T_33_mask) begin
      ram_cache[ram_cache__T_33_addr] <= ram_cache__T_33_data;
    end
    if(ram_prot__T_33_en & ram_prot__T_33_mask) begin
      ram_prot[ram_prot__T_33_addr] <= ram_prot__T_33_data;
    end
    if(ram_qos__T_33_en & ram_qos__T_33_mask) begin
      ram_qos[ram_qos__T_33_addr] <= ram_qos__T_33_data;
    end
    if(ram_user__T_33_en & ram_user__T_33_mask) begin
      ram_user[ram_user__T_33_addr] <= ram_user__T_33_data;
    end
    if(ram_wen__T_33_en & ram_wen__T_33_mask) begin
      ram_wen[ram_wen__T_33_addr] <= ram_wen__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TLToAXI4_converter(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [6:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [10:0] auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [6:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [10:0] auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [6:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [10:0] auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [6:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [10:0] auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [2:0] _T_31_a_bits_size;
  wire [6:0] _T_31_a_bits_source;
  wire [31:0] _T_31_a_bits_address;
  wire [7:0] _T_31_a_bits_mask;
  wire [63:0] _T_31_a_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [2:0] _T_31_d_bits_size;
  wire [6:0] _T_31_d_bits_source;
  wire [63:0] _T_31_d_bits_data;
  wire  _T_31_d_bits_error;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [6:0] _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire [10:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [6:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [10:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [6:0] _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire [10:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [6:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [10:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  _T_206_0;
  wire  _T_206_1;
  wire  _T_206_2;
  wire  _T_206_3;
  wire  _T_206_4;
  wire  _T_206_5;
  wire  _T_206_6;
  wire  _T_206_7;
  wire  _T_206_8;
  wire  _T_206_9;
  wire  _T_206_10;
  wire  _T_206_11;
  wire  _T_206_12;
  wire  _T_206_13;
  wire  _T_206_14;
  wire  _T_206_15;
  wire  _T_206_16;
  wire  _T_206_17;
  wire  _T_206_18;
  wire  _T_206_19;
  wire  _T_206_20;
  wire  _T_206_21;
  wire  _T_206_22;
  wire  _T_206_23;
  wire  _T_206_24;
  wire  _T_206_25;
  wire  _T_206_26;
  wire  _T_206_27;
  wire  _T_206_28;
  wire  _T_206_29;
  wire  _T_206_30;
  wire  _T_206_31;
  wire  _T_206_32;
  wire  _T_206_33;
  wire  _T_206_34;
  wire  _T_206_35;
  wire  _T_206_36;
  wire  _T_206_37;
  wire  _T_206_38;
  wire  _T_206_39;
  wire  _T_206_40;
  wire  _T_206_41;
  wire  _T_206_42;
  wire  _T_206_43;
  wire  _T_206_44;
  wire  _T_206_45;
  wire  _T_206_46;
  wire  _T_206_47;
  wire  _T_206_48;
  wire  _T_206_49;
  wire  _T_206_50;
  wire  _T_206_51;
  wire  _T_206_52;
  wire  _T_206_53;
  wire  _T_206_54;
  wire  _T_206_55;
  wire  _T_206_56;
  wire  _T_206_57;
  wire  _T_206_58;
  wire  _T_206_59;
  wire  _T_206_60;
  wire  _T_206_61;
  wire  _T_206_62;
  wire  _T_206_63;
  wire  _T_206_64;
  wire  _T_206_65;
  wire  _T_206_66;
  wire  _T_206_67;
  wire  _T_206_68;
  wire  _T_206_69;
  wire  _T_206_70;
  wire  _T_206_71;
  wire  _T_206_72;
  wire  _T_206_73;
  wire  _T_206_74;
  wire  _T_206_75;
  wire  _T_206_76;
  wire  _T_206_77;
  wire  _T_206_78;
  wire  _T_206_79;
  wire  _T_206_80;
  wire  _T_206_81;
  wire  _T_206_82;
  wire  _T_206_83;
  wire  _T_206_84;
  wire  _T_206_85;
  wire  _T_206_86;
  wire  _T_206_87;
  wire  _T_206_88;
  wire  _T_206_89;
  wire  _T_206_90;
  wire  _T_206_91;
  wire  _T_206_92;
  wire  _T_206_93;
  wire  _T_206_94;
  wire  _T_206_95;
  wire  _T_206_96;
  wire  _T_206_97;
  wire  _T_206_98;
  wire  _T_206_99;
  wire  _T_206_100;
  wire  _T_206_101;
  wire  _T_206_102;
  wire  _T_206_103;
  wire  _T_206_104;
  wire  _T_206_105;
  wire  _T_206_106;
  wire  _T_206_107;
  wire  _T_206_108;
  wire  _T_206_109;
  wire  _T_206_110;
  wire  _T_206_111;
  wire  _T_206_112;
  wire  _T_206_113;
  wire  _T_206_114;
  wire  _T_206_115;
  wire  _T_206_116;
  wire  _T_206_117;
  wire  _T_206_118;
  wire  _T_206_119;
  wire  _T_206_120;
  wire  _T_206_121;
  wire  _T_206_122;
  wire  _T_206_123;
  wire  _T_206_124;
  wire  _T_206_125;
  wire  _T_206_126;
  wire  _T_206_127;
  wire  _T_991_0;
  wire  _T_991_1;
  wire  _T_991_2;
  wire  _T_991_3;
  wire  _T_991_4;
  wire  _T_991_5;
  wire  _T_991_6;
  wire  _T_991_7;
  wire  _T_991_8;
  wire  _T_991_9;
  wire  _T_991_10;
  wire  _T_991_11;
  wire  _T_991_12;
  wire  _T_991_13;
  wire  _T_991_14;
  wire  _T_991_15;
  wire  _T_991_16;
  wire  _T_991_17;
  wire  _T_991_18;
  wire  _T_991_19;
  wire  _T_991_20;
  wire  _T_991_21;
  wire  _T_991_22;
  wire  _T_991_23;
  wire  _T_991_24;
  wire  _T_991_25;
  wire  _T_991_26;
  wire  _T_991_27;
  wire  _T_991_28;
  wire  _T_991_29;
  wire  _T_991_30;
  wire  _T_991_31;
  wire  _T_991_32;
  wire  _T_991_33;
  wire  _T_991_34;
  wire  _T_991_35;
  wire  _T_991_36;
  wire  _T_991_37;
  wire  _T_991_38;
  wire  _T_991_39;
  wire  _T_991_40;
  wire  _T_991_41;
  wire  _T_991_42;
  wire  _T_991_43;
  wire  _T_991_44;
  wire  _T_991_45;
  wire  _T_991_46;
  wire  _T_991_47;
  wire  _T_991_48;
  wire  _T_991_49;
  wire  _T_991_50;
  wire  _T_991_51;
  wire  _T_991_52;
  wire  _T_991_53;
  wire  _T_991_54;
  wire  _T_991_55;
  wire  _T_991_56;
  wire  _T_991_57;
  wire  _T_991_58;
  wire  _T_991_59;
  wire  _T_991_60;
  wire  _T_991_61;
  wire  _T_991_62;
  wire  _T_991_63;
  wire  _T_991_64;
  wire  _T_991_65;
  wire  _T_991_66;
  wire  _T_991_67;
  wire  _T_991_68;
  wire  _T_991_69;
  wire  _T_991_70;
  wire  _T_991_71;
  wire  _T_991_72;
  wire  _T_991_73;
  wire  _T_991_74;
  wire  _T_991_75;
  wire  _T_991_76;
  wire  _T_991_77;
  wire  _T_991_78;
  wire  _T_991_79;
  wire  _T_991_80;
  wire  _T_991_81;
  wire  _T_991_82;
  wire  _T_991_83;
  wire  _T_991_84;
  wire  _T_991_85;
  wire  _T_991_86;
  wire  _T_991_87;
  wire  _T_991_88;
  wire  _T_991_89;
  wire  _T_991_90;
  wire  _T_991_91;
  wire  _T_991_92;
  wire  _T_991_93;
  wire  _T_991_94;
  wire  _T_991_95;
  wire  _T_991_96;
  wire  _T_991_97;
  wire  _T_991_98;
  wire  _T_991_99;
  wire  _T_991_100;
  wire  _T_991_101;
  wire  _T_991_102;
  wire  _T_991_103;
  wire  _T_991_104;
  wire  _T_991_105;
  wire  _T_991_106;
  wire  _T_991_107;
  wire  _T_991_108;
  wire  _T_991_109;
  wire  _T_991_110;
  wire  _T_991_111;
  wire  _T_991_112;
  wire  _T_991_113;
  wire  _T_991_114;
  wire  _T_991_115;
  wire  _T_991_116;
  wire  _T_991_117;
  wire  _T_991_118;
  wire  _T_991_119;
  wire  _T_991_120;
  wire  _T_991_121;
  wire  _T_991_122;
  wire  _T_991_123;
  wire  _T_991_124;
  wire  _T_991_125;
  wire  _T_991_126;
  wire  _T_991_127;
  wire  _T_1508;
  wire  _T_1510;
  wire  _T_1511;
  wire [12:0] _T_1514;
  wire [5:0] _T_1515;
  wire [5:0] _T_1516;
  wire [2:0] _T_1517;
  wire [2:0] _T_1522;
  reg [2:0] _T_1525;
  reg [31:0] _RAND_0;
  wire [3:0] _T_1527;
  wire [3:0] _T_1528;
  wire [2:0] _T_1529;
  wire  _T_1531;
  wire  _T_1533;
  wire  _T_1535;
  wire  _T_1536;
  wire [2:0] _T_1540;
  wire [2:0] _GEN_2;
  wire [9:0] _GEN_388;
  wire [9:0] _T_1554;
  wire [9:0] _GEN_389;
  wire [9:0] _T_1555;
  wire [6:0] _T_1556;
  wire [2:0] _T_1557;
  wire [6:0] _T_1558;
  wire [2:0] _T_1559;
  wire  _T_1565_ready;
  wire  _T_1565_valid;
  wire [6:0] _T_1565_bits_id;
  wire [31:0] _T_1565_bits_addr;
  wire [7:0] _T_1565_bits_len;
  wire [2:0] _T_1565_bits_size;
  wire [10:0] _T_1565_bits_user;
  wire  _T_1565_bits_wen;
  wire  _T_1569_ready;
  wire  _T_1569_valid;
  wire [63:0] _T_1569_bits_data;
  wire [7:0] _T_1569_bits_strb;
  wire  _T_1569_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [63:0] Queue_io_enq_bits_data;
  wire [7:0] Queue_io_enq_bits_strb;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [63:0] Queue_io_deq_bits_data;
  wire [7:0] Queue_io_deq_bits_strb;
  wire  Queue_io_deq_bits_last;
  wire  _T_1577_ready;
  wire  _T_1577_valid;
  wire [63:0] _T_1577_bits_data;
  wire [7:0] _T_1577_bits_strb;
  wire  _T_1577_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [6:0] Queue_1_io_enq_bits_id;
  wire [31:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [10:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_enq_bits_wen;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [6:0] Queue_1_io_deq_bits_id;
  wire [31:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire  Queue_1_io_deq_bits_lock;
  wire [3:0] Queue_1_io_deq_bits_cache;
  wire [2:0] Queue_1_io_deq_bits_prot;
  wire [3:0] Queue_1_io_deq_bits_qos;
  wire [10:0] Queue_1_io_deq_bits_user;
  wire  Queue_1_io_deq_bits_wen;
  wire  _T_1585_ready;
  wire  _T_1585_valid;
  wire [6:0] _T_1585_bits_id;
  wire [31:0] _T_1585_bits_addr;
  wire [7:0] _T_1585_bits_len;
  wire [2:0] _T_1585_bits_size;
  wire [1:0] _T_1585_bits_burst;
  wire  _T_1585_bits_lock;
  wire [3:0] _T_1585_bits_cache;
  wire [2:0] _T_1585_bits_prot;
  wire [3:0] _T_1585_bits_qos;
  wire [10:0] _T_1585_bits_user;
  wire  _T_1585_bits_wen;
  wire  _T_1590;
  wire  _T_1591;
  wire  _T_1592;
  wire  _T_1593;
  reg  _T_1597;
  reg [31:0] _RAND_1;
  wire  _T_1600;
  wire  _GEN_3;
  wire [6:0] _GEN_0;
  wire [6:0] _GEN_4;
  wire [6:0] _GEN_5;
  wire [6:0] _GEN_6;
  wire [6:0] _GEN_7;
  wire [6:0] _GEN_8;
  wire [6:0] _GEN_9;
  wire [6:0] _GEN_10;
  wire [6:0] _GEN_11;
  wire [6:0] _GEN_12;
  wire [6:0] _GEN_13;
  wire [6:0] _GEN_14;
  wire [6:0] _GEN_15;
  wire [6:0] _GEN_16;
  wire [6:0] _GEN_17;
  wire [6:0] _GEN_18;
  wire [6:0] _GEN_19;
  wire [6:0] _GEN_20;
  wire [6:0] _GEN_21;
  wire [6:0] _GEN_22;
  wire [6:0] _GEN_23;
  wire [6:0] _GEN_24;
  wire [6:0] _GEN_25;
  wire [6:0] _GEN_26;
  wire [6:0] _GEN_27;
  wire [6:0] _GEN_28;
  wire [6:0] _GEN_29;
  wire [6:0] _GEN_30;
  wire [6:0] _GEN_31;
  wire [6:0] _GEN_32;
  wire [6:0] _GEN_33;
  wire [6:0] _GEN_34;
  wire [6:0] _GEN_35;
  wire [6:0] _GEN_36;
  wire [6:0] _GEN_37;
  wire [6:0] _GEN_38;
  wire [6:0] _GEN_39;
  wire [6:0] _GEN_40;
  wire [6:0] _GEN_41;
  wire [6:0] _GEN_42;
  wire [6:0] _GEN_43;
  wire [6:0] _GEN_44;
  wire [6:0] _GEN_45;
  wire [6:0] _GEN_46;
  wire [6:0] _GEN_47;
  wire [6:0] _GEN_48;
  wire [6:0] _GEN_49;
  wire [6:0] _GEN_50;
  wire [6:0] _GEN_51;
  wire [6:0] _GEN_52;
  wire [6:0] _GEN_53;
  wire [6:0] _GEN_54;
  wire [6:0] _GEN_55;
  wire [6:0] _GEN_56;
  wire [6:0] _GEN_57;
  wire [6:0] _GEN_58;
  wire [6:0] _GEN_59;
  wire [6:0] _GEN_60;
  wire [6:0] _GEN_61;
  wire [6:0] _GEN_62;
  wire [6:0] _GEN_63;
  wire [6:0] _GEN_64;
  wire [6:0] _GEN_65;
  wire [6:0] _GEN_66;
  wire [6:0] _GEN_67;
  wire [6:0] _GEN_68;
  wire [6:0] _GEN_69;
  wire [6:0] _GEN_70;
  wire [6:0] _GEN_71;
  wire [6:0] _GEN_72;
  wire [6:0] _GEN_73;
  wire [6:0] _GEN_74;
  wire [6:0] _GEN_75;
  wire [6:0] _GEN_76;
  wire [6:0] _GEN_77;
  wire [6:0] _GEN_78;
  wire [6:0] _GEN_79;
  wire [6:0] _GEN_80;
  wire [6:0] _GEN_81;
  wire [6:0] _GEN_82;
  wire [6:0] _GEN_83;
  wire [6:0] _GEN_84;
  wire [6:0] _GEN_85;
  wire [6:0] _GEN_86;
  wire [6:0] _GEN_87;
  wire [6:0] _GEN_88;
  wire [6:0] _GEN_89;
  wire [6:0] _GEN_90;
  wire [6:0] _GEN_91;
  wire [6:0] _GEN_92;
  wire [6:0] _GEN_93;
  wire [6:0] _GEN_94;
  wire [6:0] _GEN_95;
  wire [6:0] _GEN_96;
  wire [6:0] _GEN_97;
  wire [6:0] _GEN_98;
  wire [6:0] _GEN_99;
  wire [6:0] _GEN_100;
  wire [6:0] _GEN_101;
  wire [6:0] _GEN_102;
  wire [6:0] _GEN_103;
  wire [6:0] _GEN_104;
  wire [6:0] _GEN_105;
  wire [6:0] _GEN_106;
  wire [6:0] _GEN_107;
  wire [6:0] _GEN_108;
  wire [6:0] _GEN_109;
  wire [6:0] _GEN_110;
  wire [6:0] _GEN_111;
  wire [6:0] _GEN_112;
  wire [6:0] _GEN_113;
  wire [6:0] _GEN_114;
  wire [6:0] _GEN_115;
  wire [6:0] _GEN_116;
  wire [6:0] _GEN_117;
  wire [6:0] _GEN_118;
  wire [6:0] _GEN_119;
  wire [6:0] _GEN_120;
  wire [6:0] _GEN_121;
  wire [6:0] _GEN_122;
  wire [6:0] _GEN_123;
  wire [6:0] _GEN_124;
  wire [6:0] _GEN_125;
  wire [6:0] _GEN_126;
  wire [6:0] _GEN_127;
  wire [6:0] _GEN_128;
  wire [6:0] _GEN_129;
  wire [6:0] _GEN_130;
  wire [17:0] _T_1604;
  wire [10:0] _T_1605;
  wire [10:0] _T_1606;
  wire [7:0] _T_1607;
  wire  _T_1608;
  wire [2:0] _T_1609;
  wire  _GEN_1;
  wire  _GEN_131;
  wire  _GEN_132;
  wire  _GEN_133;
  wire  _GEN_134;
  wire  _GEN_135;
  wire  _GEN_136;
  wire  _GEN_137;
  wire  _GEN_138;
  wire  _GEN_139;
  wire  _GEN_140;
  wire  _GEN_141;
  wire  _GEN_142;
  wire  _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire  _GEN_147;
  wire  _GEN_148;
  wire  _GEN_149;
  wire  _GEN_150;
  wire  _GEN_151;
  wire  _GEN_152;
  wire  _GEN_153;
  wire  _GEN_154;
  wire  _GEN_155;
  wire  _GEN_156;
  wire  _GEN_157;
  wire  _GEN_158;
  wire  _GEN_159;
  wire  _GEN_160;
  wire  _GEN_161;
  wire  _GEN_162;
  wire  _GEN_163;
  wire  _GEN_164;
  wire  _GEN_165;
  wire  _GEN_166;
  wire  _GEN_167;
  wire  _GEN_168;
  wire  _GEN_169;
  wire  _GEN_170;
  wire  _GEN_171;
  wire  _GEN_172;
  wire  _GEN_173;
  wire  _GEN_174;
  wire  _GEN_175;
  wire  _GEN_176;
  wire  _GEN_177;
  wire  _GEN_178;
  wire  _GEN_179;
  wire  _GEN_180;
  wire  _GEN_181;
  wire  _GEN_182;
  wire  _GEN_183;
  wire  _GEN_184;
  wire  _GEN_185;
  wire  _GEN_186;
  wire  _GEN_187;
  wire  _GEN_188;
  wire  _GEN_189;
  wire  _GEN_190;
  wire  _GEN_191;
  wire  _GEN_192;
  wire  _GEN_193;
  wire  _GEN_194;
  wire  _GEN_195;
  wire  _GEN_196;
  wire  _GEN_197;
  wire  _GEN_198;
  wire  _GEN_199;
  wire  _GEN_200;
  wire  _GEN_201;
  wire  _GEN_202;
  wire  _GEN_203;
  wire  _GEN_204;
  wire  _GEN_205;
  wire  _GEN_206;
  wire  _GEN_207;
  wire  _GEN_208;
  wire  _GEN_209;
  wire  _GEN_210;
  wire  _GEN_211;
  wire  _GEN_212;
  wire  _GEN_213;
  wire  _GEN_214;
  wire  _GEN_215;
  wire  _GEN_216;
  wire  _GEN_217;
  wire  _GEN_218;
  wire  _GEN_219;
  wire  _GEN_220;
  wire  _GEN_221;
  wire  _GEN_222;
  wire  _GEN_223;
  wire  _GEN_224;
  wire  _GEN_225;
  wire  _GEN_226;
  wire  _GEN_227;
  wire  _GEN_228;
  wire  _GEN_229;
  wire  _GEN_230;
  wire  _GEN_231;
  wire  _GEN_232;
  wire  _GEN_233;
  wire  _GEN_234;
  wire  _GEN_235;
  wire  _GEN_236;
  wire  _GEN_237;
  wire  _GEN_238;
  wire  _GEN_239;
  wire  _GEN_240;
  wire  _GEN_241;
  wire  _GEN_242;
  wire  _GEN_243;
  wire  _GEN_244;
  wire  _GEN_245;
  wire  _GEN_246;
  wire  _GEN_247;
  wire  _GEN_248;
  wire  _GEN_249;
  wire  _GEN_250;
  wire  _GEN_251;
  wire  _GEN_252;
  wire  _GEN_253;
  wire  _GEN_254;
  wire  _GEN_255;
  wire  _GEN_256;
  wire  _GEN_257;
  wire  _T_1616;
  wire  _T_1618;
  wire  _T_1619;
  wire  _T_1620;
  wire  _T_1621;
  wire  _T_1622;
  wire  _T_1625;
  wire  _T_1627;
  wire  _T_1628;
  wire  _T_1630;
  wire  _T_1631;
  wire  _T_1635;
  wire  _T_1637;
  reg  _T_1640;
  reg [31:0] _RAND_2;
  wire  _T_1641;
  wire  _T_1643;
  wire  _GEN_258;
  wire  _T_1644;
  wire  _T_1646;
  wire  _T_1647;
  wire  _T_1648;
  wire  _T_1650;
  wire  _T_1652;
  reg  _T_1655;
  reg [31:0] _RAND_3;
  wire  _T_1659;
  wire  _T_1660;
  wire  _GEN_259;
  wire [2:0] _T_1664_size;
  wire [6:0] _T_1664_source;
  wire  _T_1664_error;
  wire [2:0] _T_1669_size;
  wire [6:0] _T_1669_source;
  wire  _T_1669_error;
  wire [2:0] _T_1674_opcode;
  wire [2:0] _T_1674_size;
  wire [6:0] _T_1674_source;
  wire  _T_1674_error;
  wire [127:0] _T_1677;
  wire  _T_1679;
  wire  _T_1680;
  wire  _T_1681;
  wire  _T_1682;
  wire  _T_1683;
  wire  _T_1684;
  wire  _T_1685;
  wire  _T_1686;
  wire  _T_1687;
  wire  _T_1688;
  wire  _T_1689;
  wire  _T_1690;
  wire  _T_1691;
  wire  _T_1692;
  wire  _T_1693;
  wire  _T_1694;
  wire  _T_1695;
  wire  _T_1696;
  wire  _T_1697;
  wire  _T_1698;
  wire  _T_1699;
  wire  _T_1700;
  wire  _T_1701;
  wire  _T_1702;
  wire  _T_1703;
  wire  _T_1704;
  wire  _T_1705;
  wire  _T_1706;
  wire  _T_1707;
  wire  _T_1708;
  wire  _T_1709;
  wire  _T_1710;
  wire  _T_1711;
  wire  _T_1712;
  wire  _T_1713;
  wire  _T_1714;
  wire  _T_1715;
  wire  _T_1716;
  wire  _T_1717;
  wire  _T_1718;
  wire  _T_1719;
  wire  _T_1720;
  wire  _T_1721;
  wire  _T_1722;
  wire  _T_1723;
  wire  _T_1724;
  wire  _T_1725;
  wire  _T_1726;
  wire  _T_1727;
  wire  _T_1728;
  wire  _T_1729;
  wire  _T_1730;
  wire  _T_1731;
  wire  _T_1732;
  wire  _T_1733;
  wire  _T_1734;
  wire  _T_1735;
  wire  _T_1736;
  wire  _T_1737;
  wire  _T_1738;
  wire  _T_1739;
  wire  _T_1740;
  wire  _T_1741;
  wire  _T_1742;
  wire  _T_1743;
  wire  _T_1744;
  wire  _T_1745;
  wire  _T_1746;
  wire  _T_1747;
  wire  _T_1748;
  wire  _T_1749;
  wire  _T_1750;
  wire  _T_1751;
  wire  _T_1752;
  wire  _T_1753;
  wire  _T_1754;
  wire  _T_1755;
  wire  _T_1756;
  wire  _T_1757;
  wire  _T_1758;
  wire  _T_1759;
  wire  _T_1760;
  wire  _T_1761;
  wire  _T_1762;
  wire  _T_1763;
  wire  _T_1764;
  wire  _T_1765;
  wire  _T_1766;
  wire  _T_1767;
  wire  _T_1768;
  wire  _T_1769;
  wire  _T_1770;
  wire  _T_1771;
  wire  _T_1772;
  wire  _T_1773;
  wire  _T_1774;
  wire  _T_1775;
  wire  _T_1776;
  wire  _T_1777;
  wire  _T_1778;
  wire  _T_1779;
  wire  _T_1780;
  wire  _T_1781;
  wire  _T_1782;
  wire  _T_1783;
  wire  _T_1784;
  wire  _T_1785;
  wire  _T_1786;
  wire  _T_1787;
  wire  _T_1788;
  wire  _T_1789;
  wire  _T_1790;
  wire  _T_1791;
  wire  _T_1792;
  wire  _T_1793;
  wire  _T_1794;
  wire  _T_1795;
  wire  _T_1796;
  wire  _T_1797;
  wire  _T_1798;
  wire  _T_1799;
  wire  _T_1800;
  wire  _T_1801;
  wire  _T_1802;
  wire  _T_1803;
  wire  _T_1804;
  wire  _T_1805;
  wire  _T_1806;
  wire [6:0] _T_1807;
  wire [127:0] _T_1810;
  wire  _T_1812;
  wire  _T_1813;
  wire  _T_1814;
  wire  _T_1815;
  wire  _T_1816;
  wire  _T_1817;
  wire  _T_1818;
  wire  _T_1819;
  wire  _T_1820;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1823;
  wire  _T_1824;
  wire  _T_1825;
  wire  _T_1826;
  wire  _T_1827;
  wire  _T_1828;
  wire  _T_1829;
  wire  _T_1830;
  wire  _T_1831;
  wire  _T_1832;
  wire  _T_1833;
  wire  _T_1834;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1837;
  wire  _T_1838;
  wire  _T_1839;
  wire  _T_1840;
  wire  _T_1841;
  wire  _T_1842;
  wire  _T_1843;
  wire  _T_1844;
  wire  _T_1845;
  wire  _T_1846;
  wire  _T_1847;
  wire  _T_1848;
  wire  _T_1849;
  wire  _T_1850;
  wire  _T_1851;
  wire  _T_1852;
  wire  _T_1853;
  wire  _T_1854;
  wire  _T_1855;
  wire  _T_1856;
  wire  _T_1857;
  wire  _T_1858;
  wire  _T_1859;
  wire  _T_1860;
  wire  _T_1861;
  wire  _T_1862;
  wire  _T_1863;
  wire  _T_1864;
  wire  _T_1865;
  wire  _T_1866;
  wire  _T_1867;
  wire  _T_1868;
  wire  _T_1869;
  wire  _T_1870;
  wire  _T_1871;
  wire  _T_1872;
  wire  _T_1873;
  wire  _T_1874;
  wire  _T_1875;
  wire  _T_1876;
  wire  _T_1877;
  wire  _T_1878;
  wire  _T_1879;
  wire  _T_1880;
  wire  _T_1881;
  wire  _T_1882;
  wire  _T_1883;
  wire  _T_1884;
  wire  _T_1885;
  wire  _T_1886;
  wire  _T_1887;
  wire  _T_1888;
  wire  _T_1889;
  wire  _T_1890;
  wire  _T_1891;
  wire  _T_1892;
  wire  _T_1893;
  wire  _T_1894;
  wire  _T_1895;
  wire  _T_1896;
  wire  _T_1897;
  wire  _T_1898;
  wire  _T_1899;
  wire  _T_1900;
  wire  _T_1901;
  wire  _T_1902;
  wire  _T_1903;
  wire  _T_1904;
  wire  _T_1905;
  wire  _T_1906;
  wire  _T_1907;
  wire  _T_1908;
  wire  _T_1909;
  wire  _T_1910;
  wire  _T_1911;
  wire  _T_1912;
  wire  _T_1913;
  wire  _T_1914;
  wire  _T_1915;
  wire  _T_1916;
  wire  _T_1917;
  wire  _T_1918;
  wire  _T_1919;
  wire  _T_1920;
  wire  _T_1921;
  wire  _T_1922;
  wire  _T_1923;
  wire  _T_1924;
  wire  _T_1925;
  wire  _T_1926;
  wire  _T_1927;
  wire  _T_1928;
  wire  _T_1929;
  wire  _T_1930;
  wire  _T_1931;
  wire  _T_1932;
  wire  _T_1933;
  wire  _T_1934;
  wire  _T_1935;
  wire  _T_1936;
  wire  _T_1937;
  wire  _T_1938;
  wire  _T_1939;
  wire  _T_1941;
  reg  _T_1944;
  reg [31:0] _RAND_4;
  wire  _T_1949;
  wire  _T_1950;
  wire  _T_1951;
  wire  _T_1952;
  wire  _T_1953;
  wire [1:0] _T_1954;
  wire  _T_1955;
  wire [1:0] _T_1956;
  wire [1:0] _T_1957;
  wire  _T_1958;
  wire  _T_1960;
  wire  _T_1963;
  wire  _T_1965;
  wire  _T_1967;
  wire  _T_1969;
  wire  _T_1971;
  wire  _T_1972;
  wire  _T_1974;
  wire  _T_1976;
  reg  _T_1986;
  reg [31:0] _RAND_5;
  wire  _T_1992;
  wire  _T_1993;
  wire  _T_1995;
  wire [1:0] _T_1996;
  wire  _T_1997;
  wire [1:0] _T_1998;
  wire [1:0] _T_1999;
  wire  _T_2000;
  wire  _T_2002;
  wire  _T_2005;
  wire  _T_2007;
  wire  _T_2009;
  wire  _T_2011;
  wire  _T_2013;
  wire  _T_2014;
  wire  _T_2016;
  wire  _T_2018;
  reg  _T_2028;
  reg [31:0] _RAND_6;
  wire  _T_2034;
  wire  _T_2035;
  wire  _T_2037;
  wire [1:0] _T_2038;
  wire  _T_2039;
  wire [1:0] _T_2040;
  wire [1:0] _T_2041;
  wire  _T_2042;
  wire  _T_2044;
  wire  _T_2047;
  wire  _T_2049;
  wire  _T_2051;
  wire  _T_2053;
  wire  _T_2055;
  wire  _T_2056;
  wire  _T_2058;
  wire  _T_2060;
  reg  _T_2070;
  reg [31:0] _RAND_7;
  wire  _T_2076;
  wire  _T_2077;
  wire  _T_2079;
  wire [1:0] _T_2080;
  wire  _T_2081;
  wire [1:0] _T_2082;
  wire [1:0] _T_2083;
  wire  _T_2084;
  wire  _T_2086;
  wire  _T_2089;
  wire  _T_2091;
  wire  _T_2093;
  wire  _T_2095;
  wire  _T_2097;
  wire  _T_2098;
  wire  _T_2100;
  wire  _T_2102;
  reg  _T_2112;
  reg [31:0] _RAND_8;
  wire  _T_2118;
  wire  _T_2119;
  wire  _T_2121;
  wire [1:0] _T_2122;
  wire  _T_2123;
  wire [1:0] _T_2124;
  wire [1:0] _T_2125;
  wire  _T_2126;
  wire  _T_2128;
  wire  _T_2131;
  wire  _T_2133;
  wire  _T_2135;
  wire  _T_2137;
  wire  _T_2139;
  wire  _T_2140;
  wire  _T_2142;
  wire  _T_2144;
  reg  _T_2154;
  reg [31:0] _RAND_9;
  wire  _T_2160;
  wire  _T_2161;
  wire  _T_2163;
  wire [1:0] _T_2164;
  wire  _T_2165;
  wire [1:0] _T_2166;
  wire [1:0] _T_2167;
  wire  _T_2168;
  wire  _T_2170;
  wire  _T_2173;
  wire  _T_2175;
  wire  _T_2177;
  wire  _T_2179;
  wire  _T_2181;
  wire  _T_2182;
  wire  _T_2184;
  wire  _T_2186;
  reg  _T_2196;
  reg [31:0] _RAND_10;
  wire  _T_2202;
  wire  _T_2203;
  wire  _T_2205;
  wire [1:0] _T_2206;
  wire  _T_2207;
  wire [1:0] _T_2208;
  wire [1:0] _T_2209;
  wire  _T_2210;
  wire  _T_2212;
  wire  _T_2215;
  wire  _T_2217;
  wire  _T_2219;
  wire  _T_2221;
  wire  _T_2223;
  wire  _T_2224;
  wire  _T_2226;
  wire  _T_2228;
  reg  _T_2238;
  reg [31:0] _RAND_11;
  wire  _T_2244;
  wire  _T_2245;
  wire  _T_2247;
  wire [1:0] _T_2248;
  wire  _T_2249;
  wire [1:0] _T_2250;
  wire [1:0] _T_2251;
  wire  _T_2252;
  wire  _T_2254;
  wire  _T_2257;
  wire  _T_2259;
  wire  _T_2261;
  wire  _T_2263;
  wire  _T_2265;
  wire  _T_2266;
  wire  _T_2268;
  wire  _T_2270;
  reg  _T_2280;
  reg [31:0] _RAND_12;
  wire  _T_2286;
  wire  _T_2287;
  wire  _T_2289;
  wire [1:0] _T_2290;
  wire  _T_2291;
  wire [1:0] _T_2292;
  wire [1:0] _T_2293;
  wire  _T_2294;
  wire  _T_2296;
  wire  _T_2299;
  wire  _T_2301;
  wire  _T_2303;
  wire  _T_2305;
  wire  _T_2307;
  wire  _T_2308;
  wire  _T_2310;
  wire  _T_2312;
  reg  _T_2322;
  reg [31:0] _RAND_13;
  wire  _T_2328;
  wire  _T_2329;
  wire  _T_2331;
  wire [1:0] _T_2332;
  wire  _T_2333;
  wire [1:0] _T_2334;
  wire [1:0] _T_2335;
  wire  _T_2336;
  wire  _T_2338;
  wire  _T_2341;
  wire  _T_2343;
  wire  _T_2345;
  wire  _T_2347;
  wire  _T_2349;
  wire  _T_2350;
  wire  _T_2352;
  wire  _T_2354;
  reg  _T_2364;
  reg [31:0] _RAND_14;
  wire  _T_2370;
  wire  _T_2371;
  wire  _T_2373;
  wire [1:0] _T_2374;
  wire  _T_2375;
  wire [1:0] _T_2376;
  wire [1:0] _T_2377;
  wire  _T_2378;
  wire  _T_2380;
  wire  _T_2383;
  wire  _T_2385;
  wire  _T_2387;
  wire  _T_2389;
  wire  _T_2391;
  wire  _T_2392;
  wire  _T_2394;
  wire  _T_2396;
  reg  _T_2406;
  reg [31:0] _RAND_15;
  wire  _T_2412;
  wire  _T_2413;
  wire  _T_2415;
  wire [1:0] _T_2416;
  wire  _T_2417;
  wire [1:0] _T_2418;
  wire [1:0] _T_2419;
  wire  _T_2420;
  wire  _T_2422;
  wire  _T_2425;
  wire  _T_2427;
  wire  _T_2429;
  wire  _T_2431;
  wire  _T_2433;
  wire  _T_2434;
  wire  _T_2436;
  wire  _T_2438;
  reg  _T_2448;
  reg [31:0] _RAND_16;
  wire  _T_2454;
  wire  _T_2455;
  wire  _T_2457;
  wire [1:0] _T_2458;
  wire  _T_2459;
  wire [1:0] _T_2460;
  wire [1:0] _T_2461;
  wire  _T_2462;
  wire  _T_2464;
  wire  _T_2467;
  wire  _T_2469;
  wire  _T_2471;
  wire  _T_2473;
  wire  _T_2475;
  wire  _T_2476;
  wire  _T_2478;
  wire  _T_2480;
  reg  _T_2490;
  reg [31:0] _RAND_17;
  wire  _T_2496;
  wire  _T_2497;
  wire  _T_2499;
  wire [1:0] _T_2500;
  wire  _T_2501;
  wire [1:0] _T_2502;
  wire [1:0] _T_2503;
  wire  _T_2504;
  wire  _T_2506;
  wire  _T_2509;
  wire  _T_2511;
  wire  _T_2513;
  wire  _T_2515;
  wire  _T_2517;
  wire  _T_2518;
  wire  _T_2520;
  wire  _T_2522;
  reg  _T_2532;
  reg [31:0] _RAND_18;
  wire  _T_2538;
  wire  _T_2539;
  wire  _T_2541;
  wire [1:0] _T_2542;
  wire  _T_2543;
  wire [1:0] _T_2544;
  wire [1:0] _T_2545;
  wire  _T_2546;
  wire  _T_2548;
  wire  _T_2551;
  wire  _T_2553;
  wire  _T_2555;
  wire  _T_2557;
  wire  _T_2559;
  wire  _T_2560;
  wire  _T_2562;
  wire  _T_2564;
  reg  _T_2574;
  reg [31:0] _RAND_19;
  wire  _T_2580;
  wire  _T_2581;
  wire  _T_2583;
  wire [1:0] _T_2584;
  wire  _T_2585;
  wire [1:0] _T_2586;
  wire [1:0] _T_2587;
  wire  _T_2588;
  wire  _T_2590;
  wire  _T_2593;
  wire  _T_2595;
  wire  _T_2597;
  wire  _T_2599;
  wire  _T_2601;
  wire  _T_2602;
  wire  _T_2604;
  wire  _T_2606;
  reg  _T_2616;
  reg [31:0] _RAND_20;
  wire  _T_2622;
  wire  _T_2623;
  wire  _T_2625;
  wire [1:0] _T_2626;
  wire  _T_2627;
  wire [1:0] _T_2628;
  wire [1:0] _T_2629;
  wire  _T_2630;
  wire  _T_2632;
  wire  _T_2635;
  wire  _T_2637;
  wire  _T_2639;
  wire  _T_2641;
  wire  _T_2643;
  wire  _T_2644;
  wire  _T_2646;
  wire  _T_2648;
  reg  _T_2658;
  reg [31:0] _RAND_21;
  wire  _T_2664;
  wire  _T_2665;
  wire  _T_2667;
  wire [1:0] _T_2668;
  wire  _T_2669;
  wire [1:0] _T_2670;
  wire [1:0] _T_2671;
  wire  _T_2672;
  wire  _T_2674;
  wire  _T_2677;
  wire  _T_2679;
  wire  _T_2681;
  wire  _T_2683;
  wire  _T_2685;
  wire  _T_2686;
  wire  _T_2688;
  wire  _T_2690;
  reg  _T_2700;
  reg [31:0] _RAND_22;
  wire  _T_2706;
  wire  _T_2707;
  wire  _T_2709;
  wire [1:0] _T_2710;
  wire  _T_2711;
  wire [1:0] _T_2712;
  wire [1:0] _T_2713;
  wire  _T_2714;
  wire  _T_2716;
  wire  _T_2719;
  wire  _T_2721;
  wire  _T_2723;
  wire  _T_2725;
  wire  _T_2727;
  wire  _T_2728;
  wire  _T_2730;
  wire  _T_2732;
  reg  _T_2742;
  reg [31:0] _RAND_23;
  wire  _T_2748;
  wire  _T_2749;
  wire  _T_2751;
  wire [1:0] _T_2752;
  wire  _T_2753;
  wire [1:0] _T_2754;
  wire [1:0] _T_2755;
  wire  _T_2756;
  wire  _T_2758;
  wire  _T_2761;
  wire  _T_2763;
  wire  _T_2765;
  wire  _T_2767;
  wire  _T_2769;
  wire  _T_2770;
  wire  _T_2772;
  wire  _T_2774;
  reg  _T_2784;
  reg [31:0] _RAND_24;
  wire  _T_2790;
  wire  _T_2791;
  wire  _T_2793;
  wire [1:0] _T_2794;
  wire  _T_2795;
  wire [1:0] _T_2796;
  wire [1:0] _T_2797;
  wire  _T_2798;
  wire  _T_2800;
  wire  _T_2803;
  wire  _T_2805;
  wire  _T_2807;
  wire  _T_2809;
  wire  _T_2811;
  wire  _T_2812;
  wire  _T_2814;
  wire  _T_2816;
  reg  _T_2826;
  reg [31:0] _RAND_25;
  wire  _T_2832;
  wire  _T_2833;
  wire  _T_2835;
  wire [1:0] _T_2836;
  wire  _T_2837;
  wire [1:0] _T_2838;
  wire [1:0] _T_2839;
  wire  _T_2840;
  wire  _T_2842;
  wire  _T_2845;
  wire  _T_2847;
  wire  _T_2849;
  wire  _T_2851;
  wire  _T_2853;
  wire  _T_2854;
  wire  _T_2856;
  wire  _T_2858;
  reg  _T_2868;
  reg [31:0] _RAND_26;
  wire  _T_2874;
  wire  _T_2875;
  wire  _T_2877;
  wire [1:0] _T_2878;
  wire  _T_2879;
  wire [1:0] _T_2880;
  wire [1:0] _T_2881;
  wire  _T_2882;
  wire  _T_2884;
  wire  _T_2887;
  wire  _T_2889;
  wire  _T_2891;
  wire  _T_2893;
  wire  _T_2895;
  wire  _T_2896;
  wire  _T_2898;
  wire  _T_2900;
  reg  _T_2910;
  reg [31:0] _RAND_27;
  wire  _T_2916;
  wire  _T_2917;
  wire  _T_2919;
  wire [1:0] _T_2920;
  wire  _T_2921;
  wire [1:0] _T_2922;
  wire [1:0] _T_2923;
  wire  _T_2924;
  wire  _T_2926;
  wire  _T_2929;
  wire  _T_2931;
  wire  _T_2933;
  wire  _T_2935;
  wire  _T_2937;
  wire  _T_2938;
  wire  _T_2940;
  wire  _T_2942;
  reg  _T_2952;
  reg [31:0] _RAND_28;
  wire  _T_2958;
  wire  _T_2959;
  wire  _T_2961;
  wire [1:0] _T_2962;
  wire  _T_2963;
  wire [1:0] _T_2964;
  wire [1:0] _T_2965;
  wire  _T_2966;
  wire  _T_2968;
  wire  _T_2971;
  wire  _T_2973;
  wire  _T_2975;
  wire  _T_2977;
  wire  _T_2979;
  wire  _T_2980;
  wire  _T_2982;
  wire  _T_2984;
  reg  _T_2994;
  reg [31:0] _RAND_29;
  wire  _T_3000;
  wire  _T_3001;
  wire  _T_3003;
  wire [1:0] _T_3004;
  wire  _T_3005;
  wire [1:0] _T_3006;
  wire [1:0] _T_3007;
  wire  _T_3008;
  wire  _T_3010;
  wire  _T_3013;
  wire  _T_3015;
  wire  _T_3017;
  wire  _T_3019;
  wire  _T_3021;
  wire  _T_3022;
  wire  _T_3024;
  wire  _T_3026;
  reg  _T_3036;
  reg [31:0] _RAND_30;
  wire  _T_3042;
  wire  _T_3043;
  wire  _T_3045;
  wire [1:0] _T_3046;
  wire  _T_3047;
  wire [1:0] _T_3048;
  wire [1:0] _T_3049;
  wire  _T_3050;
  wire  _T_3052;
  wire  _T_3055;
  wire  _T_3057;
  wire  _T_3059;
  wire  _T_3061;
  wire  _T_3063;
  wire  _T_3064;
  wire  _T_3066;
  wire  _T_3068;
  reg  _T_3078;
  reg [31:0] _RAND_31;
  wire  _T_3084;
  wire  _T_3085;
  wire  _T_3087;
  wire [1:0] _T_3088;
  wire  _T_3089;
  wire [1:0] _T_3090;
  wire [1:0] _T_3091;
  wire  _T_3092;
  wire  _T_3094;
  wire  _T_3097;
  wire  _T_3099;
  wire  _T_3101;
  wire  _T_3103;
  wire  _T_3105;
  wire  _T_3106;
  wire  _T_3108;
  wire  _T_3110;
  reg  _T_3120;
  reg [31:0] _RAND_32;
  wire  _T_3126;
  wire  _T_3127;
  wire  _T_3129;
  wire [1:0] _T_3130;
  wire  _T_3131;
  wire [1:0] _T_3132;
  wire [1:0] _T_3133;
  wire  _T_3134;
  wire  _T_3136;
  wire  _T_3139;
  wire  _T_3141;
  wire  _T_3143;
  wire  _T_3145;
  wire  _T_3147;
  wire  _T_3148;
  wire  _T_3150;
  wire  _T_3152;
  reg  _T_3162;
  reg [31:0] _RAND_33;
  wire  _T_3168;
  wire  _T_3169;
  wire  _T_3171;
  wire [1:0] _T_3172;
  wire  _T_3173;
  wire [1:0] _T_3174;
  wire [1:0] _T_3175;
  wire  _T_3176;
  wire  _T_3178;
  wire  _T_3181;
  wire  _T_3183;
  wire  _T_3185;
  wire  _T_3187;
  wire  _T_3189;
  wire  _T_3190;
  wire  _T_3192;
  wire  _T_3194;
  reg  _T_3204;
  reg [31:0] _RAND_34;
  wire  _T_3210;
  wire  _T_3211;
  wire  _T_3213;
  wire [1:0] _T_3214;
  wire  _T_3215;
  wire [1:0] _T_3216;
  wire [1:0] _T_3217;
  wire  _T_3218;
  wire  _T_3220;
  wire  _T_3223;
  wire  _T_3225;
  wire  _T_3227;
  wire  _T_3229;
  wire  _T_3231;
  wire  _T_3232;
  wire  _T_3234;
  wire  _T_3236;
  reg  _T_3246;
  reg [31:0] _RAND_35;
  wire  _T_3252;
  wire  _T_3253;
  wire  _T_3255;
  wire [1:0] _T_3256;
  wire  _T_3257;
  wire [1:0] _T_3258;
  wire [1:0] _T_3259;
  wire  _T_3260;
  wire  _T_3262;
  wire  _T_3265;
  wire  _T_3267;
  wire  _T_3269;
  wire  _T_3271;
  wire  _T_3273;
  wire  _T_3274;
  wire  _T_3276;
  wire  _T_3278;
  reg  _T_3288;
  reg [31:0] _RAND_36;
  wire  _T_3294;
  wire  _T_3295;
  wire  _T_3297;
  wire [1:0] _T_3298;
  wire  _T_3299;
  wire [1:0] _T_3300;
  wire [1:0] _T_3301;
  wire  _T_3302;
  wire  _T_3304;
  wire  _T_3307;
  wire  _T_3309;
  wire  _T_3311;
  wire  _T_3313;
  wire  _T_3315;
  wire  _T_3316;
  wire  _T_3318;
  wire  _T_3320;
  reg  _T_3330;
  reg [31:0] _RAND_37;
  wire  _T_3336;
  wire  _T_3337;
  wire  _T_3339;
  wire [1:0] _T_3340;
  wire  _T_3341;
  wire [1:0] _T_3342;
  wire [1:0] _T_3343;
  wire  _T_3344;
  wire  _T_3346;
  wire  _T_3349;
  wire  _T_3351;
  wire  _T_3353;
  wire  _T_3355;
  wire  _T_3357;
  wire  _T_3358;
  wire  _T_3360;
  wire  _T_3362;
  reg  _T_3372;
  reg [31:0] _RAND_38;
  wire  _T_3378;
  wire  _T_3379;
  wire  _T_3381;
  wire [1:0] _T_3382;
  wire  _T_3383;
  wire [1:0] _T_3384;
  wire [1:0] _T_3385;
  wire  _T_3386;
  wire  _T_3388;
  wire  _T_3391;
  wire  _T_3393;
  wire  _T_3395;
  wire  _T_3397;
  wire  _T_3399;
  wire  _T_3400;
  wire  _T_3402;
  wire  _T_3404;
  reg  _T_3414;
  reg [31:0] _RAND_39;
  wire  _T_3420;
  wire  _T_3421;
  wire  _T_3423;
  wire [1:0] _T_3424;
  wire  _T_3425;
  wire [1:0] _T_3426;
  wire [1:0] _T_3427;
  wire  _T_3428;
  wire  _T_3430;
  wire  _T_3433;
  wire  _T_3435;
  wire  _T_3437;
  wire  _T_3439;
  wire  _T_3441;
  wire  _T_3442;
  wire  _T_3444;
  wire  _T_3446;
  reg  _T_3456;
  reg [31:0] _RAND_40;
  wire  _T_3462;
  wire  _T_3463;
  wire  _T_3465;
  wire [1:0] _T_3466;
  wire  _T_3467;
  wire [1:0] _T_3468;
  wire [1:0] _T_3469;
  wire  _T_3470;
  wire  _T_3472;
  wire  _T_3475;
  wire  _T_3477;
  wire  _T_3479;
  wire  _T_3481;
  wire  _T_3483;
  wire  _T_3484;
  wire  _T_3486;
  wire  _T_3488;
  reg  _T_3498;
  reg [31:0] _RAND_41;
  wire  _T_3504;
  wire  _T_3505;
  wire  _T_3507;
  wire [1:0] _T_3508;
  wire  _T_3509;
  wire [1:0] _T_3510;
  wire [1:0] _T_3511;
  wire  _T_3512;
  wire  _T_3514;
  wire  _T_3517;
  wire  _T_3519;
  wire  _T_3521;
  wire  _T_3523;
  wire  _T_3525;
  wire  _T_3526;
  wire  _T_3528;
  wire  _T_3530;
  reg  _T_3540;
  reg [31:0] _RAND_42;
  wire  _T_3546;
  wire  _T_3547;
  wire  _T_3549;
  wire [1:0] _T_3550;
  wire  _T_3551;
  wire [1:0] _T_3552;
  wire [1:0] _T_3553;
  wire  _T_3554;
  wire  _T_3556;
  wire  _T_3559;
  wire  _T_3561;
  wire  _T_3563;
  wire  _T_3565;
  wire  _T_3567;
  wire  _T_3568;
  wire  _T_3570;
  wire  _T_3572;
  reg  _T_3582;
  reg [31:0] _RAND_43;
  wire  _T_3588;
  wire  _T_3589;
  wire  _T_3591;
  wire [1:0] _T_3592;
  wire  _T_3593;
  wire [1:0] _T_3594;
  wire [1:0] _T_3595;
  wire  _T_3596;
  wire  _T_3598;
  wire  _T_3601;
  wire  _T_3603;
  wire  _T_3605;
  wire  _T_3607;
  wire  _T_3609;
  wire  _T_3610;
  wire  _T_3612;
  wire  _T_3614;
  reg  _T_3624;
  reg [31:0] _RAND_44;
  wire  _T_3630;
  wire  _T_3631;
  wire  _T_3633;
  wire [1:0] _T_3634;
  wire  _T_3635;
  wire [1:0] _T_3636;
  wire [1:0] _T_3637;
  wire  _T_3638;
  wire  _T_3640;
  wire  _T_3643;
  wire  _T_3645;
  wire  _T_3647;
  wire  _T_3649;
  wire  _T_3651;
  wire  _T_3652;
  wire  _T_3654;
  wire  _T_3656;
  reg  _T_3666;
  reg [31:0] _RAND_45;
  wire  _T_3672;
  wire  _T_3673;
  wire  _T_3675;
  wire [1:0] _T_3676;
  wire  _T_3677;
  wire [1:0] _T_3678;
  wire [1:0] _T_3679;
  wire  _T_3680;
  wire  _T_3682;
  wire  _T_3685;
  wire  _T_3687;
  wire  _T_3689;
  wire  _T_3691;
  wire  _T_3693;
  wire  _T_3694;
  wire  _T_3696;
  wire  _T_3698;
  reg  _T_3708;
  reg [31:0] _RAND_46;
  wire  _T_3714;
  wire  _T_3715;
  wire  _T_3717;
  wire [1:0] _T_3718;
  wire  _T_3719;
  wire [1:0] _T_3720;
  wire [1:0] _T_3721;
  wire  _T_3722;
  wire  _T_3724;
  wire  _T_3727;
  wire  _T_3729;
  wire  _T_3731;
  wire  _T_3733;
  wire  _T_3735;
  wire  _T_3736;
  wire  _T_3738;
  wire  _T_3740;
  reg  _T_3750;
  reg [31:0] _RAND_47;
  wire  _T_3756;
  wire  _T_3757;
  wire  _T_3759;
  wire [1:0] _T_3760;
  wire  _T_3761;
  wire [1:0] _T_3762;
  wire [1:0] _T_3763;
  wire  _T_3764;
  wire  _T_3766;
  wire  _T_3769;
  wire  _T_3771;
  wire  _T_3773;
  wire  _T_3775;
  wire  _T_3777;
  wire  _T_3778;
  wire  _T_3780;
  wire  _T_3782;
  reg  _T_3792;
  reg [31:0] _RAND_48;
  wire  _T_3798;
  wire  _T_3799;
  wire  _T_3801;
  wire [1:0] _T_3802;
  wire  _T_3803;
  wire [1:0] _T_3804;
  wire [1:0] _T_3805;
  wire  _T_3806;
  wire  _T_3808;
  wire  _T_3811;
  wire  _T_3813;
  wire  _T_3815;
  wire  _T_3817;
  wire  _T_3819;
  wire  _T_3820;
  wire  _T_3822;
  wire  _T_3824;
  reg  _T_3834;
  reg [31:0] _RAND_49;
  wire  _T_3840;
  wire  _T_3841;
  wire  _T_3843;
  wire [1:0] _T_3844;
  wire  _T_3845;
  wire [1:0] _T_3846;
  wire [1:0] _T_3847;
  wire  _T_3848;
  wire  _T_3850;
  wire  _T_3853;
  wire  _T_3855;
  wire  _T_3857;
  wire  _T_3859;
  wire  _T_3861;
  wire  _T_3862;
  wire  _T_3864;
  wire  _T_3866;
  reg  _T_3876;
  reg [31:0] _RAND_50;
  wire  _T_3882;
  wire  _T_3883;
  wire  _T_3885;
  wire [1:0] _T_3886;
  wire  _T_3887;
  wire [1:0] _T_3888;
  wire [1:0] _T_3889;
  wire  _T_3890;
  wire  _T_3892;
  wire  _T_3895;
  wire  _T_3897;
  wire  _T_3899;
  wire  _T_3901;
  wire  _T_3903;
  wire  _T_3904;
  wire  _T_3906;
  wire  _T_3908;
  reg  _T_3918;
  reg [31:0] _RAND_51;
  wire  _T_3924;
  wire  _T_3925;
  wire  _T_3927;
  wire [1:0] _T_3928;
  wire  _T_3929;
  wire [1:0] _T_3930;
  wire [1:0] _T_3931;
  wire  _T_3932;
  wire  _T_3934;
  wire  _T_3937;
  wire  _T_3939;
  wire  _T_3941;
  wire  _T_3943;
  wire  _T_3945;
  wire  _T_3946;
  wire  _T_3948;
  wire  _T_3950;
  reg  _T_3960;
  reg [31:0] _RAND_52;
  wire  _T_3966;
  wire  _T_3967;
  wire  _T_3969;
  wire [1:0] _T_3970;
  wire  _T_3971;
  wire [1:0] _T_3972;
  wire [1:0] _T_3973;
  wire  _T_3974;
  wire  _T_3976;
  wire  _T_3979;
  wire  _T_3981;
  wire  _T_3983;
  wire  _T_3985;
  wire  _T_3987;
  wire  _T_3988;
  wire  _T_3990;
  wire  _T_3992;
  reg  _T_4002;
  reg [31:0] _RAND_53;
  wire  _T_4008;
  wire  _T_4009;
  wire  _T_4011;
  wire [1:0] _T_4012;
  wire  _T_4013;
  wire [1:0] _T_4014;
  wire [1:0] _T_4015;
  wire  _T_4016;
  wire  _T_4018;
  wire  _T_4021;
  wire  _T_4023;
  wire  _T_4025;
  wire  _T_4027;
  wire  _T_4029;
  wire  _T_4030;
  wire  _T_4032;
  wire  _T_4034;
  reg  _T_4044;
  reg [31:0] _RAND_54;
  wire  _T_4050;
  wire  _T_4051;
  wire  _T_4053;
  wire [1:0] _T_4054;
  wire  _T_4055;
  wire [1:0] _T_4056;
  wire [1:0] _T_4057;
  wire  _T_4058;
  wire  _T_4060;
  wire  _T_4063;
  wire  _T_4065;
  wire  _T_4067;
  wire  _T_4069;
  wire  _T_4071;
  wire  _T_4072;
  wire  _T_4074;
  wire  _T_4076;
  reg  _T_4086;
  reg [31:0] _RAND_55;
  wire  _T_4092;
  wire  _T_4093;
  wire  _T_4095;
  wire [1:0] _T_4096;
  wire  _T_4097;
  wire [1:0] _T_4098;
  wire [1:0] _T_4099;
  wire  _T_4100;
  wire  _T_4102;
  wire  _T_4105;
  wire  _T_4107;
  wire  _T_4109;
  wire  _T_4111;
  wire  _T_4113;
  wire  _T_4114;
  wire  _T_4116;
  wire  _T_4118;
  reg  _T_4128;
  reg [31:0] _RAND_56;
  wire  _T_4134;
  wire  _T_4135;
  wire  _T_4137;
  wire [1:0] _T_4138;
  wire  _T_4139;
  wire [1:0] _T_4140;
  wire [1:0] _T_4141;
  wire  _T_4142;
  wire  _T_4144;
  wire  _T_4147;
  wire  _T_4149;
  wire  _T_4151;
  wire  _T_4153;
  wire  _T_4155;
  wire  _T_4156;
  wire  _T_4158;
  wire  _T_4160;
  reg  _T_4170;
  reg [31:0] _RAND_57;
  wire  _T_4176;
  wire  _T_4177;
  wire  _T_4179;
  wire [1:0] _T_4180;
  wire  _T_4181;
  wire [1:0] _T_4182;
  wire [1:0] _T_4183;
  wire  _T_4184;
  wire  _T_4186;
  wire  _T_4189;
  wire  _T_4191;
  wire  _T_4193;
  wire  _T_4195;
  wire  _T_4197;
  wire  _T_4198;
  wire  _T_4200;
  wire  _T_4202;
  reg  _T_4212;
  reg [31:0] _RAND_58;
  wire  _T_4218;
  wire  _T_4219;
  wire  _T_4221;
  wire [1:0] _T_4222;
  wire  _T_4223;
  wire [1:0] _T_4224;
  wire [1:0] _T_4225;
  wire  _T_4226;
  wire  _T_4228;
  wire  _T_4231;
  wire  _T_4233;
  wire  _T_4235;
  wire  _T_4237;
  wire  _T_4239;
  wire  _T_4240;
  wire  _T_4242;
  wire  _T_4244;
  reg  _T_4254;
  reg [31:0] _RAND_59;
  wire  _T_4260;
  wire  _T_4261;
  wire  _T_4263;
  wire [1:0] _T_4264;
  wire  _T_4265;
  wire [1:0] _T_4266;
  wire [1:0] _T_4267;
  wire  _T_4268;
  wire  _T_4270;
  wire  _T_4273;
  wire  _T_4275;
  wire  _T_4277;
  wire  _T_4279;
  wire  _T_4281;
  wire  _T_4282;
  wire  _T_4284;
  wire  _T_4286;
  reg  _T_4296;
  reg [31:0] _RAND_60;
  wire  _T_4302;
  wire  _T_4303;
  wire  _T_4305;
  wire [1:0] _T_4306;
  wire  _T_4307;
  wire [1:0] _T_4308;
  wire [1:0] _T_4309;
  wire  _T_4310;
  wire  _T_4312;
  wire  _T_4315;
  wire  _T_4317;
  wire  _T_4319;
  wire  _T_4321;
  wire  _T_4323;
  wire  _T_4324;
  wire  _T_4326;
  wire  _T_4328;
  reg  _T_4338;
  reg [31:0] _RAND_61;
  wire  _T_4344;
  wire  _T_4345;
  wire  _T_4347;
  wire [1:0] _T_4348;
  wire  _T_4349;
  wire [1:0] _T_4350;
  wire [1:0] _T_4351;
  wire  _T_4352;
  wire  _T_4354;
  wire  _T_4357;
  wire  _T_4359;
  wire  _T_4361;
  wire  _T_4363;
  wire  _T_4365;
  wire  _T_4366;
  wire  _T_4368;
  wire  _T_4370;
  reg  _T_4380;
  reg [31:0] _RAND_62;
  wire  _T_4386;
  wire  _T_4387;
  wire  _T_4389;
  wire [1:0] _T_4390;
  wire  _T_4391;
  wire [1:0] _T_4392;
  wire [1:0] _T_4393;
  wire  _T_4394;
  wire  _T_4396;
  wire  _T_4399;
  wire  _T_4401;
  wire  _T_4403;
  wire  _T_4405;
  wire  _T_4407;
  wire  _T_4408;
  wire  _T_4410;
  wire  _T_4412;
  reg  _T_4422;
  reg [31:0] _RAND_63;
  wire  _T_4428;
  wire  _T_4429;
  wire  _T_4431;
  wire [1:0] _T_4432;
  wire  _T_4433;
  wire [1:0] _T_4434;
  wire [1:0] _T_4435;
  wire  _T_4436;
  wire  _T_4438;
  wire  _T_4441;
  wire  _T_4443;
  wire  _T_4445;
  wire  _T_4447;
  wire  _T_4449;
  wire  _T_4450;
  wire  _T_4452;
  wire  _T_4454;
  reg  _T_4464;
  reg [31:0] _RAND_64;
  wire  _T_4470;
  wire  _T_4471;
  wire  _T_4473;
  wire [1:0] _T_4474;
  wire  _T_4475;
  wire [1:0] _T_4476;
  wire [1:0] _T_4477;
  wire  _T_4478;
  wire  _T_4480;
  wire  _T_4483;
  wire  _T_4485;
  wire  _T_4487;
  wire  _T_4489;
  wire  _T_4491;
  wire  _T_4492;
  wire  _T_4494;
  wire  _T_4496;
  reg  _T_4506;
  reg [31:0] _RAND_65;
  wire  _T_4512;
  wire  _T_4513;
  wire  _T_4515;
  wire [1:0] _T_4516;
  wire  _T_4517;
  wire [1:0] _T_4518;
  wire [1:0] _T_4519;
  wire  _T_4520;
  wire  _T_4522;
  wire  _T_4525;
  wire  _T_4527;
  wire  _T_4529;
  wire  _T_4531;
  wire  _T_4533;
  wire  _T_4534;
  wire  _T_4536;
  wire  _T_4538;
  reg  _T_4548;
  reg [31:0] _RAND_66;
  wire  _T_4554;
  wire  _T_4555;
  wire  _T_4557;
  wire [1:0] _T_4558;
  wire  _T_4559;
  wire [1:0] _T_4560;
  wire [1:0] _T_4561;
  wire  _T_4562;
  wire  _T_4564;
  wire  _T_4567;
  wire  _T_4569;
  wire  _T_4571;
  wire  _T_4573;
  wire  _T_4575;
  wire  _T_4576;
  wire  _T_4578;
  wire  _T_4580;
  reg  _T_4590;
  reg [31:0] _RAND_67;
  wire  _T_4596;
  wire  _T_4597;
  wire  _T_4599;
  wire [1:0] _T_4600;
  wire  _T_4601;
  wire [1:0] _T_4602;
  wire [1:0] _T_4603;
  wire  _T_4604;
  wire  _T_4606;
  wire  _T_4609;
  wire  _T_4611;
  wire  _T_4613;
  wire  _T_4615;
  wire  _T_4617;
  wire  _T_4618;
  wire  _T_4620;
  wire  _T_4622;
  reg  _T_4632;
  reg [31:0] _RAND_68;
  wire  _T_4638;
  wire  _T_4639;
  wire  _T_4641;
  wire [1:0] _T_4642;
  wire  _T_4643;
  wire [1:0] _T_4644;
  wire [1:0] _T_4645;
  wire  _T_4646;
  wire  _T_4648;
  wire  _T_4651;
  wire  _T_4653;
  wire  _T_4655;
  wire  _T_4657;
  wire  _T_4659;
  wire  _T_4660;
  wire  _T_4662;
  wire  _T_4664;
  reg  _T_4674;
  reg [31:0] _RAND_69;
  wire  _T_4680;
  wire  _T_4681;
  wire  _T_4683;
  wire [1:0] _T_4684;
  wire  _T_4685;
  wire [1:0] _T_4686;
  wire [1:0] _T_4687;
  wire  _T_4688;
  wire  _T_4690;
  wire  _T_4693;
  wire  _T_4695;
  wire  _T_4697;
  wire  _T_4699;
  wire  _T_4701;
  wire  _T_4702;
  wire  _T_4704;
  wire  _T_4706;
  reg  _T_4716;
  reg [31:0] _RAND_70;
  wire  _T_4722;
  wire  _T_4723;
  wire  _T_4725;
  wire [1:0] _T_4726;
  wire  _T_4727;
  wire [1:0] _T_4728;
  wire [1:0] _T_4729;
  wire  _T_4730;
  wire  _T_4732;
  wire  _T_4735;
  wire  _T_4737;
  wire  _T_4739;
  wire  _T_4741;
  wire  _T_4743;
  wire  _T_4744;
  wire  _T_4746;
  wire  _T_4748;
  reg  _T_4758;
  reg [31:0] _RAND_71;
  wire  _T_4764;
  wire  _T_4765;
  wire  _T_4767;
  wire [1:0] _T_4768;
  wire  _T_4769;
  wire [1:0] _T_4770;
  wire [1:0] _T_4771;
  wire  _T_4772;
  wire  _T_4774;
  wire  _T_4777;
  wire  _T_4779;
  wire  _T_4781;
  wire  _T_4783;
  wire  _T_4785;
  wire  _T_4786;
  wire  _T_4788;
  wire  _T_4790;
  reg  _T_4800;
  reg [31:0] _RAND_72;
  wire  _T_4806;
  wire  _T_4807;
  wire  _T_4809;
  wire [1:0] _T_4810;
  wire  _T_4811;
  wire [1:0] _T_4812;
  wire [1:0] _T_4813;
  wire  _T_4814;
  wire  _T_4816;
  wire  _T_4819;
  wire  _T_4821;
  wire  _T_4823;
  wire  _T_4825;
  wire  _T_4827;
  wire  _T_4828;
  wire  _T_4830;
  wire  _T_4832;
  reg  _T_4842;
  reg [31:0] _RAND_73;
  wire  _T_4848;
  wire  _T_4849;
  wire  _T_4851;
  wire [1:0] _T_4852;
  wire  _T_4853;
  wire [1:0] _T_4854;
  wire [1:0] _T_4855;
  wire  _T_4856;
  wire  _T_4858;
  wire  _T_4861;
  wire  _T_4863;
  wire  _T_4865;
  wire  _T_4867;
  wire  _T_4869;
  wire  _T_4870;
  wire  _T_4872;
  wire  _T_4874;
  reg  _T_4884;
  reg [31:0] _RAND_74;
  wire  _T_4890;
  wire  _T_4891;
  wire  _T_4893;
  wire [1:0] _T_4894;
  wire  _T_4895;
  wire [1:0] _T_4896;
  wire [1:0] _T_4897;
  wire  _T_4898;
  wire  _T_4900;
  wire  _T_4903;
  wire  _T_4905;
  wire  _T_4907;
  wire  _T_4909;
  wire  _T_4911;
  wire  _T_4912;
  wire  _T_4914;
  wire  _T_4916;
  reg  _T_4926;
  reg [31:0] _RAND_75;
  wire  _T_4932;
  wire  _T_4933;
  wire  _T_4935;
  wire [1:0] _T_4936;
  wire  _T_4937;
  wire [1:0] _T_4938;
  wire [1:0] _T_4939;
  wire  _T_4940;
  wire  _T_4942;
  wire  _T_4945;
  wire  _T_4947;
  wire  _T_4949;
  wire  _T_4951;
  wire  _T_4953;
  wire  _T_4954;
  wire  _T_4956;
  wire  _T_4958;
  reg  _T_4968;
  reg [31:0] _RAND_76;
  wire  _T_4974;
  wire  _T_4975;
  wire  _T_4977;
  wire [1:0] _T_4978;
  wire  _T_4979;
  wire [1:0] _T_4980;
  wire [1:0] _T_4981;
  wire  _T_4982;
  wire  _T_4984;
  wire  _T_4987;
  wire  _T_4989;
  wire  _T_4991;
  wire  _T_4993;
  wire  _T_4995;
  wire  _T_4996;
  wire  _T_4998;
  wire  _T_5000;
  reg  _T_5010;
  reg [31:0] _RAND_77;
  wire  _T_5016;
  wire  _T_5017;
  wire  _T_5019;
  wire [1:0] _T_5020;
  wire  _T_5021;
  wire [1:0] _T_5022;
  wire [1:0] _T_5023;
  wire  _T_5024;
  wire  _T_5026;
  wire  _T_5029;
  wire  _T_5031;
  wire  _T_5033;
  wire  _T_5035;
  wire  _T_5037;
  wire  _T_5038;
  wire  _T_5040;
  wire  _T_5042;
  reg  _T_5052;
  reg [31:0] _RAND_78;
  wire  _T_5058;
  wire  _T_5059;
  wire  _T_5061;
  wire [1:0] _T_5062;
  wire  _T_5063;
  wire [1:0] _T_5064;
  wire [1:0] _T_5065;
  wire  _T_5066;
  wire  _T_5068;
  wire  _T_5071;
  wire  _T_5073;
  wire  _T_5075;
  wire  _T_5077;
  wire  _T_5079;
  wire  _T_5080;
  wire  _T_5082;
  wire  _T_5084;
  reg  _T_5094;
  reg [31:0] _RAND_79;
  wire  _T_5100;
  wire  _T_5101;
  wire  _T_5103;
  wire [1:0] _T_5104;
  wire  _T_5105;
  wire [1:0] _T_5106;
  wire [1:0] _T_5107;
  wire  _T_5108;
  wire  _T_5110;
  wire  _T_5113;
  wire  _T_5115;
  wire  _T_5117;
  wire  _T_5119;
  wire  _T_5121;
  wire  _T_5122;
  wire  _T_5124;
  wire  _T_5126;
  reg  _T_5136;
  reg [31:0] _RAND_80;
  wire  _T_5142;
  wire  _T_5143;
  wire  _T_5145;
  wire [1:0] _T_5146;
  wire  _T_5147;
  wire [1:0] _T_5148;
  wire [1:0] _T_5149;
  wire  _T_5150;
  wire  _T_5152;
  wire  _T_5155;
  wire  _T_5157;
  wire  _T_5159;
  wire  _T_5161;
  wire  _T_5163;
  wire  _T_5164;
  wire  _T_5166;
  wire  _T_5168;
  reg  _T_5178;
  reg [31:0] _RAND_81;
  wire  _T_5184;
  wire  _T_5185;
  wire  _T_5187;
  wire [1:0] _T_5188;
  wire  _T_5189;
  wire [1:0] _T_5190;
  wire [1:0] _T_5191;
  wire  _T_5192;
  wire  _T_5194;
  wire  _T_5197;
  wire  _T_5199;
  wire  _T_5201;
  wire  _T_5203;
  wire  _T_5205;
  wire  _T_5206;
  wire  _T_5208;
  wire  _T_5210;
  reg  _T_5220;
  reg [31:0] _RAND_82;
  wire  _T_5226;
  wire  _T_5227;
  wire  _T_5229;
  wire [1:0] _T_5230;
  wire  _T_5231;
  wire [1:0] _T_5232;
  wire [1:0] _T_5233;
  wire  _T_5234;
  wire  _T_5236;
  wire  _T_5239;
  wire  _T_5241;
  wire  _T_5243;
  wire  _T_5245;
  wire  _T_5247;
  wire  _T_5248;
  wire  _T_5250;
  wire  _T_5252;
  reg  _T_5262;
  reg [31:0] _RAND_83;
  wire  _T_5268;
  wire  _T_5269;
  wire  _T_5271;
  wire [1:0] _T_5272;
  wire  _T_5273;
  wire [1:0] _T_5274;
  wire [1:0] _T_5275;
  wire  _T_5276;
  wire  _T_5278;
  wire  _T_5281;
  wire  _T_5283;
  wire  _T_5285;
  wire  _T_5287;
  wire  _T_5289;
  wire  _T_5290;
  wire  _T_5292;
  wire  _T_5294;
  reg  _T_5304;
  reg [31:0] _RAND_84;
  wire  _T_5310;
  wire  _T_5311;
  wire  _T_5313;
  wire [1:0] _T_5314;
  wire  _T_5315;
  wire [1:0] _T_5316;
  wire [1:0] _T_5317;
  wire  _T_5318;
  wire  _T_5320;
  wire  _T_5323;
  wire  _T_5325;
  wire  _T_5327;
  wire  _T_5329;
  wire  _T_5331;
  wire  _T_5332;
  wire  _T_5334;
  wire  _T_5336;
  reg  _T_5346;
  reg [31:0] _RAND_85;
  wire  _T_5352;
  wire  _T_5353;
  wire  _T_5355;
  wire [1:0] _T_5356;
  wire  _T_5357;
  wire [1:0] _T_5358;
  wire [1:0] _T_5359;
  wire  _T_5360;
  wire  _T_5362;
  wire  _T_5365;
  wire  _T_5367;
  wire  _T_5369;
  wire  _T_5371;
  wire  _T_5373;
  wire  _T_5374;
  wire  _T_5376;
  wire  _T_5378;
  reg  _T_5388;
  reg [31:0] _RAND_86;
  wire  _T_5394;
  wire  _T_5395;
  wire  _T_5397;
  wire [1:0] _T_5398;
  wire  _T_5399;
  wire [1:0] _T_5400;
  wire [1:0] _T_5401;
  wire  _T_5402;
  wire  _T_5404;
  wire  _T_5407;
  wire  _T_5409;
  wire  _T_5411;
  wire  _T_5413;
  wire  _T_5415;
  wire  _T_5416;
  wire  _T_5418;
  wire  _T_5420;
  reg  _T_5430;
  reg [31:0] _RAND_87;
  wire  _T_5436;
  wire  _T_5437;
  wire  _T_5439;
  wire [1:0] _T_5440;
  wire  _T_5441;
  wire [1:0] _T_5442;
  wire [1:0] _T_5443;
  wire  _T_5444;
  wire  _T_5446;
  wire  _T_5449;
  wire  _T_5451;
  wire  _T_5453;
  wire  _T_5455;
  wire  _T_5457;
  wire  _T_5458;
  wire  _T_5460;
  wire  _T_5462;
  reg  _T_5472;
  reg [31:0] _RAND_88;
  wire  _T_5478;
  wire  _T_5479;
  wire  _T_5481;
  wire [1:0] _T_5482;
  wire  _T_5483;
  wire [1:0] _T_5484;
  wire [1:0] _T_5485;
  wire  _T_5486;
  wire  _T_5488;
  wire  _T_5491;
  wire  _T_5493;
  wire  _T_5495;
  wire  _T_5497;
  wire  _T_5499;
  wire  _T_5500;
  wire  _T_5502;
  wire  _T_5504;
  reg  _T_5514;
  reg [31:0] _RAND_89;
  wire  _T_5520;
  wire  _T_5521;
  wire  _T_5523;
  wire [1:0] _T_5524;
  wire  _T_5525;
  wire [1:0] _T_5526;
  wire [1:0] _T_5527;
  wire  _T_5528;
  wire  _T_5530;
  wire  _T_5533;
  wire  _T_5535;
  wire  _T_5537;
  wire  _T_5539;
  wire  _T_5541;
  wire  _T_5542;
  wire  _T_5544;
  wire  _T_5546;
  reg  _T_5556;
  reg [31:0] _RAND_90;
  wire  _T_5562;
  wire  _T_5563;
  wire  _T_5565;
  wire [1:0] _T_5566;
  wire  _T_5567;
  wire [1:0] _T_5568;
  wire [1:0] _T_5569;
  wire  _T_5570;
  wire  _T_5572;
  wire  _T_5575;
  wire  _T_5577;
  wire  _T_5579;
  wire  _T_5581;
  wire  _T_5583;
  wire  _T_5584;
  wire  _T_5586;
  wire  _T_5588;
  reg  _T_5598;
  reg [31:0] _RAND_91;
  wire  _T_5604;
  wire  _T_5605;
  wire  _T_5607;
  wire [1:0] _T_5608;
  wire  _T_5609;
  wire [1:0] _T_5610;
  wire [1:0] _T_5611;
  wire  _T_5612;
  wire  _T_5614;
  wire  _T_5617;
  wire  _T_5619;
  wire  _T_5621;
  wire  _T_5623;
  wire  _T_5625;
  wire  _T_5626;
  wire  _T_5628;
  wire  _T_5630;
  reg  _T_5640;
  reg [31:0] _RAND_92;
  wire  _T_5646;
  wire  _T_5647;
  wire  _T_5649;
  wire [1:0] _T_5650;
  wire  _T_5651;
  wire [1:0] _T_5652;
  wire [1:0] _T_5653;
  wire  _T_5654;
  wire  _T_5656;
  wire  _T_5659;
  wire  _T_5661;
  wire  _T_5663;
  wire  _T_5665;
  wire  _T_5667;
  wire  _T_5668;
  wire  _T_5670;
  wire  _T_5672;
  reg  _T_5682;
  reg [31:0] _RAND_93;
  wire  _T_5688;
  wire  _T_5689;
  wire  _T_5691;
  wire [1:0] _T_5692;
  wire  _T_5693;
  wire [1:0] _T_5694;
  wire [1:0] _T_5695;
  wire  _T_5696;
  wire  _T_5698;
  wire  _T_5701;
  wire  _T_5703;
  wire  _T_5705;
  wire  _T_5707;
  wire  _T_5709;
  wire  _T_5710;
  wire  _T_5712;
  wire  _T_5714;
  reg  _T_5724;
  reg [31:0] _RAND_94;
  wire  _T_5730;
  wire  _T_5731;
  wire  _T_5733;
  wire [1:0] _T_5734;
  wire  _T_5735;
  wire [1:0] _T_5736;
  wire [1:0] _T_5737;
  wire  _T_5738;
  wire  _T_5740;
  wire  _T_5743;
  wire  _T_5745;
  wire  _T_5747;
  wire  _T_5749;
  wire  _T_5751;
  wire  _T_5752;
  wire  _T_5754;
  wire  _T_5756;
  reg  _T_5766;
  reg [31:0] _RAND_95;
  wire  _T_5772;
  wire  _T_5773;
  wire  _T_5775;
  wire [1:0] _T_5776;
  wire  _T_5777;
  wire [1:0] _T_5778;
  wire [1:0] _T_5779;
  wire  _T_5780;
  wire  _T_5782;
  wire  _T_5785;
  wire  _T_5787;
  wire  _T_5789;
  wire  _T_5791;
  wire  _T_5793;
  wire  _T_5794;
  wire  _T_5796;
  wire  _T_5798;
  reg  _T_5808;
  reg [31:0] _RAND_96;
  wire  _T_5814;
  wire  _T_5815;
  wire  _T_5817;
  wire [1:0] _T_5818;
  wire  _T_5819;
  wire [1:0] _T_5820;
  wire [1:0] _T_5821;
  wire  _T_5822;
  wire  _T_5824;
  wire  _T_5827;
  wire  _T_5829;
  wire  _T_5831;
  wire  _T_5833;
  wire  _T_5835;
  wire  _T_5836;
  wire  _T_5838;
  wire  _T_5840;
  reg  _T_5850;
  reg [31:0] _RAND_97;
  wire  _T_5856;
  wire  _T_5857;
  wire  _T_5859;
  wire [1:0] _T_5860;
  wire  _T_5861;
  wire [1:0] _T_5862;
  wire [1:0] _T_5863;
  wire  _T_5864;
  wire  _T_5866;
  wire  _T_5869;
  wire  _T_5871;
  wire  _T_5873;
  wire  _T_5875;
  wire  _T_5877;
  wire  _T_5878;
  wire  _T_5880;
  wire  _T_5882;
  reg  _T_5892;
  reg [31:0] _RAND_98;
  wire  _T_5898;
  wire  _T_5899;
  wire  _T_5901;
  wire [1:0] _T_5902;
  wire  _T_5903;
  wire [1:0] _T_5904;
  wire [1:0] _T_5905;
  wire  _T_5906;
  wire  _T_5908;
  wire  _T_5911;
  wire  _T_5913;
  wire  _T_5915;
  wire  _T_5917;
  wire  _T_5919;
  wire  _T_5920;
  wire  _T_5922;
  wire  _T_5924;
  reg  _T_5934;
  reg [31:0] _RAND_99;
  wire  _T_5940;
  wire  _T_5941;
  wire  _T_5943;
  wire [1:0] _T_5944;
  wire  _T_5945;
  wire [1:0] _T_5946;
  wire [1:0] _T_5947;
  wire  _T_5948;
  wire  _T_5950;
  wire  _T_5953;
  wire  _T_5955;
  wire  _T_5957;
  wire  _T_5959;
  wire  _T_5961;
  wire  _T_5962;
  wire  _T_5964;
  wire  _T_5966;
  reg  _T_5976;
  reg [31:0] _RAND_100;
  wire  _T_5982;
  wire  _T_5983;
  wire  _T_5985;
  wire [1:0] _T_5986;
  wire  _T_5987;
  wire [1:0] _T_5988;
  wire [1:0] _T_5989;
  wire  _T_5990;
  wire  _T_5992;
  wire  _T_5995;
  wire  _T_5997;
  wire  _T_5999;
  wire  _T_6001;
  wire  _T_6003;
  wire  _T_6004;
  wire  _T_6006;
  wire  _T_6008;
  reg  _T_6018;
  reg [31:0] _RAND_101;
  wire  _T_6024;
  wire  _T_6025;
  wire  _T_6027;
  wire [1:0] _T_6028;
  wire  _T_6029;
  wire [1:0] _T_6030;
  wire [1:0] _T_6031;
  wire  _T_6032;
  wire  _T_6034;
  wire  _T_6037;
  wire  _T_6039;
  wire  _T_6041;
  wire  _T_6043;
  wire  _T_6045;
  wire  _T_6046;
  wire  _T_6048;
  wire  _T_6050;
  reg  _T_6060;
  reg [31:0] _RAND_102;
  wire  _T_6066;
  wire  _T_6067;
  wire  _T_6069;
  wire [1:0] _T_6070;
  wire  _T_6071;
  wire [1:0] _T_6072;
  wire [1:0] _T_6073;
  wire  _T_6074;
  wire  _T_6076;
  wire  _T_6079;
  wire  _T_6081;
  wire  _T_6083;
  wire  _T_6085;
  wire  _T_6087;
  wire  _T_6088;
  wire  _T_6090;
  wire  _T_6092;
  reg  _T_6102;
  reg [31:0] _RAND_103;
  wire  _T_6108;
  wire  _T_6109;
  wire  _T_6111;
  wire [1:0] _T_6112;
  wire  _T_6113;
  wire [1:0] _T_6114;
  wire [1:0] _T_6115;
  wire  _T_6116;
  wire  _T_6118;
  wire  _T_6121;
  wire  _T_6123;
  wire  _T_6125;
  wire  _T_6127;
  wire  _T_6129;
  wire  _T_6130;
  wire  _T_6132;
  wire  _T_6134;
  reg  _T_6144;
  reg [31:0] _RAND_104;
  wire  _T_6150;
  wire  _T_6151;
  wire  _T_6153;
  wire [1:0] _T_6154;
  wire  _T_6155;
  wire [1:0] _T_6156;
  wire [1:0] _T_6157;
  wire  _T_6158;
  wire  _T_6160;
  wire  _T_6163;
  wire  _T_6165;
  wire  _T_6167;
  wire  _T_6169;
  wire  _T_6171;
  wire  _T_6172;
  wire  _T_6174;
  wire  _T_6176;
  reg  _T_6186;
  reg [31:0] _RAND_105;
  wire  _T_6192;
  wire  _T_6193;
  wire  _T_6195;
  wire [1:0] _T_6196;
  wire  _T_6197;
  wire [1:0] _T_6198;
  wire [1:0] _T_6199;
  wire  _T_6200;
  wire  _T_6202;
  wire  _T_6205;
  wire  _T_6207;
  wire  _T_6209;
  wire  _T_6211;
  wire  _T_6213;
  wire  _T_6214;
  wire  _T_6216;
  wire  _T_6218;
  reg  _T_6228;
  reg [31:0] _RAND_106;
  wire  _T_6234;
  wire  _T_6235;
  wire  _T_6237;
  wire [1:0] _T_6238;
  wire  _T_6239;
  wire [1:0] _T_6240;
  wire [1:0] _T_6241;
  wire  _T_6242;
  wire  _T_6244;
  wire  _T_6247;
  wire  _T_6249;
  wire  _T_6251;
  wire  _T_6253;
  wire  _T_6255;
  wire  _T_6256;
  wire  _T_6258;
  wire  _T_6260;
  reg  _T_6270;
  reg [31:0] _RAND_107;
  wire  _T_6276;
  wire  _T_6277;
  wire  _T_6279;
  wire [1:0] _T_6280;
  wire  _T_6281;
  wire [1:0] _T_6282;
  wire [1:0] _T_6283;
  wire  _T_6284;
  wire  _T_6286;
  wire  _T_6289;
  wire  _T_6291;
  wire  _T_6293;
  wire  _T_6295;
  wire  _T_6297;
  wire  _T_6298;
  wire  _T_6300;
  wire  _T_6302;
  reg  _T_6312;
  reg [31:0] _RAND_108;
  wire  _T_6318;
  wire  _T_6319;
  wire  _T_6321;
  wire [1:0] _T_6322;
  wire  _T_6323;
  wire [1:0] _T_6324;
  wire [1:0] _T_6325;
  wire  _T_6326;
  wire  _T_6328;
  wire  _T_6331;
  wire  _T_6333;
  wire  _T_6335;
  wire  _T_6337;
  wire  _T_6339;
  wire  _T_6340;
  wire  _T_6342;
  wire  _T_6344;
  reg  _T_6354;
  reg [31:0] _RAND_109;
  wire  _T_6360;
  wire  _T_6361;
  wire  _T_6363;
  wire [1:0] _T_6364;
  wire  _T_6365;
  wire [1:0] _T_6366;
  wire [1:0] _T_6367;
  wire  _T_6368;
  wire  _T_6370;
  wire  _T_6373;
  wire  _T_6375;
  wire  _T_6377;
  wire  _T_6379;
  wire  _T_6381;
  wire  _T_6382;
  wire  _T_6384;
  wire  _T_6386;
  reg  _T_6396;
  reg [31:0] _RAND_110;
  wire  _T_6402;
  wire  _T_6403;
  wire  _T_6405;
  wire [1:0] _T_6406;
  wire  _T_6407;
  wire [1:0] _T_6408;
  wire [1:0] _T_6409;
  wire  _T_6410;
  wire  _T_6412;
  wire  _T_6415;
  wire  _T_6417;
  wire  _T_6419;
  wire  _T_6421;
  wire  _T_6423;
  wire  _T_6424;
  wire  _T_6426;
  wire  _T_6428;
  reg  _T_6438;
  reg [31:0] _RAND_111;
  wire  _T_6444;
  wire  _T_6445;
  wire  _T_6447;
  wire [1:0] _T_6448;
  wire  _T_6449;
  wire [1:0] _T_6450;
  wire [1:0] _T_6451;
  wire  _T_6452;
  wire  _T_6454;
  wire  _T_6457;
  wire  _T_6459;
  wire  _T_6461;
  wire  _T_6463;
  wire  _T_6465;
  wire  _T_6466;
  wire  _T_6468;
  wire  _T_6470;
  reg  _T_6480;
  reg [31:0] _RAND_112;
  wire  _T_6486;
  wire  _T_6487;
  wire  _T_6489;
  wire [1:0] _T_6490;
  wire  _T_6491;
  wire [1:0] _T_6492;
  wire [1:0] _T_6493;
  wire  _T_6494;
  wire  _T_6496;
  wire  _T_6499;
  wire  _T_6501;
  wire  _T_6503;
  wire  _T_6505;
  wire  _T_6507;
  wire  _T_6508;
  wire  _T_6510;
  wire  _T_6512;
  reg  _T_6522;
  reg [31:0] _RAND_113;
  wire  _T_6528;
  wire  _T_6529;
  wire  _T_6531;
  wire [1:0] _T_6532;
  wire  _T_6533;
  wire [1:0] _T_6534;
  wire [1:0] _T_6535;
  wire  _T_6536;
  wire  _T_6538;
  wire  _T_6541;
  wire  _T_6543;
  wire  _T_6545;
  wire  _T_6547;
  wire  _T_6549;
  wire  _T_6550;
  wire  _T_6552;
  wire  _T_6554;
  reg  _T_6564;
  reg [31:0] _RAND_114;
  wire  _T_6570;
  wire  _T_6571;
  wire  _T_6573;
  wire [1:0] _T_6574;
  wire  _T_6575;
  wire [1:0] _T_6576;
  wire [1:0] _T_6577;
  wire  _T_6578;
  wire  _T_6580;
  wire  _T_6583;
  wire  _T_6585;
  wire  _T_6587;
  wire  _T_6589;
  wire  _T_6591;
  wire  _T_6592;
  wire  _T_6594;
  wire  _T_6596;
  reg  _T_6606;
  reg [31:0] _RAND_115;
  wire  _T_6612;
  wire  _T_6613;
  wire  _T_6615;
  wire [1:0] _T_6616;
  wire  _T_6617;
  wire [1:0] _T_6618;
  wire [1:0] _T_6619;
  wire  _T_6620;
  wire  _T_6622;
  wire  _T_6625;
  wire  _T_6627;
  wire  _T_6629;
  wire  _T_6631;
  wire  _T_6633;
  wire  _T_6634;
  wire  _T_6636;
  wire  _T_6638;
  reg  _T_6648;
  reg [31:0] _RAND_116;
  wire  _T_6654;
  wire  _T_6655;
  wire  _T_6657;
  wire [1:0] _T_6658;
  wire  _T_6659;
  wire [1:0] _T_6660;
  wire [1:0] _T_6661;
  wire  _T_6662;
  wire  _T_6664;
  wire  _T_6667;
  wire  _T_6669;
  wire  _T_6671;
  wire  _T_6673;
  wire  _T_6675;
  wire  _T_6676;
  wire  _T_6678;
  wire  _T_6680;
  reg  _T_6690;
  reg [31:0] _RAND_117;
  wire  _T_6696;
  wire  _T_6697;
  wire  _T_6699;
  wire [1:0] _T_6700;
  wire  _T_6701;
  wire [1:0] _T_6702;
  wire [1:0] _T_6703;
  wire  _T_6704;
  wire  _T_6706;
  wire  _T_6709;
  wire  _T_6711;
  wire  _T_6713;
  wire  _T_6715;
  wire  _T_6717;
  wire  _T_6718;
  wire  _T_6720;
  wire  _T_6722;
  reg  _T_6732;
  reg [31:0] _RAND_118;
  wire  _T_6738;
  wire  _T_6739;
  wire  _T_6741;
  wire [1:0] _T_6742;
  wire  _T_6743;
  wire [1:0] _T_6744;
  wire [1:0] _T_6745;
  wire  _T_6746;
  wire  _T_6748;
  wire  _T_6751;
  wire  _T_6753;
  wire  _T_6755;
  wire  _T_6757;
  wire  _T_6759;
  wire  _T_6760;
  wire  _T_6762;
  wire  _T_6764;
  reg  _T_6774;
  reg [31:0] _RAND_119;
  wire  _T_6780;
  wire  _T_6781;
  wire  _T_6783;
  wire [1:0] _T_6784;
  wire  _T_6785;
  wire [1:0] _T_6786;
  wire [1:0] _T_6787;
  wire  _T_6788;
  wire  _T_6790;
  wire  _T_6793;
  wire  _T_6795;
  wire  _T_6797;
  wire  _T_6799;
  wire  _T_6801;
  wire  _T_6802;
  wire  _T_6804;
  wire  _T_6806;
  reg  _T_6816;
  reg [31:0] _RAND_120;
  wire  _T_6822;
  wire  _T_6823;
  wire  _T_6825;
  wire [1:0] _T_6826;
  wire  _T_6827;
  wire [1:0] _T_6828;
  wire [1:0] _T_6829;
  wire  _T_6830;
  wire  _T_6832;
  wire  _T_6835;
  wire  _T_6837;
  wire  _T_6839;
  wire  _T_6841;
  wire  _T_6843;
  wire  _T_6844;
  wire  _T_6846;
  wire  _T_6848;
  reg  _T_6858;
  reg [31:0] _RAND_121;
  wire  _T_6864;
  wire  _T_6865;
  wire  _T_6867;
  wire [1:0] _T_6868;
  wire  _T_6869;
  wire [1:0] _T_6870;
  wire [1:0] _T_6871;
  wire  _T_6872;
  wire  _T_6874;
  wire  _T_6877;
  wire  _T_6879;
  wire  _T_6881;
  wire  _T_6883;
  wire  _T_6885;
  wire  _T_6886;
  wire  _T_6888;
  wire  _T_6890;
  reg  _T_6900;
  reg [31:0] _RAND_122;
  wire  _T_6906;
  wire  _T_6907;
  wire  _T_6909;
  wire [1:0] _T_6910;
  wire  _T_6911;
  wire [1:0] _T_6912;
  wire [1:0] _T_6913;
  wire  _T_6914;
  wire  _T_6916;
  wire  _T_6919;
  wire  _T_6921;
  wire  _T_6923;
  wire  _T_6925;
  wire  _T_6927;
  wire  _T_6928;
  wire  _T_6930;
  wire  _T_6932;
  reg  _T_6942;
  reg [31:0] _RAND_123;
  wire  _T_6948;
  wire  _T_6949;
  wire  _T_6951;
  wire [1:0] _T_6952;
  wire  _T_6953;
  wire [1:0] _T_6954;
  wire [1:0] _T_6955;
  wire  _T_6956;
  wire  _T_6958;
  wire  _T_6961;
  wire  _T_6963;
  wire  _T_6965;
  wire  _T_6967;
  wire  _T_6969;
  wire  _T_6970;
  wire  _T_6972;
  wire  _T_6974;
  reg  _T_6984;
  reg [31:0] _RAND_124;
  wire  _T_6990;
  wire  _T_6991;
  wire  _T_6993;
  wire [1:0] _T_6994;
  wire  _T_6995;
  wire [1:0] _T_6996;
  wire [1:0] _T_6997;
  wire  _T_6998;
  wire  _T_7000;
  wire  _T_7003;
  wire  _T_7005;
  wire  _T_7007;
  wire  _T_7009;
  wire  _T_7011;
  wire  _T_7012;
  wire  _T_7014;
  wire  _T_7016;
  reg  _T_7026;
  reg [31:0] _RAND_125;
  wire  _T_7032;
  wire  _T_7033;
  wire  _T_7035;
  wire [1:0] _T_7036;
  wire  _T_7037;
  wire [1:0] _T_7038;
  wire [1:0] _T_7039;
  wire  _T_7040;
  wire  _T_7042;
  wire  _T_7045;
  wire  _T_7047;
  wire  _T_7049;
  wire  _T_7051;
  wire  _T_7053;
  wire  _T_7054;
  wire  _T_7056;
  wire  _T_7058;
  reg  _T_7068;
  reg [31:0] _RAND_126;
  wire  _T_7074;
  wire  _T_7075;
  wire  _T_7077;
  wire [1:0] _T_7078;
  wire  _T_7079;
  wire [1:0] _T_7080;
  wire [1:0] _T_7081;
  wire  _T_7082;
  wire  _T_7084;
  wire  _T_7087;
  wire  _T_7089;
  wire  _T_7091;
  wire  _T_7093;
  wire  _T_7095;
  wire  _T_7096;
  wire  _T_7098;
  wire  _T_7100;
  reg  _T_7110;
  reg [31:0] _RAND_127;
  wire  _T_7116;
  wire  _T_7117;
  wire  _T_7119;
  wire [1:0] _T_7120;
  wire  _T_7121;
  wire [1:0] _T_7122;
  wire [1:0] _T_7123;
  wire  _T_7124;
  wire  _T_7126;
  wire  _T_7129;
  wire  _T_7131;
  wire  _T_7133;
  wire  _T_7135;
  wire  _T_7137;
  wire  _T_7138;
  wire  _T_7140;
  wire  _T_7142;
  reg  _T_7152;
  reg [31:0] _RAND_128;
  wire  _T_7158;
  wire  _T_7159;
  wire  _T_7161;
  wire [1:0] _T_7162;
  wire  _T_7163;
  wire [1:0] _T_7164;
  wire [1:0] _T_7165;
  wire  _T_7166;
  wire  _T_7168;
  wire  _T_7171;
  wire  _T_7173;
  wire  _T_7175;
  wire  _T_7177;
  wire  _T_7179;
  wire  _T_7180;
  wire  _T_7182;
  wire  _T_7184;
  reg  _T_7194;
  reg [31:0] _RAND_129;
  wire  _T_7200;
  wire  _T_7201;
  wire  _T_7203;
  wire [1:0] _T_7204;
  wire  _T_7205;
  wire [1:0] _T_7206;
  wire [1:0] _T_7207;
  wire  _T_7208;
  wire  _T_7210;
  wire  _T_7213;
  wire  _T_7215;
  wire  _T_7217;
  wire  _T_7219;
  wire  _T_7221;
  wire  _T_7222;
  wire  _T_7224;
  wire  _T_7226;
  reg  _T_7236;
  reg [31:0] _RAND_130;
  wire  _T_7242;
  wire  _T_7243;
  wire  _T_7245;
  wire [1:0] _T_7246;
  wire  _T_7247;
  wire [1:0] _T_7248;
  wire [1:0] _T_7249;
  wire  _T_7250;
  wire  _T_7252;
  wire  _T_7255;
  wire  _T_7257;
  wire  _T_7259;
  wire  _T_7261;
  wire  _T_7263;
  wire  _T_7264;
  wire  _T_7266;
  wire  _T_7268;
  reg  _T_7278;
  reg [31:0] _RAND_131;
  wire  _T_7284;
  wire  _T_7285;
  wire  _T_7287;
  wire [1:0] _T_7288;
  wire  _T_7289;
  wire [1:0] _T_7290;
  wire [1:0] _T_7291;
  wire  _T_7292;
  wire  _T_7294;
  wire  _T_7297;
  wire  _T_7299;
  wire  _T_7301;
  wire  _T_7303;
  wire  _T_7305;
  wire  _T_7306;
  wire  _T_7308;
  wire  _T_7310;
  Queue_32 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_33 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_1508 = _T_31_a_bits_opcode[2];
  assign _T_1510 = _T_1508 == 1'h0;
  assign _T_1511 = _T_31_a_ready & _T_31_a_valid;
  assign _T_1514 = 13'h3f << _T_31_a_bits_size;
  assign _T_1515 = _T_1514[5:0];
  assign _T_1516 = ~ _T_1515;
  assign _T_1517 = _T_1516[5:3];
  assign _T_1522 = _T_1510 ? _T_1517 : 3'h0;
  assign _T_1527 = _T_1525 - 3'h1;
  assign _T_1528 = $unsigned(_T_1527);
  assign _T_1529 = _T_1528[2:0];
  assign _T_1531 = _T_1525 == 3'h0;
  assign _T_1533 = _T_1525 == 3'h1;
  assign _T_1535 = _T_1522 == 3'h0;
  assign _T_1536 = _T_1533 | _T_1535;
  assign _T_1540 = _T_1531 ? _T_1522 : _T_1529;
  assign _GEN_2 = _T_1511 ? _T_1540 : _T_1525;
  assign _GEN_388 = {{7'd0}, _T_31_a_bits_size};
  assign _T_1554 = _GEN_388 << 7;
  assign _GEN_389 = {{3'd0}, _T_31_a_bits_source};
  assign _T_1555 = _GEN_389 | _T_1554;
  assign _T_1556 = _T_89_r_bits_user[6:0];
  assign _T_1557 = _T_89_r_bits_user[9:7];
  assign _T_1558 = _T_89_b_bits_user[6:0];
  assign _T_1559 = _T_89_b_bits_user[9:7];
  assign _T_1590 = _T_1585_bits_wen == 1'h0;
  assign _T_1591 = _T_1585_valid & _T_1590;
  assign _T_1592 = _T_1585_valid & _T_1585_bits_wen;
  assign _T_1593 = _T_1585_bits_wen ? _T_89_aw_ready : _T_89_ar_ready;
  assign _T_1600 = _T_1536 == 1'h0;
  assign _GEN_3 = _T_1511 ? _T_1600 : _T_1597;
  assign _GEN_4 = 7'h1 == _T_31_a_bits_source ? 7'h1 : 7'h0;
  assign _GEN_5 = 7'h2 == _T_31_a_bits_source ? 7'h2 : _GEN_4;
  assign _GEN_6 = 7'h3 == _T_31_a_bits_source ? 7'h3 : _GEN_5;
  assign _GEN_7 = 7'h4 == _T_31_a_bits_source ? 7'h4 : _GEN_6;
  assign _GEN_8 = 7'h5 == _T_31_a_bits_source ? 7'h5 : _GEN_7;
  assign _GEN_9 = 7'h6 == _T_31_a_bits_source ? 7'h6 : _GEN_8;
  assign _GEN_10 = 7'h7 == _T_31_a_bits_source ? 7'h7 : _GEN_9;
  assign _GEN_11 = 7'h8 == _T_31_a_bits_source ? 7'h8 : _GEN_10;
  assign _GEN_12 = 7'h9 == _T_31_a_bits_source ? 7'h9 : _GEN_11;
  assign _GEN_13 = 7'ha == _T_31_a_bits_source ? 7'ha : _GEN_12;
  assign _GEN_14 = 7'hb == _T_31_a_bits_source ? 7'hb : _GEN_13;
  assign _GEN_15 = 7'hc == _T_31_a_bits_source ? 7'hc : _GEN_14;
  assign _GEN_16 = 7'hd == _T_31_a_bits_source ? 7'hd : _GEN_15;
  assign _GEN_17 = 7'he == _T_31_a_bits_source ? 7'he : _GEN_16;
  assign _GEN_18 = 7'hf == _T_31_a_bits_source ? 7'hf : _GEN_17;
  assign _GEN_19 = 7'h10 == _T_31_a_bits_source ? 7'h10 : _GEN_18;
  assign _GEN_20 = 7'h11 == _T_31_a_bits_source ? 7'h11 : _GEN_19;
  assign _GEN_21 = 7'h12 == _T_31_a_bits_source ? 7'h12 : _GEN_20;
  assign _GEN_22 = 7'h13 == _T_31_a_bits_source ? 7'h13 : _GEN_21;
  assign _GEN_23 = 7'h14 == _T_31_a_bits_source ? 7'h14 : _GEN_22;
  assign _GEN_24 = 7'h15 == _T_31_a_bits_source ? 7'h15 : _GEN_23;
  assign _GEN_25 = 7'h16 == _T_31_a_bits_source ? 7'h16 : _GEN_24;
  assign _GEN_26 = 7'h17 == _T_31_a_bits_source ? 7'h17 : _GEN_25;
  assign _GEN_27 = 7'h18 == _T_31_a_bits_source ? 7'h18 : _GEN_26;
  assign _GEN_28 = 7'h19 == _T_31_a_bits_source ? 7'h19 : _GEN_27;
  assign _GEN_29 = 7'h1a == _T_31_a_bits_source ? 7'h1a : _GEN_28;
  assign _GEN_30 = 7'h1b == _T_31_a_bits_source ? 7'h1b : _GEN_29;
  assign _GEN_31 = 7'h1c == _T_31_a_bits_source ? 7'h1c : _GEN_30;
  assign _GEN_32 = 7'h1d == _T_31_a_bits_source ? 7'h1d : _GEN_31;
  assign _GEN_33 = 7'h1e == _T_31_a_bits_source ? 7'h1e : _GEN_32;
  assign _GEN_34 = 7'h1f == _T_31_a_bits_source ? 7'h1f : _GEN_33;
  assign _GEN_35 = 7'h20 == _T_31_a_bits_source ? 7'h20 : _GEN_34;
  assign _GEN_36 = 7'h21 == _T_31_a_bits_source ? 7'h21 : _GEN_35;
  assign _GEN_37 = 7'h22 == _T_31_a_bits_source ? 7'h22 : _GEN_36;
  assign _GEN_38 = 7'h23 == _T_31_a_bits_source ? 7'h23 : _GEN_37;
  assign _GEN_39 = 7'h24 == _T_31_a_bits_source ? 7'h24 : _GEN_38;
  assign _GEN_40 = 7'h25 == _T_31_a_bits_source ? 7'h25 : _GEN_39;
  assign _GEN_41 = 7'h26 == _T_31_a_bits_source ? 7'h26 : _GEN_40;
  assign _GEN_42 = 7'h27 == _T_31_a_bits_source ? 7'h27 : _GEN_41;
  assign _GEN_43 = 7'h28 == _T_31_a_bits_source ? 7'h28 : _GEN_42;
  assign _GEN_44 = 7'h29 == _T_31_a_bits_source ? 7'h29 : _GEN_43;
  assign _GEN_45 = 7'h2a == _T_31_a_bits_source ? 7'h2a : _GEN_44;
  assign _GEN_46 = 7'h2b == _T_31_a_bits_source ? 7'h2b : _GEN_45;
  assign _GEN_47 = 7'h2c == _T_31_a_bits_source ? 7'h2c : _GEN_46;
  assign _GEN_48 = 7'h2d == _T_31_a_bits_source ? 7'h2d : _GEN_47;
  assign _GEN_49 = 7'h2e == _T_31_a_bits_source ? 7'h2e : _GEN_48;
  assign _GEN_50 = 7'h2f == _T_31_a_bits_source ? 7'h2f : _GEN_49;
  assign _GEN_51 = 7'h30 == _T_31_a_bits_source ? 7'h30 : _GEN_50;
  assign _GEN_52 = 7'h31 == _T_31_a_bits_source ? 7'h31 : _GEN_51;
  assign _GEN_53 = 7'h32 == _T_31_a_bits_source ? 7'h32 : _GEN_52;
  assign _GEN_54 = 7'h33 == _T_31_a_bits_source ? 7'h33 : _GEN_53;
  assign _GEN_55 = 7'h34 == _T_31_a_bits_source ? 7'h34 : _GEN_54;
  assign _GEN_56 = 7'h35 == _T_31_a_bits_source ? 7'h35 : _GEN_55;
  assign _GEN_57 = 7'h36 == _T_31_a_bits_source ? 7'h36 : _GEN_56;
  assign _GEN_58 = 7'h37 == _T_31_a_bits_source ? 7'h37 : _GEN_57;
  assign _GEN_59 = 7'h38 == _T_31_a_bits_source ? 7'h38 : _GEN_58;
  assign _GEN_60 = 7'h39 == _T_31_a_bits_source ? 7'h39 : _GEN_59;
  assign _GEN_61 = 7'h3a == _T_31_a_bits_source ? 7'h3a : _GEN_60;
  assign _GEN_62 = 7'h3b == _T_31_a_bits_source ? 7'h3b : _GEN_61;
  assign _GEN_63 = 7'h3c == _T_31_a_bits_source ? 7'h3c : _GEN_62;
  assign _GEN_64 = 7'h3d == _T_31_a_bits_source ? 7'h3d : _GEN_63;
  assign _GEN_65 = 7'h3e == _T_31_a_bits_source ? 7'h3e : _GEN_64;
  assign _GEN_66 = 7'h3f == _T_31_a_bits_source ? 7'h3f : _GEN_65;
  assign _GEN_67 = 7'h40 == _T_31_a_bits_source ? 7'h40 : _GEN_66;
  assign _GEN_68 = 7'h41 == _T_31_a_bits_source ? 7'h41 : _GEN_67;
  assign _GEN_69 = 7'h42 == _T_31_a_bits_source ? 7'h42 : _GEN_68;
  assign _GEN_70 = 7'h43 == _T_31_a_bits_source ? 7'h43 : _GEN_69;
  assign _GEN_71 = 7'h44 == _T_31_a_bits_source ? 7'h44 : _GEN_70;
  assign _GEN_72 = 7'h45 == _T_31_a_bits_source ? 7'h45 : _GEN_71;
  assign _GEN_73 = 7'h46 == _T_31_a_bits_source ? 7'h46 : _GEN_72;
  assign _GEN_74 = 7'h47 == _T_31_a_bits_source ? 7'h47 : _GEN_73;
  assign _GEN_75 = 7'h48 == _T_31_a_bits_source ? 7'h48 : _GEN_74;
  assign _GEN_76 = 7'h49 == _T_31_a_bits_source ? 7'h49 : _GEN_75;
  assign _GEN_77 = 7'h4a == _T_31_a_bits_source ? 7'h4a : _GEN_76;
  assign _GEN_78 = 7'h4b == _T_31_a_bits_source ? 7'h4b : _GEN_77;
  assign _GEN_79 = 7'h4c == _T_31_a_bits_source ? 7'h4c : _GEN_78;
  assign _GEN_80 = 7'h4d == _T_31_a_bits_source ? 7'h4d : _GEN_79;
  assign _GEN_81 = 7'h4e == _T_31_a_bits_source ? 7'h4e : _GEN_80;
  assign _GEN_82 = 7'h4f == _T_31_a_bits_source ? 7'h4f : _GEN_81;
  assign _GEN_83 = 7'h50 == _T_31_a_bits_source ? 7'h50 : _GEN_82;
  assign _GEN_84 = 7'h51 == _T_31_a_bits_source ? 7'h51 : _GEN_83;
  assign _GEN_85 = 7'h52 == _T_31_a_bits_source ? 7'h52 : _GEN_84;
  assign _GEN_86 = 7'h53 == _T_31_a_bits_source ? 7'h53 : _GEN_85;
  assign _GEN_87 = 7'h54 == _T_31_a_bits_source ? 7'h54 : _GEN_86;
  assign _GEN_88 = 7'h55 == _T_31_a_bits_source ? 7'h55 : _GEN_87;
  assign _GEN_89 = 7'h56 == _T_31_a_bits_source ? 7'h56 : _GEN_88;
  assign _GEN_90 = 7'h57 == _T_31_a_bits_source ? 7'h57 : _GEN_89;
  assign _GEN_91 = 7'h58 == _T_31_a_bits_source ? 7'h58 : _GEN_90;
  assign _GEN_92 = 7'h59 == _T_31_a_bits_source ? 7'h59 : _GEN_91;
  assign _GEN_93 = 7'h5a == _T_31_a_bits_source ? 7'h5a : _GEN_92;
  assign _GEN_94 = 7'h5b == _T_31_a_bits_source ? 7'h5b : _GEN_93;
  assign _GEN_95 = 7'h5c == _T_31_a_bits_source ? 7'h5c : _GEN_94;
  assign _GEN_96 = 7'h5d == _T_31_a_bits_source ? 7'h5d : _GEN_95;
  assign _GEN_97 = 7'h5e == _T_31_a_bits_source ? 7'h5e : _GEN_96;
  assign _GEN_98 = 7'h5f == _T_31_a_bits_source ? 7'h5f : _GEN_97;
  assign _GEN_99 = 7'h60 == _T_31_a_bits_source ? 7'h60 : _GEN_98;
  assign _GEN_100 = 7'h61 == _T_31_a_bits_source ? 7'h61 : _GEN_99;
  assign _GEN_101 = 7'h62 == _T_31_a_bits_source ? 7'h62 : _GEN_100;
  assign _GEN_102 = 7'h63 == _T_31_a_bits_source ? 7'h63 : _GEN_101;
  assign _GEN_103 = 7'h64 == _T_31_a_bits_source ? 7'h64 : _GEN_102;
  assign _GEN_104 = 7'h65 == _T_31_a_bits_source ? 7'h65 : _GEN_103;
  assign _GEN_105 = 7'h66 == _T_31_a_bits_source ? 7'h66 : _GEN_104;
  assign _GEN_106 = 7'h67 == _T_31_a_bits_source ? 7'h67 : _GEN_105;
  assign _GEN_107 = 7'h68 == _T_31_a_bits_source ? 7'h68 : _GEN_106;
  assign _GEN_108 = 7'h69 == _T_31_a_bits_source ? 7'h69 : _GEN_107;
  assign _GEN_109 = 7'h6a == _T_31_a_bits_source ? 7'h6a : _GEN_108;
  assign _GEN_110 = 7'h6b == _T_31_a_bits_source ? 7'h6b : _GEN_109;
  assign _GEN_111 = 7'h6c == _T_31_a_bits_source ? 7'h6c : _GEN_110;
  assign _GEN_112 = 7'h6d == _T_31_a_bits_source ? 7'h6d : _GEN_111;
  assign _GEN_113 = 7'h6e == _T_31_a_bits_source ? 7'h6e : _GEN_112;
  assign _GEN_114 = 7'h6f == _T_31_a_bits_source ? 7'h6f : _GEN_113;
  assign _GEN_115 = 7'h70 == _T_31_a_bits_source ? 7'h70 : _GEN_114;
  assign _GEN_116 = 7'h71 == _T_31_a_bits_source ? 7'h71 : _GEN_115;
  assign _GEN_117 = 7'h72 == _T_31_a_bits_source ? 7'h72 : _GEN_116;
  assign _GEN_118 = 7'h73 == _T_31_a_bits_source ? 7'h73 : _GEN_117;
  assign _GEN_119 = 7'h74 == _T_31_a_bits_source ? 7'h74 : _GEN_118;
  assign _GEN_120 = 7'h75 == _T_31_a_bits_source ? 7'h75 : _GEN_119;
  assign _GEN_121 = 7'h76 == _T_31_a_bits_source ? 7'h76 : _GEN_120;
  assign _GEN_122 = 7'h77 == _T_31_a_bits_source ? 7'h77 : _GEN_121;
  assign _GEN_123 = 7'h78 == _T_31_a_bits_source ? 7'h78 : _GEN_122;
  assign _GEN_124 = 7'h79 == _T_31_a_bits_source ? 7'h79 : _GEN_123;
  assign _GEN_125 = 7'h7a == _T_31_a_bits_source ? 7'h7a : _GEN_124;
  assign _GEN_126 = 7'h7b == _T_31_a_bits_source ? 7'h7b : _GEN_125;
  assign _GEN_127 = 7'h7c == _T_31_a_bits_source ? 7'h7c : _GEN_126;
  assign _GEN_128 = 7'h7d == _T_31_a_bits_source ? 7'h7d : _GEN_127;
  assign _GEN_129 = 7'h7e == _T_31_a_bits_source ? 7'h7e : _GEN_128;
  assign _GEN_130 = 7'h7f == _T_31_a_bits_source ? 7'h7f : _GEN_129;
  assign _T_1604 = 18'h7ff << _T_31_a_bits_size;
  assign _T_1605 = _T_1604[10:0];
  assign _T_1606 = ~ _T_1605;
  assign _T_1607 = _T_1606[10:3];
  assign _T_1608 = _T_31_a_bits_size >= 3'h3;
  assign _T_1609 = _T_1608 ? 3'h3 : _T_31_a_bits_size;
  assign _GEN_131 = 7'h1 == _T_31_a_bits_source ? _T_206_1 : _T_206_0;
  assign _GEN_132 = 7'h2 == _T_31_a_bits_source ? _T_206_2 : _GEN_131;
  assign _GEN_133 = 7'h3 == _T_31_a_bits_source ? _T_206_3 : _GEN_132;
  assign _GEN_134 = 7'h4 == _T_31_a_bits_source ? _T_206_4 : _GEN_133;
  assign _GEN_135 = 7'h5 == _T_31_a_bits_source ? _T_206_5 : _GEN_134;
  assign _GEN_136 = 7'h6 == _T_31_a_bits_source ? _T_206_6 : _GEN_135;
  assign _GEN_137 = 7'h7 == _T_31_a_bits_source ? _T_206_7 : _GEN_136;
  assign _GEN_138 = 7'h8 == _T_31_a_bits_source ? _T_206_8 : _GEN_137;
  assign _GEN_139 = 7'h9 == _T_31_a_bits_source ? _T_206_9 : _GEN_138;
  assign _GEN_140 = 7'ha == _T_31_a_bits_source ? _T_206_10 : _GEN_139;
  assign _GEN_141 = 7'hb == _T_31_a_bits_source ? _T_206_11 : _GEN_140;
  assign _GEN_142 = 7'hc == _T_31_a_bits_source ? _T_206_12 : _GEN_141;
  assign _GEN_143 = 7'hd == _T_31_a_bits_source ? _T_206_13 : _GEN_142;
  assign _GEN_144 = 7'he == _T_31_a_bits_source ? _T_206_14 : _GEN_143;
  assign _GEN_145 = 7'hf == _T_31_a_bits_source ? _T_206_15 : _GEN_144;
  assign _GEN_146 = 7'h10 == _T_31_a_bits_source ? _T_206_16 : _GEN_145;
  assign _GEN_147 = 7'h11 == _T_31_a_bits_source ? _T_206_17 : _GEN_146;
  assign _GEN_148 = 7'h12 == _T_31_a_bits_source ? _T_206_18 : _GEN_147;
  assign _GEN_149 = 7'h13 == _T_31_a_bits_source ? _T_206_19 : _GEN_148;
  assign _GEN_150 = 7'h14 == _T_31_a_bits_source ? _T_206_20 : _GEN_149;
  assign _GEN_151 = 7'h15 == _T_31_a_bits_source ? _T_206_21 : _GEN_150;
  assign _GEN_152 = 7'h16 == _T_31_a_bits_source ? _T_206_22 : _GEN_151;
  assign _GEN_153 = 7'h17 == _T_31_a_bits_source ? _T_206_23 : _GEN_152;
  assign _GEN_154 = 7'h18 == _T_31_a_bits_source ? _T_206_24 : _GEN_153;
  assign _GEN_155 = 7'h19 == _T_31_a_bits_source ? _T_206_25 : _GEN_154;
  assign _GEN_156 = 7'h1a == _T_31_a_bits_source ? _T_206_26 : _GEN_155;
  assign _GEN_157 = 7'h1b == _T_31_a_bits_source ? _T_206_27 : _GEN_156;
  assign _GEN_158 = 7'h1c == _T_31_a_bits_source ? _T_206_28 : _GEN_157;
  assign _GEN_159 = 7'h1d == _T_31_a_bits_source ? _T_206_29 : _GEN_158;
  assign _GEN_160 = 7'h1e == _T_31_a_bits_source ? _T_206_30 : _GEN_159;
  assign _GEN_161 = 7'h1f == _T_31_a_bits_source ? _T_206_31 : _GEN_160;
  assign _GEN_162 = 7'h20 == _T_31_a_bits_source ? _T_206_32 : _GEN_161;
  assign _GEN_163 = 7'h21 == _T_31_a_bits_source ? _T_206_33 : _GEN_162;
  assign _GEN_164 = 7'h22 == _T_31_a_bits_source ? _T_206_34 : _GEN_163;
  assign _GEN_165 = 7'h23 == _T_31_a_bits_source ? _T_206_35 : _GEN_164;
  assign _GEN_166 = 7'h24 == _T_31_a_bits_source ? _T_206_36 : _GEN_165;
  assign _GEN_167 = 7'h25 == _T_31_a_bits_source ? _T_206_37 : _GEN_166;
  assign _GEN_168 = 7'h26 == _T_31_a_bits_source ? _T_206_38 : _GEN_167;
  assign _GEN_169 = 7'h27 == _T_31_a_bits_source ? _T_206_39 : _GEN_168;
  assign _GEN_170 = 7'h28 == _T_31_a_bits_source ? _T_206_40 : _GEN_169;
  assign _GEN_171 = 7'h29 == _T_31_a_bits_source ? _T_206_41 : _GEN_170;
  assign _GEN_172 = 7'h2a == _T_31_a_bits_source ? _T_206_42 : _GEN_171;
  assign _GEN_173 = 7'h2b == _T_31_a_bits_source ? _T_206_43 : _GEN_172;
  assign _GEN_174 = 7'h2c == _T_31_a_bits_source ? _T_206_44 : _GEN_173;
  assign _GEN_175 = 7'h2d == _T_31_a_bits_source ? _T_206_45 : _GEN_174;
  assign _GEN_176 = 7'h2e == _T_31_a_bits_source ? _T_206_46 : _GEN_175;
  assign _GEN_177 = 7'h2f == _T_31_a_bits_source ? _T_206_47 : _GEN_176;
  assign _GEN_178 = 7'h30 == _T_31_a_bits_source ? _T_206_48 : _GEN_177;
  assign _GEN_179 = 7'h31 == _T_31_a_bits_source ? _T_206_49 : _GEN_178;
  assign _GEN_180 = 7'h32 == _T_31_a_bits_source ? _T_206_50 : _GEN_179;
  assign _GEN_181 = 7'h33 == _T_31_a_bits_source ? _T_206_51 : _GEN_180;
  assign _GEN_182 = 7'h34 == _T_31_a_bits_source ? _T_206_52 : _GEN_181;
  assign _GEN_183 = 7'h35 == _T_31_a_bits_source ? _T_206_53 : _GEN_182;
  assign _GEN_184 = 7'h36 == _T_31_a_bits_source ? _T_206_54 : _GEN_183;
  assign _GEN_185 = 7'h37 == _T_31_a_bits_source ? _T_206_55 : _GEN_184;
  assign _GEN_186 = 7'h38 == _T_31_a_bits_source ? _T_206_56 : _GEN_185;
  assign _GEN_187 = 7'h39 == _T_31_a_bits_source ? _T_206_57 : _GEN_186;
  assign _GEN_188 = 7'h3a == _T_31_a_bits_source ? _T_206_58 : _GEN_187;
  assign _GEN_189 = 7'h3b == _T_31_a_bits_source ? _T_206_59 : _GEN_188;
  assign _GEN_190 = 7'h3c == _T_31_a_bits_source ? _T_206_60 : _GEN_189;
  assign _GEN_191 = 7'h3d == _T_31_a_bits_source ? _T_206_61 : _GEN_190;
  assign _GEN_192 = 7'h3e == _T_31_a_bits_source ? _T_206_62 : _GEN_191;
  assign _GEN_193 = 7'h3f == _T_31_a_bits_source ? _T_206_63 : _GEN_192;
  assign _GEN_194 = 7'h40 == _T_31_a_bits_source ? _T_206_64 : _GEN_193;
  assign _GEN_195 = 7'h41 == _T_31_a_bits_source ? _T_206_65 : _GEN_194;
  assign _GEN_196 = 7'h42 == _T_31_a_bits_source ? _T_206_66 : _GEN_195;
  assign _GEN_197 = 7'h43 == _T_31_a_bits_source ? _T_206_67 : _GEN_196;
  assign _GEN_198 = 7'h44 == _T_31_a_bits_source ? _T_206_68 : _GEN_197;
  assign _GEN_199 = 7'h45 == _T_31_a_bits_source ? _T_206_69 : _GEN_198;
  assign _GEN_200 = 7'h46 == _T_31_a_bits_source ? _T_206_70 : _GEN_199;
  assign _GEN_201 = 7'h47 == _T_31_a_bits_source ? _T_206_71 : _GEN_200;
  assign _GEN_202 = 7'h48 == _T_31_a_bits_source ? _T_206_72 : _GEN_201;
  assign _GEN_203 = 7'h49 == _T_31_a_bits_source ? _T_206_73 : _GEN_202;
  assign _GEN_204 = 7'h4a == _T_31_a_bits_source ? _T_206_74 : _GEN_203;
  assign _GEN_205 = 7'h4b == _T_31_a_bits_source ? _T_206_75 : _GEN_204;
  assign _GEN_206 = 7'h4c == _T_31_a_bits_source ? _T_206_76 : _GEN_205;
  assign _GEN_207 = 7'h4d == _T_31_a_bits_source ? _T_206_77 : _GEN_206;
  assign _GEN_208 = 7'h4e == _T_31_a_bits_source ? _T_206_78 : _GEN_207;
  assign _GEN_209 = 7'h4f == _T_31_a_bits_source ? _T_206_79 : _GEN_208;
  assign _GEN_210 = 7'h50 == _T_31_a_bits_source ? _T_206_80 : _GEN_209;
  assign _GEN_211 = 7'h51 == _T_31_a_bits_source ? _T_206_81 : _GEN_210;
  assign _GEN_212 = 7'h52 == _T_31_a_bits_source ? _T_206_82 : _GEN_211;
  assign _GEN_213 = 7'h53 == _T_31_a_bits_source ? _T_206_83 : _GEN_212;
  assign _GEN_214 = 7'h54 == _T_31_a_bits_source ? _T_206_84 : _GEN_213;
  assign _GEN_215 = 7'h55 == _T_31_a_bits_source ? _T_206_85 : _GEN_214;
  assign _GEN_216 = 7'h56 == _T_31_a_bits_source ? _T_206_86 : _GEN_215;
  assign _GEN_217 = 7'h57 == _T_31_a_bits_source ? _T_206_87 : _GEN_216;
  assign _GEN_218 = 7'h58 == _T_31_a_bits_source ? _T_206_88 : _GEN_217;
  assign _GEN_219 = 7'h59 == _T_31_a_bits_source ? _T_206_89 : _GEN_218;
  assign _GEN_220 = 7'h5a == _T_31_a_bits_source ? _T_206_90 : _GEN_219;
  assign _GEN_221 = 7'h5b == _T_31_a_bits_source ? _T_206_91 : _GEN_220;
  assign _GEN_222 = 7'h5c == _T_31_a_bits_source ? _T_206_92 : _GEN_221;
  assign _GEN_223 = 7'h5d == _T_31_a_bits_source ? _T_206_93 : _GEN_222;
  assign _GEN_224 = 7'h5e == _T_31_a_bits_source ? _T_206_94 : _GEN_223;
  assign _GEN_225 = 7'h5f == _T_31_a_bits_source ? _T_206_95 : _GEN_224;
  assign _GEN_226 = 7'h60 == _T_31_a_bits_source ? _T_206_96 : _GEN_225;
  assign _GEN_227 = 7'h61 == _T_31_a_bits_source ? _T_206_97 : _GEN_226;
  assign _GEN_228 = 7'h62 == _T_31_a_bits_source ? _T_206_98 : _GEN_227;
  assign _GEN_229 = 7'h63 == _T_31_a_bits_source ? _T_206_99 : _GEN_228;
  assign _GEN_230 = 7'h64 == _T_31_a_bits_source ? _T_206_100 : _GEN_229;
  assign _GEN_231 = 7'h65 == _T_31_a_bits_source ? _T_206_101 : _GEN_230;
  assign _GEN_232 = 7'h66 == _T_31_a_bits_source ? _T_206_102 : _GEN_231;
  assign _GEN_233 = 7'h67 == _T_31_a_bits_source ? _T_206_103 : _GEN_232;
  assign _GEN_234 = 7'h68 == _T_31_a_bits_source ? _T_206_104 : _GEN_233;
  assign _GEN_235 = 7'h69 == _T_31_a_bits_source ? _T_206_105 : _GEN_234;
  assign _GEN_236 = 7'h6a == _T_31_a_bits_source ? _T_206_106 : _GEN_235;
  assign _GEN_237 = 7'h6b == _T_31_a_bits_source ? _T_206_107 : _GEN_236;
  assign _GEN_238 = 7'h6c == _T_31_a_bits_source ? _T_206_108 : _GEN_237;
  assign _GEN_239 = 7'h6d == _T_31_a_bits_source ? _T_206_109 : _GEN_238;
  assign _GEN_240 = 7'h6e == _T_31_a_bits_source ? _T_206_110 : _GEN_239;
  assign _GEN_241 = 7'h6f == _T_31_a_bits_source ? _T_206_111 : _GEN_240;
  assign _GEN_242 = 7'h70 == _T_31_a_bits_source ? _T_206_112 : _GEN_241;
  assign _GEN_243 = 7'h71 == _T_31_a_bits_source ? _T_206_113 : _GEN_242;
  assign _GEN_244 = 7'h72 == _T_31_a_bits_source ? _T_206_114 : _GEN_243;
  assign _GEN_245 = 7'h73 == _T_31_a_bits_source ? _T_206_115 : _GEN_244;
  assign _GEN_246 = 7'h74 == _T_31_a_bits_source ? _T_206_116 : _GEN_245;
  assign _GEN_247 = 7'h75 == _T_31_a_bits_source ? _T_206_117 : _GEN_246;
  assign _GEN_248 = 7'h76 == _T_31_a_bits_source ? _T_206_118 : _GEN_247;
  assign _GEN_249 = 7'h77 == _T_31_a_bits_source ? _T_206_119 : _GEN_248;
  assign _GEN_250 = 7'h78 == _T_31_a_bits_source ? _T_206_120 : _GEN_249;
  assign _GEN_251 = 7'h79 == _T_31_a_bits_source ? _T_206_121 : _GEN_250;
  assign _GEN_252 = 7'h7a == _T_31_a_bits_source ? _T_206_122 : _GEN_251;
  assign _GEN_253 = 7'h7b == _T_31_a_bits_source ? _T_206_123 : _GEN_252;
  assign _GEN_254 = 7'h7c == _T_31_a_bits_source ? _T_206_124 : _GEN_253;
  assign _GEN_255 = 7'h7d == _T_31_a_bits_source ? _T_206_125 : _GEN_254;
  assign _GEN_256 = 7'h7e == _T_31_a_bits_source ? _T_206_126 : _GEN_255;
  assign _GEN_257 = 7'h7f == _T_31_a_bits_source ? _T_206_127 : _GEN_256;
  assign _T_1616 = _GEN_1 & _T_1531;
  assign _T_1618 = _T_1616 == 1'h0;
  assign _T_1619 = _T_1597 | _T_1565_ready;
  assign _T_1620 = _T_1619 & _T_1569_ready;
  assign _T_1621 = _T_1510 ? _T_1620 : _T_1565_ready;
  assign _T_1622 = _T_1618 & _T_1621;
  assign _T_1625 = _T_1618 & _T_31_a_valid;
  assign _T_1627 = _T_1597 == 1'h0;
  assign _T_1628 = _T_1627 & _T_1569_ready;
  assign _T_1630 = _T_1510 ? _T_1628 : 1'h1;
  assign _T_1631 = _T_1625 & _T_1630;
  assign _T_1635 = _T_1625 & _T_1510;
  assign _T_1637 = _T_1635 & _T_1619;
  assign _T_1641 = _T_89_r_ready & _T_89_r_valid;
  assign _T_1643 = _T_89_r_bits_last == 1'h0;
  assign _GEN_258 = _T_1641 ? _T_1643 : _T_1640;
  assign _T_1644 = _T_89_r_valid | _T_1640;
  assign _T_1646 = _T_1644 == 1'h0;
  assign _T_1647 = _T_31_d_ready & _T_1646;
  assign _T_1648 = _T_1644 ? _T_89_r_valid : _T_89_b_valid;
  assign _T_1650 = _T_89_r_bits_resp != 2'h0;
  assign _T_1652 = _T_89_b_bits_resp != 2'h0;
  assign _T_1659 = _T_1655 | _T_1650;
  assign _T_1660 = _T_1643 & _T_1659;
  assign _GEN_259 = _T_1641 ? _T_1660 : _T_1655;
  assign _T_1674_opcode = _T_1644 ? 3'h1 : 3'h0;
  assign _T_1674_size = _T_1644 ? _T_1664_size : _T_1669_size;
  assign _T_1674_source = _T_1644 ? _T_1664_source : _T_1669_source;
  assign _T_1674_error = _T_1644 ? _T_1664_error : _T_1669_error;
  assign _T_1677 = 128'h1 << _T_1565_bits_id;
  assign _T_1679 = _T_1677[0];
  assign _T_1680 = _T_1677[1];
  assign _T_1681 = _T_1677[2];
  assign _T_1682 = _T_1677[3];
  assign _T_1683 = _T_1677[4];
  assign _T_1684 = _T_1677[5];
  assign _T_1685 = _T_1677[6];
  assign _T_1686 = _T_1677[7];
  assign _T_1687 = _T_1677[8];
  assign _T_1688 = _T_1677[9];
  assign _T_1689 = _T_1677[10];
  assign _T_1690 = _T_1677[11];
  assign _T_1691 = _T_1677[12];
  assign _T_1692 = _T_1677[13];
  assign _T_1693 = _T_1677[14];
  assign _T_1694 = _T_1677[15];
  assign _T_1695 = _T_1677[16];
  assign _T_1696 = _T_1677[17];
  assign _T_1697 = _T_1677[18];
  assign _T_1698 = _T_1677[19];
  assign _T_1699 = _T_1677[20];
  assign _T_1700 = _T_1677[21];
  assign _T_1701 = _T_1677[22];
  assign _T_1702 = _T_1677[23];
  assign _T_1703 = _T_1677[24];
  assign _T_1704 = _T_1677[25];
  assign _T_1705 = _T_1677[26];
  assign _T_1706 = _T_1677[27];
  assign _T_1707 = _T_1677[28];
  assign _T_1708 = _T_1677[29];
  assign _T_1709 = _T_1677[30];
  assign _T_1710 = _T_1677[31];
  assign _T_1711 = _T_1677[32];
  assign _T_1712 = _T_1677[33];
  assign _T_1713 = _T_1677[34];
  assign _T_1714 = _T_1677[35];
  assign _T_1715 = _T_1677[36];
  assign _T_1716 = _T_1677[37];
  assign _T_1717 = _T_1677[38];
  assign _T_1718 = _T_1677[39];
  assign _T_1719 = _T_1677[40];
  assign _T_1720 = _T_1677[41];
  assign _T_1721 = _T_1677[42];
  assign _T_1722 = _T_1677[43];
  assign _T_1723 = _T_1677[44];
  assign _T_1724 = _T_1677[45];
  assign _T_1725 = _T_1677[46];
  assign _T_1726 = _T_1677[47];
  assign _T_1727 = _T_1677[48];
  assign _T_1728 = _T_1677[49];
  assign _T_1729 = _T_1677[50];
  assign _T_1730 = _T_1677[51];
  assign _T_1731 = _T_1677[52];
  assign _T_1732 = _T_1677[53];
  assign _T_1733 = _T_1677[54];
  assign _T_1734 = _T_1677[55];
  assign _T_1735 = _T_1677[56];
  assign _T_1736 = _T_1677[57];
  assign _T_1737 = _T_1677[58];
  assign _T_1738 = _T_1677[59];
  assign _T_1739 = _T_1677[60];
  assign _T_1740 = _T_1677[61];
  assign _T_1741 = _T_1677[62];
  assign _T_1742 = _T_1677[63];
  assign _T_1743 = _T_1677[64];
  assign _T_1744 = _T_1677[65];
  assign _T_1745 = _T_1677[66];
  assign _T_1746 = _T_1677[67];
  assign _T_1747 = _T_1677[68];
  assign _T_1748 = _T_1677[69];
  assign _T_1749 = _T_1677[70];
  assign _T_1750 = _T_1677[71];
  assign _T_1751 = _T_1677[72];
  assign _T_1752 = _T_1677[73];
  assign _T_1753 = _T_1677[74];
  assign _T_1754 = _T_1677[75];
  assign _T_1755 = _T_1677[76];
  assign _T_1756 = _T_1677[77];
  assign _T_1757 = _T_1677[78];
  assign _T_1758 = _T_1677[79];
  assign _T_1759 = _T_1677[80];
  assign _T_1760 = _T_1677[81];
  assign _T_1761 = _T_1677[82];
  assign _T_1762 = _T_1677[83];
  assign _T_1763 = _T_1677[84];
  assign _T_1764 = _T_1677[85];
  assign _T_1765 = _T_1677[86];
  assign _T_1766 = _T_1677[87];
  assign _T_1767 = _T_1677[88];
  assign _T_1768 = _T_1677[89];
  assign _T_1769 = _T_1677[90];
  assign _T_1770 = _T_1677[91];
  assign _T_1771 = _T_1677[92];
  assign _T_1772 = _T_1677[93];
  assign _T_1773 = _T_1677[94];
  assign _T_1774 = _T_1677[95];
  assign _T_1775 = _T_1677[96];
  assign _T_1776 = _T_1677[97];
  assign _T_1777 = _T_1677[98];
  assign _T_1778 = _T_1677[99];
  assign _T_1779 = _T_1677[100];
  assign _T_1780 = _T_1677[101];
  assign _T_1781 = _T_1677[102];
  assign _T_1782 = _T_1677[103];
  assign _T_1783 = _T_1677[104];
  assign _T_1784 = _T_1677[105];
  assign _T_1785 = _T_1677[106];
  assign _T_1786 = _T_1677[107];
  assign _T_1787 = _T_1677[108];
  assign _T_1788 = _T_1677[109];
  assign _T_1789 = _T_1677[110];
  assign _T_1790 = _T_1677[111];
  assign _T_1791 = _T_1677[112];
  assign _T_1792 = _T_1677[113];
  assign _T_1793 = _T_1677[114];
  assign _T_1794 = _T_1677[115];
  assign _T_1795 = _T_1677[116];
  assign _T_1796 = _T_1677[117];
  assign _T_1797 = _T_1677[118];
  assign _T_1798 = _T_1677[119];
  assign _T_1799 = _T_1677[120];
  assign _T_1800 = _T_1677[121];
  assign _T_1801 = _T_1677[122];
  assign _T_1802 = _T_1677[123];
  assign _T_1803 = _T_1677[124];
  assign _T_1804 = _T_1677[125];
  assign _T_1805 = _T_1677[126];
  assign _T_1806 = _T_1677[127];
  assign _T_1807 = _T_1644 ? _T_89_r_bits_id : _T_89_b_bits_id;
  assign _T_1810 = 128'h1 << _T_1807;
  assign _T_1812 = _T_1810[0];
  assign _T_1813 = _T_1810[1];
  assign _T_1814 = _T_1810[2];
  assign _T_1815 = _T_1810[3];
  assign _T_1816 = _T_1810[4];
  assign _T_1817 = _T_1810[5];
  assign _T_1818 = _T_1810[6];
  assign _T_1819 = _T_1810[7];
  assign _T_1820 = _T_1810[8];
  assign _T_1821 = _T_1810[9];
  assign _T_1822 = _T_1810[10];
  assign _T_1823 = _T_1810[11];
  assign _T_1824 = _T_1810[12];
  assign _T_1825 = _T_1810[13];
  assign _T_1826 = _T_1810[14];
  assign _T_1827 = _T_1810[15];
  assign _T_1828 = _T_1810[16];
  assign _T_1829 = _T_1810[17];
  assign _T_1830 = _T_1810[18];
  assign _T_1831 = _T_1810[19];
  assign _T_1832 = _T_1810[20];
  assign _T_1833 = _T_1810[21];
  assign _T_1834 = _T_1810[22];
  assign _T_1835 = _T_1810[23];
  assign _T_1836 = _T_1810[24];
  assign _T_1837 = _T_1810[25];
  assign _T_1838 = _T_1810[26];
  assign _T_1839 = _T_1810[27];
  assign _T_1840 = _T_1810[28];
  assign _T_1841 = _T_1810[29];
  assign _T_1842 = _T_1810[30];
  assign _T_1843 = _T_1810[31];
  assign _T_1844 = _T_1810[32];
  assign _T_1845 = _T_1810[33];
  assign _T_1846 = _T_1810[34];
  assign _T_1847 = _T_1810[35];
  assign _T_1848 = _T_1810[36];
  assign _T_1849 = _T_1810[37];
  assign _T_1850 = _T_1810[38];
  assign _T_1851 = _T_1810[39];
  assign _T_1852 = _T_1810[40];
  assign _T_1853 = _T_1810[41];
  assign _T_1854 = _T_1810[42];
  assign _T_1855 = _T_1810[43];
  assign _T_1856 = _T_1810[44];
  assign _T_1857 = _T_1810[45];
  assign _T_1858 = _T_1810[46];
  assign _T_1859 = _T_1810[47];
  assign _T_1860 = _T_1810[48];
  assign _T_1861 = _T_1810[49];
  assign _T_1862 = _T_1810[50];
  assign _T_1863 = _T_1810[51];
  assign _T_1864 = _T_1810[52];
  assign _T_1865 = _T_1810[53];
  assign _T_1866 = _T_1810[54];
  assign _T_1867 = _T_1810[55];
  assign _T_1868 = _T_1810[56];
  assign _T_1869 = _T_1810[57];
  assign _T_1870 = _T_1810[58];
  assign _T_1871 = _T_1810[59];
  assign _T_1872 = _T_1810[60];
  assign _T_1873 = _T_1810[61];
  assign _T_1874 = _T_1810[62];
  assign _T_1875 = _T_1810[63];
  assign _T_1876 = _T_1810[64];
  assign _T_1877 = _T_1810[65];
  assign _T_1878 = _T_1810[66];
  assign _T_1879 = _T_1810[67];
  assign _T_1880 = _T_1810[68];
  assign _T_1881 = _T_1810[69];
  assign _T_1882 = _T_1810[70];
  assign _T_1883 = _T_1810[71];
  assign _T_1884 = _T_1810[72];
  assign _T_1885 = _T_1810[73];
  assign _T_1886 = _T_1810[74];
  assign _T_1887 = _T_1810[75];
  assign _T_1888 = _T_1810[76];
  assign _T_1889 = _T_1810[77];
  assign _T_1890 = _T_1810[78];
  assign _T_1891 = _T_1810[79];
  assign _T_1892 = _T_1810[80];
  assign _T_1893 = _T_1810[81];
  assign _T_1894 = _T_1810[82];
  assign _T_1895 = _T_1810[83];
  assign _T_1896 = _T_1810[84];
  assign _T_1897 = _T_1810[85];
  assign _T_1898 = _T_1810[86];
  assign _T_1899 = _T_1810[87];
  assign _T_1900 = _T_1810[88];
  assign _T_1901 = _T_1810[89];
  assign _T_1902 = _T_1810[90];
  assign _T_1903 = _T_1810[91];
  assign _T_1904 = _T_1810[92];
  assign _T_1905 = _T_1810[93];
  assign _T_1906 = _T_1810[94];
  assign _T_1907 = _T_1810[95];
  assign _T_1908 = _T_1810[96];
  assign _T_1909 = _T_1810[97];
  assign _T_1910 = _T_1810[98];
  assign _T_1911 = _T_1810[99];
  assign _T_1912 = _T_1810[100];
  assign _T_1913 = _T_1810[101];
  assign _T_1914 = _T_1810[102];
  assign _T_1915 = _T_1810[103];
  assign _T_1916 = _T_1810[104];
  assign _T_1917 = _T_1810[105];
  assign _T_1918 = _T_1810[106];
  assign _T_1919 = _T_1810[107];
  assign _T_1920 = _T_1810[108];
  assign _T_1921 = _T_1810[109];
  assign _T_1922 = _T_1810[110];
  assign _T_1923 = _T_1810[111];
  assign _T_1924 = _T_1810[112];
  assign _T_1925 = _T_1810[113];
  assign _T_1926 = _T_1810[114];
  assign _T_1927 = _T_1810[115];
  assign _T_1928 = _T_1810[116];
  assign _T_1929 = _T_1810[117];
  assign _T_1930 = _T_1810[118];
  assign _T_1931 = _T_1810[119];
  assign _T_1932 = _T_1810[120];
  assign _T_1933 = _T_1810[121];
  assign _T_1934 = _T_1810[122];
  assign _T_1935 = _T_1810[123];
  assign _T_1936 = _T_1810[124];
  assign _T_1937 = _T_1810[125];
  assign _T_1938 = _T_1810[126];
  assign _T_1939 = _T_1810[127];
  assign _T_1941 = _T_1644 ? _T_89_r_bits_last : 1'h1;
  assign _T_1949 = _T_1565_ready & _T_1565_valid;
  assign _T_1950 = _T_1679 & _T_1949;
  assign _T_1951 = _T_1812 & _T_1941;
  assign _T_1952 = _T_31_d_ready & _T_31_d_valid;
  assign _T_1953 = _T_1951 & _T_1952;
  assign _T_1954 = _T_1944 + _T_1950;
  assign _T_1955 = _T_1954[0:0];
  assign _T_1956 = _T_1955 - _T_1953;
  assign _T_1957 = $unsigned(_T_1956);
  assign _T_1958 = _T_1957[0:0];
  assign _T_1960 = _T_1953 == 1'h0;
  assign _T_1963 = _T_1960 | _T_1944;
  assign _T_1965 = _T_1963 | reset;
  assign _T_1967 = _T_1965 == 1'h0;
  assign _T_1969 = _T_1950 == 1'h0;
  assign _T_1971 = _T_1944 != 1'h1;
  assign _T_1972 = _T_1969 | _T_1971;
  assign _T_1974 = _T_1972 | reset;
  assign _T_1976 = _T_1974 == 1'h0;
  assign _T_1992 = _T_1680 & _T_1949;
  assign _T_1993 = _T_1813 & _T_1941;
  assign _T_1995 = _T_1993 & _T_1952;
  assign _T_1996 = _T_1986 + _T_1992;
  assign _T_1997 = _T_1996[0:0];
  assign _T_1998 = _T_1997 - _T_1995;
  assign _T_1999 = $unsigned(_T_1998);
  assign _T_2000 = _T_1999[0:0];
  assign _T_2002 = _T_1995 == 1'h0;
  assign _T_2005 = _T_2002 | _T_1986;
  assign _T_2007 = _T_2005 | reset;
  assign _T_2009 = _T_2007 == 1'h0;
  assign _T_2011 = _T_1992 == 1'h0;
  assign _T_2013 = _T_1986 != 1'h1;
  assign _T_2014 = _T_2011 | _T_2013;
  assign _T_2016 = _T_2014 | reset;
  assign _T_2018 = _T_2016 == 1'h0;
  assign _T_2034 = _T_1681 & _T_1949;
  assign _T_2035 = _T_1814 & _T_1941;
  assign _T_2037 = _T_2035 & _T_1952;
  assign _T_2038 = _T_2028 + _T_2034;
  assign _T_2039 = _T_2038[0:0];
  assign _T_2040 = _T_2039 - _T_2037;
  assign _T_2041 = $unsigned(_T_2040);
  assign _T_2042 = _T_2041[0:0];
  assign _T_2044 = _T_2037 == 1'h0;
  assign _T_2047 = _T_2044 | _T_2028;
  assign _T_2049 = _T_2047 | reset;
  assign _T_2051 = _T_2049 == 1'h0;
  assign _T_2053 = _T_2034 == 1'h0;
  assign _T_2055 = _T_2028 != 1'h1;
  assign _T_2056 = _T_2053 | _T_2055;
  assign _T_2058 = _T_2056 | reset;
  assign _T_2060 = _T_2058 == 1'h0;
  assign _T_2076 = _T_1682 & _T_1949;
  assign _T_2077 = _T_1815 & _T_1941;
  assign _T_2079 = _T_2077 & _T_1952;
  assign _T_2080 = _T_2070 + _T_2076;
  assign _T_2081 = _T_2080[0:0];
  assign _T_2082 = _T_2081 - _T_2079;
  assign _T_2083 = $unsigned(_T_2082);
  assign _T_2084 = _T_2083[0:0];
  assign _T_2086 = _T_2079 == 1'h0;
  assign _T_2089 = _T_2086 | _T_2070;
  assign _T_2091 = _T_2089 | reset;
  assign _T_2093 = _T_2091 == 1'h0;
  assign _T_2095 = _T_2076 == 1'h0;
  assign _T_2097 = _T_2070 != 1'h1;
  assign _T_2098 = _T_2095 | _T_2097;
  assign _T_2100 = _T_2098 | reset;
  assign _T_2102 = _T_2100 == 1'h0;
  assign _T_2118 = _T_1683 & _T_1949;
  assign _T_2119 = _T_1816 & _T_1941;
  assign _T_2121 = _T_2119 & _T_1952;
  assign _T_2122 = _T_2112 + _T_2118;
  assign _T_2123 = _T_2122[0:0];
  assign _T_2124 = _T_2123 - _T_2121;
  assign _T_2125 = $unsigned(_T_2124);
  assign _T_2126 = _T_2125[0:0];
  assign _T_2128 = _T_2121 == 1'h0;
  assign _T_2131 = _T_2128 | _T_2112;
  assign _T_2133 = _T_2131 | reset;
  assign _T_2135 = _T_2133 == 1'h0;
  assign _T_2137 = _T_2118 == 1'h0;
  assign _T_2139 = _T_2112 != 1'h1;
  assign _T_2140 = _T_2137 | _T_2139;
  assign _T_2142 = _T_2140 | reset;
  assign _T_2144 = _T_2142 == 1'h0;
  assign _T_2160 = _T_1684 & _T_1949;
  assign _T_2161 = _T_1817 & _T_1941;
  assign _T_2163 = _T_2161 & _T_1952;
  assign _T_2164 = _T_2154 + _T_2160;
  assign _T_2165 = _T_2164[0:0];
  assign _T_2166 = _T_2165 - _T_2163;
  assign _T_2167 = $unsigned(_T_2166);
  assign _T_2168 = _T_2167[0:0];
  assign _T_2170 = _T_2163 == 1'h0;
  assign _T_2173 = _T_2170 | _T_2154;
  assign _T_2175 = _T_2173 | reset;
  assign _T_2177 = _T_2175 == 1'h0;
  assign _T_2179 = _T_2160 == 1'h0;
  assign _T_2181 = _T_2154 != 1'h1;
  assign _T_2182 = _T_2179 | _T_2181;
  assign _T_2184 = _T_2182 | reset;
  assign _T_2186 = _T_2184 == 1'h0;
  assign _T_2202 = _T_1685 & _T_1949;
  assign _T_2203 = _T_1818 & _T_1941;
  assign _T_2205 = _T_2203 & _T_1952;
  assign _T_2206 = _T_2196 + _T_2202;
  assign _T_2207 = _T_2206[0:0];
  assign _T_2208 = _T_2207 - _T_2205;
  assign _T_2209 = $unsigned(_T_2208);
  assign _T_2210 = _T_2209[0:0];
  assign _T_2212 = _T_2205 == 1'h0;
  assign _T_2215 = _T_2212 | _T_2196;
  assign _T_2217 = _T_2215 | reset;
  assign _T_2219 = _T_2217 == 1'h0;
  assign _T_2221 = _T_2202 == 1'h0;
  assign _T_2223 = _T_2196 != 1'h1;
  assign _T_2224 = _T_2221 | _T_2223;
  assign _T_2226 = _T_2224 | reset;
  assign _T_2228 = _T_2226 == 1'h0;
  assign _T_2244 = _T_1686 & _T_1949;
  assign _T_2245 = _T_1819 & _T_1941;
  assign _T_2247 = _T_2245 & _T_1952;
  assign _T_2248 = _T_2238 + _T_2244;
  assign _T_2249 = _T_2248[0:0];
  assign _T_2250 = _T_2249 - _T_2247;
  assign _T_2251 = $unsigned(_T_2250);
  assign _T_2252 = _T_2251[0:0];
  assign _T_2254 = _T_2247 == 1'h0;
  assign _T_2257 = _T_2254 | _T_2238;
  assign _T_2259 = _T_2257 | reset;
  assign _T_2261 = _T_2259 == 1'h0;
  assign _T_2263 = _T_2244 == 1'h0;
  assign _T_2265 = _T_2238 != 1'h1;
  assign _T_2266 = _T_2263 | _T_2265;
  assign _T_2268 = _T_2266 | reset;
  assign _T_2270 = _T_2268 == 1'h0;
  assign _T_2286 = _T_1687 & _T_1949;
  assign _T_2287 = _T_1820 & _T_1941;
  assign _T_2289 = _T_2287 & _T_1952;
  assign _T_2290 = _T_2280 + _T_2286;
  assign _T_2291 = _T_2290[0:0];
  assign _T_2292 = _T_2291 - _T_2289;
  assign _T_2293 = $unsigned(_T_2292);
  assign _T_2294 = _T_2293[0:0];
  assign _T_2296 = _T_2289 == 1'h0;
  assign _T_2299 = _T_2296 | _T_2280;
  assign _T_2301 = _T_2299 | reset;
  assign _T_2303 = _T_2301 == 1'h0;
  assign _T_2305 = _T_2286 == 1'h0;
  assign _T_2307 = _T_2280 != 1'h1;
  assign _T_2308 = _T_2305 | _T_2307;
  assign _T_2310 = _T_2308 | reset;
  assign _T_2312 = _T_2310 == 1'h0;
  assign _T_2328 = _T_1688 & _T_1949;
  assign _T_2329 = _T_1821 & _T_1941;
  assign _T_2331 = _T_2329 & _T_1952;
  assign _T_2332 = _T_2322 + _T_2328;
  assign _T_2333 = _T_2332[0:0];
  assign _T_2334 = _T_2333 - _T_2331;
  assign _T_2335 = $unsigned(_T_2334);
  assign _T_2336 = _T_2335[0:0];
  assign _T_2338 = _T_2331 == 1'h0;
  assign _T_2341 = _T_2338 | _T_2322;
  assign _T_2343 = _T_2341 | reset;
  assign _T_2345 = _T_2343 == 1'h0;
  assign _T_2347 = _T_2328 == 1'h0;
  assign _T_2349 = _T_2322 != 1'h1;
  assign _T_2350 = _T_2347 | _T_2349;
  assign _T_2352 = _T_2350 | reset;
  assign _T_2354 = _T_2352 == 1'h0;
  assign _T_2370 = _T_1689 & _T_1949;
  assign _T_2371 = _T_1822 & _T_1941;
  assign _T_2373 = _T_2371 & _T_1952;
  assign _T_2374 = _T_2364 + _T_2370;
  assign _T_2375 = _T_2374[0:0];
  assign _T_2376 = _T_2375 - _T_2373;
  assign _T_2377 = $unsigned(_T_2376);
  assign _T_2378 = _T_2377[0:0];
  assign _T_2380 = _T_2373 == 1'h0;
  assign _T_2383 = _T_2380 | _T_2364;
  assign _T_2385 = _T_2383 | reset;
  assign _T_2387 = _T_2385 == 1'h0;
  assign _T_2389 = _T_2370 == 1'h0;
  assign _T_2391 = _T_2364 != 1'h1;
  assign _T_2392 = _T_2389 | _T_2391;
  assign _T_2394 = _T_2392 | reset;
  assign _T_2396 = _T_2394 == 1'h0;
  assign _T_2412 = _T_1690 & _T_1949;
  assign _T_2413 = _T_1823 & _T_1941;
  assign _T_2415 = _T_2413 & _T_1952;
  assign _T_2416 = _T_2406 + _T_2412;
  assign _T_2417 = _T_2416[0:0];
  assign _T_2418 = _T_2417 - _T_2415;
  assign _T_2419 = $unsigned(_T_2418);
  assign _T_2420 = _T_2419[0:0];
  assign _T_2422 = _T_2415 == 1'h0;
  assign _T_2425 = _T_2422 | _T_2406;
  assign _T_2427 = _T_2425 | reset;
  assign _T_2429 = _T_2427 == 1'h0;
  assign _T_2431 = _T_2412 == 1'h0;
  assign _T_2433 = _T_2406 != 1'h1;
  assign _T_2434 = _T_2431 | _T_2433;
  assign _T_2436 = _T_2434 | reset;
  assign _T_2438 = _T_2436 == 1'h0;
  assign _T_2454 = _T_1691 & _T_1949;
  assign _T_2455 = _T_1824 & _T_1941;
  assign _T_2457 = _T_2455 & _T_1952;
  assign _T_2458 = _T_2448 + _T_2454;
  assign _T_2459 = _T_2458[0:0];
  assign _T_2460 = _T_2459 - _T_2457;
  assign _T_2461 = $unsigned(_T_2460);
  assign _T_2462 = _T_2461[0:0];
  assign _T_2464 = _T_2457 == 1'h0;
  assign _T_2467 = _T_2464 | _T_2448;
  assign _T_2469 = _T_2467 | reset;
  assign _T_2471 = _T_2469 == 1'h0;
  assign _T_2473 = _T_2454 == 1'h0;
  assign _T_2475 = _T_2448 != 1'h1;
  assign _T_2476 = _T_2473 | _T_2475;
  assign _T_2478 = _T_2476 | reset;
  assign _T_2480 = _T_2478 == 1'h0;
  assign _T_2496 = _T_1692 & _T_1949;
  assign _T_2497 = _T_1825 & _T_1941;
  assign _T_2499 = _T_2497 & _T_1952;
  assign _T_2500 = _T_2490 + _T_2496;
  assign _T_2501 = _T_2500[0:0];
  assign _T_2502 = _T_2501 - _T_2499;
  assign _T_2503 = $unsigned(_T_2502);
  assign _T_2504 = _T_2503[0:0];
  assign _T_2506 = _T_2499 == 1'h0;
  assign _T_2509 = _T_2506 | _T_2490;
  assign _T_2511 = _T_2509 | reset;
  assign _T_2513 = _T_2511 == 1'h0;
  assign _T_2515 = _T_2496 == 1'h0;
  assign _T_2517 = _T_2490 != 1'h1;
  assign _T_2518 = _T_2515 | _T_2517;
  assign _T_2520 = _T_2518 | reset;
  assign _T_2522 = _T_2520 == 1'h0;
  assign _T_2538 = _T_1693 & _T_1949;
  assign _T_2539 = _T_1826 & _T_1941;
  assign _T_2541 = _T_2539 & _T_1952;
  assign _T_2542 = _T_2532 + _T_2538;
  assign _T_2543 = _T_2542[0:0];
  assign _T_2544 = _T_2543 - _T_2541;
  assign _T_2545 = $unsigned(_T_2544);
  assign _T_2546 = _T_2545[0:0];
  assign _T_2548 = _T_2541 == 1'h0;
  assign _T_2551 = _T_2548 | _T_2532;
  assign _T_2553 = _T_2551 | reset;
  assign _T_2555 = _T_2553 == 1'h0;
  assign _T_2557 = _T_2538 == 1'h0;
  assign _T_2559 = _T_2532 != 1'h1;
  assign _T_2560 = _T_2557 | _T_2559;
  assign _T_2562 = _T_2560 | reset;
  assign _T_2564 = _T_2562 == 1'h0;
  assign _T_2580 = _T_1694 & _T_1949;
  assign _T_2581 = _T_1827 & _T_1941;
  assign _T_2583 = _T_2581 & _T_1952;
  assign _T_2584 = _T_2574 + _T_2580;
  assign _T_2585 = _T_2584[0:0];
  assign _T_2586 = _T_2585 - _T_2583;
  assign _T_2587 = $unsigned(_T_2586);
  assign _T_2588 = _T_2587[0:0];
  assign _T_2590 = _T_2583 == 1'h0;
  assign _T_2593 = _T_2590 | _T_2574;
  assign _T_2595 = _T_2593 | reset;
  assign _T_2597 = _T_2595 == 1'h0;
  assign _T_2599 = _T_2580 == 1'h0;
  assign _T_2601 = _T_2574 != 1'h1;
  assign _T_2602 = _T_2599 | _T_2601;
  assign _T_2604 = _T_2602 | reset;
  assign _T_2606 = _T_2604 == 1'h0;
  assign _T_2622 = _T_1695 & _T_1949;
  assign _T_2623 = _T_1828 & _T_1941;
  assign _T_2625 = _T_2623 & _T_1952;
  assign _T_2626 = _T_2616 + _T_2622;
  assign _T_2627 = _T_2626[0:0];
  assign _T_2628 = _T_2627 - _T_2625;
  assign _T_2629 = $unsigned(_T_2628);
  assign _T_2630 = _T_2629[0:0];
  assign _T_2632 = _T_2625 == 1'h0;
  assign _T_2635 = _T_2632 | _T_2616;
  assign _T_2637 = _T_2635 | reset;
  assign _T_2639 = _T_2637 == 1'h0;
  assign _T_2641 = _T_2622 == 1'h0;
  assign _T_2643 = _T_2616 != 1'h1;
  assign _T_2644 = _T_2641 | _T_2643;
  assign _T_2646 = _T_2644 | reset;
  assign _T_2648 = _T_2646 == 1'h0;
  assign _T_2664 = _T_1696 & _T_1949;
  assign _T_2665 = _T_1829 & _T_1941;
  assign _T_2667 = _T_2665 & _T_1952;
  assign _T_2668 = _T_2658 + _T_2664;
  assign _T_2669 = _T_2668[0:0];
  assign _T_2670 = _T_2669 - _T_2667;
  assign _T_2671 = $unsigned(_T_2670);
  assign _T_2672 = _T_2671[0:0];
  assign _T_2674 = _T_2667 == 1'h0;
  assign _T_2677 = _T_2674 | _T_2658;
  assign _T_2679 = _T_2677 | reset;
  assign _T_2681 = _T_2679 == 1'h0;
  assign _T_2683 = _T_2664 == 1'h0;
  assign _T_2685 = _T_2658 != 1'h1;
  assign _T_2686 = _T_2683 | _T_2685;
  assign _T_2688 = _T_2686 | reset;
  assign _T_2690 = _T_2688 == 1'h0;
  assign _T_2706 = _T_1697 & _T_1949;
  assign _T_2707 = _T_1830 & _T_1941;
  assign _T_2709 = _T_2707 & _T_1952;
  assign _T_2710 = _T_2700 + _T_2706;
  assign _T_2711 = _T_2710[0:0];
  assign _T_2712 = _T_2711 - _T_2709;
  assign _T_2713 = $unsigned(_T_2712);
  assign _T_2714 = _T_2713[0:0];
  assign _T_2716 = _T_2709 == 1'h0;
  assign _T_2719 = _T_2716 | _T_2700;
  assign _T_2721 = _T_2719 | reset;
  assign _T_2723 = _T_2721 == 1'h0;
  assign _T_2725 = _T_2706 == 1'h0;
  assign _T_2727 = _T_2700 != 1'h1;
  assign _T_2728 = _T_2725 | _T_2727;
  assign _T_2730 = _T_2728 | reset;
  assign _T_2732 = _T_2730 == 1'h0;
  assign _T_2748 = _T_1698 & _T_1949;
  assign _T_2749 = _T_1831 & _T_1941;
  assign _T_2751 = _T_2749 & _T_1952;
  assign _T_2752 = _T_2742 + _T_2748;
  assign _T_2753 = _T_2752[0:0];
  assign _T_2754 = _T_2753 - _T_2751;
  assign _T_2755 = $unsigned(_T_2754);
  assign _T_2756 = _T_2755[0:0];
  assign _T_2758 = _T_2751 == 1'h0;
  assign _T_2761 = _T_2758 | _T_2742;
  assign _T_2763 = _T_2761 | reset;
  assign _T_2765 = _T_2763 == 1'h0;
  assign _T_2767 = _T_2748 == 1'h0;
  assign _T_2769 = _T_2742 != 1'h1;
  assign _T_2770 = _T_2767 | _T_2769;
  assign _T_2772 = _T_2770 | reset;
  assign _T_2774 = _T_2772 == 1'h0;
  assign _T_2790 = _T_1699 & _T_1949;
  assign _T_2791 = _T_1832 & _T_1941;
  assign _T_2793 = _T_2791 & _T_1952;
  assign _T_2794 = _T_2784 + _T_2790;
  assign _T_2795 = _T_2794[0:0];
  assign _T_2796 = _T_2795 - _T_2793;
  assign _T_2797 = $unsigned(_T_2796);
  assign _T_2798 = _T_2797[0:0];
  assign _T_2800 = _T_2793 == 1'h0;
  assign _T_2803 = _T_2800 | _T_2784;
  assign _T_2805 = _T_2803 | reset;
  assign _T_2807 = _T_2805 == 1'h0;
  assign _T_2809 = _T_2790 == 1'h0;
  assign _T_2811 = _T_2784 != 1'h1;
  assign _T_2812 = _T_2809 | _T_2811;
  assign _T_2814 = _T_2812 | reset;
  assign _T_2816 = _T_2814 == 1'h0;
  assign _T_2832 = _T_1700 & _T_1949;
  assign _T_2833 = _T_1833 & _T_1941;
  assign _T_2835 = _T_2833 & _T_1952;
  assign _T_2836 = _T_2826 + _T_2832;
  assign _T_2837 = _T_2836[0:0];
  assign _T_2838 = _T_2837 - _T_2835;
  assign _T_2839 = $unsigned(_T_2838);
  assign _T_2840 = _T_2839[0:0];
  assign _T_2842 = _T_2835 == 1'h0;
  assign _T_2845 = _T_2842 | _T_2826;
  assign _T_2847 = _T_2845 | reset;
  assign _T_2849 = _T_2847 == 1'h0;
  assign _T_2851 = _T_2832 == 1'h0;
  assign _T_2853 = _T_2826 != 1'h1;
  assign _T_2854 = _T_2851 | _T_2853;
  assign _T_2856 = _T_2854 | reset;
  assign _T_2858 = _T_2856 == 1'h0;
  assign _T_2874 = _T_1701 & _T_1949;
  assign _T_2875 = _T_1834 & _T_1941;
  assign _T_2877 = _T_2875 & _T_1952;
  assign _T_2878 = _T_2868 + _T_2874;
  assign _T_2879 = _T_2878[0:0];
  assign _T_2880 = _T_2879 - _T_2877;
  assign _T_2881 = $unsigned(_T_2880);
  assign _T_2882 = _T_2881[0:0];
  assign _T_2884 = _T_2877 == 1'h0;
  assign _T_2887 = _T_2884 | _T_2868;
  assign _T_2889 = _T_2887 | reset;
  assign _T_2891 = _T_2889 == 1'h0;
  assign _T_2893 = _T_2874 == 1'h0;
  assign _T_2895 = _T_2868 != 1'h1;
  assign _T_2896 = _T_2893 | _T_2895;
  assign _T_2898 = _T_2896 | reset;
  assign _T_2900 = _T_2898 == 1'h0;
  assign _T_2916 = _T_1702 & _T_1949;
  assign _T_2917 = _T_1835 & _T_1941;
  assign _T_2919 = _T_2917 & _T_1952;
  assign _T_2920 = _T_2910 + _T_2916;
  assign _T_2921 = _T_2920[0:0];
  assign _T_2922 = _T_2921 - _T_2919;
  assign _T_2923 = $unsigned(_T_2922);
  assign _T_2924 = _T_2923[0:0];
  assign _T_2926 = _T_2919 == 1'h0;
  assign _T_2929 = _T_2926 | _T_2910;
  assign _T_2931 = _T_2929 | reset;
  assign _T_2933 = _T_2931 == 1'h0;
  assign _T_2935 = _T_2916 == 1'h0;
  assign _T_2937 = _T_2910 != 1'h1;
  assign _T_2938 = _T_2935 | _T_2937;
  assign _T_2940 = _T_2938 | reset;
  assign _T_2942 = _T_2940 == 1'h0;
  assign _T_2958 = _T_1703 & _T_1949;
  assign _T_2959 = _T_1836 & _T_1941;
  assign _T_2961 = _T_2959 & _T_1952;
  assign _T_2962 = _T_2952 + _T_2958;
  assign _T_2963 = _T_2962[0:0];
  assign _T_2964 = _T_2963 - _T_2961;
  assign _T_2965 = $unsigned(_T_2964);
  assign _T_2966 = _T_2965[0:0];
  assign _T_2968 = _T_2961 == 1'h0;
  assign _T_2971 = _T_2968 | _T_2952;
  assign _T_2973 = _T_2971 | reset;
  assign _T_2975 = _T_2973 == 1'h0;
  assign _T_2977 = _T_2958 == 1'h0;
  assign _T_2979 = _T_2952 != 1'h1;
  assign _T_2980 = _T_2977 | _T_2979;
  assign _T_2982 = _T_2980 | reset;
  assign _T_2984 = _T_2982 == 1'h0;
  assign _T_3000 = _T_1704 & _T_1949;
  assign _T_3001 = _T_1837 & _T_1941;
  assign _T_3003 = _T_3001 & _T_1952;
  assign _T_3004 = _T_2994 + _T_3000;
  assign _T_3005 = _T_3004[0:0];
  assign _T_3006 = _T_3005 - _T_3003;
  assign _T_3007 = $unsigned(_T_3006);
  assign _T_3008 = _T_3007[0:0];
  assign _T_3010 = _T_3003 == 1'h0;
  assign _T_3013 = _T_3010 | _T_2994;
  assign _T_3015 = _T_3013 | reset;
  assign _T_3017 = _T_3015 == 1'h0;
  assign _T_3019 = _T_3000 == 1'h0;
  assign _T_3021 = _T_2994 != 1'h1;
  assign _T_3022 = _T_3019 | _T_3021;
  assign _T_3024 = _T_3022 | reset;
  assign _T_3026 = _T_3024 == 1'h0;
  assign _T_3042 = _T_1705 & _T_1949;
  assign _T_3043 = _T_1838 & _T_1941;
  assign _T_3045 = _T_3043 & _T_1952;
  assign _T_3046 = _T_3036 + _T_3042;
  assign _T_3047 = _T_3046[0:0];
  assign _T_3048 = _T_3047 - _T_3045;
  assign _T_3049 = $unsigned(_T_3048);
  assign _T_3050 = _T_3049[0:0];
  assign _T_3052 = _T_3045 == 1'h0;
  assign _T_3055 = _T_3052 | _T_3036;
  assign _T_3057 = _T_3055 | reset;
  assign _T_3059 = _T_3057 == 1'h0;
  assign _T_3061 = _T_3042 == 1'h0;
  assign _T_3063 = _T_3036 != 1'h1;
  assign _T_3064 = _T_3061 | _T_3063;
  assign _T_3066 = _T_3064 | reset;
  assign _T_3068 = _T_3066 == 1'h0;
  assign _T_3084 = _T_1706 & _T_1949;
  assign _T_3085 = _T_1839 & _T_1941;
  assign _T_3087 = _T_3085 & _T_1952;
  assign _T_3088 = _T_3078 + _T_3084;
  assign _T_3089 = _T_3088[0:0];
  assign _T_3090 = _T_3089 - _T_3087;
  assign _T_3091 = $unsigned(_T_3090);
  assign _T_3092 = _T_3091[0:0];
  assign _T_3094 = _T_3087 == 1'h0;
  assign _T_3097 = _T_3094 | _T_3078;
  assign _T_3099 = _T_3097 | reset;
  assign _T_3101 = _T_3099 == 1'h0;
  assign _T_3103 = _T_3084 == 1'h0;
  assign _T_3105 = _T_3078 != 1'h1;
  assign _T_3106 = _T_3103 | _T_3105;
  assign _T_3108 = _T_3106 | reset;
  assign _T_3110 = _T_3108 == 1'h0;
  assign _T_3126 = _T_1707 & _T_1949;
  assign _T_3127 = _T_1840 & _T_1941;
  assign _T_3129 = _T_3127 & _T_1952;
  assign _T_3130 = _T_3120 + _T_3126;
  assign _T_3131 = _T_3130[0:0];
  assign _T_3132 = _T_3131 - _T_3129;
  assign _T_3133 = $unsigned(_T_3132);
  assign _T_3134 = _T_3133[0:0];
  assign _T_3136 = _T_3129 == 1'h0;
  assign _T_3139 = _T_3136 | _T_3120;
  assign _T_3141 = _T_3139 | reset;
  assign _T_3143 = _T_3141 == 1'h0;
  assign _T_3145 = _T_3126 == 1'h0;
  assign _T_3147 = _T_3120 != 1'h1;
  assign _T_3148 = _T_3145 | _T_3147;
  assign _T_3150 = _T_3148 | reset;
  assign _T_3152 = _T_3150 == 1'h0;
  assign _T_3168 = _T_1708 & _T_1949;
  assign _T_3169 = _T_1841 & _T_1941;
  assign _T_3171 = _T_3169 & _T_1952;
  assign _T_3172 = _T_3162 + _T_3168;
  assign _T_3173 = _T_3172[0:0];
  assign _T_3174 = _T_3173 - _T_3171;
  assign _T_3175 = $unsigned(_T_3174);
  assign _T_3176 = _T_3175[0:0];
  assign _T_3178 = _T_3171 == 1'h0;
  assign _T_3181 = _T_3178 | _T_3162;
  assign _T_3183 = _T_3181 | reset;
  assign _T_3185 = _T_3183 == 1'h0;
  assign _T_3187 = _T_3168 == 1'h0;
  assign _T_3189 = _T_3162 != 1'h1;
  assign _T_3190 = _T_3187 | _T_3189;
  assign _T_3192 = _T_3190 | reset;
  assign _T_3194 = _T_3192 == 1'h0;
  assign _T_3210 = _T_1709 & _T_1949;
  assign _T_3211 = _T_1842 & _T_1941;
  assign _T_3213 = _T_3211 & _T_1952;
  assign _T_3214 = _T_3204 + _T_3210;
  assign _T_3215 = _T_3214[0:0];
  assign _T_3216 = _T_3215 - _T_3213;
  assign _T_3217 = $unsigned(_T_3216);
  assign _T_3218 = _T_3217[0:0];
  assign _T_3220 = _T_3213 == 1'h0;
  assign _T_3223 = _T_3220 | _T_3204;
  assign _T_3225 = _T_3223 | reset;
  assign _T_3227 = _T_3225 == 1'h0;
  assign _T_3229 = _T_3210 == 1'h0;
  assign _T_3231 = _T_3204 != 1'h1;
  assign _T_3232 = _T_3229 | _T_3231;
  assign _T_3234 = _T_3232 | reset;
  assign _T_3236 = _T_3234 == 1'h0;
  assign _T_3252 = _T_1710 & _T_1949;
  assign _T_3253 = _T_1843 & _T_1941;
  assign _T_3255 = _T_3253 & _T_1952;
  assign _T_3256 = _T_3246 + _T_3252;
  assign _T_3257 = _T_3256[0:0];
  assign _T_3258 = _T_3257 - _T_3255;
  assign _T_3259 = $unsigned(_T_3258);
  assign _T_3260 = _T_3259[0:0];
  assign _T_3262 = _T_3255 == 1'h0;
  assign _T_3265 = _T_3262 | _T_3246;
  assign _T_3267 = _T_3265 | reset;
  assign _T_3269 = _T_3267 == 1'h0;
  assign _T_3271 = _T_3252 == 1'h0;
  assign _T_3273 = _T_3246 != 1'h1;
  assign _T_3274 = _T_3271 | _T_3273;
  assign _T_3276 = _T_3274 | reset;
  assign _T_3278 = _T_3276 == 1'h0;
  assign _T_3294 = _T_1711 & _T_1949;
  assign _T_3295 = _T_1844 & _T_1941;
  assign _T_3297 = _T_3295 & _T_1952;
  assign _T_3298 = _T_3288 + _T_3294;
  assign _T_3299 = _T_3298[0:0];
  assign _T_3300 = _T_3299 - _T_3297;
  assign _T_3301 = $unsigned(_T_3300);
  assign _T_3302 = _T_3301[0:0];
  assign _T_3304 = _T_3297 == 1'h0;
  assign _T_3307 = _T_3304 | _T_3288;
  assign _T_3309 = _T_3307 | reset;
  assign _T_3311 = _T_3309 == 1'h0;
  assign _T_3313 = _T_3294 == 1'h0;
  assign _T_3315 = _T_3288 != 1'h1;
  assign _T_3316 = _T_3313 | _T_3315;
  assign _T_3318 = _T_3316 | reset;
  assign _T_3320 = _T_3318 == 1'h0;
  assign _T_3336 = _T_1712 & _T_1949;
  assign _T_3337 = _T_1845 & _T_1941;
  assign _T_3339 = _T_3337 & _T_1952;
  assign _T_3340 = _T_3330 + _T_3336;
  assign _T_3341 = _T_3340[0:0];
  assign _T_3342 = _T_3341 - _T_3339;
  assign _T_3343 = $unsigned(_T_3342);
  assign _T_3344 = _T_3343[0:0];
  assign _T_3346 = _T_3339 == 1'h0;
  assign _T_3349 = _T_3346 | _T_3330;
  assign _T_3351 = _T_3349 | reset;
  assign _T_3353 = _T_3351 == 1'h0;
  assign _T_3355 = _T_3336 == 1'h0;
  assign _T_3357 = _T_3330 != 1'h1;
  assign _T_3358 = _T_3355 | _T_3357;
  assign _T_3360 = _T_3358 | reset;
  assign _T_3362 = _T_3360 == 1'h0;
  assign _T_3378 = _T_1713 & _T_1949;
  assign _T_3379 = _T_1846 & _T_1941;
  assign _T_3381 = _T_3379 & _T_1952;
  assign _T_3382 = _T_3372 + _T_3378;
  assign _T_3383 = _T_3382[0:0];
  assign _T_3384 = _T_3383 - _T_3381;
  assign _T_3385 = $unsigned(_T_3384);
  assign _T_3386 = _T_3385[0:0];
  assign _T_3388 = _T_3381 == 1'h0;
  assign _T_3391 = _T_3388 | _T_3372;
  assign _T_3393 = _T_3391 | reset;
  assign _T_3395 = _T_3393 == 1'h0;
  assign _T_3397 = _T_3378 == 1'h0;
  assign _T_3399 = _T_3372 != 1'h1;
  assign _T_3400 = _T_3397 | _T_3399;
  assign _T_3402 = _T_3400 | reset;
  assign _T_3404 = _T_3402 == 1'h0;
  assign _T_3420 = _T_1714 & _T_1949;
  assign _T_3421 = _T_1847 & _T_1941;
  assign _T_3423 = _T_3421 & _T_1952;
  assign _T_3424 = _T_3414 + _T_3420;
  assign _T_3425 = _T_3424[0:0];
  assign _T_3426 = _T_3425 - _T_3423;
  assign _T_3427 = $unsigned(_T_3426);
  assign _T_3428 = _T_3427[0:0];
  assign _T_3430 = _T_3423 == 1'h0;
  assign _T_3433 = _T_3430 | _T_3414;
  assign _T_3435 = _T_3433 | reset;
  assign _T_3437 = _T_3435 == 1'h0;
  assign _T_3439 = _T_3420 == 1'h0;
  assign _T_3441 = _T_3414 != 1'h1;
  assign _T_3442 = _T_3439 | _T_3441;
  assign _T_3444 = _T_3442 | reset;
  assign _T_3446 = _T_3444 == 1'h0;
  assign _T_3462 = _T_1715 & _T_1949;
  assign _T_3463 = _T_1848 & _T_1941;
  assign _T_3465 = _T_3463 & _T_1952;
  assign _T_3466 = _T_3456 + _T_3462;
  assign _T_3467 = _T_3466[0:0];
  assign _T_3468 = _T_3467 - _T_3465;
  assign _T_3469 = $unsigned(_T_3468);
  assign _T_3470 = _T_3469[0:0];
  assign _T_3472 = _T_3465 == 1'h0;
  assign _T_3475 = _T_3472 | _T_3456;
  assign _T_3477 = _T_3475 | reset;
  assign _T_3479 = _T_3477 == 1'h0;
  assign _T_3481 = _T_3462 == 1'h0;
  assign _T_3483 = _T_3456 != 1'h1;
  assign _T_3484 = _T_3481 | _T_3483;
  assign _T_3486 = _T_3484 | reset;
  assign _T_3488 = _T_3486 == 1'h0;
  assign _T_3504 = _T_1716 & _T_1949;
  assign _T_3505 = _T_1849 & _T_1941;
  assign _T_3507 = _T_3505 & _T_1952;
  assign _T_3508 = _T_3498 + _T_3504;
  assign _T_3509 = _T_3508[0:0];
  assign _T_3510 = _T_3509 - _T_3507;
  assign _T_3511 = $unsigned(_T_3510);
  assign _T_3512 = _T_3511[0:0];
  assign _T_3514 = _T_3507 == 1'h0;
  assign _T_3517 = _T_3514 | _T_3498;
  assign _T_3519 = _T_3517 | reset;
  assign _T_3521 = _T_3519 == 1'h0;
  assign _T_3523 = _T_3504 == 1'h0;
  assign _T_3525 = _T_3498 != 1'h1;
  assign _T_3526 = _T_3523 | _T_3525;
  assign _T_3528 = _T_3526 | reset;
  assign _T_3530 = _T_3528 == 1'h0;
  assign _T_3546 = _T_1717 & _T_1949;
  assign _T_3547 = _T_1850 & _T_1941;
  assign _T_3549 = _T_3547 & _T_1952;
  assign _T_3550 = _T_3540 + _T_3546;
  assign _T_3551 = _T_3550[0:0];
  assign _T_3552 = _T_3551 - _T_3549;
  assign _T_3553 = $unsigned(_T_3552);
  assign _T_3554 = _T_3553[0:0];
  assign _T_3556 = _T_3549 == 1'h0;
  assign _T_3559 = _T_3556 | _T_3540;
  assign _T_3561 = _T_3559 | reset;
  assign _T_3563 = _T_3561 == 1'h0;
  assign _T_3565 = _T_3546 == 1'h0;
  assign _T_3567 = _T_3540 != 1'h1;
  assign _T_3568 = _T_3565 | _T_3567;
  assign _T_3570 = _T_3568 | reset;
  assign _T_3572 = _T_3570 == 1'h0;
  assign _T_3588 = _T_1718 & _T_1949;
  assign _T_3589 = _T_1851 & _T_1941;
  assign _T_3591 = _T_3589 & _T_1952;
  assign _T_3592 = _T_3582 + _T_3588;
  assign _T_3593 = _T_3592[0:0];
  assign _T_3594 = _T_3593 - _T_3591;
  assign _T_3595 = $unsigned(_T_3594);
  assign _T_3596 = _T_3595[0:0];
  assign _T_3598 = _T_3591 == 1'h0;
  assign _T_3601 = _T_3598 | _T_3582;
  assign _T_3603 = _T_3601 | reset;
  assign _T_3605 = _T_3603 == 1'h0;
  assign _T_3607 = _T_3588 == 1'h0;
  assign _T_3609 = _T_3582 != 1'h1;
  assign _T_3610 = _T_3607 | _T_3609;
  assign _T_3612 = _T_3610 | reset;
  assign _T_3614 = _T_3612 == 1'h0;
  assign _T_3630 = _T_1719 & _T_1949;
  assign _T_3631 = _T_1852 & _T_1941;
  assign _T_3633 = _T_3631 & _T_1952;
  assign _T_3634 = _T_3624 + _T_3630;
  assign _T_3635 = _T_3634[0:0];
  assign _T_3636 = _T_3635 - _T_3633;
  assign _T_3637 = $unsigned(_T_3636);
  assign _T_3638 = _T_3637[0:0];
  assign _T_3640 = _T_3633 == 1'h0;
  assign _T_3643 = _T_3640 | _T_3624;
  assign _T_3645 = _T_3643 | reset;
  assign _T_3647 = _T_3645 == 1'h0;
  assign _T_3649 = _T_3630 == 1'h0;
  assign _T_3651 = _T_3624 != 1'h1;
  assign _T_3652 = _T_3649 | _T_3651;
  assign _T_3654 = _T_3652 | reset;
  assign _T_3656 = _T_3654 == 1'h0;
  assign _T_3672 = _T_1720 & _T_1949;
  assign _T_3673 = _T_1853 & _T_1941;
  assign _T_3675 = _T_3673 & _T_1952;
  assign _T_3676 = _T_3666 + _T_3672;
  assign _T_3677 = _T_3676[0:0];
  assign _T_3678 = _T_3677 - _T_3675;
  assign _T_3679 = $unsigned(_T_3678);
  assign _T_3680 = _T_3679[0:0];
  assign _T_3682 = _T_3675 == 1'h0;
  assign _T_3685 = _T_3682 | _T_3666;
  assign _T_3687 = _T_3685 | reset;
  assign _T_3689 = _T_3687 == 1'h0;
  assign _T_3691 = _T_3672 == 1'h0;
  assign _T_3693 = _T_3666 != 1'h1;
  assign _T_3694 = _T_3691 | _T_3693;
  assign _T_3696 = _T_3694 | reset;
  assign _T_3698 = _T_3696 == 1'h0;
  assign _T_3714 = _T_1721 & _T_1949;
  assign _T_3715 = _T_1854 & _T_1941;
  assign _T_3717 = _T_3715 & _T_1952;
  assign _T_3718 = _T_3708 + _T_3714;
  assign _T_3719 = _T_3718[0:0];
  assign _T_3720 = _T_3719 - _T_3717;
  assign _T_3721 = $unsigned(_T_3720);
  assign _T_3722 = _T_3721[0:0];
  assign _T_3724 = _T_3717 == 1'h0;
  assign _T_3727 = _T_3724 | _T_3708;
  assign _T_3729 = _T_3727 | reset;
  assign _T_3731 = _T_3729 == 1'h0;
  assign _T_3733 = _T_3714 == 1'h0;
  assign _T_3735 = _T_3708 != 1'h1;
  assign _T_3736 = _T_3733 | _T_3735;
  assign _T_3738 = _T_3736 | reset;
  assign _T_3740 = _T_3738 == 1'h0;
  assign _T_3756 = _T_1722 & _T_1949;
  assign _T_3757 = _T_1855 & _T_1941;
  assign _T_3759 = _T_3757 & _T_1952;
  assign _T_3760 = _T_3750 + _T_3756;
  assign _T_3761 = _T_3760[0:0];
  assign _T_3762 = _T_3761 - _T_3759;
  assign _T_3763 = $unsigned(_T_3762);
  assign _T_3764 = _T_3763[0:0];
  assign _T_3766 = _T_3759 == 1'h0;
  assign _T_3769 = _T_3766 | _T_3750;
  assign _T_3771 = _T_3769 | reset;
  assign _T_3773 = _T_3771 == 1'h0;
  assign _T_3775 = _T_3756 == 1'h0;
  assign _T_3777 = _T_3750 != 1'h1;
  assign _T_3778 = _T_3775 | _T_3777;
  assign _T_3780 = _T_3778 | reset;
  assign _T_3782 = _T_3780 == 1'h0;
  assign _T_3798 = _T_1723 & _T_1949;
  assign _T_3799 = _T_1856 & _T_1941;
  assign _T_3801 = _T_3799 & _T_1952;
  assign _T_3802 = _T_3792 + _T_3798;
  assign _T_3803 = _T_3802[0:0];
  assign _T_3804 = _T_3803 - _T_3801;
  assign _T_3805 = $unsigned(_T_3804);
  assign _T_3806 = _T_3805[0:0];
  assign _T_3808 = _T_3801 == 1'h0;
  assign _T_3811 = _T_3808 | _T_3792;
  assign _T_3813 = _T_3811 | reset;
  assign _T_3815 = _T_3813 == 1'h0;
  assign _T_3817 = _T_3798 == 1'h0;
  assign _T_3819 = _T_3792 != 1'h1;
  assign _T_3820 = _T_3817 | _T_3819;
  assign _T_3822 = _T_3820 | reset;
  assign _T_3824 = _T_3822 == 1'h0;
  assign _T_3840 = _T_1724 & _T_1949;
  assign _T_3841 = _T_1857 & _T_1941;
  assign _T_3843 = _T_3841 & _T_1952;
  assign _T_3844 = _T_3834 + _T_3840;
  assign _T_3845 = _T_3844[0:0];
  assign _T_3846 = _T_3845 - _T_3843;
  assign _T_3847 = $unsigned(_T_3846);
  assign _T_3848 = _T_3847[0:0];
  assign _T_3850 = _T_3843 == 1'h0;
  assign _T_3853 = _T_3850 | _T_3834;
  assign _T_3855 = _T_3853 | reset;
  assign _T_3857 = _T_3855 == 1'h0;
  assign _T_3859 = _T_3840 == 1'h0;
  assign _T_3861 = _T_3834 != 1'h1;
  assign _T_3862 = _T_3859 | _T_3861;
  assign _T_3864 = _T_3862 | reset;
  assign _T_3866 = _T_3864 == 1'h0;
  assign _T_3882 = _T_1725 & _T_1949;
  assign _T_3883 = _T_1858 & _T_1941;
  assign _T_3885 = _T_3883 & _T_1952;
  assign _T_3886 = _T_3876 + _T_3882;
  assign _T_3887 = _T_3886[0:0];
  assign _T_3888 = _T_3887 - _T_3885;
  assign _T_3889 = $unsigned(_T_3888);
  assign _T_3890 = _T_3889[0:0];
  assign _T_3892 = _T_3885 == 1'h0;
  assign _T_3895 = _T_3892 | _T_3876;
  assign _T_3897 = _T_3895 | reset;
  assign _T_3899 = _T_3897 == 1'h0;
  assign _T_3901 = _T_3882 == 1'h0;
  assign _T_3903 = _T_3876 != 1'h1;
  assign _T_3904 = _T_3901 | _T_3903;
  assign _T_3906 = _T_3904 | reset;
  assign _T_3908 = _T_3906 == 1'h0;
  assign _T_3924 = _T_1726 & _T_1949;
  assign _T_3925 = _T_1859 & _T_1941;
  assign _T_3927 = _T_3925 & _T_1952;
  assign _T_3928 = _T_3918 + _T_3924;
  assign _T_3929 = _T_3928[0:0];
  assign _T_3930 = _T_3929 - _T_3927;
  assign _T_3931 = $unsigned(_T_3930);
  assign _T_3932 = _T_3931[0:0];
  assign _T_3934 = _T_3927 == 1'h0;
  assign _T_3937 = _T_3934 | _T_3918;
  assign _T_3939 = _T_3937 | reset;
  assign _T_3941 = _T_3939 == 1'h0;
  assign _T_3943 = _T_3924 == 1'h0;
  assign _T_3945 = _T_3918 != 1'h1;
  assign _T_3946 = _T_3943 | _T_3945;
  assign _T_3948 = _T_3946 | reset;
  assign _T_3950 = _T_3948 == 1'h0;
  assign _T_3966 = _T_1727 & _T_1949;
  assign _T_3967 = _T_1860 & _T_1941;
  assign _T_3969 = _T_3967 & _T_1952;
  assign _T_3970 = _T_3960 + _T_3966;
  assign _T_3971 = _T_3970[0:0];
  assign _T_3972 = _T_3971 - _T_3969;
  assign _T_3973 = $unsigned(_T_3972);
  assign _T_3974 = _T_3973[0:0];
  assign _T_3976 = _T_3969 == 1'h0;
  assign _T_3979 = _T_3976 | _T_3960;
  assign _T_3981 = _T_3979 | reset;
  assign _T_3983 = _T_3981 == 1'h0;
  assign _T_3985 = _T_3966 == 1'h0;
  assign _T_3987 = _T_3960 != 1'h1;
  assign _T_3988 = _T_3985 | _T_3987;
  assign _T_3990 = _T_3988 | reset;
  assign _T_3992 = _T_3990 == 1'h0;
  assign _T_4008 = _T_1728 & _T_1949;
  assign _T_4009 = _T_1861 & _T_1941;
  assign _T_4011 = _T_4009 & _T_1952;
  assign _T_4012 = _T_4002 + _T_4008;
  assign _T_4013 = _T_4012[0:0];
  assign _T_4014 = _T_4013 - _T_4011;
  assign _T_4015 = $unsigned(_T_4014);
  assign _T_4016 = _T_4015[0:0];
  assign _T_4018 = _T_4011 == 1'h0;
  assign _T_4021 = _T_4018 | _T_4002;
  assign _T_4023 = _T_4021 | reset;
  assign _T_4025 = _T_4023 == 1'h0;
  assign _T_4027 = _T_4008 == 1'h0;
  assign _T_4029 = _T_4002 != 1'h1;
  assign _T_4030 = _T_4027 | _T_4029;
  assign _T_4032 = _T_4030 | reset;
  assign _T_4034 = _T_4032 == 1'h0;
  assign _T_4050 = _T_1729 & _T_1949;
  assign _T_4051 = _T_1862 & _T_1941;
  assign _T_4053 = _T_4051 & _T_1952;
  assign _T_4054 = _T_4044 + _T_4050;
  assign _T_4055 = _T_4054[0:0];
  assign _T_4056 = _T_4055 - _T_4053;
  assign _T_4057 = $unsigned(_T_4056);
  assign _T_4058 = _T_4057[0:0];
  assign _T_4060 = _T_4053 == 1'h0;
  assign _T_4063 = _T_4060 | _T_4044;
  assign _T_4065 = _T_4063 | reset;
  assign _T_4067 = _T_4065 == 1'h0;
  assign _T_4069 = _T_4050 == 1'h0;
  assign _T_4071 = _T_4044 != 1'h1;
  assign _T_4072 = _T_4069 | _T_4071;
  assign _T_4074 = _T_4072 | reset;
  assign _T_4076 = _T_4074 == 1'h0;
  assign _T_4092 = _T_1730 & _T_1949;
  assign _T_4093 = _T_1863 & _T_1941;
  assign _T_4095 = _T_4093 & _T_1952;
  assign _T_4096 = _T_4086 + _T_4092;
  assign _T_4097 = _T_4096[0:0];
  assign _T_4098 = _T_4097 - _T_4095;
  assign _T_4099 = $unsigned(_T_4098);
  assign _T_4100 = _T_4099[0:0];
  assign _T_4102 = _T_4095 == 1'h0;
  assign _T_4105 = _T_4102 | _T_4086;
  assign _T_4107 = _T_4105 | reset;
  assign _T_4109 = _T_4107 == 1'h0;
  assign _T_4111 = _T_4092 == 1'h0;
  assign _T_4113 = _T_4086 != 1'h1;
  assign _T_4114 = _T_4111 | _T_4113;
  assign _T_4116 = _T_4114 | reset;
  assign _T_4118 = _T_4116 == 1'h0;
  assign _T_4134 = _T_1731 & _T_1949;
  assign _T_4135 = _T_1864 & _T_1941;
  assign _T_4137 = _T_4135 & _T_1952;
  assign _T_4138 = _T_4128 + _T_4134;
  assign _T_4139 = _T_4138[0:0];
  assign _T_4140 = _T_4139 - _T_4137;
  assign _T_4141 = $unsigned(_T_4140);
  assign _T_4142 = _T_4141[0:0];
  assign _T_4144 = _T_4137 == 1'h0;
  assign _T_4147 = _T_4144 | _T_4128;
  assign _T_4149 = _T_4147 | reset;
  assign _T_4151 = _T_4149 == 1'h0;
  assign _T_4153 = _T_4134 == 1'h0;
  assign _T_4155 = _T_4128 != 1'h1;
  assign _T_4156 = _T_4153 | _T_4155;
  assign _T_4158 = _T_4156 | reset;
  assign _T_4160 = _T_4158 == 1'h0;
  assign _T_4176 = _T_1732 & _T_1949;
  assign _T_4177 = _T_1865 & _T_1941;
  assign _T_4179 = _T_4177 & _T_1952;
  assign _T_4180 = _T_4170 + _T_4176;
  assign _T_4181 = _T_4180[0:0];
  assign _T_4182 = _T_4181 - _T_4179;
  assign _T_4183 = $unsigned(_T_4182);
  assign _T_4184 = _T_4183[0:0];
  assign _T_4186 = _T_4179 == 1'h0;
  assign _T_4189 = _T_4186 | _T_4170;
  assign _T_4191 = _T_4189 | reset;
  assign _T_4193 = _T_4191 == 1'h0;
  assign _T_4195 = _T_4176 == 1'h0;
  assign _T_4197 = _T_4170 != 1'h1;
  assign _T_4198 = _T_4195 | _T_4197;
  assign _T_4200 = _T_4198 | reset;
  assign _T_4202 = _T_4200 == 1'h0;
  assign _T_4218 = _T_1733 & _T_1949;
  assign _T_4219 = _T_1866 & _T_1941;
  assign _T_4221 = _T_4219 & _T_1952;
  assign _T_4222 = _T_4212 + _T_4218;
  assign _T_4223 = _T_4222[0:0];
  assign _T_4224 = _T_4223 - _T_4221;
  assign _T_4225 = $unsigned(_T_4224);
  assign _T_4226 = _T_4225[0:0];
  assign _T_4228 = _T_4221 == 1'h0;
  assign _T_4231 = _T_4228 | _T_4212;
  assign _T_4233 = _T_4231 | reset;
  assign _T_4235 = _T_4233 == 1'h0;
  assign _T_4237 = _T_4218 == 1'h0;
  assign _T_4239 = _T_4212 != 1'h1;
  assign _T_4240 = _T_4237 | _T_4239;
  assign _T_4242 = _T_4240 | reset;
  assign _T_4244 = _T_4242 == 1'h0;
  assign _T_4260 = _T_1734 & _T_1949;
  assign _T_4261 = _T_1867 & _T_1941;
  assign _T_4263 = _T_4261 & _T_1952;
  assign _T_4264 = _T_4254 + _T_4260;
  assign _T_4265 = _T_4264[0:0];
  assign _T_4266 = _T_4265 - _T_4263;
  assign _T_4267 = $unsigned(_T_4266);
  assign _T_4268 = _T_4267[0:0];
  assign _T_4270 = _T_4263 == 1'h0;
  assign _T_4273 = _T_4270 | _T_4254;
  assign _T_4275 = _T_4273 | reset;
  assign _T_4277 = _T_4275 == 1'h0;
  assign _T_4279 = _T_4260 == 1'h0;
  assign _T_4281 = _T_4254 != 1'h1;
  assign _T_4282 = _T_4279 | _T_4281;
  assign _T_4284 = _T_4282 | reset;
  assign _T_4286 = _T_4284 == 1'h0;
  assign _T_4302 = _T_1735 & _T_1949;
  assign _T_4303 = _T_1868 & _T_1941;
  assign _T_4305 = _T_4303 & _T_1952;
  assign _T_4306 = _T_4296 + _T_4302;
  assign _T_4307 = _T_4306[0:0];
  assign _T_4308 = _T_4307 - _T_4305;
  assign _T_4309 = $unsigned(_T_4308);
  assign _T_4310 = _T_4309[0:0];
  assign _T_4312 = _T_4305 == 1'h0;
  assign _T_4315 = _T_4312 | _T_4296;
  assign _T_4317 = _T_4315 | reset;
  assign _T_4319 = _T_4317 == 1'h0;
  assign _T_4321 = _T_4302 == 1'h0;
  assign _T_4323 = _T_4296 != 1'h1;
  assign _T_4324 = _T_4321 | _T_4323;
  assign _T_4326 = _T_4324 | reset;
  assign _T_4328 = _T_4326 == 1'h0;
  assign _T_4344 = _T_1736 & _T_1949;
  assign _T_4345 = _T_1869 & _T_1941;
  assign _T_4347 = _T_4345 & _T_1952;
  assign _T_4348 = _T_4338 + _T_4344;
  assign _T_4349 = _T_4348[0:0];
  assign _T_4350 = _T_4349 - _T_4347;
  assign _T_4351 = $unsigned(_T_4350);
  assign _T_4352 = _T_4351[0:0];
  assign _T_4354 = _T_4347 == 1'h0;
  assign _T_4357 = _T_4354 | _T_4338;
  assign _T_4359 = _T_4357 | reset;
  assign _T_4361 = _T_4359 == 1'h0;
  assign _T_4363 = _T_4344 == 1'h0;
  assign _T_4365 = _T_4338 != 1'h1;
  assign _T_4366 = _T_4363 | _T_4365;
  assign _T_4368 = _T_4366 | reset;
  assign _T_4370 = _T_4368 == 1'h0;
  assign _T_4386 = _T_1737 & _T_1949;
  assign _T_4387 = _T_1870 & _T_1941;
  assign _T_4389 = _T_4387 & _T_1952;
  assign _T_4390 = _T_4380 + _T_4386;
  assign _T_4391 = _T_4390[0:0];
  assign _T_4392 = _T_4391 - _T_4389;
  assign _T_4393 = $unsigned(_T_4392);
  assign _T_4394 = _T_4393[0:0];
  assign _T_4396 = _T_4389 == 1'h0;
  assign _T_4399 = _T_4396 | _T_4380;
  assign _T_4401 = _T_4399 | reset;
  assign _T_4403 = _T_4401 == 1'h0;
  assign _T_4405 = _T_4386 == 1'h0;
  assign _T_4407 = _T_4380 != 1'h1;
  assign _T_4408 = _T_4405 | _T_4407;
  assign _T_4410 = _T_4408 | reset;
  assign _T_4412 = _T_4410 == 1'h0;
  assign _T_4428 = _T_1738 & _T_1949;
  assign _T_4429 = _T_1871 & _T_1941;
  assign _T_4431 = _T_4429 & _T_1952;
  assign _T_4432 = _T_4422 + _T_4428;
  assign _T_4433 = _T_4432[0:0];
  assign _T_4434 = _T_4433 - _T_4431;
  assign _T_4435 = $unsigned(_T_4434);
  assign _T_4436 = _T_4435[0:0];
  assign _T_4438 = _T_4431 == 1'h0;
  assign _T_4441 = _T_4438 | _T_4422;
  assign _T_4443 = _T_4441 | reset;
  assign _T_4445 = _T_4443 == 1'h0;
  assign _T_4447 = _T_4428 == 1'h0;
  assign _T_4449 = _T_4422 != 1'h1;
  assign _T_4450 = _T_4447 | _T_4449;
  assign _T_4452 = _T_4450 | reset;
  assign _T_4454 = _T_4452 == 1'h0;
  assign _T_4470 = _T_1739 & _T_1949;
  assign _T_4471 = _T_1872 & _T_1941;
  assign _T_4473 = _T_4471 & _T_1952;
  assign _T_4474 = _T_4464 + _T_4470;
  assign _T_4475 = _T_4474[0:0];
  assign _T_4476 = _T_4475 - _T_4473;
  assign _T_4477 = $unsigned(_T_4476);
  assign _T_4478 = _T_4477[0:0];
  assign _T_4480 = _T_4473 == 1'h0;
  assign _T_4483 = _T_4480 | _T_4464;
  assign _T_4485 = _T_4483 | reset;
  assign _T_4487 = _T_4485 == 1'h0;
  assign _T_4489 = _T_4470 == 1'h0;
  assign _T_4491 = _T_4464 != 1'h1;
  assign _T_4492 = _T_4489 | _T_4491;
  assign _T_4494 = _T_4492 | reset;
  assign _T_4496 = _T_4494 == 1'h0;
  assign _T_4512 = _T_1740 & _T_1949;
  assign _T_4513 = _T_1873 & _T_1941;
  assign _T_4515 = _T_4513 & _T_1952;
  assign _T_4516 = _T_4506 + _T_4512;
  assign _T_4517 = _T_4516[0:0];
  assign _T_4518 = _T_4517 - _T_4515;
  assign _T_4519 = $unsigned(_T_4518);
  assign _T_4520 = _T_4519[0:0];
  assign _T_4522 = _T_4515 == 1'h0;
  assign _T_4525 = _T_4522 | _T_4506;
  assign _T_4527 = _T_4525 | reset;
  assign _T_4529 = _T_4527 == 1'h0;
  assign _T_4531 = _T_4512 == 1'h0;
  assign _T_4533 = _T_4506 != 1'h1;
  assign _T_4534 = _T_4531 | _T_4533;
  assign _T_4536 = _T_4534 | reset;
  assign _T_4538 = _T_4536 == 1'h0;
  assign _T_4554 = _T_1741 & _T_1949;
  assign _T_4555 = _T_1874 & _T_1941;
  assign _T_4557 = _T_4555 & _T_1952;
  assign _T_4558 = _T_4548 + _T_4554;
  assign _T_4559 = _T_4558[0:0];
  assign _T_4560 = _T_4559 - _T_4557;
  assign _T_4561 = $unsigned(_T_4560);
  assign _T_4562 = _T_4561[0:0];
  assign _T_4564 = _T_4557 == 1'h0;
  assign _T_4567 = _T_4564 | _T_4548;
  assign _T_4569 = _T_4567 | reset;
  assign _T_4571 = _T_4569 == 1'h0;
  assign _T_4573 = _T_4554 == 1'h0;
  assign _T_4575 = _T_4548 != 1'h1;
  assign _T_4576 = _T_4573 | _T_4575;
  assign _T_4578 = _T_4576 | reset;
  assign _T_4580 = _T_4578 == 1'h0;
  assign _T_4596 = _T_1742 & _T_1949;
  assign _T_4597 = _T_1875 & _T_1941;
  assign _T_4599 = _T_4597 & _T_1952;
  assign _T_4600 = _T_4590 + _T_4596;
  assign _T_4601 = _T_4600[0:0];
  assign _T_4602 = _T_4601 - _T_4599;
  assign _T_4603 = $unsigned(_T_4602);
  assign _T_4604 = _T_4603[0:0];
  assign _T_4606 = _T_4599 == 1'h0;
  assign _T_4609 = _T_4606 | _T_4590;
  assign _T_4611 = _T_4609 | reset;
  assign _T_4613 = _T_4611 == 1'h0;
  assign _T_4615 = _T_4596 == 1'h0;
  assign _T_4617 = _T_4590 != 1'h1;
  assign _T_4618 = _T_4615 | _T_4617;
  assign _T_4620 = _T_4618 | reset;
  assign _T_4622 = _T_4620 == 1'h0;
  assign _T_4638 = _T_1743 & _T_1949;
  assign _T_4639 = _T_1876 & _T_1941;
  assign _T_4641 = _T_4639 & _T_1952;
  assign _T_4642 = _T_4632 + _T_4638;
  assign _T_4643 = _T_4642[0:0];
  assign _T_4644 = _T_4643 - _T_4641;
  assign _T_4645 = $unsigned(_T_4644);
  assign _T_4646 = _T_4645[0:0];
  assign _T_4648 = _T_4641 == 1'h0;
  assign _T_4651 = _T_4648 | _T_4632;
  assign _T_4653 = _T_4651 | reset;
  assign _T_4655 = _T_4653 == 1'h0;
  assign _T_4657 = _T_4638 == 1'h0;
  assign _T_4659 = _T_4632 != 1'h1;
  assign _T_4660 = _T_4657 | _T_4659;
  assign _T_4662 = _T_4660 | reset;
  assign _T_4664 = _T_4662 == 1'h0;
  assign _T_4680 = _T_1744 & _T_1949;
  assign _T_4681 = _T_1877 & _T_1941;
  assign _T_4683 = _T_4681 & _T_1952;
  assign _T_4684 = _T_4674 + _T_4680;
  assign _T_4685 = _T_4684[0:0];
  assign _T_4686 = _T_4685 - _T_4683;
  assign _T_4687 = $unsigned(_T_4686);
  assign _T_4688 = _T_4687[0:0];
  assign _T_4690 = _T_4683 == 1'h0;
  assign _T_4693 = _T_4690 | _T_4674;
  assign _T_4695 = _T_4693 | reset;
  assign _T_4697 = _T_4695 == 1'h0;
  assign _T_4699 = _T_4680 == 1'h0;
  assign _T_4701 = _T_4674 != 1'h1;
  assign _T_4702 = _T_4699 | _T_4701;
  assign _T_4704 = _T_4702 | reset;
  assign _T_4706 = _T_4704 == 1'h0;
  assign _T_4722 = _T_1745 & _T_1949;
  assign _T_4723 = _T_1878 & _T_1941;
  assign _T_4725 = _T_4723 & _T_1952;
  assign _T_4726 = _T_4716 + _T_4722;
  assign _T_4727 = _T_4726[0:0];
  assign _T_4728 = _T_4727 - _T_4725;
  assign _T_4729 = $unsigned(_T_4728);
  assign _T_4730 = _T_4729[0:0];
  assign _T_4732 = _T_4725 == 1'h0;
  assign _T_4735 = _T_4732 | _T_4716;
  assign _T_4737 = _T_4735 | reset;
  assign _T_4739 = _T_4737 == 1'h0;
  assign _T_4741 = _T_4722 == 1'h0;
  assign _T_4743 = _T_4716 != 1'h1;
  assign _T_4744 = _T_4741 | _T_4743;
  assign _T_4746 = _T_4744 | reset;
  assign _T_4748 = _T_4746 == 1'h0;
  assign _T_4764 = _T_1746 & _T_1949;
  assign _T_4765 = _T_1879 & _T_1941;
  assign _T_4767 = _T_4765 & _T_1952;
  assign _T_4768 = _T_4758 + _T_4764;
  assign _T_4769 = _T_4768[0:0];
  assign _T_4770 = _T_4769 - _T_4767;
  assign _T_4771 = $unsigned(_T_4770);
  assign _T_4772 = _T_4771[0:0];
  assign _T_4774 = _T_4767 == 1'h0;
  assign _T_4777 = _T_4774 | _T_4758;
  assign _T_4779 = _T_4777 | reset;
  assign _T_4781 = _T_4779 == 1'h0;
  assign _T_4783 = _T_4764 == 1'h0;
  assign _T_4785 = _T_4758 != 1'h1;
  assign _T_4786 = _T_4783 | _T_4785;
  assign _T_4788 = _T_4786 | reset;
  assign _T_4790 = _T_4788 == 1'h0;
  assign _T_4806 = _T_1747 & _T_1949;
  assign _T_4807 = _T_1880 & _T_1941;
  assign _T_4809 = _T_4807 & _T_1952;
  assign _T_4810 = _T_4800 + _T_4806;
  assign _T_4811 = _T_4810[0:0];
  assign _T_4812 = _T_4811 - _T_4809;
  assign _T_4813 = $unsigned(_T_4812);
  assign _T_4814 = _T_4813[0:0];
  assign _T_4816 = _T_4809 == 1'h0;
  assign _T_4819 = _T_4816 | _T_4800;
  assign _T_4821 = _T_4819 | reset;
  assign _T_4823 = _T_4821 == 1'h0;
  assign _T_4825 = _T_4806 == 1'h0;
  assign _T_4827 = _T_4800 != 1'h1;
  assign _T_4828 = _T_4825 | _T_4827;
  assign _T_4830 = _T_4828 | reset;
  assign _T_4832 = _T_4830 == 1'h0;
  assign _T_4848 = _T_1748 & _T_1949;
  assign _T_4849 = _T_1881 & _T_1941;
  assign _T_4851 = _T_4849 & _T_1952;
  assign _T_4852 = _T_4842 + _T_4848;
  assign _T_4853 = _T_4852[0:0];
  assign _T_4854 = _T_4853 - _T_4851;
  assign _T_4855 = $unsigned(_T_4854);
  assign _T_4856 = _T_4855[0:0];
  assign _T_4858 = _T_4851 == 1'h0;
  assign _T_4861 = _T_4858 | _T_4842;
  assign _T_4863 = _T_4861 | reset;
  assign _T_4865 = _T_4863 == 1'h0;
  assign _T_4867 = _T_4848 == 1'h0;
  assign _T_4869 = _T_4842 != 1'h1;
  assign _T_4870 = _T_4867 | _T_4869;
  assign _T_4872 = _T_4870 | reset;
  assign _T_4874 = _T_4872 == 1'h0;
  assign _T_4890 = _T_1749 & _T_1949;
  assign _T_4891 = _T_1882 & _T_1941;
  assign _T_4893 = _T_4891 & _T_1952;
  assign _T_4894 = _T_4884 + _T_4890;
  assign _T_4895 = _T_4894[0:0];
  assign _T_4896 = _T_4895 - _T_4893;
  assign _T_4897 = $unsigned(_T_4896);
  assign _T_4898 = _T_4897[0:0];
  assign _T_4900 = _T_4893 == 1'h0;
  assign _T_4903 = _T_4900 | _T_4884;
  assign _T_4905 = _T_4903 | reset;
  assign _T_4907 = _T_4905 == 1'h0;
  assign _T_4909 = _T_4890 == 1'h0;
  assign _T_4911 = _T_4884 != 1'h1;
  assign _T_4912 = _T_4909 | _T_4911;
  assign _T_4914 = _T_4912 | reset;
  assign _T_4916 = _T_4914 == 1'h0;
  assign _T_4932 = _T_1750 & _T_1949;
  assign _T_4933 = _T_1883 & _T_1941;
  assign _T_4935 = _T_4933 & _T_1952;
  assign _T_4936 = _T_4926 + _T_4932;
  assign _T_4937 = _T_4936[0:0];
  assign _T_4938 = _T_4937 - _T_4935;
  assign _T_4939 = $unsigned(_T_4938);
  assign _T_4940 = _T_4939[0:0];
  assign _T_4942 = _T_4935 == 1'h0;
  assign _T_4945 = _T_4942 | _T_4926;
  assign _T_4947 = _T_4945 | reset;
  assign _T_4949 = _T_4947 == 1'h0;
  assign _T_4951 = _T_4932 == 1'h0;
  assign _T_4953 = _T_4926 != 1'h1;
  assign _T_4954 = _T_4951 | _T_4953;
  assign _T_4956 = _T_4954 | reset;
  assign _T_4958 = _T_4956 == 1'h0;
  assign _T_4974 = _T_1751 & _T_1949;
  assign _T_4975 = _T_1884 & _T_1941;
  assign _T_4977 = _T_4975 & _T_1952;
  assign _T_4978 = _T_4968 + _T_4974;
  assign _T_4979 = _T_4978[0:0];
  assign _T_4980 = _T_4979 - _T_4977;
  assign _T_4981 = $unsigned(_T_4980);
  assign _T_4982 = _T_4981[0:0];
  assign _T_4984 = _T_4977 == 1'h0;
  assign _T_4987 = _T_4984 | _T_4968;
  assign _T_4989 = _T_4987 | reset;
  assign _T_4991 = _T_4989 == 1'h0;
  assign _T_4993 = _T_4974 == 1'h0;
  assign _T_4995 = _T_4968 != 1'h1;
  assign _T_4996 = _T_4993 | _T_4995;
  assign _T_4998 = _T_4996 | reset;
  assign _T_5000 = _T_4998 == 1'h0;
  assign _T_5016 = _T_1752 & _T_1949;
  assign _T_5017 = _T_1885 & _T_1941;
  assign _T_5019 = _T_5017 & _T_1952;
  assign _T_5020 = _T_5010 + _T_5016;
  assign _T_5021 = _T_5020[0:0];
  assign _T_5022 = _T_5021 - _T_5019;
  assign _T_5023 = $unsigned(_T_5022);
  assign _T_5024 = _T_5023[0:0];
  assign _T_5026 = _T_5019 == 1'h0;
  assign _T_5029 = _T_5026 | _T_5010;
  assign _T_5031 = _T_5029 | reset;
  assign _T_5033 = _T_5031 == 1'h0;
  assign _T_5035 = _T_5016 == 1'h0;
  assign _T_5037 = _T_5010 != 1'h1;
  assign _T_5038 = _T_5035 | _T_5037;
  assign _T_5040 = _T_5038 | reset;
  assign _T_5042 = _T_5040 == 1'h0;
  assign _T_5058 = _T_1753 & _T_1949;
  assign _T_5059 = _T_1886 & _T_1941;
  assign _T_5061 = _T_5059 & _T_1952;
  assign _T_5062 = _T_5052 + _T_5058;
  assign _T_5063 = _T_5062[0:0];
  assign _T_5064 = _T_5063 - _T_5061;
  assign _T_5065 = $unsigned(_T_5064);
  assign _T_5066 = _T_5065[0:0];
  assign _T_5068 = _T_5061 == 1'h0;
  assign _T_5071 = _T_5068 | _T_5052;
  assign _T_5073 = _T_5071 | reset;
  assign _T_5075 = _T_5073 == 1'h0;
  assign _T_5077 = _T_5058 == 1'h0;
  assign _T_5079 = _T_5052 != 1'h1;
  assign _T_5080 = _T_5077 | _T_5079;
  assign _T_5082 = _T_5080 | reset;
  assign _T_5084 = _T_5082 == 1'h0;
  assign _T_5100 = _T_1754 & _T_1949;
  assign _T_5101 = _T_1887 & _T_1941;
  assign _T_5103 = _T_5101 & _T_1952;
  assign _T_5104 = _T_5094 + _T_5100;
  assign _T_5105 = _T_5104[0:0];
  assign _T_5106 = _T_5105 - _T_5103;
  assign _T_5107 = $unsigned(_T_5106);
  assign _T_5108 = _T_5107[0:0];
  assign _T_5110 = _T_5103 == 1'h0;
  assign _T_5113 = _T_5110 | _T_5094;
  assign _T_5115 = _T_5113 | reset;
  assign _T_5117 = _T_5115 == 1'h0;
  assign _T_5119 = _T_5100 == 1'h0;
  assign _T_5121 = _T_5094 != 1'h1;
  assign _T_5122 = _T_5119 | _T_5121;
  assign _T_5124 = _T_5122 | reset;
  assign _T_5126 = _T_5124 == 1'h0;
  assign _T_5142 = _T_1755 & _T_1949;
  assign _T_5143 = _T_1888 & _T_1941;
  assign _T_5145 = _T_5143 & _T_1952;
  assign _T_5146 = _T_5136 + _T_5142;
  assign _T_5147 = _T_5146[0:0];
  assign _T_5148 = _T_5147 - _T_5145;
  assign _T_5149 = $unsigned(_T_5148);
  assign _T_5150 = _T_5149[0:0];
  assign _T_5152 = _T_5145 == 1'h0;
  assign _T_5155 = _T_5152 | _T_5136;
  assign _T_5157 = _T_5155 | reset;
  assign _T_5159 = _T_5157 == 1'h0;
  assign _T_5161 = _T_5142 == 1'h0;
  assign _T_5163 = _T_5136 != 1'h1;
  assign _T_5164 = _T_5161 | _T_5163;
  assign _T_5166 = _T_5164 | reset;
  assign _T_5168 = _T_5166 == 1'h0;
  assign _T_5184 = _T_1756 & _T_1949;
  assign _T_5185 = _T_1889 & _T_1941;
  assign _T_5187 = _T_5185 & _T_1952;
  assign _T_5188 = _T_5178 + _T_5184;
  assign _T_5189 = _T_5188[0:0];
  assign _T_5190 = _T_5189 - _T_5187;
  assign _T_5191 = $unsigned(_T_5190);
  assign _T_5192 = _T_5191[0:0];
  assign _T_5194 = _T_5187 == 1'h0;
  assign _T_5197 = _T_5194 | _T_5178;
  assign _T_5199 = _T_5197 | reset;
  assign _T_5201 = _T_5199 == 1'h0;
  assign _T_5203 = _T_5184 == 1'h0;
  assign _T_5205 = _T_5178 != 1'h1;
  assign _T_5206 = _T_5203 | _T_5205;
  assign _T_5208 = _T_5206 | reset;
  assign _T_5210 = _T_5208 == 1'h0;
  assign _T_5226 = _T_1757 & _T_1949;
  assign _T_5227 = _T_1890 & _T_1941;
  assign _T_5229 = _T_5227 & _T_1952;
  assign _T_5230 = _T_5220 + _T_5226;
  assign _T_5231 = _T_5230[0:0];
  assign _T_5232 = _T_5231 - _T_5229;
  assign _T_5233 = $unsigned(_T_5232);
  assign _T_5234 = _T_5233[0:0];
  assign _T_5236 = _T_5229 == 1'h0;
  assign _T_5239 = _T_5236 | _T_5220;
  assign _T_5241 = _T_5239 | reset;
  assign _T_5243 = _T_5241 == 1'h0;
  assign _T_5245 = _T_5226 == 1'h0;
  assign _T_5247 = _T_5220 != 1'h1;
  assign _T_5248 = _T_5245 | _T_5247;
  assign _T_5250 = _T_5248 | reset;
  assign _T_5252 = _T_5250 == 1'h0;
  assign _T_5268 = _T_1758 & _T_1949;
  assign _T_5269 = _T_1891 & _T_1941;
  assign _T_5271 = _T_5269 & _T_1952;
  assign _T_5272 = _T_5262 + _T_5268;
  assign _T_5273 = _T_5272[0:0];
  assign _T_5274 = _T_5273 - _T_5271;
  assign _T_5275 = $unsigned(_T_5274);
  assign _T_5276 = _T_5275[0:0];
  assign _T_5278 = _T_5271 == 1'h0;
  assign _T_5281 = _T_5278 | _T_5262;
  assign _T_5283 = _T_5281 | reset;
  assign _T_5285 = _T_5283 == 1'h0;
  assign _T_5287 = _T_5268 == 1'h0;
  assign _T_5289 = _T_5262 != 1'h1;
  assign _T_5290 = _T_5287 | _T_5289;
  assign _T_5292 = _T_5290 | reset;
  assign _T_5294 = _T_5292 == 1'h0;
  assign _T_5310 = _T_1759 & _T_1949;
  assign _T_5311 = _T_1892 & _T_1941;
  assign _T_5313 = _T_5311 & _T_1952;
  assign _T_5314 = _T_5304 + _T_5310;
  assign _T_5315 = _T_5314[0:0];
  assign _T_5316 = _T_5315 - _T_5313;
  assign _T_5317 = $unsigned(_T_5316);
  assign _T_5318 = _T_5317[0:0];
  assign _T_5320 = _T_5313 == 1'h0;
  assign _T_5323 = _T_5320 | _T_5304;
  assign _T_5325 = _T_5323 | reset;
  assign _T_5327 = _T_5325 == 1'h0;
  assign _T_5329 = _T_5310 == 1'h0;
  assign _T_5331 = _T_5304 != 1'h1;
  assign _T_5332 = _T_5329 | _T_5331;
  assign _T_5334 = _T_5332 | reset;
  assign _T_5336 = _T_5334 == 1'h0;
  assign _T_5352 = _T_1760 & _T_1949;
  assign _T_5353 = _T_1893 & _T_1941;
  assign _T_5355 = _T_5353 & _T_1952;
  assign _T_5356 = _T_5346 + _T_5352;
  assign _T_5357 = _T_5356[0:0];
  assign _T_5358 = _T_5357 - _T_5355;
  assign _T_5359 = $unsigned(_T_5358);
  assign _T_5360 = _T_5359[0:0];
  assign _T_5362 = _T_5355 == 1'h0;
  assign _T_5365 = _T_5362 | _T_5346;
  assign _T_5367 = _T_5365 | reset;
  assign _T_5369 = _T_5367 == 1'h0;
  assign _T_5371 = _T_5352 == 1'h0;
  assign _T_5373 = _T_5346 != 1'h1;
  assign _T_5374 = _T_5371 | _T_5373;
  assign _T_5376 = _T_5374 | reset;
  assign _T_5378 = _T_5376 == 1'h0;
  assign _T_5394 = _T_1761 & _T_1949;
  assign _T_5395 = _T_1894 & _T_1941;
  assign _T_5397 = _T_5395 & _T_1952;
  assign _T_5398 = _T_5388 + _T_5394;
  assign _T_5399 = _T_5398[0:0];
  assign _T_5400 = _T_5399 - _T_5397;
  assign _T_5401 = $unsigned(_T_5400);
  assign _T_5402 = _T_5401[0:0];
  assign _T_5404 = _T_5397 == 1'h0;
  assign _T_5407 = _T_5404 | _T_5388;
  assign _T_5409 = _T_5407 | reset;
  assign _T_5411 = _T_5409 == 1'h0;
  assign _T_5413 = _T_5394 == 1'h0;
  assign _T_5415 = _T_5388 != 1'h1;
  assign _T_5416 = _T_5413 | _T_5415;
  assign _T_5418 = _T_5416 | reset;
  assign _T_5420 = _T_5418 == 1'h0;
  assign _T_5436 = _T_1762 & _T_1949;
  assign _T_5437 = _T_1895 & _T_1941;
  assign _T_5439 = _T_5437 & _T_1952;
  assign _T_5440 = _T_5430 + _T_5436;
  assign _T_5441 = _T_5440[0:0];
  assign _T_5442 = _T_5441 - _T_5439;
  assign _T_5443 = $unsigned(_T_5442);
  assign _T_5444 = _T_5443[0:0];
  assign _T_5446 = _T_5439 == 1'h0;
  assign _T_5449 = _T_5446 | _T_5430;
  assign _T_5451 = _T_5449 | reset;
  assign _T_5453 = _T_5451 == 1'h0;
  assign _T_5455 = _T_5436 == 1'h0;
  assign _T_5457 = _T_5430 != 1'h1;
  assign _T_5458 = _T_5455 | _T_5457;
  assign _T_5460 = _T_5458 | reset;
  assign _T_5462 = _T_5460 == 1'h0;
  assign _T_5478 = _T_1763 & _T_1949;
  assign _T_5479 = _T_1896 & _T_1941;
  assign _T_5481 = _T_5479 & _T_1952;
  assign _T_5482 = _T_5472 + _T_5478;
  assign _T_5483 = _T_5482[0:0];
  assign _T_5484 = _T_5483 - _T_5481;
  assign _T_5485 = $unsigned(_T_5484);
  assign _T_5486 = _T_5485[0:0];
  assign _T_5488 = _T_5481 == 1'h0;
  assign _T_5491 = _T_5488 | _T_5472;
  assign _T_5493 = _T_5491 | reset;
  assign _T_5495 = _T_5493 == 1'h0;
  assign _T_5497 = _T_5478 == 1'h0;
  assign _T_5499 = _T_5472 != 1'h1;
  assign _T_5500 = _T_5497 | _T_5499;
  assign _T_5502 = _T_5500 | reset;
  assign _T_5504 = _T_5502 == 1'h0;
  assign _T_5520 = _T_1764 & _T_1949;
  assign _T_5521 = _T_1897 & _T_1941;
  assign _T_5523 = _T_5521 & _T_1952;
  assign _T_5524 = _T_5514 + _T_5520;
  assign _T_5525 = _T_5524[0:0];
  assign _T_5526 = _T_5525 - _T_5523;
  assign _T_5527 = $unsigned(_T_5526);
  assign _T_5528 = _T_5527[0:0];
  assign _T_5530 = _T_5523 == 1'h0;
  assign _T_5533 = _T_5530 | _T_5514;
  assign _T_5535 = _T_5533 | reset;
  assign _T_5537 = _T_5535 == 1'h0;
  assign _T_5539 = _T_5520 == 1'h0;
  assign _T_5541 = _T_5514 != 1'h1;
  assign _T_5542 = _T_5539 | _T_5541;
  assign _T_5544 = _T_5542 | reset;
  assign _T_5546 = _T_5544 == 1'h0;
  assign _T_5562 = _T_1765 & _T_1949;
  assign _T_5563 = _T_1898 & _T_1941;
  assign _T_5565 = _T_5563 & _T_1952;
  assign _T_5566 = _T_5556 + _T_5562;
  assign _T_5567 = _T_5566[0:0];
  assign _T_5568 = _T_5567 - _T_5565;
  assign _T_5569 = $unsigned(_T_5568);
  assign _T_5570 = _T_5569[0:0];
  assign _T_5572 = _T_5565 == 1'h0;
  assign _T_5575 = _T_5572 | _T_5556;
  assign _T_5577 = _T_5575 | reset;
  assign _T_5579 = _T_5577 == 1'h0;
  assign _T_5581 = _T_5562 == 1'h0;
  assign _T_5583 = _T_5556 != 1'h1;
  assign _T_5584 = _T_5581 | _T_5583;
  assign _T_5586 = _T_5584 | reset;
  assign _T_5588 = _T_5586 == 1'h0;
  assign _T_5604 = _T_1766 & _T_1949;
  assign _T_5605 = _T_1899 & _T_1941;
  assign _T_5607 = _T_5605 & _T_1952;
  assign _T_5608 = _T_5598 + _T_5604;
  assign _T_5609 = _T_5608[0:0];
  assign _T_5610 = _T_5609 - _T_5607;
  assign _T_5611 = $unsigned(_T_5610);
  assign _T_5612 = _T_5611[0:0];
  assign _T_5614 = _T_5607 == 1'h0;
  assign _T_5617 = _T_5614 | _T_5598;
  assign _T_5619 = _T_5617 | reset;
  assign _T_5621 = _T_5619 == 1'h0;
  assign _T_5623 = _T_5604 == 1'h0;
  assign _T_5625 = _T_5598 != 1'h1;
  assign _T_5626 = _T_5623 | _T_5625;
  assign _T_5628 = _T_5626 | reset;
  assign _T_5630 = _T_5628 == 1'h0;
  assign _T_5646 = _T_1767 & _T_1949;
  assign _T_5647 = _T_1900 & _T_1941;
  assign _T_5649 = _T_5647 & _T_1952;
  assign _T_5650 = _T_5640 + _T_5646;
  assign _T_5651 = _T_5650[0:0];
  assign _T_5652 = _T_5651 - _T_5649;
  assign _T_5653 = $unsigned(_T_5652);
  assign _T_5654 = _T_5653[0:0];
  assign _T_5656 = _T_5649 == 1'h0;
  assign _T_5659 = _T_5656 | _T_5640;
  assign _T_5661 = _T_5659 | reset;
  assign _T_5663 = _T_5661 == 1'h0;
  assign _T_5665 = _T_5646 == 1'h0;
  assign _T_5667 = _T_5640 != 1'h1;
  assign _T_5668 = _T_5665 | _T_5667;
  assign _T_5670 = _T_5668 | reset;
  assign _T_5672 = _T_5670 == 1'h0;
  assign _T_5688 = _T_1768 & _T_1949;
  assign _T_5689 = _T_1901 & _T_1941;
  assign _T_5691 = _T_5689 & _T_1952;
  assign _T_5692 = _T_5682 + _T_5688;
  assign _T_5693 = _T_5692[0:0];
  assign _T_5694 = _T_5693 - _T_5691;
  assign _T_5695 = $unsigned(_T_5694);
  assign _T_5696 = _T_5695[0:0];
  assign _T_5698 = _T_5691 == 1'h0;
  assign _T_5701 = _T_5698 | _T_5682;
  assign _T_5703 = _T_5701 | reset;
  assign _T_5705 = _T_5703 == 1'h0;
  assign _T_5707 = _T_5688 == 1'h0;
  assign _T_5709 = _T_5682 != 1'h1;
  assign _T_5710 = _T_5707 | _T_5709;
  assign _T_5712 = _T_5710 | reset;
  assign _T_5714 = _T_5712 == 1'h0;
  assign _T_5730 = _T_1769 & _T_1949;
  assign _T_5731 = _T_1902 & _T_1941;
  assign _T_5733 = _T_5731 & _T_1952;
  assign _T_5734 = _T_5724 + _T_5730;
  assign _T_5735 = _T_5734[0:0];
  assign _T_5736 = _T_5735 - _T_5733;
  assign _T_5737 = $unsigned(_T_5736);
  assign _T_5738 = _T_5737[0:0];
  assign _T_5740 = _T_5733 == 1'h0;
  assign _T_5743 = _T_5740 | _T_5724;
  assign _T_5745 = _T_5743 | reset;
  assign _T_5747 = _T_5745 == 1'h0;
  assign _T_5749 = _T_5730 == 1'h0;
  assign _T_5751 = _T_5724 != 1'h1;
  assign _T_5752 = _T_5749 | _T_5751;
  assign _T_5754 = _T_5752 | reset;
  assign _T_5756 = _T_5754 == 1'h0;
  assign _T_5772 = _T_1770 & _T_1949;
  assign _T_5773 = _T_1903 & _T_1941;
  assign _T_5775 = _T_5773 & _T_1952;
  assign _T_5776 = _T_5766 + _T_5772;
  assign _T_5777 = _T_5776[0:0];
  assign _T_5778 = _T_5777 - _T_5775;
  assign _T_5779 = $unsigned(_T_5778);
  assign _T_5780 = _T_5779[0:0];
  assign _T_5782 = _T_5775 == 1'h0;
  assign _T_5785 = _T_5782 | _T_5766;
  assign _T_5787 = _T_5785 | reset;
  assign _T_5789 = _T_5787 == 1'h0;
  assign _T_5791 = _T_5772 == 1'h0;
  assign _T_5793 = _T_5766 != 1'h1;
  assign _T_5794 = _T_5791 | _T_5793;
  assign _T_5796 = _T_5794 | reset;
  assign _T_5798 = _T_5796 == 1'h0;
  assign _T_5814 = _T_1771 & _T_1949;
  assign _T_5815 = _T_1904 & _T_1941;
  assign _T_5817 = _T_5815 & _T_1952;
  assign _T_5818 = _T_5808 + _T_5814;
  assign _T_5819 = _T_5818[0:0];
  assign _T_5820 = _T_5819 - _T_5817;
  assign _T_5821 = $unsigned(_T_5820);
  assign _T_5822 = _T_5821[0:0];
  assign _T_5824 = _T_5817 == 1'h0;
  assign _T_5827 = _T_5824 | _T_5808;
  assign _T_5829 = _T_5827 | reset;
  assign _T_5831 = _T_5829 == 1'h0;
  assign _T_5833 = _T_5814 == 1'h0;
  assign _T_5835 = _T_5808 != 1'h1;
  assign _T_5836 = _T_5833 | _T_5835;
  assign _T_5838 = _T_5836 | reset;
  assign _T_5840 = _T_5838 == 1'h0;
  assign _T_5856 = _T_1772 & _T_1949;
  assign _T_5857 = _T_1905 & _T_1941;
  assign _T_5859 = _T_5857 & _T_1952;
  assign _T_5860 = _T_5850 + _T_5856;
  assign _T_5861 = _T_5860[0:0];
  assign _T_5862 = _T_5861 - _T_5859;
  assign _T_5863 = $unsigned(_T_5862);
  assign _T_5864 = _T_5863[0:0];
  assign _T_5866 = _T_5859 == 1'h0;
  assign _T_5869 = _T_5866 | _T_5850;
  assign _T_5871 = _T_5869 | reset;
  assign _T_5873 = _T_5871 == 1'h0;
  assign _T_5875 = _T_5856 == 1'h0;
  assign _T_5877 = _T_5850 != 1'h1;
  assign _T_5878 = _T_5875 | _T_5877;
  assign _T_5880 = _T_5878 | reset;
  assign _T_5882 = _T_5880 == 1'h0;
  assign _T_5898 = _T_1773 & _T_1949;
  assign _T_5899 = _T_1906 & _T_1941;
  assign _T_5901 = _T_5899 & _T_1952;
  assign _T_5902 = _T_5892 + _T_5898;
  assign _T_5903 = _T_5902[0:0];
  assign _T_5904 = _T_5903 - _T_5901;
  assign _T_5905 = $unsigned(_T_5904);
  assign _T_5906 = _T_5905[0:0];
  assign _T_5908 = _T_5901 == 1'h0;
  assign _T_5911 = _T_5908 | _T_5892;
  assign _T_5913 = _T_5911 | reset;
  assign _T_5915 = _T_5913 == 1'h0;
  assign _T_5917 = _T_5898 == 1'h0;
  assign _T_5919 = _T_5892 != 1'h1;
  assign _T_5920 = _T_5917 | _T_5919;
  assign _T_5922 = _T_5920 | reset;
  assign _T_5924 = _T_5922 == 1'h0;
  assign _T_5940 = _T_1774 & _T_1949;
  assign _T_5941 = _T_1907 & _T_1941;
  assign _T_5943 = _T_5941 & _T_1952;
  assign _T_5944 = _T_5934 + _T_5940;
  assign _T_5945 = _T_5944[0:0];
  assign _T_5946 = _T_5945 - _T_5943;
  assign _T_5947 = $unsigned(_T_5946);
  assign _T_5948 = _T_5947[0:0];
  assign _T_5950 = _T_5943 == 1'h0;
  assign _T_5953 = _T_5950 | _T_5934;
  assign _T_5955 = _T_5953 | reset;
  assign _T_5957 = _T_5955 == 1'h0;
  assign _T_5959 = _T_5940 == 1'h0;
  assign _T_5961 = _T_5934 != 1'h1;
  assign _T_5962 = _T_5959 | _T_5961;
  assign _T_5964 = _T_5962 | reset;
  assign _T_5966 = _T_5964 == 1'h0;
  assign _T_5982 = _T_1775 & _T_1949;
  assign _T_5983 = _T_1908 & _T_1941;
  assign _T_5985 = _T_5983 & _T_1952;
  assign _T_5986 = _T_5976 + _T_5982;
  assign _T_5987 = _T_5986[0:0];
  assign _T_5988 = _T_5987 - _T_5985;
  assign _T_5989 = $unsigned(_T_5988);
  assign _T_5990 = _T_5989[0:0];
  assign _T_5992 = _T_5985 == 1'h0;
  assign _T_5995 = _T_5992 | _T_5976;
  assign _T_5997 = _T_5995 | reset;
  assign _T_5999 = _T_5997 == 1'h0;
  assign _T_6001 = _T_5982 == 1'h0;
  assign _T_6003 = _T_5976 != 1'h1;
  assign _T_6004 = _T_6001 | _T_6003;
  assign _T_6006 = _T_6004 | reset;
  assign _T_6008 = _T_6006 == 1'h0;
  assign _T_6024 = _T_1776 & _T_1949;
  assign _T_6025 = _T_1909 & _T_1941;
  assign _T_6027 = _T_6025 & _T_1952;
  assign _T_6028 = _T_6018 + _T_6024;
  assign _T_6029 = _T_6028[0:0];
  assign _T_6030 = _T_6029 - _T_6027;
  assign _T_6031 = $unsigned(_T_6030);
  assign _T_6032 = _T_6031[0:0];
  assign _T_6034 = _T_6027 == 1'h0;
  assign _T_6037 = _T_6034 | _T_6018;
  assign _T_6039 = _T_6037 | reset;
  assign _T_6041 = _T_6039 == 1'h0;
  assign _T_6043 = _T_6024 == 1'h0;
  assign _T_6045 = _T_6018 != 1'h1;
  assign _T_6046 = _T_6043 | _T_6045;
  assign _T_6048 = _T_6046 | reset;
  assign _T_6050 = _T_6048 == 1'h0;
  assign _T_6066 = _T_1777 & _T_1949;
  assign _T_6067 = _T_1910 & _T_1941;
  assign _T_6069 = _T_6067 & _T_1952;
  assign _T_6070 = _T_6060 + _T_6066;
  assign _T_6071 = _T_6070[0:0];
  assign _T_6072 = _T_6071 - _T_6069;
  assign _T_6073 = $unsigned(_T_6072);
  assign _T_6074 = _T_6073[0:0];
  assign _T_6076 = _T_6069 == 1'h0;
  assign _T_6079 = _T_6076 | _T_6060;
  assign _T_6081 = _T_6079 | reset;
  assign _T_6083 = _T_6081 == 1'h0;
  assign _T_6085 = _T_6066 == 1'h0;
  assign _T_6087 = _T_6060 != 1'h1;
  assign _T_6088 = _T_6085 | _T_6087;
  assign _T_6090 = _T_6088 | reset;
  assign _T_6092 = _T_6090 == 1'h0;
  assign _T_6108 = _T_1778 & _T_1949;
  assign _T_6109 = _T_1911 & _T_1941;
  assign _T_6111 = _T_6109 & _T_1952;
  assign _T_6112 = _T_6102 + _T_6108;
  assign _T_6113 = _T_6112[0:0];
  assign _T_6114 = _T_6113 - _T_6111;
  assign _T_6115 = $unsigned(_T_6114);
  assign _T_6116 = _T_6115[0:0];
  assign _T_6118 = _T_6111 == 1'h0;
  assign _T_6121 = _T_6118 | _T_6102;
  assign _T_6123 = _T_6121 | reset;
  assign _T_6125 = _T_6123 == 1'h0;
  assign _T_6127 = _T_6108 == 1'h0;
  assign _T_6129 = _T_6102 != 1'h1;
  assign _T_6130 = _T_6127 | _T_6129;
  assign _T_6132 = _T_6130 | reset;
  assign _T_6134 = _T_6132 == 1'h0;
  assign _T_6150 = _T_1779 & _T_1949;
  assign _T_6151 = _T_1912 & _T_1941;
  assign _T_6153 = _T_6151 & _T_1952;
  assign _T_6154 = _T_6144 + _T_6150;
  assign _T_6155 = _T_6154[0:0];
  assign _T_6156 = _T_6155 - _T_6153;
  assign _T_6157 = $unsigned(_T_6156);
  assign _T_6158 = _T_6157[0:0];
  assign _T_6160 = _T_6153 == 1'h0;
  assign _T_6163 = _T_6160 | _T_6144;
  assign _T_6165 = _T_6163 | reset;
  assign _T_6167 = _T_6165 == 1'h0;
  assign _T_6169 = _T_6150 == 1'h0;
  assign _T_6171 = _T_6144 != 1'h1;
  assign _T_6172 = _T_6169 | _T_6171;
  assign _T_6174 = _T_6172 | reset;
  assign _T_6176 = _T_6174 == 1'h0;
  assign _T_6192 = _T_1780 & _T_1949;
  assign _T_6193 = _T_1913 & _T_1941;
  assign _T_6195 = _T_6193 & _T_1952;
  assign _T_6196 = _T_6186 + _T_6192;
  assign _T_6197 = _T_6196[0:0];
  assign _T_6198 = _T_6197 - _T_6195;
  assign _T_6199 = $unsigned(_T_6198);
  assign _T_6200 = _T_6199[0:0];
  assign _T_6202 = _T_6195 == 1'h0;
  assign _T_6205 = _T_6202 | _T_6186;
  assign _T_6207 = _T_6205 | reset;
  assign _T_6209 = _T_6207 == 1'h0;
  assign _T_6211 = _T_6192 == 1'h0;
  assign _T_6213 = _T_6186 != 1'h1;
  assign _T_6214 = _T_6211 | _T_6213;
  assign _T_6216 = _T_6214 | reset;
  assign _T_6218 = _T_6216 == 1'h0;
  assign _T_6234 = _T_1781 & _T_1949;
  assign _T_6235 = _T_1914 & _T_1941;
  assign _T_6237 = _T_6235 & _T_1952;
  assign _T_6238 = _T_6228 + _T_6234;
  assign _T_6239 = _T_6238[0:0];
  assign _T_6240 = _T_6239 - _T_6237;
  assign _T_6241 = $unsigned(_T_6240);
  assign _T_6242 = _T_6241[0:0];
  assign _T_6244 = _T_6237 == 1'h0;
  assign _T_6247 = _T_6244 | _T_6228;
  assign _T_6249 = _T_6247 | reset;
  assign _T_6251 = _T_6249 == 1'h0;
  assign _T_6253 = _T_6234 == 1'h0;
  assign _T_6255 = _T_6228 != 1'h1;
  assign _T_6256 = _T_6253 | _T_6255;
  assign _T_6258 = _T_6256 | reset;
  assign _T_6260 = _T_6258 == 1'h0;
  assign _T_6276 = _T_1782 & _T_1949;
  assign _T_6277 = _T_1915 & _T_1941;
  assign _T_6279 = _T_6277 & _T_1952;
  assign _T_6280 = _T_6270 + _T_6276;
  assign _T_6281 = _T_6280[0:0];
  assign _T_6282 = _T_6281 - _T_6279;
  assign _T_6283 = $unsigned(_T_6282);
  assign _T_6284 = _T_6283[0:0];
  assign _T_6286 = _T_6279 == 1'h0;
  assign _T_6289 = _T_6286 | _T_6270;
  assign _T_6291 = _T_6289 | reset;
  assign _T_6293 = _T_6291 == 1'h0;
  assign _T_6295 = _T_6276 == 1'h0;
  assign _T_6297 = _T_6270 != 1'h1;
  assign _T_6298 = _T_6295 | _T_6297;
  assign _T_6300 = _T_6298 | reset;
  assign _T_6302 = _T_6300 == 1'h0;
  assign _T_6318 = _T_1783 & _T_1949;
  assign _T_6319 = _T_1916 & _T_1941;
  assign _T_6321 = _T_6319 & _T_1952;
  assign _T_6322 = _T_6312 + _T_6318;
  assign _T_6323 = _T_6322[0:0];
  assign _T_6324 = _T_6323 - _T_6321;
  assign _T_6325 = $unsigned(_T_6324);
  assign _T_6326 = _T_6325[0:0];
  assign _T_6328 = _T_6321 == 1'h0;
  assign _T_6331 = _T_6328 | _T_6312;
  assign _T_6333 = _T_6331 | reset;
  assign _T_6335 = _T_6333 == 1'h0;
  assign _T_6337 = _T_6318 == 1'h0;
  assign _T_6339 = _T_6312 != 1'h1;
  assign _T_6340 = _T_6337 | _T_6339;
  assign _T_6342 = _T_6340 | reset;
  assign _T_6344 = _T_6342 == 1'h0;
  assign _T_6360 = _T_1784 & _T_1949;
  assign _T_6361 = _T_1917 & _T_1941;
  assign _T_6363 = _T_6361 & _T_1952;
  assign _T_6364 = _T_6354 + _T_6360;
  assign _T_6365 = _T_6364[0:0];
  assign _T_6366 = _T_6365 - _T_6363;
  assign _T_6367 = $unsigned(_T_6366);
  assign _T_6368 = _T_6367[0:0];
  assign _T_6370 = _T_6363 == 1'h0;
  assign _T_6373 = _T_6370 | _T_6354;
  assign _T_6375 = _T_6373 | reset;
  assign _T_6377 = _T_6375 == 1'h0;
  assign _T_6379 = _T_6360 == 1'h0;
  assign _T_6381 = _T_6354 != 1'h1;
  assign _T_6382 = _T_6379 | _T_6381;
  assign _T_6384 = _T_6382 | reset;
  assign _T_6386 = _T_6384 == 1'h0;
  assign _T_6402 = _T_1785 & _T_1949;
  assign _T_6403 = _T_1918 & _T_1941;
  assign _T_6405 = _T_6403 & _T_1952;
  assign _T_6406 = _T_6396 + _T_6402;
  assign _T_6407 = _T_6406[0:0];
  assign _T_6408 = _T_6407 - _T_6405;
  assign _T_6409 = $unsigned(_T_6408);
  assign _T_6410 = _T_6409[0:0];
  assign _T_6412 = _T_6405 == 1'h0;
  assign _T_6415 = _T_6412 | _T_6396;
  assign _T_6417 = _T_6415 | reset;
  assign _T_6419 = _T_6417 == 1'h0;
  assign _T_6421 = _T_6402 == 1'h0;
  assign _T_6423 = _T_6396 != 1'h1;
  assign _T_6424 = _T_6421 | _T_6423;
  assign _T_6426 = _T_6424 | reset;
  assign _T_6428 = _T_6426 == 1'h0;
  assign _T_6444 = _T_1786 & _T_1949;
  assign _T_6445 = _T_1919 & _T_1941;
  assign _T_6447 = _T_6445 & _T_1952;
  assign _T_6448 = _T_6438 + _T_6444;
  assign _T_6449 = _T_6448[0:0];
  assign _T_6450 = _T_6449 - _T_6447;
  assign _T_6451 = $unsigned(_T_6450);
  assign _T_6452 = _T_6451[0:0];
  assign _T_6454 = _T_6447 == 1'h0;
  assign _T_6457 = _T_6454 | _T_6438;
  assign _T_6459 = _T_6457 | reset;
  assign _T_6461 = _T_6459 == 1'h0;
  assign _T_6463 = _T_6444 == 1'h0;
  assign _T_6465 = _T_6438 != 1'h1;
  assign _T_6466 = _T_6463 | _T_6465;
  assign _T_6468 = _T_6466 | reset;
  assign _T_6470 = _T_6468 == 1'h0;
  assign _T_6486 = _T_1787 & _T_1949;
  assign _T_6487 = _T_1920 & _T_1941;
  assign _T_6489 = _T_6487 & _T_1952;
  assign _T_6490 = _T_6480 + _T_6486;
  assign _T_6491 = _T_6490[0:0];
  assign _T_6492 = _T_6491 - _T_6489;
  assign _T_6493 = $unsigned(_T_6492);
  assign _T_6494 = _T_6493[0:0];
  assign _T_6496 = _T_6489 == 1'h0;
  assign _T_6499 = _T_6496 | _T_6480;
  assign _T_6501 = _T_6499 | reset;
  assign _T_6503 = _T_6501 == 1'h0;
  assign _T_6505 = _T_6486 == 1'h0;
  assign _T_6507 = _T_6480 != 1'h1;
  assign _T_6508 = _T_6505 | _T_6507;
  assign _T_6510 = _T_6508 | reset;
  assign _T_6512 = _T_6510 == 1'h0;
  assign _T_6528 = _T_1788 & _T_1949;
  assign _T_6529 = _T_1921 & _T_1941;
  assign _T_6531 = _T_6529 & _T_1952;
  assign _T_6532 = _T_6522 + _T_6528;
  assign _T_6533 = _T_6532[0:0];
  assign _T_6534 = _T_6533 - _T_6531;
  assign _T_6535 = $unsigned(_T_6534);
  assign _T_6536 = _T_6535[0:0];
  assign _T_6538 = _T_6531 == 1'h0;
  assign _T_6541 = _T_6538 | _T_6522;
  assign _T_6543 = _T_6541 | reset;
  assign _T_6545 = _T_6543 == 1'h0;
  assign _T_6547 = _T_6528 == 1'h0;
  assign _T_6549 = _T_6522 != 1'h1;
  assign _T_6550 = _T_6547 | _T_6549;
  assign _T_6552 = _T_6550 | reset;
  assign _T_6554 = _T_6552 == 1'h0;
  assign _T_6570 = _T_1789 & _T_1949;
  assign _T_6571 = _T_1922 & _T_1941;
  assign _T_6573 = _T_6571 & _T_1952;
  assign _T_6574 = _T_6564 + _T_6570;
  assign _T_6575 = _T_6574[0:0];
  assign _T_6576 = _T_6575 - _T_6573;
  assign _T_6577 = $unsigned(_T_6576);
  assign _T_6578 = _T_6577[0:0];
  assign _T_6580 = _T_6573 == 1'h0;
  assign _T_6583 = _T_6580 | _T_6564;
  assign _T_6585 = _T_6583 | reset;
  assign _T_6587 = _T_6585 == 1'h0;
  assign _T_6589 = _T_6570 == 1'h0;
  assign _T_6591 = _T_6564 != 1'h1;
  assign _T_6592 = _T_6589 | _T_6591;
  assign _T_6594 = _T_6592 | reset;
  assign _T_6596 = _T_6594 == 1'h0;
  assign _T_6612 = _T_1790 & _T_1949;
  assign _T_6613 = _T_1923 & _T_1941;
  assign _T_6615 = _T_6613 & _T_1952;
  assign _T_6616 = _T_6606 + _T_6612;
  assign _T_6617 = _T_6616[0:0];
  assign _T_6618 = _T_6617 - _T_6615;
  assign _T_6619 = $unsigned(_T_6618);
  assign _T_6620 = _T_6619[0:0];
  assign _T_6622 = _T_6615 == 1'h0;
  assign _T_6625 = _T_6622 | _T_6606;
  assign _T_6627 = _T_6625 | reset;
  assign _T_6629 = _T_6627 == 1'h0;
  assign _T_6631 = _T_6612 == 1'h0;
  assign _T_6633 = _T_6606 != 1'h1;
  assign _T_6634 = _T_6631 | _T_6633;
  assign _T_6636 = _T_6634 | reset;
  assign _T_6638 = _T_6636 == 1'h0;
  assign _T_6654 = _T_1791 & _T_1949;
  assign _T_6655 = _T_1924 & _T_1941;
  assign _T_6657 = _T_6655 & _T_1952;
  assign _T_6658 = _T_6648 + _T_6654;
  assign _T_6659 = _T_6658[0:0];
  assign _T_6660 = _T_6659 - _T_6657;
  assign _T_6661 = $unsigned(_T_6660);
  assign _T_6662 = _T_6661[0:0];
  assign _T_6664 = _T_6657 == 1'h0;
  assign _T_6667 = _T_6664 | _T_6648;
  assign _T_6669 = _T_6667 | reset;
  assign _T_6671 = _T_6669 == 1'h0;
  assign _T_6673 = _T_6654 == 1'h0;
  assign _T_6675 = _T_6648 != 1'h1;
  assign _T_6676 = _T_6673 | _T_6675;
  assign _T_6678 = _T_6676 | reset;
  assign _T_6680 = _T_6678 == 1'h0;
  assign _T_6696 = _T_1792 & _T_1949;
  assign _T_6697 = _T_1925 & _T_1941;
  assign _T_6699 = _T_6697 & _T_1952;
  assign _T_6700 = _T_6690 + _T_6696;
  assign _T_6701 = _T_6700[0:0];
  assign _T_6702 = _T_6701 - _T_6699;
  assign _T_6703 = $unsigned(_T_6702);
  assign _T_6704 = _T_6703[0:0];
  assign _T_6706 = _T_6699 == 1'h0;
  assign _T_6709 = _T_6706 | _T_6690;
  assign _T_6711 = _T_6709 | reset;
  assign _T_6713 = _T_6711 == 1'h0;
  assign _T_6715 = _T_6696 == 1'h0;
  assign _T_6717 = _T_6690 != 1'h1;
  assign _T_6718 = _T_6715 | _T_6717;
  assign _T_6720 = _T_6718 | reset;
  assign _T_6722 = _T_6720 == 1'h0;
  assign _T_6738 = _T_1793 & _T_1949;
  assign _T_6739 = _T_1926 & _T_1941;
  assign _T_6741 = _T_6739 & _T_1952;
  assign _T_6742 = _T_6732 + _T_6738;
  assign _T_6743 = _T_6742[0:0];
  assign _T_6744 = _T_6743 - _T_6741;
  assign _T_6745 = $unsigned(_T_6744);
  assign _T_6746 = _T_6745[0:0];
  assign _T_6748 = _T_6741 == 1'h0;
  assign _T_6751 = _T_6748 | _T_6732;
  assign _T_6753 = _T_6751 | reset;
  assign _T_6755 = _T_6753 == 1'h0;
  assign _T_6757 = _T_6738 == 1'h0;
  assign _T_6759 = _T_6732 != 1'h1;
  assign _T_6760 = _T_6757 | _T_6759;
  assign _T_6762 = _T_6760 | reset;
  assign _T_6764 = _T_6762 == 1'h0;
  assign _T_6780 = _T_1794 & _T_1949;
  assign _T_6781 = _T_1927 & _T_1941;
  assign _T_6783 = _T_6781 & _T_1952;
  assign _T_6784 = _T_6774 + _T_6780;
  assign _T_6785 = _T_6784[0:0];
  assign _T_6786 = _T_6785 - _T_6783;
  assign _T_6787 = $unsigned(_T_6786);
  assign _T_6788 = _T_6787[0:0];
  assign _T_6790 = _T_6783 == 1'h0;
  assign _T_6793 = _T_6790 | _T_6774;
  assign _T_6795 = _T_6793 | reset;
  assign _T_6797 = _T_6795 == 1'h0;
  assign _T_6799 = _T_6780 == 1'h0;
  assign _T_6801 = _T_6774 != 1'h1;
  assign _T_6802 = _T_6799 | _T_6801;
  assign _T_6804 = _T_6802 | reset;
  assign _T_6806 = _T_6804 == 1'h0;
  assign _T_6822 = _T_1795 & _T_1949;
  assign _T_6823 = _T_1928 & _T_1941;
  assign _T_6825 = _T_6823 & _T_1952;
  assign _T_6826 = _T_6816 + _T_6822;
  assign _T_6827 = _T_6826[0:0];
  assign _T_6828 = _T_6827 - _T_6825;
  assign _T_6829 = $unsigned(_T_6828);
  assign _T_6830 = _T_6829[0:0];
  assign _T_6832 = _T_6825 == 1'h0;
  assign _T_6835 = _T_6832 | _T_6816;
  assign _T_6837 = _T_6835 | reset;
  assign _T_6839 = _T_6837 == 1'h0;
  assign _T_6841 = _T_6822 == 1'h0;
  assign _T_6843 = _T_6816 != 1'h1;
  assign _T_6844 = _T_6841 | _T_6843;
  assign _T_6846 = _T_6844 | reset;
  assign _T_6848 = _T_6846 == 1'h0;
  assign _T_6864 = _T_1796 & _T_1949;
  assign _T_6865 = _T_1929 & _T_1941;
  assign _T_6867 = _T_6865 & _T_1952;
  assign _T_6868 = _T_6858 + _T_6864;
  assign _T_6869 = _T_6868[0:0];
  assign _T_6870 = _T_6869 - _T_6867;
  assign _T_6871 = $unsigned(_T_6870);
  assign _T_6872 = _T_6871[0:0];
  assign _T_6874 = _T_6867 == 1'h0;
  assign _T_6877 = _T_6874 | _T_6858;
  assign _T_6879 = _T_6877 | reset;
  assign _T_6881 = _T_6879 == 1'h0;
  assign _T_6883 = _T_6864 == 1'h0;
  assign _T_6885 = _T_6858 != 1'h1;
  assign _T_6886 = _T_6883 | _T_6885;
  assign _T_6888 = _T_6886 | reset;
  assign _T_6890 = _T_6888 == 1'h0;
  assign _T_6906 = _T_1797 & _T_1949;
  assign _T_6907 = _T_1930 & _T_1941;
  assign _T_6909 = _T_6907 & _T_1952;
  assign _T_6910 = _T_6900 + _T_6906;
  assign _T_6911 = _T_6910[0:0];
  assign _T_6912 = _T_6911 - _T_6909;
  assign _T_6913 = $unsigned(_T_6912);
  assign _T_6914 = _T_6913[0:0];
  assign _T_6916 = _T_6909 == 1'h0;
  assign _T_6919 = _T_6916 | _T_6900;
  assign _T_6921 = _T_6919 | reset;
  assign _T_6923 = _T_6921 == 1'h0;
  assign _T_6925 = _T_6906 == 1'h0;
  assign _T_6927 = _T_6900 != 1'h1;
  assign _T_6928 = _T_6925 | _T_6927;
  assign _T_6930 = _T_6928 | reset;
  assign _T_6932 = _T_6930 == 1'h0;
  assign _T_6948 = _T_1798 & _T_1949;
  assign _T_6949 = _T_1931 & _T_1941;
  assign _T_6951 = _T_6949 & _T_1952;
  assign _T_6952 = _T_6942 + _T_6948;
  assign _T_6953 = _T_6952[0:0];
  assign _T_6954 = _T_6953 - _T_6951;
  assign _T_6955 = $unsigned(_T_6954);
  assign _T_6956 = _T_6955[0:0];
  assign _T_6958 = _T_6951 == 1'h0;
  assign _T_6961 = _T_6958 | _T_6942;
  assign _T_6963 = _T_6961 | reset;
  assign _T_6965 = _T_6963 == 1'h0;
  assign _T_6967 = _T_6948 == 1'h0;
  assign _T_6969 = _T_6942 != 1'h1;
  assign _T_6970 = _T_6967 | _T_6969;
  assign _T_6972 = _T_6970 | reset;
  assign _T_6974 = _T_6972 == 1'h0;
  assign _T_6990 = _T_1799 & _T_1949;
  assign _T_6991 = _T_1932 & _T_1941;
  assign _T_6993 = _T_6991 & _T_1952;
  assign _T_6994 = _T_6984 + _T_6990;
  assign _T_6995 = _T_6994[0:0];
  assign _T_6996 = _T_6995 - _T_6993;
  assign _T_6997 = $unsigned(_T_6996);
  assign _T_6998 = _T_6997[0:0];
  assign _T_7000 = _T_6993 == 1'h0;
  assign _T_7003 = _T_7000 | _T_6984;
  assign _T_7005 = _T_7003 | reset;
  assign _T_7007 = _T_7005 == 1'h0;
  assign _T_7009 = _T_6990 == 1'h0;
  assign _T_7011 = _T_6984 != 1'h1;
  assign _T_7012 = _T_7009 | _T_7011;
  assign _T_7014 = _T_7012 | reset;
  assign _T_7016 = _T_7014 == 1'h0;
  assign _T_7032 = _T_1800 & _T_1949;
  assign _T_7033 = _T_1933 & _T_1941;
  assign _T_7035 = _T_7033 & _T_1952;
  assign _T_7036 = _T_7026 + _T_7032;
  assign _T_7037 = _T_7036[0:0];
  assign _T_7038 = _T_7037 - _T_7035;
  assign _T_7039 = $unsigned(_T_7038);
  assign _T_7040 = _T_7039[0:0];
  assign _T_7042 = _T_7035 == 1'h0;
  assign _T_7045 = _T_7042 | _T_7026;
  assign _T_7047 = _T_7045 | reset;
  assign _T_7049 = _T_7047 == 1'h0;
  assign _T_7051 = _T_7032 == 1'h0;
  assign _T_7053 = _T_7026 != 1'h1;
  assign _T_7054 = _T_7051 | _T_7053;
  assign _T_7056 = _T_7054 | reset;
  assign _T_7058 = _T_7056 == 1'h0;
  assign _T_7074 = _T_1801 & _T_1949;
  assign _T_7075 = _T_1934 & _T_1941;
  assign _T_7077 = _T_7075 & _T_1952;
  assign _T_7078 = _T_7068 + _T_7074;
  assign _T_7079 = _T_7078[0:0];
  assign _T_7080 = _T_7079 - _T_7077;
  assign _T_7081 = $unsigned(_T_7080);
  assign _T_7082 = _T_7081[0:0];
  assign _T_7084 = _T_7077 == 1'h0;
  assign _T_7087 = _T_7084 | _T_7068;
  assign _T_7089 = _T_7087 | reset;
  assign _T_7091 = _T_7089 == 1'h0;
  assign _T_7093 = _T_7074 == 1'h0;
  assign _T_7095 = _T_7068 != 1'h1;
  assign _T_7096 = _T_7093 | _T_7095;
  assign _T_7098 = _T_7096 | reset;
  assign _T_7100 = _T_7098 == 1'h0;
  assign _T_7116 = _T_1802 & _T_1949;
  assign _T_7117 = _T_1935 & _T_1941;
  assign _T_7119 = _T_7117 & _T_1952;
  assign _T_7120 = _T_7110 + _T_7116;
  assign _T_7121 = _T_7120[0:0];
  assign _T_7122 = _T_7121 - _T_7119;
  assign _T_7123 = $unsigned(_T_7122);
  assign _T_7124 = _T_7123[0:0];
  assign _T_7126 = _T_7119 == 1'h0;
  assign _T_7129 = _T_7126 | _T_7110;
  assign _T_7131 = _T_7129 | reset;
  assign _T_7133 = _T_7131 == 1'h0;
  assign _T_7135 = _T_7116 == 1'h0;
  assign _T_7137 = _T_7110 != 1'h1;
  assign _T_7138 = _T_7135 | _T_7137;
  assign _T_7140 = _T_7138 | reset;
  assign _T_7142 = _T_7140 == 1'h0;
  assign _T_7158 = _T_1803 & _T_1949;
  assign _T_7159 = _T_1936 & _T_1941;
  assign _T_7161 = _T_7159 & _T_1952;
  assign _T_7162 = _T_7152 + _T_7158;
  assign _T_7163 = _T_7162[0:0];
  assign _T_7164 = _T_7163 - _T_7161;
  assign _T_7165 = $unsigned(_T_7164);
  assign _T_7166 = _T_7165[0:0];
  assign _T_7168 = _T_7161 == 1'h0;
  assign _T_7171 = _T_7168 | _T_7152;
  assign _T_7173 = _T_7171 | reset;
  assign _T_7175 = _T_7173 == 1'h0;
  assign _T_7177 = _T_7158 == 1'h0;
  assign _T_7179 = _T_7152 != 1'h1;
  assign _T_7180 = _T_7177 | _T_7179;
  assign _T_7182 = _T_7180 | reset;
  assign _T_7184 = _T_7182 == 1'h0;
  assign _T_7200 = _T_1804 & _T_1949;
  assign _T_7201 = _T_1937 & _T_1941;
  assign _T_7203 = _T_7201 & _T_1952;
  assign _T_7204 = _T_7194 + _T_7200;
  assign _T_7205 = _T_7204[0:0];
  assign _T_7206 = _T_7205 - _T_7203;
  assign _T_7207 = $unsigned(_T_7206);
  assign _T_7208 = _T_7207[0:0];
  assign _T_7210 = _T_7203 == 1'h0;
  assign _T_7213 = _T_7210 | _T_7194;
  assign _T_7215 = _T_7213 | reset;
  assign _T_7217 = _T_7215 == 1'h0;
  assign _T_7219 = _T_7200 == 1'h0;
  assign _T_7221 = _T_7194 != 1'h1;
  assign _T_7222 = _T_7219 | _T_7221;
  assign _T_7224 = _T_7222 | reset;
  assign _T_7226 = _T_7224 == 1'h0;
  assign _T_7242 = _T_1805 & _T_1949;
  assign _T_7243 = _T_1938 & _T_1941;
  assign _T_7245 = _T_7243 & _T_1952;
  assign _T_7246 = _T_7236 + _T_7242;
  assign _T_7247 = _T_7246[0:0];
  assign _T_7248 = _T_7247 - _T_7245;
  assign _T_7249 = $unsigned(_T_7248);
  assign _T_7250 = _T_7249[0:0];
  assign _T_7252 = _T_7245 == 1'h0;
  assign _T_7255 = _T_7252 | _T_7236;
  assign _T_7257 = _T_7255 | reset;
  assign _T_7259 = _T_7257 == 1'h0;
  assign _T_7261 = _T_7242 == 1'h0;
  assign _T_7263 = _T_7236 != 1'h1;
  assign _T_7264 = _T_7261 | _T_7263;
  assign _T_7266 = _T_7264 | reset;
  assign _T_7268 = _T_7266 == 1'h0;
  assign _T_7284 = _T_1806 & _T_1949;
  assign _T_7285 = _T_1939 & _T_1941;
  assign _T_7287 = _T_7285 & _T_1952;
  assign _T_7288 = _T_7278 + _T_7284;
  assign _T_7289 = _T_7288[0:0];
  assign _T_7290 = _T_7289 - _T_7287;
  assign _T_7291 = $unsigned(_T_7290);
  assign _T_7292 = _T_7291[0:0];
  assign _T_7294 = _T_7287 == 1'h0;
  assign _T_7297 = _T_7294 | _T_7278;
  assign _T_7299 = _T_7297 | reset;
  assign _T_7301 = _T_7299 == 1'h0;
  assign _T_7303 = _T_7284 == 1'h0;
  assign _T_7305 = _T_7278 != 1'h1;
  assign _T_7306 = _T_7303 | _T_7305;
  assign _T_7308 = _T_7306 | reset;
  assign _T_7310 = _T_7308 == 1'h0;
  assign auto_in_a_ready = _T_31_a_ready;
  assign auto_in_d_valid = _T_31_d_valid;
  assign auto_in_d_bits_opcode = _T_31_d_bits_opcode;
  assign auto_in_d_bits_size = _T_31_d_bits_size;
  assign auto_in_d_bits_source = _T_31_d_bits_source;
  assign auto_in_d_bits_data = _T_31_d_bits_data;
  assign auto_in_d_bits_error = _T_31_d_bits_error;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_a_ready = _T_1622;
  assign _T_31_a_valid = auto_in_a_valid;
  assign _T_31_a_bits_opcode = auto_in_a_bits_opcode;
  assign _T_31_a_bits_size = auto_in_a_bits_size;
  assign _T_31_a_bits_source = auto_in_a_bits_source;
  assign _T_31_a_bits_address = auto_in_a_bits_address;
  assign _T_31_a_bits_mask = auto_in_a_bits_mask;
  assign _T_31_a_bits_data = auto_in_a_bits_data;
  assign _T_31_d_ready = auto_in_d_ready;
  assign _T_31_d_valid = _T_1648;
  assign _T_31_d_bits_opcode = _T_1674_opcode;
  assign _T_31_d_bits_size = _T_1674_size;
  assign _T_31_d_bits_source = _T_1674_source;
  assign _T_31_d_bits_data = _T_89_r_bits_data;
  assign _T_31_d_bits_error = _T_1674_error;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_1592;
  assign _T_89_aw_bits_id = _T_1585_bits_id;
  assign _T_89_aw_bits_addr = _T_1585_bits_addr;
  assign _T_89_aw_bits_len = _T_1585_bits_len;
  assign _T_89_aw_bits_size = _T_1585_bits_size;
  assign _T_89_aw_bits_burst = _T_1585_bits_burst;
  assign _T_89_aw_bits_lock = _T_1585_bits_lock;
  assign _T_89_aw_bits_cache = _T_1585_bits_cache;
  assign _T_89_aw_bits_prot = _T_1585_bits_prot;
  assign _T_89_aw_bits_qos = _T_1585_bits_qos;
  assign _T_89_aw_bits_user = _T_1585_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_1577_valid;
  assign _T_89_w_bits_data = _T_1577_bits_data;
  assign _T_89_w_bits_strb = _T_1577_bits_strb;
  assign _T_89_w_bits_last = _T_1577_bits_last;
  assign _T_89_b_ready = _T_1647;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_1591;
  assign _T_89_ar_bits_id = _T_1585_bits_id;
  assign _T_89_ar_bits_addr = _T_1585_bits_addr;
  assign _T_89_ar_bits_len = _T_1585_bits_len;
  assign _T_89_ar_bits_size = _T_1585_bits_size;
  assign _T_89_ar_bits_burst = _T_1585_bits_burst;
  assign _T_89_ar_bits_lock = _T_1585_bits_lock;
  assign _T_89_ar_bits_cache = _T_1585_bits_cache;
  assign _T_89_ar_bits_prot = _T_1585_bits_prot;
  assign _T_89_ar_bits_qos = _T_1585_bits_qos;
  assign _T_89_ar_bits_user = _T_1585_bits_user;
  assign _T_89_r_ready = _T_31_d_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign _T_206_0 = _T_991_0;
  assign _T_206_1 = _T_991_1;
  assign _T_206_2 = _T_991_2;
  assign _T_206_3 = _T_991_3;
  assign _T_206_4 = _T_991_4;
  assign _T_206_5 = _T_991_5;
  assign _T_206_6 = _T_991_6;
  assign _T_206_7 = _T_991_7;
  assign _T_206_8 = _T_991_8;
  assign _T_206_9 = _T_991_9;
  assign _T_206_10 = _T_991_10;
  assign _T_206_11 = _T_991_11;
  assign _T_206_12 = _T_991_12;
  assign _T_206_13 = _T_991_13;
  assign _T_206_14 = _T_991_14;
  assign _T_206_15 = _T_991_15;
  assign _T_206_16 = _T_991_16;
  assign _T_206_17 = _T_991_17;
  assign _T_206_18 = _T_991_18;
  assign _T_206_19 = _T_991_19;
  assign _T_206_20 = _T_991_20;
  assign _T_206_21 = _T_991_21;
  assign _T_206_22 = _T_991_22;
  assign _T_206_23 = _T_991_23;
  assign _T_206_24 = _T_991_24;
  assign _T_206_25 = _T_991_25;
  assign _T_206_26 = _T_991_26;
  assign _T_206_27 = _T_991_27;
  assign _T_206_28 = _T_991_28;
  assign _T_206_29 = _T_991_29;
  assign _T_206_30 = _T_991_30;
  assign _T_206_31 = _T_991_31;
  assign _T_206_32 = _T_991_32;
  assign _T_206_33 = _T_991_33;
  assign _T_206_34 = _T_991_34;
  assign _T_206_35 = _T_991_35;
  assign _T_206_36 = _T_991_36;
  assign _T_206_37 = _T_991_37;
  assign _T_206_38 = _T_991_38;
  assign _T_206_39 = _T_991_39;
  assign _T_206_40 = _T_991_40;
  assign _T_206_41 = _T_991_41;
  assign _T_206_42 = _T_991_42;
  assign _T_206_43 = _T_991_43;
  assign _T_206_44 = _T_991_44;
  assign _T_206_45 = _T_991_45;
  assign _T_206_46 = _T_991_46;
  assign _T_206_47 = _T_991_47;
  assign _T_206_48 = _T_991_48;
  assign _T_206_49 = _T_991_49;
  assign _T_206_50 = _T_991_50;
  assign _T_206_51 = _T_991_51;
  assign _T_206_52 = _T_991_52;
  assign _T_206_53 = _T_991_53;
  assign _T_206_54 = _T_991_54;
  assign _T_206_55 = _T_991_55;
  assign _T_206_56 = _T_991_56;
  assign _T_206_57 = _T_991_57;
  assign _T_206_58 = _T_991_58;
  assign _T_206_59 = _T_991_59;
  assign _T_206_60 = _T_991_60;
  assign _T_206_61 = _T_991_61;
  assign _T_206_62 = _T_991_62;
  assign _T_206_63 = _T_991_63;
  assign _T_206_64 = _T_991_64;
  assign _T_206_65 = _T_991_65;
  assign _T_206_66 = _T_991_66;
  assign _T_206_67 = _T_991_67;
  assign _T_206_68 = _T_991_68;
  assign _T_206_69 = _T_991_69;
  assign _T_206_70 = _T_991_70;
  assign _T_206_71 = _T_991_71;
  assign _T_206_72 = _T_991_72;
  assign _T_206_73 = _T_991_73;
  assign _T_206_74 = _T_991_74;
  assign _T_206_75 = _T_991_75;
  assign _T_206_76 = _T_991_76;
  assign _T_206_77 = _T_991_77;
  assign _T_206_78 = _T_991_78;
  assign _T_206_79 = _T_991_79;
  assign _T_206_80 = _T_991_80;
  assign _T_206_81 = _T_991_81;
  assign _T_206_82 = _T_991_82;
  assign _T_206_83 = _T_991_83;
  assign _T_206_84 = _T_991_84;
  assign _T_206_85 = _T_991_85;
  assign _T_206_86 = _T_991_86;
  assign _T_206_87 = _T_991_87;
  assign _T_206_88 = _T_991_88;
  assign _T_206_89 = _T_991_89;
  assign _T_206_90 = _T_991_90;
  assign _T_206_91 = _T_991_91;
  assign _T_206_92 = _T_991_92;
  assign _T_206_93 = _T_991_93;
  assign _T_206_94 = _T_991_94;
  assign _T_206_95 = _T_991_95;
  assign _T_206_96 = _T_991_96;
  assign _T_206_97 = _T_991_97;
  assign _T_206_98 = _T_991_98;
  assign _T_206_99 = _T_991_99;
  assign _T_206_100 = _T_991_100;
  assign _T_206_101 = _T_991_101;
  assign _T_206_102 = _T_991_102;
  assign _T_206_103 = _T_991_103;
  assign _T_206_104 = _T_991_104;
  assign _T_206_105 = _T_991_105;
  assign _T_206_106 = _T_991_106;
  assign _T_206_107 = _T_991_107;
  assign _T_206_108 = _T_991_108;
  assign _T_206_109 = _T_991_109;
  assign _T_206_110 = _T_991_110;
  assign _T_206_111 = _T_991_111;
  assign _T_206_112 = _T_991_112;
  assign _T_206_113 = _T_991_113;
  assign _T_206_114 = _T_991_114;
  assign _T_206_115 = _T_991_115;
  assign _T_206_116 = _T_991_116;
  assign _T_206_117 = _T_991_117;
  assign _T_206_118 = _T_991_118;
  assign _T_206_119 = _T_991_119;
  assign _T_206_120 = _T_991_120;
  assign _T_206_121 = _T_991_121;
  assign _T_206_122 = _T_991_122;
  assign _T_206_123 = _T_991_123;
  assign _T_206_124 = _T_991_124;
  assign _T_206_125 = _T_991_125;
  assign _T_206_126 = _T_991_126;
  assign _T_206_127 = _T_991_127;
  assign _T_991_0 = _T_1944;
  assign _T_991_1 = _T_1986;
  assign _T_991_2 = _T_2028;
  assign _T_991_3 = _T_2070;
  assign _T_991_4 = _T_2112;
  assign _T_991_5 = _T_2154;
  assign _T_991_6 = _T_2196;
  assign _T_991_7 = _T_2238;
  assign _T_991_8 = _T_2280;
  assign _T_991_9 = _T_2322;
  assign _T_991_10 = _T_2364;
  assign _T_991_11 = _T_2406;
  assign _T_991_12 = _T_2448;
  assign _T_991_13 = _T_2490;
  assign _T_991_14 = _T_2532;
  assign _T_991_15 = _T_2574;
  assign _T_991_16 = _T_2616;
  assign _T_991_17 = _T_2658;
  assign _T_991_18 = _T_2700;
  assign _T_991_19 = _T_2742;
  assign _T_991_20 = _T_2784;
  assign _T_991_21 = _T_2826;
  assign _T_991_22 = _T_2868;
  assign _T_991_23 = _T_2910;
  assign _T_991_24 = _T_2952;
  assign _T_991_25 = _T_2994;
  assign _T_991_26 = _T_3036;
  assign _T_991_27 = _T_3078;
  assign _T_991_28 = _T_3120;
  assign _T_991_29 = _T_3162;
  assign _T_991_30 = _T_3204;
  assign _T_991_31 = _T_3246;
  assign _T_991_32 = _T_3288;
  assign _T_991_33 = _T_3330;
  assign _T_991_34 = _T_3372;
  assign _T_991_35 = _T_3414;
  assign _T_991_36 = _T_3456;
  assign _T_991_37 = _T_3498;
  assign _T_991_38 = _T_3540;
  assign _T_991_39 = _T_3582;
  assign _T_991_40 = _T_3624;
  assign _T_991_41 = _T_3666;
  assign _T_991_42 = _T_3708;
  assign _T_991_43 = _T_3750;
  assign _T_991_44 = _T_3792;
  assign _T_991_45 = _T_3834;
  assign _T_991_46 = _T_3876;
  assign _T_991_47 = _T_3918;
  assign _T_991_48 = _T_3960;
  assign _T_991_49 = _T_4002;
  assign _T_991_50 = _T_4044;
  assign _T_991_51 = _T_4086;
  assign _T_991_52 = _T_4128;
  assign _T_991_53 = _T_4170;
  assign _T_991_54 = _T_4212;
  assign _T_991_55 = _T_4254;
  assign _T_991_56 = _T_4296;
  assign _T_991_57 = _T_4338;
  assign _T_991_58 = _T_4380;
  assign _T_991_59 = _T_4422;
  assign _T_991_60 = _T_4464;
  assign _T_991_61 = _T_4506;
  assign _T_991_62 = _T_4548;
  assign _T_991_63 = _T_4590;
  assign _T_991_64 = _T_4632;
  assign _T_991_65 = _T_4674;
  assign _T_991_66 = _T_4716;
  assign _T_991_67 = _T_4758;
  assign _T_991_68 = _T_4800;
  assign _T_991_69 = _T_4842;
  assign _T_991_70 = _T_4884;
  assign _T_991_71 = _T_4926;
  assign _T_991_72 = _T_4968;
  assign _T_991_73 = _T_5010;
  assign _T_991_74 = _T_5052;
  assign _T_991_75 = _T_5094;
  assign _T_991_76 = _T_5136;
  assign _T_991_77 = _T_5178;
  assign _T_991_78 = _T_5220;
  assign _T_991_79 = _T_5262;
  assign _T_991_80 = _T_5304;
  assign _T_991_81 = _T_5346;
  assign _T_991_82 = _T_5388;
  assign _T_991_83 = _T_5430;
  assign _T_991_84 = _T_5472;
  assign _T_991_85 = _T_5514;
  assign _T_991_86 = _T_5556;
  assign _T_991_87 = _T_5598;
  assign _T_991_88 = _T_5640;
  assign _T_991_89 = _T_5682;
  assign _T_991_90 = _T_5724;
  assign _T_991_91 = _T_5766;
  assign _T_991_92 = _T_5808;
  assign _T_991_93 = _T_5850;
  assign _T_991_94 = _T_5892;
  assign _T_991_95 = _T_5934;
  assign _T_991_96 = _T_5976;
  assign _T_991_97 = _T_6018;
  assign _T_991_98 = _T_6060;
  assign _T_991_99 = _T_6102;
  assign _T_991_100 = _T_6144;
  assign _T_991_101 = _T_6186;
  assign _T_991_102 = _T_6228;
  assign _T_991_103 = _T_6270;
  assign _T_991_104 = _T_6312;
  assign _T_991_105 = _T_6354;
  assign _T_991_106 = _T_6396;
  assign _T_991_107 = _T_6438;
  assign _T_991_108 = _T_6480;
  assign _T_991_109 = _T_6522;
  assign _T_991_110 = _T_6564;
  assign _T_991_111 = _T_6606;
  assign _T_991_112 = _T_6648;
  assign _T_991_113 = _T_6690;
  assign _T_991_114 = _T_6732;
  assign _T_991_115 = _T_6774;
  assign _T_991_116 = _T_6816;
  assign _T_991_117 = _T_6858;
  assign _T_991_118 = _T_6900;
  assign _T_991_119 = _T_6942;
  assign _T_991_120 = _T_6984;
  assign _T_991_121 = _T_7026;
  assign _T_991_122 = _T_7068;
  assign _T_991_123 = _T_7110;
  assign _T_991_124 = _T_7152;
  assign _T_991_125 = _T_7194;
  assign _T_991_126 = _T_7236;
  assign _T_991_127 = _T_7278;
  assign _T_1565_ready = Queue_1_io_enq_ready;
  assign _T_1565_valid = _T_1631;
  assign _T_1565_bits_id = _GEN_0;
  assign _T_1565_bits_addr = _T_31_a_bits_address;
  assign _T_1565_bits_len = _T_1607;
  assign _T_1565_bits_size = _T_1609;
  assign _T_1565_bits_user = {{1'd0}, _T_1555};
  assign _T_1565_bits_wen = _T_1510;
  assign _T_1569_ready = Queue_io_enq_ready;
  assign _T_1569_valid = _T_1637;
  assign _T_1569_bits_data = _T_31_a_bits_data;
  assign _T_1569_bits_strb = _T_31_a_bits_mask;
  assign _T_1569_bits_last = _T_1536;
  assign Queue_io_enq_valid = _T_1569_valid;
  assign Queue_io_enq_bits_data = _T_1569_bits_data;
  assign Queue_io_enq_bits_strb = _T_1569_bits_strb;
  assign Queue_io_enq_bits_last = _T_1569_bits_last;
  assign Queue_io_deq_ready = _T_1577_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_1577_ready = _T_89_w_ready;
  assign _T_1577_valid = Queue_io_deq_valid;
  assign _T_1577_bits_data = Queue_io_deq_bits_data;
  assign _T_1577_bits_strb = Queue_io_deq_bits_strb;
  assign _T_1577_bits_last = Queue_io_deq_bits_last;
  assign Queue_1_io_enq_valid = _T_1565_valid;
  assign Queue_1_io_enq_bits_id = _T_1565_bits_id;
  assign Queue_1_io_enq_bits_addr = _T_1565_bits_addr;
  assign Queue_1_io_enq_bits_len = _T_1565_bits_len;
  assign Queue_1_io_enq_bits_size = _T_1565_bits_size;
  assign Queue_1_io_enq_bits_user = _T_1565_bits_user;
  assign Queue_1_io_enq_bits_wen = _T_1565_bits_wen;
  assign Queue_1_io_deq_ready = _T_1585_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_1585_ready = _T_1593;
  assign _T_1585_valid = Queue_1_io_deq_valid;
  assign _T_1585_bits_id = Queue_1_io_deq_bits_id;
  assign _T_1585_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_1585_bits_len = Queue_1_io_deq_bits_len;
  assign _T_1585_bits_size = Queue_1_io_deq_bits_size;
  assign _T_1585_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_1585_bits_lock = Queue_1_io_deq_bits_lock;
  assign _T_1585_bits_cache = Queue_1_io_deq_bits_cache;
  assign _T_1585_bits_prot = Queue_1_io_deq_bits_prot;
  assign _T_1585_bits_qos = Queue_1_io_deq_bits_qos;
  assign _T_1585_bits_user = Queue_1_io_deq_bits_user;
  assign _T_1585_bits_wen = Queue_1_io_deq_bits_wen;
  assign _GEN_0 = _GEN_130;
  assign _GEN_1 = _GEN_257;
  assign _T_1664_size = _T_1557;
  assign _T_1664_source = _T_1556;
  assign _T_1664_error = _T_1659;
  assign _T_1669_size = _T_1559;
  assign _T_1669_source = _T_1558;
  assign _T_1669_error = _T_1652;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1525 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1597 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_1640 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_1655 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_1944 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_1986 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_2028 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_2070 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_2112 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_2154 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_2196 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_2238 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_2280 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_2322 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_2364 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_2406 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_2448 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_2490 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_2532 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_2574 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_2616 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_2658 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_2700 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_2742 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_2784 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_2826 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_2868 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_2910 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_2952 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_2994 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_3036 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_3078 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_3120 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_3162 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_3204 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_3246 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_3288 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_3330 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_3372 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_3414 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_3456 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_3498 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_3540 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_3582 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_3624 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_3666 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_3708 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_3750 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_3792 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_3834 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_3876 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_3918 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_3960 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_4002 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_4044 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_4086 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_4128 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_4170 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_4212 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_4254 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_4296 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_4338 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_4380 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_4422 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_4464 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_4506 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_4548 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_4590 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_4632 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_4674 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_4716 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_4758 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_4800 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_4842 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_4884 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_4926 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_4968 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_5010 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_5052 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_5094 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_5136 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_5178 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_5220 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_5262 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_5304 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_5346 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_5388 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_5430 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_5472 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_5514 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_5556 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_5598 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_5640 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_5682 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_5724 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_5766 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_5808 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_5850 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_5892 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_5934 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_5976 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_6018 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_6060 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_6102 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_6144 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_6186 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_6228 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_6270 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_6312 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_6354 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_6396 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_6438 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_6480 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_6522 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_6564 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_6606 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_6648 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_6690 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_6732 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_6774 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_6816 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_6858 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_6900 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_6942 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_6984 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_7026 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_7068 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_7110 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_7152 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_7194 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_7236 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_7278 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1525 <= 3'h0;
    end else begin
      if (_T_1511) begin
        if (_T_1531) begin
          if (_T_1510) begin
            _T_1525 <= _T_1517;
          end else begin
            _T_1525 <= 3'h0;
          end
        end else begin
          _T_1525 <= _T_1529;
        end
      end
    end
    if (reset) begin
      _T_1597 <= 1'h0;
    end else begin
      if (_T_1511) begin
        _T_1597 <= _T_1600;
      end
    end
    if (reset) begin
      _T_1640 <= 1'h0;
    end else begin
      if (_T_1641) begin
        _T_1640 <= _T_1643;
      end
    end
    if (reset) begin
      _T_1655 <= 1'h0;
    end else begin
      if (_T_1641) begin
        _T_1655 <= _T_1660;
      end
    end
    if (reset) begin
      _T_1944 <= 1'h0;
    end else begin
      _T_1944 <= _T_1958;
    end
    if (reset) begin
      _T_1986 <= 1'h0;
    end else begin
      _T_1986 <= _T_2000;
    end
    if (reset) begin
      _T_2028 <= 1'h0;
    end else begin
      _T_2028 <= _T_2042;
    end
    if (reset) begin
      _T_2070 <= 1'h0;
    end else begin
      _T_2070 <= _T_2084;
    end
    if (reset) begin
      _T_2112 <= 1'h0;
    end else begin
      _T_2112 <= _T_2126;
    end
    if (reset) begin
      _T_2154 <= 1'h0;
    end else begin
      _T_2154 <= _T_2168;
    end
    if (reset) begin
      _T_2196 <= 1'h0;
    end else begin
      _T_2196 <= _T_2210;
    end
    if (reset) begin
      _T_2238 <= 1'h0;
    end else begin
      _T_2238 <= _T_2252;
    end
    if (reset) begin
      _T_2280 <= 1'h0;
    end else begin
      _T_2280 <= _T_2294;
    end
    if (reset) begin
      _T_2322 <= 1'h0;
    end else begin
      _T_2322 <= _T_2336;
    end
    if (reset) begin
      _T_2364 <= 1'h0;
    end else begin
      _T_2364 <= _T_2378;
    end
    if (reset) begin
      _T_2406 <= 1'h0;
    end else begin
      _T_2406 <= _T_2420;
    end
    if (reset) begin
      _T_2448 <= 1'h0;
    end else begin
      _T_2448 <= _T_2462;
    end
    if (reset) begin
      _T_2490 <= 1'h0;
    end else begin
      _T_2490 <= _T_2504;
    end
    if (reset) begin
      _T_2532 <= 1'h0;
    end else begin
      _T_2532 <= _T_2546;
    end
    if (reset) begin
      _T_2574 <= 1'h0;
    end else begin
      _T_2574 <= _T_2588;
    end
    if (reset) begin
      _T_2616 <= 1'h0;
    end else begin
      _T_2616 <= _T_2630;
    end
    if (reset) begin
      _T_2658 <= 1'h0;
    end else begin
      _T_2658 <= _T_2672;
    end
    if (reset) begin
      _T_2700 <= 1'h0;
    end else begin
      _T_2700 <= _T_2714;
    end
    if (reset) begin
      _T_2742 <= 1'h0;
    end else begin
      _T_2742 <= _T_2756;
    end
    if (reset) begin
      _T_2784 <= 1'h0;
    end else begin
      _T_2784 <= _T_2798;
    end
    if (reset) begin
      _T_2826 <= 1'h0;
    end else begin
      _T_2826 <= _T_2840;
    end
    if (reset) begin
      _T_2868 <= 1'h0;
    end else begin
      _T_2868 <= _T_2882;
    end
    if (reset) begin
      _T_2910 <= 1'h0;
    end else begin
      _T_2910 <= _T_2924;
    end
    if (reset) begin
      _T_2952 <= 1'h0;
    end else begin
      _T_2952 <= _T_2966;
    end
    if (reset) begin
      _T_2994 <= 1'h0;
    end else begin
      _T_2994 <= _T_3008;
    end
    if (reset) begin
      _T_3036 <= 1'h0;
    end else begin
      _T_3036 <= _T_3050;
    end
    if (reset) begin
      _T_3078 <= 1'h0;
    end else begin
      _T_3078 <= _T_3092;
    end
    if (reset) begin
      _T_3120 <= 1'h0;
    end else begin
      _T_3120 <= _T_3134;
    end
    if (reset) begin
      _T_3162 <= 1'h0;
    end else begin
      _T_3162 <= _T_3176;
    end
    if (reset) begin
      _T_3204 <= 1'h0;
    end else begin
      _T_3204 <= _T_3218;
    end
    if (reset) begin
      _T_3246 <= 1'h0;
    end else begin
      _T_3246 <= _T_3260;
    end
    if (reset) begin
      _T_3288 <= 1'h0;
    end else begin
      _T_3288 <= _T_3302;
    end
    if (reset) begin
      _T_3330 <= 1'h0;
    end else begin
      _T_3330 <= _T_3344;
    end
    if (reset) begin
      _T_3372 <= 1'h0;
    end else begin
      _T_3372 <= _T_3386;
    end
    if (reset) begin
      _T_3414 <= 1'h0;
    end else begin
      _T_3414 <= _T_3428;
    end
    if (reset) begin
      _T_3456 <= 1'h0;
    end else begin
      _T_3456 <= _T_3470;
    end
    if (reset) begin
      _T_3498 <= 1'h0;
    end else begin
      _T_3498 <= _T_3512;
    end
    if (reset) begin
      _T_3540 <= 1'h0;
    end else begin
      _T_3540 <= _T_3554;
    end
    if (reset) begin
      _T_3582 <= 1'h0;
    end else begin
      _T_3582 <= _T_3596;
    end
    if (reset) begin
      _T_3624 <= 1'h0;
    end else begin
      _T_3624 <= _T_3638;
    end
    if (reset) begin
      _T_3666 <= 1'h0;
    end else begin
      _T_3666 <= _T_3680;
    end
    if (reset) begin
      _T_3708 <= 1'h0;
    end else begin
      _T_3708 <= _T_3722;
    end
    if (reset) begin
      _T_3750 <= 1'h0;
    end else begin
      _T_3750 <= _T_3764;
    end
    if (reset) begin
      _T_3792 <= 1'h0;
    end else begin
      _T_3792 <= _T_3806;
    end
    if (reset) begin
      _T_3834 <= 1'h0;
    end else begin
      _T_3834 <= _T_3848;
    end
    if (reset) begin
      _T_3876 <= 1'h0;
    end else begin
      _T_3876 <= _T_3890;
    end
    if (reset) begin
      _T_3918 <= 1'h0;
    end else begin
      _T_3918 <= _T_3932;
    end
    if (reset) begin
      _T_3960 <= 1'h0;
    end else begin
      _T_3960 <= _T_3974;
    end
    if (reset) begin
      _T_4002 <= 1'h0;
    end else begin
      _T_4002 <= _T_4016;
    end
    if (reset) begin
      _T_4044 <= 1'h0;
    end else begin
      _T_4044 <= _T_4058;
    end
    if (reset) begin
      _T_4086 <= 1'h0;
    end else begin
      _T_4086 <= _T_4100;
    end
    if (reset) begin
      _T_4128 <= 1'h0;
    end else begin
      _T_4128 <= _T_4142;
    end
    if (reset) begin
      _T_4170 <= 1'h0;
    end else begin
      _T_4170 <= _T_4184;
    end
    if (reset) begin
      _T_4212 <= 1'h0;
    end else begin
      _T_4212 <= _T_4226;
    end
    if (reset) begin
      _T_4254 <= 1'h0;
    end else begin
      _T_4254 <= _T_4268;
    end
    if (reset) begin
      _T_4296 <= 1'h0;
    end else begin
      _T_4296 <= _T_4310;
    end
    if (reset) begin
      _T_4338 <= 1'h0;
    end else begin
      _T_4338 <= _T_4352;
    end
    if (reset) begin
      _T_4380 <= 1'h0;
    end else begin
      _T_4380 <= _T_4394;
    end
    if (reset) begin
      _T_4422 <= 1'h0;
    end else begin
      _T_4422 <= _T_4436;
    end
    if (reset) begin
      _T_4464 <= 1'h0;
    end else begin
      _T_4464 <= _T_4478;
    end
    if (reset) begin
      _T_4506 <= 1'h0;
    end else begin
      _T_4506 <= _T_4520;
    end
    if (reset) begin
      _T_4548 <= 1'h0;
    end else begin
      _T_4548 <= _T_4562;
    end
    if (reset) begin
      _T_4590 <= 1'h0;
    end else begin
      _T_4590 <= _T_4604;
    end
    if (reset) begin
      _T_4632 <= 1'h0;
    end else begin
      _T_4632 <= _T_4646;
    end
    if (reset) begin
      _T_4674 <= 1'h0;
    end else begin
      _T_4674 <= _T_4688;
    end
    if (reset) begin
      _T_4716 <= 1'h0;
    end else begin
      _T_4716 <= _T_4730;
    end
    if (reset) begin
      _T_4758 <= 1'h0;
    end else begin
      _T_4758 <= _T_4772;
    end
    if (reset) begin
      _T_4800 <= 1'h0;
    end else begin
      _T_4800 <= _T_4814;
    end
    if (reset) begin
      _T_4842 <= 1'h0;
    end else begin
      _T_4842 <= _T_4856;
    end
    if (reset) begin
      _T_4884 <= 1'h0;
    end else begin
      _T_4884 <= _T_4898;
    end
    if (reset) begin
      _T_4926 <= 1'h0;
    end else begin
      _T_4926 <= _T_4940;
    end
    if (reset) begin
      _T_4968 <= 1'h0;
    end else begin
      _T_4968 <= _T_4982;
    end
    if (reset) begin
      _T_5010 <= 1'h0;
    end else begin
      _T_5010 <= _T_5024;
    end
    if (reset) begin
      _T_5052 <= 1'h0;
    end else begin
      _T_5052 <= _T_5066;
    end
    if (reset) begin
      _T_5094 <= 1'h0;
    end else begin
      _T_5094 <= _T_5108;
    end
    if (reset) begin
      _T_5136 <= 1'h0;
    end else begin
      _T_5136 <= _T_5150;
    end
    if (reset) begin
      _T_5178 <= 1'h0;
    end else begin
      _T_5178 <= _T_5192;
    end
    if (reset) begin
      _T_5220 <= 1'h0;
    end else begin
      _T_5220 <= _T_5234;
    end
    if (reset) begin
      _T_5262 <= 1'h0;
    end else begin
      _T_5262 <= _T_5276;
    end
    if (reset) begin
      _T_5304 <= 1'h0;
    end else begin
      _T_5304 <= _T_5318;
    end
    if (reset) begin
      _T_5346 <= 1'h0;
    end else begin
      _T_5346 <= _T_5360;
    end
    if (reset) begin
      _T_5388 <= 1'h0;
    end else begin
      _T_5388 <= _T_5402;
    end
    if (reset) begin
      _T_5430 <= 1'h0;
    end else begin
      _T_5430 <= _T_5444;
    end
    if (reset) begin
      _T_5472 <= 1'h0;
    end else begin
      _T_5472 <= _T_5486;
    end
    if (reset) begin
      _T_5514 <= 1'h0;
    end else begin
      _T_5514 <= _T_5528;
    end
    if (reset) begin
      _T_5556 <= 1'h0;
    end else begin
      _T_5556 <= _T_5570;
    end
    if (reset) begin
      _T_5598 <= 1'h0;
    end else begin
      _T_5598 <= _T_5612;
    end
    if (reset) begin
      _T_5640 <= 1'h0;
    end else begin
      _T_5640 <= _T_5654;
    end
    if (reset) begin
      _T_5682 <= 1'h0;
    end else begin
      _T_5682 <= _T_5696;
    end
    if (reset) begin
      _T_5724 <= 1'h0;
    end else begin
      _T_5724 <= _T_5738;
    end
    if (reset) begin
      _T_5766 <= 1'h0;
    end else begin
      _T_5766 <= _T_5780;
    end
    if (reset) begin
      _T_5808 <= 1'h0;
    end else begin
      _T_5808 <= _T_5822;
    end
    if (reset) begin
      _T_5850 <= 1'h0;
    end else begin
      _T_5850 <= _T_5864;
    end
    if (reset) begin
      _T_5892 <= 1'h0;
    end else begin
      _T_5892 <= _T_5906;
    end
    if (reset) begin
      _T_5934 <= 1'h0;
    end else begin
      _T_5934 <= _T_5948;
    end
    if (reset) begin
      _T_5976 <= 1'h0;
    end else begin
      _T_5976 <= _T_5990;
    end
    if (reset) begin
      _T_6018 <= 1'h0;
    end else begin
      _T_6018 <= _T_6032;
    end
    if (reset) begin
      _T_6060 <= 1'h0;
    end else begin
      _T_6060 <= _T_6074;
    end
    if (reset) begin
      _T_6102 <= 1'h0;
    end else begin
      _T_6102 <= _T_6116;
    end
    if (reset) begin
      _T_6144 <= 1'h0;
    end else begin
      _T_6144 <= _T_6158;
    end
    if (reset) begin
      _T_6186 <= 1'h0;
    end else begin
      _T_6186 <= _T_6200;
    end
    if (reset) begin
      _T_6228 <= 1'h0;
    end else begin
      _T_6228 <= _T_6242;
    end
    if (reset) begin
      _T_6270 <= 1'h0;
    end else begin
      _T_6270 <= _T_6284;
    end
    if (reset) begin
      _T_6312 <= 1'h0;
    end else begin
      _T_6312 <= _T_6326;
    end
    if (reset) begin
      _T_6354 <= 1'h0;
    end else begin
      _T_6354 <= _T_6368;
    end
    if (reset) begin
      _T_6396 <= 1'h0;
    end else begin
      _T_6396 <= _T_6410;
    end
    if (reset) begin
      _T_6438 <= 1'h0;
    end else begin
      _T_6438 <= _T_6452;
    end
    if (reset) begin
      _T_6480 <= 1'h0;
    end else begin
      _T_6480 <= _T_6494;
    end
    if (reset) begin
      _T_6522 <= 1'h0;
    end else begin
      _T_6522 <= _T_6536;
    end
    if (reset) begin
      _T_6564 <= 1'h0;
    end else begin
      _T_6564 <= _T_6578;
    end
    if (reset) begin
      _T_6606 <= 1'h0;
    end else begin
      _T_6606 <= _T_6620;
    end
    if (reset) begin
      _T_6648 <= 1'h0;
    end else begin
      _T_6648 <= _T_6662;
    end
    if (reset) begin
      _T_6690 <= 1'h0;
    end else begin
      _T_6690 <= _T_6704;
    end
    if (reset) begin
      _T_6732 <= 1'h0;
    end else begin
      _T_6732 <= _T_6746;
    end
    if (reset) begin
      _T_6774 <= 1'h0;
    end else begin
      _T_6774 <= _T_6788;
    end
    if (reset) begin
      _T_6816 <= 1'h0;
    end else begin
      _T_6816 <= _T_6830;
    end
    if (reset) begin
      _T_6858 <= 1'h0;
    end else begin
      _T_6858 <= _T_6872;
    end
    if (reset) begin
      _T_6900 <= 1'h0;
    end else begin
      _T_6900 <= _T_6914;
    end
    if (reset) begin
      _T_6942 <= 1'h0;
    end else begin
      _T_6942 <= _T_6956;
    end
    if (reset) begin
      _T_6984 <= 1'h0;
    end else begin
      _T_6984 <= _T_6998;
    end
    if (reset) begin
      _T_7026 <= 1'h0;
    end else begin
      _T_7026 <= _T_7040;
    end
    if (reset) begin
      _T_7068 <= 1'h0;
    end else begin
      _T_7068 <= _T_7082;
    end
    if (reset) begin
      _T_7110 <= 1'h0;
    end else begin
      _T_7110 <= _T_7124;
    end
    if (reset) begin
      _T_7152 <= 1'h0;
    end else begin
      _T_7152 <= _T_7166;
    end
    if (reset) begin
      _T_7194 <= 1'h0;
    end else begin
      _T_7194 <= _T_7208;
    end
    if (reset) begin
      _T_7236 <= 1'h0;
    end else begin
      _T_7236 <= _T_7250;
    end
    if (reset) begin
      _T_7278 <= 1'h0;
    end else begin
      _T_7278 <= _T_7292;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:106 assert (a_source  < UInt(BigInt(1) << sourceBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:107 assert (a_size    < UInt(BigInt(1) << sizeBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1967) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1967) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1976) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1976) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2009) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2009) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2018) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2018) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2051) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2051) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2060) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2060) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2093) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2093) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2102) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2135) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2144) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2177) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2186) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2228) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2261) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2270) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2303) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2312) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2345) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2354) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2387) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2396) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2396) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2429) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2429) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2438) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2438) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2471) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2471) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2480) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2480) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2513) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2513) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2522) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2522) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2555) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2555) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2564) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2564) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2597) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2597) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2606) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2639) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2639) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2648) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2648) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2681) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2681) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2690) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2690) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2723) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2732) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2732) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2765) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2765) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2774) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2774) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2807) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2807) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2816) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2816) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2849) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2849) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2858) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2858) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2891) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2891) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2900) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2900) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2933) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2933) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2942) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2942) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2975) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2975) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2984) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2984) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3017) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3017) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3026) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3026) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3059) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3059) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3068) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3068) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3101) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3110) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3143) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3152) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3185) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3194) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3227) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3236) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3269) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3278) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3311) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3311) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3320) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3353) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3362) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3395) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3395) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3404) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3404) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3437) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3437) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3446) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3446) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3479) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3479) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3488) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3488) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3521) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3521) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3530) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3530) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3563) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3563) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3572) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3572) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3605) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3605) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3614) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3614) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3647) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3647) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3656) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3656) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3689) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3689) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3698) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3698) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3731) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3731) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3740) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3740) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3773) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3773) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3782) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3782) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3815) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3815) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3824) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3824) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3857) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3857) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3866) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3866) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3899) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3899) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3908) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3908) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3941) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3941) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3950) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3950) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3983) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3983) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3992) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3992) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4025) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4025) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4034) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4034) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4067) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4067) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4076) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4076) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4109) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4118) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4151) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4160) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4193) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4235) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4244) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4277) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4286) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4319) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4328) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4328) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4361) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4361) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4370) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4370) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4403) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4403) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4412) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4412) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4445) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4445) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4454) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4454) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4487) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4487) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4496) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4496) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4529) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4529) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4538) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4538) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4571) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4571) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4580) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4613) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4622) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4622) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4655) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4655) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4664) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4664) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4697) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4697) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4706) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4706) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4739) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4739) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4748) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4748) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4781) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4781) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4790) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4790) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4823) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4823) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4832) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4832) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4865) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4865) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4874) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4874) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4907) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4907) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4916) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4916) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4949) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4949) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4958) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4958) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4991) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4991) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5000) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5033) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5033) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5042) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5042) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5075) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5075) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5084) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5084) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5117) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5126) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5159) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5168) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5210) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5243) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5252) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5285) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5294) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5327) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5336) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5369) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5369) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5378) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5378) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5411) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5411) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5420) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5420) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5453) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5453) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5462) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5462) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5495) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5504) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5504) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5537) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5537) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5546) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5546) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5579) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5579) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5588) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5588) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5621) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5621) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5630) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5630) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5663) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5663) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5672) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5672) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5705) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5705) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5714) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5714) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5747) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5747) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5756) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5756) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5789) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5789) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5798) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5798) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5831) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5831) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5840) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5840) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5873) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5873) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5882) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5882) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5915) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5915) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5924) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5924) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5957) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5957) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5966) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5966) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5999) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5999) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6008) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6008) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6041) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6041) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6050) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6050) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6083) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6083) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6092) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6092) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6134) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6167) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6176) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6209) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6218) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6251) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6260) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6293) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6302) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6335) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6344) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6377) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6377) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6386) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6386) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6419) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6419) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6428) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6428) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6461) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6461) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6470) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6470) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6503) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6503) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6512) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6512) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6545) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6545) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6554) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6554) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6587) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6587) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6596) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6596) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6629) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6629) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6638) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6638) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6671) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6671) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6680) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6680) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6713) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6713) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6722) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6722) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6755) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6755) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6764) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6764) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6797) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6797) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6806) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6806) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6839) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6839) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6848) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6848) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6881) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6881) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6890) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6890) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6923) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6923) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6932) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6932) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6965) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6965) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6974) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6974) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7007) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7007) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7016) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7016) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7049) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7049) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7058) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7058) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7091) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7091) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7100) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7133) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7142) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7175) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7184) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7217) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7226) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7259) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7268) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7301) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7310) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_7310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_trim(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [6:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [10:0] auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [6:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [10:0] auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [6:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [10:0] auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [6:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [10:0] auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [13:0] auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [13:0] auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [13:0] auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [13:0] auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [6:0] _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire [10:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [6:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [10:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [6:0] _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire [10:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [6:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [10:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire [13:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [13:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire [13:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [13:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire [2:0] _T_203;
  wire [13:0] _T_204;
  wire [2:0] _T_205;
  wire [13:0] _T_206;
  wire [10:0] _T_207;
  wire [10:0] _T_208;
  wire [17:0] _T_209;
  wire [17:0] _T_210;
  assign _T_203 = _T_31_ar_bits_id[6:4];
  assign _T_204 = {_T_31_ar_bits_user,_T_203};
  assign _T_205 = _T_31_aw_bits_id[6:4];
  assign _T_206 = {_T_31_aw_bits_user,_T_205};
  assign _T_207 = _T_89_r_bits_user[13:3];
  assign _T_208 = _T_89_b_bits_user[13:3];
  assign _T_209 = {_T_89_r_bits_user,_T_89_r_bits_id};
  assign _T_210 = {_T_89_b_bits_user,_T_89_b_bits_id};
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_89_aw_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_210[6:0];
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _T_208;
  assign _T_31_ar_ready = _T_89_ar_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_209[6:0];
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _T_207;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_31_aw_valid;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id[3:0];
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_lock = _T_31_aw_bits_lock;
  assign _T_89_aw_bits_cache = _T_31_aw_bits_cache;
  assign _T_89_aw_bits_prot = _T_31_aw_bits_prot;
  assign _T_89_aw_bits_qos = _T_31_aw_bits_qos;
  assign _T_89_aw_bits_user = _T_206;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_31_ar_valid;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id[3:0];
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_lock = _T_31_ar_bits_lock;
  assign _T_89_ar_bits_cache = _T_31_ar_bits_cache;
  assign _T_89_ar_bits_prot = _T_31_ar_bits_prot;
  assign _T_89_ar_bits_qos = _T_31_ar_bits_qos;
  assign _T_89_ar_bits_user = _T_204;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
endmodule
module Queue_34(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [13:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [13:0] io_deq_bits
);
  reg [13:0] ram [0:7];
  reg [31:0] _RAND_0;
  wire [13:0] ram__T_50_data;
  wire [2:0] ram__T_50_addr;
  wire [13:0] ram__T_36_data;
  wire [2:0] ram__T_36_addr;
  wire  ram__T_36_mask;
  wire  ram__T_36_en;
  reg [2:0] value;
  reg [31:0] _RAND_1;
  reg [2:0] value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [3:0] _T_39;
  wire [2:0] _T_40;
  wire [2:0] _GEN_4;
  wire [3:0] _T_43;
  wire [2:0] _T_44;
  wire [2:0] _GEN_5;
  wire  _T_45;
  wire  _GEN_6;
  wire  _T_47;
  wire  _T_49;
  assign ram__T_50_addr = value_1;
  assign ram__T_50_data = ram[ram__T_50_addr];
  assign ram__T_36_data = io_enq_bits;
  assign ram__T_36_addr = value;
  assign ram__T_36_mask = do_enq;
  assign ram__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 3'h1;
  assign _T_40 = _T_39[2:0];
  assign _GEN_4 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 3'h1;
  assign _T_44 = _T_43[2:0];
  assign _GEN_5 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_6 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits = ram__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[13:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_36_en & ram__T_36_mask) begin
      ram[ram__T_36_addr] <= ram__T_36_data;
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4UserYanker_yank(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [13:0] auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [13:0] auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [13:0] auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [13:0] auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire [13:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [13:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire [13:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [13:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [13:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [13:0] Queue_io_deq_bits;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [13:0] Queue_1_io_enq_bits;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [13:0] Queue_1_io_deq_bits;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [13:0] Queue_2_io_enq_bits;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [13:0] Queue_2_io_deq_bits;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [13:0] Queue_3_io_enq_bits;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [13:0] Queue_3_io_deq_bits;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [13:0] Queue_4_io_enq_bits;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [13:0] Queue_4_io_deq_bits;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [13:0] Queue_5_io_enq_bits;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [13:0] Queue_5_io_deq_bits;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [13:0] Queue_6_io_enq_bits;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [13:0] Queue_6_io_deq_bits;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [13:0] Queue_7_io_enq_bits;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [13:0] Queue_7_io_deq_bits;
  wire  Queue_8_clock;
  wire  Queue_8_reset;
  wire  Queue_8_io_enq_ready;
  wire  Queue_8_io_enq_valid;
  wire [13:0] Queue_8_io_enq_bits;
  wire  Queue_8_io_deq_ready;
  wire  Queue_8_io_deq_valid;
  wire [13:0] Queue_8_io_deq_bits;
  wire  Queue_9_clock;
  wire  Queue_9_reset;
  wire  Queue_9_io_enq_ready;
  wire  Queue_9_io_enq_valid;
  wire [13:0] Queue_9_io_enq_bits;
  wire  Queue_9_io_deq_ready;
  wire  Queue_9_io_deq_valid;
  wire [13:0] Queue_9_io_deq_bits;
  wire  Queue_10_clock;
  wire  Queue_10_reset;
  wire  Queue_10_io_enq_ready;
  wire  Queue_10_io_enq_valid;
  wire [13:0] Queue_10_io_enq_bits;
  wire  Queue_10_io_deq_ready;
  wire  Queue_10_io_deq_valid;
  wire [13:0] Queue_10_io_deq_bits;
  wire  Queue_11_clock;
  wire  Queue_11_reset;
  wire  Queue_11_io_enq_ready;
  wire  Queue_11_io_enq_valid;
  wire [13:0] Queue_11_io_enq_bits;
  wire  Queue_11_io_deq_ready;
  wire  Queue_11_io_deq_valid;
  wire [13:0] Queue_11_io_deq_bits;
  wire  Queue_12_clock;
  wire  Queue_12_reset;
  wire  Queue_12_io_enq_ready;
  wire  Queue_12_io_enq_valid;
  wire [13:0] Queue_12_io_enq_bits;
  wire  Queue_12_io_deq_ready;
  wire  Queue_12_io_deq_valid;
  wire [13:0] Queue_12_io_deq_bits;
  wire  Queue_13_clock;
  wire  Queue_13_reset;
  wire  Queue_13_io_enq_ready;
  wire  Queue_13_io_enq_valid;
  wire [13:0] Queue_13_io_enq_bits;
  wire  Queue_13_io_deq_ready;
  wire  Queue_13_io_deq_valid;
  wire [13:0] Queue_13_io_deq_bits;
  wire  Queue_14_clock;
  wire  Queue_14_reset;
  wire  Queue_14_io_enq_ready;
  wire  Queue_14_io_enq_valid;
  wire [13:0] Queue_14_io_enq_bits;
  wire  Queue_14_io_deq_ready;
  wire  Queue_14_io_deq_valid;
  wire [13:0] Queue_14_io_deq_bits;
  wire  Queue_15_clock;
  wire  Queue_15_reset;
  wire  Queue_15_io_enq_ready;
  wire  Queue_15_io_enq_valid;
  wire [13:0] Queue_15_io_enq_bits;
  wire  Queue_15_io_deq_ready;
  wire  Queue_15_io_deq_valid;
  wire [13:0] Queue_15_io_deq_bits;
  wire  Queue_16_clock;
  wire  Queue_16_reset;
  wire  Queue_16_io_enq_ready;
  wire  Queue_16_io_enq_valid;
  wire [13:0] Queue_16_io_enq_bits;
  wire  Queue_16_io_deq_ready;
  wire  Queue_16_io_deq_valid;
  wire [13:0] Queue_16_io_deq_bits;
  wire  Queue_17_clock;
  wire  Queue_17_reset;
  wire  Queue_17_io_enq_ready;
  wire  Queue_17_io_enq_valid;
  wire [13:0] Queue_17_io_enq_bits;
  wire  Queue_17_io_deq_ready;
  wire  Queue_17_io_deq_valid;
  wire [13:0] Queue_17_io_deq_bits;
  wire  Queue_18_clock;
  wire  Queue_18_reset;
  wire  Queue_18_io_enq_ready;
  wire  Queue_18_io_enq_valid;
  wire [13:0] Queue_18_io_enq_bits;
  wire  Queue_18_io_deq_ready;
  wire  Queue_18_io_deq_valid;
  wire [13:0] Queue_18_io_deq_bits;
  wire  Queue_19_clock;
  wire  Queue_19_reset;
  wire  Queue_19_io_enq_ready;
  wire  Queue_19_io_enq_valid;
  wire [13:0] Queue_19_io_enq_bits;
  wire  Queue_19_io_deq_ready;
  wire  Queue_19_io_deq_valid;
  wire [13:0] Queue_19_io_deq_bits;
  wire  Queue_20_clock;
  wire  Queue_20_reset;
  wire  Queue_20_io_enq_ready;
  wire  Queue_20_io_enq_valid;
  wire [13:0] Queue_20_io_enq_bits;
  wire  Queue_20_io_deq_ready;
  wire  Queue_20_io_deq_valid;
  wire [13:0] Queue_20_io_deq_bits;
  wire  Queue_21_clock;
  wire  Queue_21_reset;
  wire  Queue_21_io_enq_ready;
  wire  Queue_21_io_enq_valid;
  wire [13:0] Queue_21_io_enq_bits;
  wire  Queue_21_io_deq_ready;
  wire  Queue_21_io_deq_valid;
  wire [13:0] Queue_21_io_deq_bits;
  wire  Queue_22_clock;
  wire  Queue_22_reset;
  wire  Queue_22_io_enq_ready;
  wire  Queue_22_io_enq_valid;
  wire [13:0] Queue_22_io_enq_bits;
  wire  Queue_22_io_deq_ready;
  wire  Queue_22_io_deq_valid;
  wire [13:0] Queue_22_io_deq_bits;
  wire  Queue_23_clock;
  wire  Queue_23_reset;
  wire  Queue_23_io_enq_ready;
  wire  Queue_23_io_enq_valid;
  wire [13:0] Queue_23_io_enq_bits;
  wire  Queue_23_io_deq_ready;
  wire  Queue_23_io_deq_valid;
  wire [13:0] Queue_23_io_deq_bits;
  wire  Queue_24_clock;
  wire  Queue_24_reset;
  wire  Queue_24_io_enq_ready;
  wire  Queue_24_io_enq_valid;
  wire [13:0] Queue_24_io_enq_bits;
  wire  Queue_24_io_deq_ready;
  wire  Queue_24_io_deq_valid;
  wire [13:0] Queue_24_io_deq_bits;
  wire  Queue_25_clock;
  wire  Queue_25_reset;
  wire  Queue_25_io_enq_ready;
  wire  Queue_25_io_enq_valid;
  wire [13:0] Queue_25_io_enq_bits;
  wire  Queue_25_io_deq_ready;
  wire  Queue_25_io_deq_valid;
  wire [13:0] Queue_25_io_deq_bits;
  wire  Queue_26_clock;
  wire  Queue_26_reset;
  wire  Queue_26_io_enq_ready;
  wire  Queue_26_io_enq_valid;
  wire [13:0] Queue_26_io_enq_bits;
  wire  Queue_26_io_deq_ready;
  wire  Queue_26_io_deq_valid;
  wire [13:0] Queue_26_io_deq_bits;
  wire  Queue_27_clock;
  wire  Queue_27_reset;
  wire  Queue_27_io_enq_ready;
  wire  Queue_27_io_enq_valid;
  wire [13:0] Queue_27_io_enq_bits;
  wire  Queue_27_io_deq_ready;
  wire  Queue_27_io_deq_valid;
  wire [13:0] Queue_27_io_deq_bits;
  wire  Queue_28_clock;
  wire  Queue_28_reset;
  wire  Queue_28_io_enq_ready;
  wire  Queue_28_io_enq_valid;
  wire [13:0] Queue_28_io_enq_bits;
  wire  Queue_28_io_deq_ready;
  wire  Queue_28_io_deq_valid;
  wire [13:0] Queue_28_io_deq_bits;
  wire  Queue_29_clock;
  wire  Queue_29_reset;
  wire  Queue_29_io_enq_ready;
  wire  Queue_29_io_enq_valid;
  wire [13:0] Queue_29_io_enq_bits;
  wire  Queue_29_io_deq_ready;
  wire  Queue_29_io_deq_valid;
  wire [13:0] Queue_29_io_deq_bits;
  wire  Queue_30_clock;
  wire  Queue_30_reset;
  wire  Queue_30_io_enq_ready;
  wire  Queue_30_io_enq_valid;
  wire [13:0] Queue_30_io_enq_bits;
  wire  Queue_30_io_deq_ready;
  wire  Queue_30_io_deq_valid;
  wire [13:0] Queue_30_io_deq_bits;
  wire  Queue_31_clock;
  wire  Queue_31_reset;
  wire  Queue_31_io_enq_ready;
  wire  Queue_31_io_enq_valid;
  wire [13:0] Queue_31_io_enq_bits;
  wire  Queue_31_io_deq_ready;
  wire  Queue_31_io_deq_valid;
  wire [13:0] Queue_31_io_deq_bits;
  wire  _T_205_0;
  wire  _T_205_1;
  wire  _T_205_2;
  wire  _T_205_3;
  wire  _T_205_4;
  wire  _T_205_5;
  wire  _T_205_6;
  wire  _T_205_7;
  wire  _T_205_8;
  wire  _T_205_9;
  wire  _T_205_10;
  wire  _T_205_11;
  wire  _T_205_12;
  wire  _T_205_13;
  wire  _T_205_14;
  wire  _T_205_15;
  wire  _GEN_0;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _T_225;
  wire  _GEN_1;
  wire  _T_226;
  wire  _T_229_0;
  wire  _T_229_1;
  wire  _T_229_2;
  wire  _T_229_3;
  wire  _T_229_4;
  wire  _T_229_5;
  wire  _T_229_6;
  wire  _T_229_7;
  wire  _T_229_8;
  wire  _T_229_9;
  wire  _T_229_10;
  wire  _T_229_11;
  wire  _T_229_12;
  wire  _T_229_13;
  wire  _T_229_14;
  wire  _T_229_15;
  wire [13:0] _T_251_0;
  wire [13:0] _T_251_1;
  wire [13:0] _T_251_2;
  wire [13:0] _T_251_3;
  wire [13:0] _T_251_4;
  wire [13:0] _T_251_5;
  wire [13:0] _T_251_6;
  wire [13:0] _T_251_7;
  wire [13:0] _T_251_8;
  wire [13:0] _T_251_9;
  wire [13:0] _T_251_10;
  wire [13:0] _T_251_11;
  wire [13:0] _T_251_12;
  wire [13:0] _T_251_13;
  wire [13:0] _T_251_14;
  wire [13:0] _T_251_15;
  wire  _T_272;
  wire  _GEN_2;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _T_273;
  wire  _T_275;
  wire  _T_277;
  wire [13:0] _GEN_3;
  wire [13:0] _GEN_38;
  wire [13:0] _GEN_39;
  wire [13:0] _GEN_40;
  wire [13:0] _GEN_41;
  wire [13:0] _GEN_42;
  wire [13:0] _GEN_43;
  wire [13:0] _GEN_44;
  wire [13:0] _GEN_45;
  wire [13:0] _GEN_46;
  wire [13:0] _GEN_47;
  wire [13:0] _GEN_48;
  wire [13:0] _GEN_49;
  wire [13:0] _GEN_50;
  wire [13:0] _GEN_51;
  wire [13:0] _GEN_52;
  wire [15:0] _T_280;
  wire  _T_282;
  wire  _T_283;
  wire  _T_284;
  wire  _T_285;
  wire  _T_286;
  wire  _T_287;
  wire  _T_288;
  wire  _T_289;
  wire  _T_290;
  wire  _T_291;
  wire  _T_292;
  wire  _T_293;
  wire  _T_294;
  wire  _T_295;
  wire  _T_296;
  wire  _T_297;
  wire [15:0] _T_300;
  wire  _T_302;
  wire  _T_303;
  wire  _T_304;
  wire  _T_305;
  wire  _T_306;
  wire  _T_307;
  wire  _T_308;
  wire  _T_309;
  wire  _T_310;
  wire  _T_311;
  wire  _T_312;
  wire  _T_313;
  wire  _T_314;
  wire  _T_315;
  wire  _T_316;
  wire  _T_317;
  wire  _T_318;
  wire  _T_319;
  wire  _T_320;
  wire  _T_321;
  wire  _T_322;
  wire  _T_324;
  wire  _T_325;
  wire  _T_327;
  wire  _T_329;
  wire  _T_330;
  wire  _T_332;
  wire  _T_334;
  wire  _T_335;
  wire  _T_337;
  wire  _T_339;
  wire  _T_340;
  wire  _T_342;
  wire  _T_344;
  wire  _T_345;
  wire  _T_347;
  wire  _T_349;
  wire  _T_350;
  wire  _T_352;
  wire  _T_354;
  wire  _T_355;
  wire  _T_357;
  wire  _T_359;
  wire  _T_360;
  wire  _T_362;
  wire  _T_364;
  wire  _T_365;
  wire  _T_367;
  wire  _T_369;
  wire  _T_370;
  wire  _T_372;
  wire  _T_374;
  wire  _T_375;
  wire  _T_377;
  wire  _T_379;
  wire  _T_380;
  wire  _T_382;
  wire  _T_384;
  wire  _T_385;
  wire  _T_387;
  wire  _T_389;
  wire  _T_390;
  wire  _T_392;
  wire  _T_394;
  wire  _T_395;
  wire  _T_397;
  wire  _T_400_0;
  wire  _T_400_1;
  wire  _T_400_2;
  wire  _T_400_3;
  wire  _T_400_4;
  wire  _T_400_5;
  wire  _T_400_6;
  wire  _T_400_7;
  wire  _T_400_8;
  wire  _T_400_9;
  wire  _T_400_10;
  wire  _T_400_11;
  wire  _T_400_12;
  wire  _T_400_13;
  wire  _T_400_14;
  wire  _T_400_15;
  wire  _GEN_4;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _T_420;
  wire  _GEN_5;
  wire  _T_421;
  wire  _T_424_0;
  wire  _T_424_1;
  wire  _T_424_2;
  wire  _T_424_3;
  wire  _T_424_4;
  wire  _T_424_5;
  wire  _T_424_6;
  wire  _T_424_7;
  wire  _T_424_8;
  wire  _T_424_9;
  wire  _T_424_10;
  wire  _T_424_11;
  wire  _T_424_12;
  wire  _T_424_13;
  wire  _T_424_14;
  wire  _T_424_15;
  wire [13:0] _T_446_0;
  wire [13:0] _T_446_1;
  wire [13:0] _T_446_2;
  wire [13:0] _T_446_3;
  wire [13:0] _T_446_4;
  wire [13:0] _T_446_5;
  wire [13:0] _T_446_6;
  wire [13:0] _T_446_7;
  wire [13:0] _T_446_8;
  wire [13:0] _T_446_9;
  wire [13:0] _T_446_10;
  wire [13:0] _T_446_11;
  wire [13:0] _T_446_12;
  wire [13:0] _T_446_13;
  wire [13:0] _T_446_14;
  wire [13:0] _T_446_15;
  wire  _T_467;
  wire  _GEN_6;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _T_468;
  wire  _T_470;
  wire  _T_472;
  wire [13:0] _GEN_7;
  wire [13:0] _GEN_83;
  wire [13:0] _GEN_84;
  wire [13:0] _GEN_85;
  wire [13:0] _GEN_86;
  wire [13:0] _GEN_87;
  wire [13:0] _GEN_88;
  wire [13:0] _GEN_89;
  wire [13:0] _GEN_90;
  wire [13:0] _GEN_91;
  wire [13:0] _GEN_92;
  wire [13:0] _GEN_93;
  wire [13:0] _GEN_94;
  wire [13:0] _GEN_95;
  wire [13:0] _GEN_96;
  wire [13:0] _GEN_97;
  wire [15:0] _T_475;
  wire  _T_477;
  wire  _T_478;
  wire  _T_479;
  wire  _T_480;
  wire  _T_481;
  wire  _T_482;
  wire  _T_483;
  wire  _T_484;
  wire  _T_485;
  wire  _T_486;
  wire  _T_487;
  wire  _T_488;
  wire  _T_489;
  wire  _T_490;
  wire  _T_491;
  wire  _T_492;
  wire [15:0] _T_495;
  wire  _T_497;
  wire  _T_498;
  wire  _T_499;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire  _T_507;
  wire  _T_508;
  wire  _T_509;
  wire  _T_510;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_515;
  wire  _T_516;
  wire  _T_518;
  wire  _T_520;
  wire  _T_522;
  wire  _T_524;
  wire  _T_526;
  wire  _T_528;
  wire  _T_530;
  wire  _T_532;
  wire  _T_534;
  wire  _T_536;
  wire  _T_538;
  wire  _T_540;
  wire  _T_542;
  wire  _T_544;
  wire  _T_546;
  wire  _T_548;
  wire  _T_550;
  wire  _T_552;
  wire  _T_554;
  wire  _T_556;
  wire  _T_558;
  wire  _T_560;
  wire  _T_562;
  wire  _T_564;
  wire  _T_566;
  wire  _T_568;
  wire  _T_570;
  wire  _T_572;
  wire  _T_574;
  wire  _T_576;
  Queue_34 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_34 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_34 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_34 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  Queue_34 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_34 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  Queue_34 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  Queue_34 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  Queue_34 Queue_8 (
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits(Queue_8_io_enq_bits),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits(Queue_8_io_deq_bits)
  );
  Queue_34 Queue_9 (
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits(Queue_9_io_enq_bits),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits(Queue_9_io_deq_bits)
  );
  Queue_34 Queue_10 (
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  Queue_34 Queue_11 (
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits(Queue_11_io_enq_bits),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits(Queue_11_io_deq_bits)
  );
  Queue_34 Queue_12 (
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits(Queue_12_io_enq_bits),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits(Queue_12_io_deq_bits)
  );
  Queue_34 Queue_13 (
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits(Queue_13_io_enq_bits),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits(Queue_13_io_deq_bits)
  );
  Queue_34 Queue_14 (
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits(Queue_14_io_enq_bits),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits(Queue_14_io_deq_bits)
  );
  Queue_34 Queue_15 (
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits(Queue_15_io_enq_bits),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits(Queue_15_io_deq_bits)
  );
  Queue_34 Queue_16 (
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits(Queue_16_io_enq_bits),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits(Queue_16_io_deq_bits)
  );
  Queue_34 Queue_17 (
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits(Queue_17_io_enq_bits),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits(Queue_17_io_deq_bits)
  );
  Queue_34 Queue_18 (
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits(Queue_18_io_enq_bits),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits(Queue_18_io_deq_bits)
  );
  Queue_34 Queue_19 (
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits(Queue_19_io_enq_bits),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits(Queue_19_io_deq_bits)
  );
  Queue_34 Queue_20 (
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits(Queue_20_io_enq_bits),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits(Queue_20_io_deq_bits)
  );
  Queue_34 Queue_21 (
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits(Queue_21_io_enq_bits),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits(Queue_21_io_deq_bits)
  );
  Queue_34 Queue_22 (
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits(Queue_22_io_enq_bits),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits(Queue_22_io_deq_bits)
  );
  Queue_34 Queue_23 (
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits(Queue_23_io_enq_bits),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits(Queue_23_io_deq_bits)
  );
  Queue_34 Queue_24 (
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits(Queue_24_io_enq_bits),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits(Queue_24_io_deq_bits)
  );
  Queue_34 Queue_25 (
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits(Queue_25_io_enq_bits),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits(Queue_25_io_deq_bits)
  );
  Queue_34 Queue_26 (
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits(Queue_26_io_enq_bits),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits(Queue_26_io_deq_bits)
  );
  Queue_34 Queue_27 (
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits(Queue_27_io_enq_bits),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits(Queue_27_io_deq_bits)
  );
  Queue_34 Queue_28 (
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits(Queue_28_io_enq_bits),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits(Queue_28_io_deq_bits)
  );
  Queue_34 Queue_29 (
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits(Queue_29_io_enq_bits),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits(Queue_29_io_deq_bits)
  );
  Queue_34 Queue_30 (
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits(Queue_30_io_enq_bits),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits(Queue_30_io_deq_bits)
  );
  Queue_34 Queue_31 (
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits(Queue_31_io_enq_bits),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits(Queue_31_io_deq_bits)
  );
  assign _GEN_8 = 4'h1 == _T_31_ar_bits_id ? _T_205_1 : _T_205_0;
  assign _GEN_9 = 4'h2 == _T_31_ar_bits_id ? _T_205_2 : _GEN_8;
  assign _GEN_10 = 4'h3 == _T_31_ar_bits_id ? _T_205_3 : _GEN_9;
  assign _GEN_11 = 4'h4 == _T_31_ar_bits_id ? _T_205_4 : _GEN_10;
  assign _GEN_12 = 4'h5 == _T_31_ar_bits_id ? _T_205_5 : _GEN_11;
  assign _GEN_13 = 4'h6 == _T_31_ar_bits_id ? _T_205_6 : _GEN_12;
  assign _GEN_14 = 4'h7 == _T_31_ar_bits_id ? _T_205_7 : _GEN_13;
  assign _GEN_15 = 4'h8 == _T_31_ar_bits_id ? _T_205_8 : _GEN_14;
  assign _GEN_16 = 4'h9 == _T_31_ar_bits_id ? _T_205_9 : _GEN_15;
  assign _GEN_17 = 4'ha == _T_31_ar_bits_id ? _T_205_10 : _GEN_16;
  assign _GEN_18 = 4'hb == _T_31_ar_bits_id ? _T_205_11 : _GEN_17;
  assign _GEN_19 = 4'hc == _T_31_ar_bits_id ? _T_205_12 : _GEN_18;
  assign _GEN_20 = 4'hd == _T_31_ar_bits_id ? _T_205_13 : _GEN_19;
  assign _GEN_21 = 4'he == _T_31_ar_bits_id ? _T_205_14 : _GEN_20;
  assign _GEN_22 = 4'hf == _T_31_ar_bits_id ? _T_205_15 : _GEN_21;
  assign _T_225 = _T_89_ar_ready & _GEN_0;
  assign _T_226 = _T_31_ar_valid & _GEN_1;
  assign _T_272 = _T_89_r_valid == 1'h0;
  assign _GEN_23 = 4'h1 == _T_89_r_bits_id ? _T_229_1 : _T_229_0;
  assign _GEN_24 = 4'h2 == _T_89_r_bits_id ? _T_229_2 : _GEN_23;
  assign _GEN_25 = 4'h3 == _T_89_r_bits_id ? _T_229_3 : _GEN_24;
  assign _GEN_26 = 4'h4 == _T_89_r_bits_id ? _T_229_4 : _GEN_25;
  assign _GEN_27 = 4'h5 == _T_89_r_bits_id ? _T_229_5 : _GEN_26;
  assign _GEN_28 = 4'h6 == _T_89_r_bits_id ? _T_229_6 : _GEN_27;
  assign _GEN_29 = 4'h7 == _T_89_r_bits_id ? _T_229_7 : _GEN_28;
  assign _GEN_30 = 4'h8 == _T_89_r_bits_id ? _T_229_8 : _GEN_29;
  assign _GEN_31 = 4'h9 == _T_89_r_bits_id ? _T_229_9 : _GEN_30;
  assign _GEN_32 = 4'ha == _T_89_r_bits_id ? _T_229_10 : _GEN_31;
  assign _GEN_33 = 4'hb == _T_89_r_bits_id ? _T_229_11 : _GEN_32;
  assign _GEN_34 = 4'hc == _T_89_r_bits_id ? _T_229_12 : _GEN_33;
  assign _GEN_35 = 4'hd == _T_89_r_bits_id ? _T_229_13 : _GEN_34;
  assign _GEN_36 = 4'he == _T_89_r_bits_id ? _T_229_14 : _GEN_35;
  assign _GEN_37 = 4'hf == _T_89_r_bits_id ? _T_229_15 : _GEN_36;
  assign _T_273 = _T_272 | _GEN_2;
  assign _T_275 = _T_273 | reset;
  assign _T_277 = _T_275 == 1'h0;
  assign _GEN_38 = 4'h1 == _T_89_r_bits_id ? _T_251_1 : _T_251_0;
  assign _GEN_39 = 4'h2 == _T_89_r_bits_id ? _T_251_2 : _GEN_38;
  assign _GEN_40 = 4'h3 == _T_89_r_bits_id ? _T_251_3 : _GEN_39;
  assign _GEN_41 = 4'h4 == _T_89_r_bits_id ? _T_251_4 : _GEN_40;
  assign _GEN_42 = 4'h5 == _T_89_r_bits_id ? _T_251_5 : _GEN_41;
  assign _GEN_43 = 4'h6 == _T_89_r_bits_id ? _T_251_6 : _GEN_42;
  assign _GEN_44 = 4'h7 == _T_89_r_bits_id ? _T_251_7 : _GEN_43;
  assign _GEN_45 = 4'h8 == _T_89_r_bits_id ? _T_251_8 : _GEN_44;
  assign _GEN_46 = 4'h9 == _T_89_r_bits_id ? _T_251_9 : _GEN_45;
  assign _GEN_47 = 4'ha == _T_89_r_bits_id ? _T_251_10 : _GEN_46;
  assign _GEN_48 = 4'hb == _T_89_r_bits_id ? _T_251_11 : _GEN_47;
  assign _GEN_49 = 4'hc == _T_89_r_bits_id ? _T_251_12 : _GEN_48;
  assign _GEN_50 = 4'hd == _T_89_r_bits_id ? _T_251_13 : _GEN_49;
  assign _GEN_51 = 4'he == _T_89_r_bits_id ? _T_251_14 : _GEN_50;
  assign _GEN_52 = 4'hf == _T_89_r_bits_id ? _T_251_15 : _GEN_51;
  assign _T_280 = 16'h1 << _T_31_ar_bits_id;
  assign _T_282 = _T_280[0];
  assign _T_283 = _T_280[1];
  assign _T_284 = _T_280[2];
  assign _T_285 = _T_280[3];
  assign _T_286 = _T_280[4];
  assign _T_287 = _T_280[5];
  assign _T_288 = _T_280[6];
  assign _T_289 = _T_280[7];
  assign _T_290 = _T_280[8];
  assign _T_291 = _T_280[9];
  assign _T_292 = _T_280[10];
  assign _T_293 = _T_280[11];
  assign _T_294 = _T_280[12];
  assign _T_295 = _T_280[13];
  assign _T_296 = _T_280[14];
  assign _T_297 = _T_280[15];
  assign _T_300 = 16'h1 << _T_89_r_bits_id;
  assign _T_302 = _T_300[0];
  assign _T_303 = _T_300[1];
  assign _T_304 = _T_300[2];
  assign _T_305 = _T_300[3];
  assign _T_306 = _T_300[4];
  assign _T_307 = _T_300[5];
  assign _T_308 = _T_300[6];
  assign _T_309 = _T_300[7];
  assign _T_310 = _T_300[8];
  assign _T_311 = _T_300[9];
  assign _T_312 = _T_300[10];
  assign _T_313 = _T_300[11];
  assign _T_314 = _T_300[12];
  assign _T_315 = _T_300[13];
  assign _T_316 = _T_300[14];
  assign _T_317 = _T_300[15];
  assign _T_318 = _T_89_r_valid & _T_31_r_ready;
  assign _T_319 = _T_318 & _T_302;
  assign _T_320 = _T_319 & _T_89_r_bits_last;
  assign _T_321 = _T_31_ar_valid & _T_89_ar_ready;
  assign _T_322 = _T_321 & _T_282;
  assign _T_324 = _T_318 & _T_303;
  assign _T_325 = _T_324 & _T_89_r_bits_last;
  assign _T_327 = _T_321 & _T_283;
  assign _T_329 = _T_318 & _T_304;
  assign _T_330 = _T_329 & _T_89_r_bits_last;
  assign _T_332 = _T_321 & _T_284;
  assign _T_334 = _T_318 & _T_305;
  assign _T_335 = _T_334 & _T_89_r_bits_last;
  assign _T_337 = _T_321 & _T_285;
  assign _T_339 = _T_318 & _T_306;
  assign _T_340 = _T_339 & _T_89_r_bits_last;
  assign _T_342 = _T_321 & _T_286;
  assign _T_344 = _T_318 & _T_307;
  assign _T_345 = _T_344 & _T_89_r_bits_last;
  assign _T_347 = _T_321 & _T_287;
  assign _T_349 = _T_318 & _T_308;
  assign _T_350 = _T_349 & _T_89_r_bits_last;
  assign _T_352 = _T_321 & _T_288;
  assign _T_354 = _T_318 & _T_309;
  assign _T_355 = _T_354 & _T_89_r_bits_last;
  assign _T_357 = _T_321 & _T_289;
  assign _T_359 = _T_318 & _T_310;
  assign _T_360 = _T_359 & _T_89_r_bits_last;
  assign _T_362 = _T_321 & _T_290;
  assign _T_364 = _T_318 & _T_311;
  assign _T_365 = _T_364 & _T_89_r_bits_last;
  assign _T_367 = _T_321 & _T_291;
  assign _T_369 = _T_318 & _T_312;
  assign _T_370 = _T_369 & _T_89_r_bits_last;
  assign _T_372 = _T_321 & _T_292;
  assign _T_374 = _T_318 & _T_313;
  assign _T_375 = _T_374 & _T_89_r_bits_last;
  assign _T_377 = _T_321 & _T_293;
  assign _T_379 = _T_318 & _T_314;
  assign _T_380 = _T_379 & _T_89_r_bits_last;
  assign _T_382 = _T_321 & _T_294;
  assign _T_384 = _T_318 & _T_315;
  assign _T_385 = _T_384 & _T_89_r_bits_last;
  assign _T_387 = _T_321 & _T_295;
  assign _T_389 = _T_318 & _T_316;
  assign _T_390 = _T_389 & _T_89_r_bits_last;
  assign _T_392 = _T_321 & _T_296;
  assign _T_394 = _T_318 & _T_317;
  assign _T_395 = _T_394 & _T_89_r_bits_last;
  assign _T_397 = _T_321 & _T_297;
  assign _GEN_53 = 4'h1 == _T_31_aw_bits_id ? _T_400_1 : _T_400_0;
  assign _GEN_54 = 4'h2 == _T_31_aw_bits_id ? _T_400_2 : _GEN_53;
  assign _GEN_55 = 4'h3 == _T_31_aw_bits_id ? _T_400_3 : _GEN_54;
  assign _GEN_56 = 4'h4 == _T_31_aw_bits_id ? _T_400_4 : _GEN_55;
  assign _GEN_57 = 4'h5 == _T_31_aw_bits_id ? _T_400_5 : _GEN_56;
  assign _GEN_58 = 4'h6 == _T_31_aw_bits_id ? _T_400_6 : _GEN_57;
  assign _GEN_59 = 4'h7 == _T_31_aw_bits_id ? _T_400_7 : _GEN_58;
  assign _GEN_60 = 4'h8 == _T_31_aw_bits_id ? _T_400_8 : _GEN_59;
  assign _GEN_61 = 4'h9 == _T_31_aw_bits_id ? _T_400_9 : _GEN_60;
  assign _GEN_62 = 4'ha == _T_31_aw_bits_id ? _T_400_10 : _GEN_61;
  assign _GEN_63 = 4'hb == _T_31_aw_bits_id ? _T_400_11 : _GEN_62;
  assign _GEN_64 = 4'hc == _T_31_aw_bits_id ? _T_400_12 : _GEN_63;
  assign _GEN_65 = 4'hd == _T_31_aw_bits_id ? _T_400_13 : _GEN_64;
  assign _GEN_66 = 4'he == _T_31_aw_bits_id ? _T_400_14 : _GEN_65;
  assign _GEN_67 = 4'hf == _T_31_aw_bits_id ? _T_400_15 : _GEN_66;
  assign _T_420 = _T_89_aw_ready & _GEN_4;
  assign _T_421 = _T_31_aw_valid & _GEN_5;
  assign _T_467 = _T_89_b_valid == 1'h0;
  assign _GEN_68 = 4'h1 == _T_89_b_bits_id ? _T_424_1 : _T_424_0;
  assign _GEN_69 = 4'h2 == _T_89_b_bits_id ? _T_424_2 : _GEN_68;
  assign _GEN_70 = 4'h3 == _T_89_b_bits_id ? _T_424_3 : _GEN_69;
  assign _GEN_71 = 4'h4 == _T_89_b_bits_id ? _T_424_4 : _GEN_70;
  assign _GEN_72 = 4'h5 == _T_89_b_bits_id ? _T_424_5 : _GEN_71;
  assign _GEN_73 = 4'h6 == _T_89_b_bits_id ? _T_424_6 : _GEN_72;
  assign _GEN_74 = 4'h7 == _T_89_b_bits_id ? _T_424_7 : _GEN_73;
  assign _GEN_75 = 4'h8 == _T_89_b_bits_id ? _T_424_8 : _GEN_74;
  assign _GEN_76 = 4'h9 == _T_89_b_bits_id ? _T_424_9 : _GEN_75;
  assign _GEN_77 = 4'ha == _T_89_b_bits_id ? _T_424_10 : _GEN_76;
  assign _GEN_78 = 4'hb == _T_89_b_bits_id ? _T_424_11 : _GEN_77;
  assign _GEN_79 = 4'hc == _T_89_b_bits_id ? _T_424_12 : _GEN_78;
  assign _GEN_80 = 4'hd == _T_89_b_bits_id ? _T_424_13 : _GEN_79;
  assign _GEN_81 = 4'he == _T_89_b_bits_id ? _T_424_14 : _GEN_80;
  assign _GEN_82 = 4'hf == _T_89_b_bits_id ? _T_424_15 : _GEN_81;
  assign _T_468 = _T_467 | _GEN_6;
  assign _T_470 = _T_468 | reset;
  assign _T_472 = _T_470 == 1'h0;
  assign _GEN_83 = 4'h1 == _T_89_b_bits_id ? _T_446_1 : _T_446_0;
  assign _GEN_84 = 4'h2 == _T_89_b_bits_id ? _T_446_2 : _GEN_83;
  assign _GEN_85 = 4'h3 == _T_89_b_bits_id ? _T_446_3 : _GEN_84;
  assign _GEN_86 = 4'h4 == _T_89_b_bits_id ? _T_446_4 : _GEN_85;
  assign _GEN_87 = 4'h5 == _T_89_b_bits_id ? _T_446_5 : _GEN_86;
  assign _GEN_88 = 4'h6 == _T_89_b_bits_id ? _T_446_6 : _GEN_87;
  assign _GEN_89 = 4'h7 == _T_89_b_bits_id ? _T_446_7 : _GEN_88;
  assign _GEN_90 = 4'h8 == _T_89_b_bits_id ? _T_446_8 : _GEN_89;
  assign _GEN_91 = 4'h9 == _T_89_b_bits_id ? _T_446_9 : _GEN_90;
  assign _GEN_92 = 4'ha == _T_89_b_bits_id ? _T_446_10 : _GEN_91;
  assign _GEN_93 = 4'hb == _T_89_b_bits_id ? _T_446_11 : _GEN_92;
  assign _GEN_94 = 4'hc == _T_89_b_bits_id ? _T_446_12 : _GEN_93;
  assign _GEN_95 = 4'hd == _T_89_b_bits_id ? _T_446_13 : _GEN_94;
  assign _GEN_96 = 4'he == _T_89_b_bits_id ? _T_446_14 : _GEN_95;
  assign _GEN_97 = 4'hf == _T_89_b_bits_id ? _T_446_15 : _GEN_96;
  assign _T_475 = 16'h1 << _T_31_aw_bits_id;
  assign _T_477 = _T_475[0];
  assign _T_478 = _T_475[1];
  assign _T_479 = _T_475[2];
  assign _T_480 = _T_475[3];
  assign _T_481 = _T_475[4];
  assign _T_482 = _T_475[5];
  assign _T_483 = _T_475[6];
  assign _T_484 = _T_475[7];
  assign _T_485 = _T_475[8];
  assign _T_486 = _T_475[9];
  assign _T_487 = _T_475[10];
  assign _T_488 = _T_475[11];
  assign _T_489 = _T_475[12];
  assign _T_490 = _T_475[13];
  assign _T_491 = _T_475[14];
  assign _T_492 = _T_475[15];
  assign _T_495 = 16'h1 << _T_89_b_bits_id;
  assign _T_497 = _T_495[0];
  assign _T_498 = _T_495[1];
  assign _T_499 = _T_495[2];
  assign _T_500 = _T_495[3];
  assign _T_501 = _T_495[4];
  assign _T_502 = _T_495[5];
  assign _T_503 = _T_495[6];
  assign _T_504 = _T_495[7];
  assign _T_505 = _T_495[8];
  assign _T_506 = _T_495[9];
  assign _T_507 = _T_495[10];
  assign _T_508 = _T_495[11];
  assign _T_509 = _T_495[12];
  assign _T_510 = _T_495[13];
  assign _T_511 = _T_495[14];
  assign _T_512 = _T_495[15];
  assign _T_513 = _T_89_b_valid & _T_31_b_ready;
  assign _T_514 = _T_513 & _T_497;
  assign _T_515 = _T_31_aw_valid & _T_89_aw_ready;
  assign _T_516 = _T_515 & _T_477;
  assign _T_518 = _T_513 & _T_498;
  assign _T_520 = _T_515 & _T_478;
  assign _T_522 = _T_513 & _T_499;
  assign _T_524 = _T_515 & _T_479;
  assign _T_526 = _T_513 & _T_500;
  assign _T_528 = _T_515 & _T_480;
  assign _T_530 = _T_513 & _T_501;
  assign _T_532 = _T_515 & _T_481;
  assign _T_534 = _T_513 & _T_502;
  assign _T_536 = _T_515 & _T_482;
  assign _T_538 = _T_513 & _T_503;
  assign _T_540 = _T_515 & _T_483;
  assign _T_542 = _T_513 & _T_504;
  assign _T_544 = _T_515 & _T_484;
  assign _T_546 = _T_513 & _T_505;
  assign _T_548 = _T_515 & _T_485;
  assign _T_550 = _T_513 & _T_506;
  assign _T_552 = _T_515 & _T_486;
  assign _T_554 = _T_513 & _T_507;
  assign _T_556 = _T_515 & _T_487;
  assign _T_558 = _T_513 & _T_508;
  assign _T_560 = _T_515 & _T_488;
  assign _T_562 = _T_513 & _T_509;
  assign _T_564 = _T_515 & _T_489;
  assign _T_566 = _T_513 & _T_510;
  assign _T_568 = _T_515 & _T_490;
  assign _T_570 = _T_513 & _T_511;
  assign _T_572 = _T_515 & _T_491;
  assign _T_574 = _T_513 & _T_512;
  assign _T_576 = _T_515 & _T_492;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_420;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _GEN_7;
  assign _T_31_ar_ready = _T_225;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _GEN_3;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_421;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id;
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_lock = _T_31_aw_bits_lock;
  assign _T_89_aw_bits_cache = _T_31_aw_bits_cache;
  assign _T_89_aw_bits_prot = _T_31_aw_bits_prot;
  assign _T_89_aw_bits_qos = _T_31_aw_bits_qos;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_226;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id;
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_lock = _T_31_ar_bits_lock;
  assign _T_89_ar_bits_cache = _T_31_ar_bits_cache;
  assign _T_89_ar_bits_prot = _T_31_ar_bits_prot;
  assign _T_89_ar_bits_qos = _T_31_ar_bits_qos;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_322;
  assign Queue_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_io_deq_ready = _T_320;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_327;
  assign Queue_1_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_1_io_deq_ready = _T_325;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_2_io_enq_valid = _T_332;
  assign Queue_2_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_2_io_deq_ready = _T_330;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_3_io_enq_valid = _T_337;
  assign Queue_3_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_3_io_deq_ready = _T_335;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_4_io_enq_valid = _T_342;
  assign Queue_4_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_4_io_deq_ready = _T_340;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_5_io_enq_valid = _T_347;
  assign Queue_5_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_5_io_deq_ready = _T_345;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_6_io_enq_valid = _T_352;
  assign Queue_6_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_6_io_deq_ready = _T_350;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_7_io_enq_valid = _T_357;
  assign Queue_7_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_7_io_deq_ready = _T_355;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_8_io_enq_valid = _T_362;
  assign Queue_8_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_8_io_deq_ready = _T_360;
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_9_io_enq_valid = _T_367;
  assign Queue_9_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_9_io_deq_ready = _T_365;
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_10_io_enq_valid = _T_372;
  assign Queue_10_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_10_io_deq_ready = _T_370;
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_11_io_enq_valid = _T_377;
  assign Queue_11_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_11_io_deq_ready = _T_375;
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_12_io_enq_valid = _T_382;
  assign Queue_12_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_12_io_deq_ready = _T_380;
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_13_io_enq_valid = _T_387;
  assign Queue_13_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_13_io_deq_ready = _T_385;
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_14_io_enq_valid = _T_392;
  assign Queue_14_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_14_io_deq_ready = _T_390;
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_15_io_enq_valid = _T_397;
  assign Queue_15_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_15_io_deq_ready = _T_395;
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign Queue_16_io_enq_valid = _T_516;
  assign Queue_16_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_16_io_deq_ready = _T_514;
  assign Queue_16_clock = clock;
  assign Queue_16_reset = reset;
  assign Queue_17_io_enq_valid = _T_520;
  assign Queue_17_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_17_io_deq_ready = _T_518;
  assign Queue_17_clock = clock;
  assign Queue_17_reset = reset;
  assign Queue_18_io_enq_valid = _T_524;
  assign Queue_18_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_18_io_deq_ready = _T_522;
  assign Queue_18_clock = clock;
  assign Queue_18_reset = reset;
  assign Queue_19_io_enq_valid = _T_528;
  assign Queue_19_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_19_io_deq_ready = _T_526;
  assign Queue_19_clock = clock;
  assign Queue_19_reset = reset;
  assign Queue_20_io_enq_valid = _T_532;
  assign Queue_20_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_20_io_deq_ready = _T_530;
  assign Queue_20_clock = clock;
  assign Queue_20_reset = reset;
  assign Queue_21_io_enq_valid = _T_536;
  assign Queue_21_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_21_io_deq_ready = _T_534;
  assign Queue_21_clock = clock;
  assign Queue_21_reset = reset;
  assign Queue_22_io_enq_valid = _T_540;
  assign Queue_22_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_22_io_deq_ready = _T_538;
  assign Queue_22_clock = clock;
  assign Queue_22_reset = reset;
  assign Queue_23_io_enq_valid = _T_544;
  assign Queue_23_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_23_io_deq_ready = _T_542;
  assign Queue_23_clock = clock;
  assign Queue_23_reset = reset;
  assign Queue_24_io_enq_valid = _T_548;
  assign Queue_24_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_24_io_deq_ready = _T_546;
  assign Queue_24_clock = clock;
  assign Queue_24_reset = reset;
  assign Queue_25_io_enq_valid = _T_552;
  assign Queue_25_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_25_io_deq_ready = _T_550;
  assign Queue_25_clock = clock;
  assign Queue_25_reset = reset;
  assign Queue_26_io_enq_valid = _T_556;
  assign Queue_26_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_26_io_deq_ready = _T_554;
  assign Queue_26_clock = clock;
  assign Queue_26_reset = reset;
  assign Queue_27_io_enq_valid = _T_560;
  assign Queue_27_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_27_io_deq_ready = _T_558;
  assign Queue_27_clock = clock;
  assign Queue_27_reset = reset;
  assign Queue_28_io_enq_valid = _T_564;
  assign Queue_28_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_28_io_deq_ready = _T_562;
  assign Queue_28_clock = clock;
  assign Queue_28_reset = reset;
  assign Queue_29_io_enq_valid = _T_568;
  assign Queue_29_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_29_io_deq_ready = _T_566;
  assign Queue_29_clock = clock;
  assign Queue_29_reset = reset;
  assign Queue_30_io_enq_valid = _T_572;
  assign Queue_30_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_30_io_deq_ready = _T_570;
  assign Queue_30_clock = clock;
  assign Queue_30_reset = reset;
  assign Queue_31_io_enq_valid = _T_576;
  assign Queue_31_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_31_io_deq_ready = _T_574;
  assign Queue_31_clock = clock;
  assign Queue_31_reset = reset;
  assign _T_205_0 = Queue_io_enq_ready;
  assign _T_205_1 = Queue_1_io_enq_ready;
  assign _T_205_2 = Queue_2_io_enq_ready;
  assign _T_205_3 = Queue_3_io_enq_ready;
  assign _T_205_4 = Queue_4_io_enq_ready;
  assign _T_205_5 = Queue_5_io_enq_ready;
  assign _T_205_6 = Queue_6_io_enq_ready;
  assign _T_205_7 = Queue_7_io_enq_ready;
  assign _T_205_8 = Queue_8_io_enq_ready;
  assign _T_205_9 = Queue_9_io_enq_ready;
  assign _T_205_10 = Queue_10_io_enq_ready;
  assign _T_205_11 = Queue_11_io_enq_ready;
  assign _T_205_12 = Queue_12_io_enq_ready;
  assign _T_205_13 = Queue_13_io_enq_ready;
  assign _T_205_14 = Queue_14_io_enq_ready;
  assign _T_205_15 = Queue_15_io_enq_ready;
  assign _GEN_0 = _GEN_22;
  assign _GEN_1 = _GEN_22;
  assign _T_229_0 = Queue_io_deq_valid;
  assign _T_229_1 = Queue_1_io_deq_valid;
  assign _T_229_2 = Queue_2_io_deq_valid;
  assign _T_229_3 = Queue_3_io_deq_valid;
  assign _T_229_4 = Queue_4_io_deq_valid;
  assign _T_229_5 = Queue_5_io_deq_valid;
  assign _T_229_6 = Queue_6_io_deq_valid;
  assign _T_229_7 = Queue_7_io_deq_valid;
  assign _T_229_8 = Queue_8_io_deq_valid;
  assign _T_229_9 = Queue_9_io_deq_valid;
  assign _T_229_10 = Queue_10_io_deq_valid;
  assign _T_229_11 = Queue_11_io_deq_valid;
  assign _T_229_12 = Queue_12_io_deq_valid;
  assign _T_229_13 = Queue_13_io_deq_valid;
  assign _T_229_14 = Queue_14_io_deq_valid;
  assign _T_229_15 = Queue_15_io_deq_valid;
  assign _T_251_0 = Queue_io_deq_bits;
  assign _T_251_1 = Queue_1_io_deq_bits;
  assign _T_251_2 = Queue_2_io_deq_bits;
  assign _T_251_3 = Queue_3_io_deq_bits;
  assign _T_251_4 = Queue_4_io_deq_bits;
  assign _T_251_5 = Queue_5_io_deq_bits;
  assign _T_251_6 = Queue_6_io_deq_bits;
  assign _T_251_7 = Queue_7_io_deq_bits;
  assign _T_251_8 = Queue_8_io_deq_bits;
  assign _T_251_9 = Queue_9_io_deq_bits;
  assign _T_251_10 = Queue_10_io_deq_bits;
  assign _T_251_11 = Queue_11_io_deq_bits;
  assign _T_251_12 = Queue_12_io_deq_bits;
  assign _T_251_13 = Queue_13_io_deq_bits;
  assign _T_251_14 = Queue_14_io_deq_bits;
  assign _T_251_15 = Queue_15_io_deq_bits;
  assign _GEN_2 = _GEN_37;
  assign _GEN_3 = _GEN_52;
  assign _T_400_0 = Queue_16_io_enq_ready;
  assign _T_400_1 = Queue_17_io_enq_ready;
  assign _T_400_2 = Queue_18_io_enq_ready;
  assign _T_400_3 = Queue_19_io_enq_ready;
  assign _T_400_4 = Queue_20_io_enq_ready;
  assign _T_400_5 = Queue_21_io_enq_ready;
  assign _T_400_6 = Queue_22_io_enq_ready;
  assign _T_400_7 = Queue_23_io_enq_ready;
  assign _T_400_8 = Queue_24_io_enq_ready;
  assign _T_400_9 = Queue_25_io_enq_ready;
  assign _T_400_10 = Queue_26_io_enq_ready;
  assign _T_400_11 = Queue_27_io_enq_ready;
  assign _T_400_12 = Queue_28_io_enq_ready;
  assign _T_400_13 = Queue_29_io_enq_ready;
  assign _T_400_14 = Queue_30_io_enq_ready;
  assign _T_400_15 = Queue_31_io_enq_ready;
  assign _GEN_4 = _GEN_67;
  assign _GEN_5 = _GEN_67;
  assign _T_424_0 = Queue_16_io_deq_valid;
  assign _T_424_1 = Queue_17_io_deq_valid;
  assign _T_424_2 = Queue_18_io_deq_valid;
  assign _T_424_3 = Queue_19_io_deq_valid;
  assign _T_424_4 = Queue_20_io_deq_valid;
  assign _T_424_5 = Queue_21_io_deq_valid;
  assign _T_424_6 = Queue_22_io_deq_valid;
  assign _T_424_7 = Queue_23_io_deq_valid;
  assign _T_424_8 = Queue_24_io_deq_valid;
  assign _T_424_9 = Queue_25_io_deq_valid;
  assign _T_424_10 = Queue_26_io_deq_valid;
  assign _T_424_11 = Queue_27_io_deq_valid;
  assign _T_424_12 = Queue_28_io_deq_valid;
  assign _T_424_13 = Queue_29_io_deq_valid;
  assign _T_424_14 = Queue_30_io_deq_valid;
  assign _T_424_15 = Queue_31_io_deq_valid;
  assign _T_446_0 = Queue_16_io_deq_bits;
  assign _T_446_1 = Queue_17_io_deq_bits;
  assign _T_446_2 = Queue_18_io_deq_bits;
  assign _T_446_3 = Queue_19_io_deq_bits;
  assign _T_446_4 = Queue_20_io_deq_bits;
  assign _T_446_5 = Queue_21_io_deq_bits;
  assign _T_446_6 = Queue_22_io_deq_bits;
  assign _T_446_7 = Queue_23_io_deq_bits;
  assign _T_446_8 = Queue_24_io_deq_bits;
  assign _T_446_9 = Queue_25_io_deq_bits;
  assign _T_446_10 = Queue_26_io_deq_bits;
  assign _T_446_11 = Queue_27_io_deq_bits;
  assign _T_446_12 = Queue_28_io_deq_bits;
  assign _T_446_13 = Queue_29_io_deq_bits;
  assign _T_446_14 = Queue_30_io_deq_bits;
  assign _T_446_15 = Queue_31_io_deq_bits;
  assign _GEN_6 = _GEN_82;
  assign _GEN_7 = _GEN_97;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_277) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_472) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_472) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_66(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [31:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [31:0] ram_addr__T_50_data;
  wire  ram_addr__T_50_addr;
  wire [31:0] ram_addr__T_36_data;
  wire  ram_addr__T_36_addr;
  wire  ram_addr__T_36_mask;
  wire  ram_addr__T_36_en;
  reg [7:0] ram_len [0:1];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_50_data;
  wire  ram_len__T_50_addr;
  wire [7:0] ram_len__T_36_data;
  wire  ram_len__T_36_addr;
  wire  ram_len__T_36_mask;
  wire  ram_len__T_36_en;
  reg [2:0] ram_size [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [2:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [1:0] ram_burst [0:1];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_50_data;
  wire  ram_burst__T_50_addr;
  wire [1:0] ram_burst__T_36_data;
  wire  ram_burst__T_36_addr;
  wire  ram_burst__T_36_mask;
  wire  ram_burst__T_36_en;
  reg  ram_lock [0:1];
  reg [31:0] _RAND_5;
  wire  ram_lock__T_50_data;
  wire  ram_lock__T_50_addr;
  wire  ram_lock__T_36_data;
  wire  ram_lock__T_36_addr;
  wire  ram_lock__T_36_mask;
  wire  ram_lock__T_36_en;
  reg [3:0] ram_cache [0:1];
  reg [31:0] _RAND_6;
  wire [3:0] ram_cache__T_50_data;
  wire  ram_cache__T_50_addr;
  wire [3:0] ram_cache__T_36_data;
  wire  ram_cache__T_36_addr;
  wire  ram_cache__T_36_mask;
  wire  ram_cache__T_36_en;
  reg [2:0] ram_prot [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] ram_prot__T_50_data;
  wire  ram_prot__T_50_addr;
  wire [2:0] ram_prot__T_36_data;
  wire  ram_prot__T_36_addr;
  wire  ram_prot__T_36_mask;
  wire  ram_prot__T_36_en;
  reg [3:0] ram_qos [0:1];
  reg [31:0] _RAND_8;
  wire [3:0] ram_qos__T_50_data;
  wire  ram_qos__T_50_addr;
  wire [3:0] ram_qos__T_36_data;
  wire  ram_qos__T_36_addr;
  wire  ram_qos__T_36_mask;
  wire  ram_qos__T_36_en;
  reg  value;
  reg [31:0] _RAND_9;
  reg  value_1;
  reg [31:0] _RAND_10;
  reg  maybe_full;
  reg [31:0] _RAND_11;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_12;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_13;
  wire  _T_45;
  wire  _GEN_14;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_addr__T_50_addr = value_1;
  assign ram_addr__T_50_data = ram_addr[ram_addr__T_50_addr];
  assign ram_addr__T_36_data = io_enq_bits_addr;
  assign ram_addr__T_36_addr = value;
  assign ram_addr__T_36_mask = do_enq;
  assign ram_addr__T_36_en = do_enq;
  assign ram_len__T_50_addr = value_1;
  assign ram_len__T_50_data = ram_len[ram_len__T_50_addr];
  assign ram_len__T_36_data = io_enq_bits_len;
  assign ram_len__T_36_addr = value;
  assign ram_len__T_36_mask = do_enq;
  assign ram_len__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_burst__T_50_addr = value_1;
  assign ram_burst__T_50_data = ram_burst[ram_burst__T_50_addr];
  assign ram_burst__T_36_data = io_enq_bits_burst;
  assign ram_burst__T_36_addr = value;
  assign ram_burst__T_36_mask = do_enq;
  assign ram_burst__T_36_en = do_enq;
  assign ram_lock__T_50_addr = value_1;
  assign ram_lock__T_50_data = ram_lock[ram_lock__T_50_addr];
  assign ram_lock__T_36_data = io_enq_bits_lock;
  assign ram_lock__T_36_addr = value;
  assign ram_lock__T_36_mask = do_enq;
  assign ram_lock__T_36_en = do_enq;
  assign ram_cache__T_50_addr = value_1;
  assign ram_cache__T_50_data = ram_cache[ram_cache__T_50_addr];
  assign ram_cache__T_36_data = io_enq_bits_cache;
  assign ram_cache__T_36_addr = value;
  assign ram_cache__T_36_mask = do_enq;
  assign ram_cache__T_36_en = do_enq;
  assign ram_prot__T_50_addr = value_1;
  assign ram_prot__T_50_data = ram_prot[ram_prot__T_50_addr];
  assign ram_prot__T_36_data = io_enq_bits_prot;
  assign ram_prot__T_36_addr = value;
  assign ram_prot__T_36_mask = do_enq;
  assign ram_prot__T_36_en = do_enq;
  assign ram_qos__T_50_addr = value_1;
  assign ram_qos__T_50_data = ram_qos[ram_qos__T_50_addr];
  assign ram_qos__T_36_data = io_enq_bits_qos;
  assign ram_qos__T_36_addr = value;
  assign ram_qos__T_36_mask = do_enq;
  assign ram_qos__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_12 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_13 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_14 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_addr = ram_addr__T_50_data;
  assign io_deq_bits_len = ram_len__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_burst = ram_burst__T_50_data;
  assign io_deq_bits_lock = ram_lock__T_50_data;
  assign io_deq_bits_cache = ram_cache__T_50_data;
  assign io_deq_bits_prot = ram_prot__T_50_data;
  assign io_deq_bits_qos = ram_qos__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  value = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  value_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  maybe_full = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_addr__T_36_en & ram_addr__T_36_mask) begin
      ram_addr[ram_addr__T_36_addr] <= ram_addr__T_36_data;
    end
    if(ram_len__T_36_en & ram_len__T_36_mask) begin
      ram_len[ram_len__T_36_addr] <= ram_len__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_burst__T_36_en & ram_burst__T_36_mask) begin
      ram_burst[ram_burst__T_36_addr] <= ram_burst__T_36_data;
    end
    if(ram_lock__T_36_en & ram_lock__T_36_mask) begin
      ram_lock[ram_lock__T_36_addr] <= ram_lock__T_36_data;
    end
    if(ram_cache__T_36_en & ram_cache__T_36_mask) begin
      ram_cache[ram_cache__T_36_addr] <= ram_cache__T_36_data;
    end
    if(ram_prot__T_36_en & ram_prot__T_36_mask) begin
      ram_prot[ram_prot__T_36_addr] <= ram_prot__T_36_data;
    end
    if(ram_qos__T_36_en & ram_qos__T_36_mask) begin
      ram_qos[ram_qos__T_36_addr] <= ram_qos__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_67(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_0;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] _RAND_1;
  wire [7:0] ram_strb__T_50_data;
  wire  ram_strb__T_50_addr;
  wire [7:0] ram_strb__T_36_data;
  wire  ram_strb__T_36_addr;
  wire  ram_strb__T_36_mask;
  wire  ram_strb__T_36_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_2;
  wire  ram_last__T_50_data;
  wire  ram_last__T_50_addr;
  wire  ram_last__T_36_data;
  wire  ram_last__T_36_addr;
  wire  ram_last__T_36_mask;
  wire  ram_last__T_36_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_6;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_7;
  wire  _T_45;
  wire  _GEN_8;
  wire  _T_47;
  wire  _T_49;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign ram_strb__T_50_addr = value_1;
  assign ram_strb__T_50_data = ram_strb[ram_strb__T_50_addr];
  assign ram_strb__T_36_data = io_enq_bits_strb;
  assign ram_strb__T_36_addr = value;
  assign ram_strb__T_36_mask = do_enq;
  assign ram_strb__T_36_en = do_enq;
  assign ram_last__T_50_addr = value_1;
  assign ram_last__T_50_data = ram_last[ram_last__T_50_addr];
  assign ram_last__T_36_data = io_enq_bits_last;
  assign ram_last__T_36_addr = value;
  assign ram_last__T_36_mask = do_enq;
  assign ram_last__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_6 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_7 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_8 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign io_deq_bits_strb = ram_strb__T_50_data;
  assign io_deq_bits_last = ram_last__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if(ram_strb__T_36_en & ram_strb__T_36_mask) begin
      ram_strb[ram_strb__T_36_addr] <= ram_strb__T_36_data;
    end
    if(ram_last__T_36_en & ram_last__T_36_mask) begin
      ram_last[ram_last__T_36_addr] <= ram_last__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_68(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_resp__T_50_data;
  wire  ram_resp__T_50_addr;
  wire [1:0] ram_resp__T_36_data;
  wire  ram_resp__T_36_addr;
  wire  ram_resp__T_36_mask;
  wire  ram_resp__T_36_en;
  reg  value;
  reg [31:0] _RAND_2;
  reg  value_1;
  reg [31:0] _RAND_3;
  reg  maybe_full;
  reg [31:0] _RAND_4;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_5;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_6;
  wire  _T_45;
  wire  _GEN_7;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_resp__T_50_addr = value_1;
  assign ram_resp__T_50_data = ram_resp[ram_resp__T_50_addr];
  assign ram_resp__T_36_data = io_enq_bits_resp;
  assign ram_resp__T_36_addr = value;
  assign ram_resp__T_36_mask = do_enq;
  assign ram_resp__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_5 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_6 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_7 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_resp = ram_resp__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  maybe_full = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_resp__T_36_en & ram_resp__T_36_mask) begin
      ram_resp[ram_resp__T_36_addr] <= ram_resp__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_70(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_50_data;
  wire  ram_resp__T_50_addr;
  wire [1:0] ram_resp__T_36_data;
  wire  ram_resp__T_36_addr;
  wire  ram_resp__T_36_mask;
  wire  ram_resp__T_36_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_3;
  wire  ram_last__T_50_data;
  wire  ram_last__T_50_addr;
  wire  ram_last__T_36_data;
  wire  ram_last__T_36_addr;
  wire  ram_last__T_36_mask;
  wire  ram_last__T_36_en;
  reg  value;
  reg [31:0] _RAND_4;
  reg  value_1;
  reg [31:0] _RAND_5;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_7;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_8;
  wire  _T_45;
  wire  _GEN_9;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign ram_resp__T_50_addr = value_1;
  assign ram_resp__T_50_data = ram_resp[ram_resp__T_50_addr];
  assign ram_resp__T_36_data = io_enq_bits_resp;
  assign ram_resp__T_36_addr = value;
  assign ram_resp__T_36_mask = do_enq;
  assign ram_resp__T_36_en = do_enq;
  assign ram_last__T_50_addr = value_1;
  assign ram_last__T_50_data = ram_last[ram_last__T_50_addr];
  assign ram_last__T_36_data = io_enq_bits_last;
  assign ram_last__T_36_addr = value;
  assign ram_last__T_36_mask = do_enq;
  assign ram_last__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_7 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_8 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_9 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign io_deq_bits_resp = ram_resp__T_50_data;
  assign io_deq_bits_last = ram_last__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if(ram_resp__T_36_en & ram_resp__T_36_mask) begin
      ram_resp[ram_resp__T_36_addr] <= ram_resp__T_36_data;
    end
    if(ram_last__T_36_en & ram_last__T_36_mask) begin
      ram_last[ram_last__T_36_addr] <= ram_last__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Buffer_buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [31:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_enq_bits_lock;
  wire [3:0] Queue_io_enq_bits_cache;
  wire [2:0] Queue_io_enq_bits_prot;
  wire [3:0] Queue_io_enq_bits_qos;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [31:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  Queue_io_deq_bits_lock;
  wire [3:0] Queue_io_deq_bits_cache;
  wire [2:0] Queue_io_deq_bits_prot;
  wire [3:0] Queue_io_deq_bits_qos;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [31:0] _T_207_bits_addr;
  wire [7:0] _T_207_bits_len;
  wire [2:0] _T_207_bits_size;
  wire [1:0] _T_207_bits_burst;
  wire  _T_207_bits_lock;
  wire [3:0] _T_207_bits_cache;
  wire [2:0] _T_207_bits_prot;
  wire [3:0] _T_207_bits_qos;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_215_ready;
  wire  _T_215_valid;
  wire [63:0] _T_215_bits_data;
  wire [7:0] _T_215_bits_strb;
  wire  _T_215_bits_last;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  _T_223_ready;
  wire  _T_223_valid;
  wire [3:0] _T_223_bits_id;
  wire [1:0] _T_223_bits_resp;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [31:0] Queue_3_io_enq_bits_addr;
  wire [7:0] Queue_3_io_enq_bits_len;
  wire [2:0] Queue_3_io_enq_bits_size;
  wire [1:0] Queue_3_io_enq_bits_burst;
  wire  Queue_3_io_enq_bits_lock;
  wire [3:0] Queue_3_io_enq_bits_cache;
  wire [2:0] Queue_3_io_enq_bits_prot;
  wire [3:0] Queue_3_io_enq_bits_qos;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [31:0] Queue_3_io_deq_bits_addr;
  wire [7:0] Queue_3_io_deq_bits_len;
  wire [2:0] Queue_3_io_deq_bits_size;
  wire [1:0] Queue_3_io_deq_bits_burst;
  wire  Queue_3_io_deq_bits_lock;
  wire [3:0] Queue_3_io_deq_bits_cache;
  wire [2:0] Queue_3_io_deq_bits_prot;
  wire [3:0] Queue_3_io_deq_bits_qos;
  wire  _T_231_ready;
  wire  _T_231_valid;
  wire [3:0] _T_231_bits_id;
  wire [31:0] _T_231_bits_addr;
  wire [7:0] _T_231_bits_len;
  wire [2:0] _T_231_bits_size;
  wire [1:0] _T_231_bits_burst;
  wire  _T_231_bits_lock;
  wire [3:0] _T_231_bits_cache;
  wire [2:0] _T_231_bits_prot;
  wire [3:0] _T_231_bits_qos;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_last;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_239_ready;
  wire  _T_239_valid;
  wire [3:0] _T_239_bits_id;
  wire [63:0] _T_239_bits_data;
  wire [1:0] _T_239_bits_resp;
  wire  _T_239_bits_last;
  Queue_66 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_io_enq_bits_qos),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_io_deq_bits_qos)
  );
  Queue_67 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_68 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_66 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_len(Queue_3_io_enq_bits_len),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_burst(Queue_3_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_3_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_3_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_3_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_3_io_enq_bits_qos),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_len(Queue_3_io_deq_bits_len),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_burst(Queue_3_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_3_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_3_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_3_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_3_io_deq_bits_qos)
  );
  Queue_70 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_w_ready = Queue_1_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_223_valid;
  assign _T_31_b_bits_id = _T_223_bits_id;
  assign _T_31_b_bits_resp = _T_223_bits_resp;
  assign _T_31_ar_ready = Queue_3_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_239_valid;
  assign _T_31_r_bits_id = _T_239_bits_id;
  assign _T_31_r_bits_data = _T_239_bits_data;
  assign _T_31_r_bits_resp = _T_239_bits_resp;
  assign _T_31_r_bits_last = _T_239_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_207_valid;
  assign _T_89_aw_bits_id = _T_207_bits_id;
  assign _T_89_aw_bits_addr = _T_207_bits_addr;
  assign _T_89_aw_bits_len = _T_207_bits_len;
  assign _T_89_aw_bits_size = _T_207_bits_size;
  assign _T_89_aw_bits_burst = _T_207_bits_burst;
  assign _T_89_aw_bits_lock = _T_207_bits_lock;
  assign _T_89_aw_bits_cache = _T_207_bits_cache;
  assign _T_89_aw_bits_prot = _T_207_bits_prot;
  assign _T_89_aw_bits_qos = _T_207_bits_qos;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_215_valid;
  assign _T_89_w_bits_data = _T_215_bits_data;
  assign _T_89_w_bits_strb = _T_215_bits_strb;
  assign _T_89_w_bits_last = _T_215_bits_last;
  assign _T_89_b_ready = Queue_2_io_enq_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_231_valid;
  assign _T_89_ar_bits_id = _T_231_bits_id;
  assign _T_89_ar_bits_addr = _T_231_bits_addr;
  assign _T_89_ar_bits_len = _T_231_bits_len;
  assign _T_89_ar_bits_size = _T_231_bits_size;
  assign _T_89_ar_bits_burst = _T_231_bits_burst;
  assign _T_89_ar_bits_lock = _T_231_bits_lock;
  assign _T_89_ar_bits_cache = _T_231_bits_cache;
  assign _T_89_ar_bits_prot = _T_231_bits_prot;
  assign _T_89_ar_bits_qos = _T_231_bits_qos;
  assign _T_89_r_ready = Queue_4_io_enq_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_31_aw_valid;
  assign Queue_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_io_enq_bits_len = _T_31_aw_bits_len;
  assign Queue_io_enq_bits_size = _T_31_aw_bits_size;
  assign Queue_io_enq_bits_burst = _T_31_aw_bits_burst;
  assign Queue_io_enq_bits_lock = _T_31_aw_bits_lock;
  assign Queue_io_enq_bits_cache = _T_31_aw_bits_cache;
  assign Queue_io_enq_bits_prot = _T_31_aw_bits_prot;
  assign Queue_io_enq_bits_qos = _T_31_aw_bits_qos;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_89_aw_ready;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_len = Queue_io_deq_bits_len;
  assign _T_207_bits_size = Queue_io_deq_bits_size;
  assign _T_207_bits_burst = Queue_io_deq_bits_burst;
  assign _T_207_bits_lock = Queue_io_deq_bits_lock;
  assign _T_207_bits_cache = Queue_io_deq_bits_cache;
  assign _T_207_bits_prot = Queue_io_deq_bits_prot;
  assign _T_207_bits_qos = Queue_io_deq_bits_qos;
  assign Queue_1_io_enq_valid = _T_31_w_valid;
  assign Queue_1_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_1_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_1_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_1_io_deq_ready = _T_215_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_215_ready = _T_89_w_ready;
  assign _T_215_valid = Queue_1_io_deq_valid;
  assign _T_215_bits_data = Queue_1_io_deq_bits_data;
  assign _T_215_bits_strb = Queue_1_io_deq_bits_strb;
  assign _T_215_bits_last = Queue_1_io_deq_bits_last;
  assign Queue_2_io_enq_valid = _T_89_b_valid;
  assign Queue_2_io_enq_bits_id = _T_89_b_bits_id;
  assign Queue_2_io_enq_bits_resp = _T_89_b_bits_resp;
  assign Queue_2_io_deq_ready = _T_223_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_223_ready = _T_31_b_ready;
  assign _T_223_valid = Queue_2_io_deq_valid;
  assign _T_223_bits_id = Queue_2_io_deq_bits_id;
  assign _T_223_bits_resp = Queue_2_io_deq_bits_resp;
  assign Queue_3_io_enq_valid = _T_31_ar_valid;
  assign Queue_3_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_3_io_enq_bits_len = _T_31_ar_bits_len;
  assign Queue_3_io_enq_bits_size = _T_31_ar_bits_size;
  assign Queue_3_io_enq_bits_burst = _T_31_ar_bits_burst;
  assign Queue_3_io_enq_bits_lock = _T_31_ar_bits_lock;
  assign Queue_3_io_enq_bits_cache = _T_31_ar_bits_cache;
  assign Queue_3_io_enq_bits_prot = _T_31_ar_bits_prot;
  assign Queue_3_io_enq_bits_qos = _T_31_ar_bits_qos;
  assign Queue_3_io_deq_ready = _T_231_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign _T_231_ready = _T_89_ar_ready;
  assign _T_231_valid = Queue_3_io_deq_valid;
  assign _T_231_bits_id = Queue_3_io_deq_bits_id;
  assign _T_231_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_231_bits_len = Queue_3_io_deq_bits_len;
  assign _T_231_bits_size = Queue_3_io_deq_bits_size;
  assign _T_231_bits_burst = Queue_3_io_deq_bits_burst;
  assign _T_231_bits_lock = Queue_3_io_deq_bits_lock;
  assign _T_231_bits_cache = Queue_3_io_deq_bits_cache;
  assign _T_231_bits_prot = Queue_3_io_deq_bits_prot;
  assign _T_231_bits_qos = Queue_3_io_deq_bits_qos;
  assign Queue_4_io_enq_valid = _T_89_r_valid;
  assign Queue_4_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_4_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_4_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_4_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_4_io_deq_ready = _T_239_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign _T_239_ready = _T_31_r_ready;
  assign _T_239_valid = Queue_4_io_deq_valid;
  assign _T_239_bits_id = Queue_4_io_deq_bits_id;
  assign _T_239_bits_data = Queue_4_io_deq_bits_data;
  assign _T_239_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_239_bits_last = Queue_4_io_deq_bits_last;
endmodule
module Queue_71(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [30:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_enq_bits_lock,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_qos,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [30:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [30:0] ram_addr__T_50_data;
  wire  ram_addr__T_50_addr;
  wire [30:0] ram_addr__T_36_data;
  wire  ram_addr__T_36_addr;
  wire  ram_addr__T_36_mask;
  wire  ram_addr__T_36_en;
  reg [7:0] ram_len [0:1];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_50_data;
  wire  ram_len__T_50_addr;
  wire [7:0] ram_len__T_36_data;
  wire  ram_len__T_36_addr;
  wire  ram_len__T_36_mask;
  wire  ram_len__T_36_en;
  reg [2:0] ram_size [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_50_data;
  wire  ram_size__T_50_addr;
  wire [2:0] ram_size__T_36_data;
  wire  ram_size__T_36_addr;
  wire  ram_size__T_36_mask;
  wire  ram_size__T_36_en;
  reg [1:0] ram_burst [0:1];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_50_data;
  wire  ram_burst__T_50_addr;
  wire [1:0] ram_burst__T_36_data;
  wire  ram_burst__T_36_addr;
  wire  ram_burst__T_36_mask;
  wire  ram_burst__T_36_en;
  reg  ram_lock [0:1];
  reg [31:0] _RAND_5;
  wire  ram_lock__T_50_data;
  wire  ram_lock__T_50_addr;
  wire  ram_lock__T_36_data;
  wire  ram_lock__T_36_addr;
  wire  ram_lock__T_36_mask;
  wire  ram_lock__T_36_en;
  reg [3:0] ram_cache [0:1];
  reg [31:0] _RAND_6;
  wire [3:0] ram_cache__T_50_data;
  wire  ram_cache__T_50_addr;
  wire [3:0] ram_cache__T_36_data;
  wire  ram_cache__T_36_addr;
  wire  ram_cache__T_36_mask;
  wire  ram_cache__T_36_en;
  reg [2:0] ram_prot [0:1];
  reg [31:0] _RAND_7;
  wire [2:0] ram_prot__T_50_data;
  wire  ram_prot__T_50_addr;
  wire [2:0] ram_prot__T_36_data;
  wire  ram_prot__T_36_addr;
  wire  ram_prot__T_36_mask;
  wire  ram_prot__T_36_en;
  reg [3:0] ram_qos [0:1];
  reg [31:0] _RAND_8;
  wire [3:0] ram_qos__T_50_data;
  wire  ram_qos__T_50_addr;
  wire [3:0] ram_qos__T_36_data;
  wire  ram_qos__T_36_addr;
  wire  ram_qos__T_36_mask;
  wire  ram_qos__T_36_en;
  reg  value;
  reg [31:0] _RAND_9;
  reg  value_1;
  reg [31:0] _RAND_10;
  reg  maybe_full;
  reg [31:0] _RAND_11;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_12;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_13;
  wire  _T_45;
  wire  _GEN_14;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_addr__T_50_addr = value_1;
  assign ram_addr__T_50_data = ram_addr[ram_addr__T_50_addr];
  assign ram_addr__T_36_data = io_enq_bits_addr;
  assign ram_addr__T_36_addr = value;
  assign ram_addr__T_36_mask = do_enq;
  assign ram_addr__T_36_en = do_enq;
  assign ram_len__T_50_addr = value_1;
  assign ram_len__T_50_data = ram_len[ram_len__T_50_addr];
  assign ram_len__T_36_data = io_enq_bits_len;
  assign ram_len__T_36_addr = value;
  assign ram_len__T_36_mask = do_enq;
  assign ram_len__T_36_en = do_enq;
  assign ram_size__T_50_addr = value_1;
  assign ram_size__T_50_data = ram_size[ram_size__T_50_addr];
  assign ram_size__T_36_data = io_enq_bits_size;
  assign ram_size__T_36_addr = value;
  assign ram_size__T_36_mask = do_enq;
  assign ram_size__T_36_en = do_enq;
  assign ram_burst__T_50_addr = value_1;
  assign ram_burst__T_50_data = ram_burst[ram_burst__T_50_addr];
  assign ram_burst__T_36_data = io_enq_bits_burst;
  assign ram_burst__T_36_addr = value;
  assign ram_burst__T_36_mask = do_enq;
  assign ram_burst__T_36_en = do_enq;
  assign ram_lock__T_50_addr = value_1;
  assign ram_lock__T_50_data = ram_lock[ram_lock__T_50_addr];
  assign ram_lock__T_36_data = io_enq_bits_lock;
  assign ram_lock__T_36_addr = value;
  assign ram_lock__T_36_mask = do_enq;
  assign ram_lock__T_36_en = do_enq;
  assign ram_cache__T_50_addr = value_1;
  assign ram_cache__T_50_data = ram_cache[ram_cache__T_50_addr];
  assign ram_cache__T_36_data = io_enq_bits_cache;
  assign ram_cache__T_36_addr = value;
  assign ram_cache__T_36_mask = do_enq;
  assign ram_cache__T_36_en = do_enq;
  assign ram_prot__T_50_addr = value_1;
  assign ram_prot__T_50_data = ram_prot[ram_prot__T_50_addr];
  assign ram_prot__T_36_data = io_enq_bits_prot;
  assign ram_prot__T_36_addr = value;
  assign ram_prot__T_36_mask = do_enq;
  assign ram_prot__T_36_en = do_enq;
  assign ram_qos__T_50_addr = value_1;
  assign ram_qos__T_50_data = ram_qos[ram_qos__T_50_addr];
  assign ram_qos__T_36_data = io_enq_bits_qos;
  assign ram_qos__T_36_addr = value;
  assign ram_qos__T_36_mask = do_enq;
  assign ram_qos__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_12 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_13 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_14 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_addr = ram_addr__T_50_data;
  assign io_deq_bits_len = ram_len__T_50_data;
  assign io_deq_bits_size = ram_size__T_50_data;
  assign io_deq_bits_burst = ram_burst__T_50_data;
  assign io_deq_bits_lock = ram_lock__T_50_data;
  assign io_deq_bits_cache = ram_cache__T_50_data;
  assign io_deq_bits_prot = ram_prot__T_50_data;
  assign io_deq_bits_qos = ram_qos__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  value = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  value_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  maybe_full = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_addr__T_36_en & ram_addr__T_36_mask) begin
      ram_addr[ram_addr__T_36_addr] <= ram_addr__T_36_data;
    end
    if(ram_len__T_36_en & ram_len__T_36_mask) begin
      ram_len[ram_len__T_36_addr] <= ram_len__T_36_data;
    end
    if(ram_size__T_36_en & ram_size__T_36_mask) begin
      ram_size[ram_size__T_36_addr] <= ram_size__T_36_data;
    end
    if(ram_burst__T_36_en & ram_burst__T_36_mask) begin
      ram_burst[ram_burst__T_36_addr] <= ram_burst__T_36_data;
    end
    if(ram_lock__T_36_en & ram_lock__T_36_mask) begin
      ram_lock[ram_lock__T_36_addr] <= ram_lock__T_36_data;
    end
    if(ram_cache__T_36_en & ram_cache__T_36_mask) begin
      ram_cache[ram_cache__T_36_addr] <= ram_cache__T_36_data;
    end
    if(ram_prot__T_36_en & ram_prot__T_36_mask) begin
      ram_prot[ram_prot__T_36_addr] <= ram_prot__T_36_data;
    end
    if(ram_qos__T_36_en & ram_qos__T_36_mask) begin
      ram_qos[ram_qos__T_36_addr] <= ram_qos__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [30:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [30:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [30:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [30:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [30:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [30:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [30:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_enq_bits_lock;
  wire [3:0] Queue_io_enq_bits_cache;
  wire [2:0] Queue_io_enq_bits_prot;
  wire [3:0] Queue_io_enq_bits_qos;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [30:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  Queue_io_deq_bits_lock;
  wire [3:0] Queue_io_deq_bits_cache;
  wire [2:0] Queue_io_deq_bits_prot;
  wire [3:0] Queue_io_deq_bits_qos;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [30:0] _T_207_bits_addr;
  wire [7:0] _T_207_bits_len;
  wire [2:0] _T_207_bits_size;
  wire [1:0] _T_207_bits_burst;
  wire  _T_207_bits_lock;
  wire [3:0] _T_207_bits_cache;
  wire [2:0] _T_207_bits_prot;
  wire [3:0] _T_207_bits_qos;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_215_ready;
  wire  _T_215_valid;
  wire [63:0] _T_215_bits_data;
  wire [7:0] _T_215_bits_strb;
  wire  _T_215_bits_last;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  _T_223_ready;
  wire  _T_223_valid;
  wire [3:0] _T_223_bits_id;
  wire [1:0] _T_223_bits_resp;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [30:0] Queue_3_io_enq_bits_addr;
  wire [7:0] Queue_3_io_enq_bits_len;
  wire [2:0] Queue_3_io_enq_bits_size;
  wire [1:0] Queue_3_io_enq_bits_burst;
  wire  Queue_3_io_enq_bits_lock;
  wire [3:0] Queue_3_io_enq_bits_cache;
  wire [2:0] Queue_3_io_enq_bits_prot;
  wire [3:0] Queue_3_io_enq_bits_qos;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [30:0] Queue_3_io_deq_bits_addr;
  wire [7:0] Queue_3_io_deq_bits_len;
  wire [2:0] Queue_3_io_deq_bits_size;
  wire [1:0] Queue_3_io_deq_bits_burst;
  wire  Queue_3_io_deq_bits_lock;
  wire [3:0] Queue_3_io_deq_bits_cache;
  wire [2:0] Queue_3_io_deq_bits_prot;
  wire [3:0] Queue_3_io_deq_bits_qos;
  wire  _T_231_ready;
  wire  _T_231_valid;
  wire [3:0] _T_231_bits_id;
  wire [30:0] _T_231_bits_addr;
  wire [7:0] _T_231_bits_len;
  wire [2:0] _T_231_bits_size;
  wire [1:0] _T_231_bits_burst;
  wire  _T_231_bits_lock;
  wire [3:0] _T_231_bits_cache;
  wire [2:0] _T_231_bits_prot;
  wire [3:0] _T_231_bits_qos;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_last;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_239_ready;
  wire  _T_239_valid;
  wire [3:0] _T_239_bits_id;
  wire [63:0] _T_239_bits_data;
  wire [1:0] _T_239_bits_resp;
  wire  _T_239_bits_last;
  Queue_71 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_io_enq_bits_qos),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_io_deq_bits_qos)
  );
  Queue_67 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_68 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_71 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_len(Queue_3_io_enq_bits_len),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_burst(Queue_3_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_3_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_3_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_3_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_3_io_enq_bits_qos),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_len(Queue_3_io_deq_bits_len),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_burst(Queue_3_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_3_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_3_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_3_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_3_io_deq_bits_qos)
  );
  Queue_70 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_w_ready = Queue_1_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_223_valid;
  assign _T_31_b_bits_id = _T_223_bits_id;
  assign _T_31_b_bits_resp = _T_223_bits_resp;
  assign _T_31_ar_ready = Queue_3_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_239_valid;
  assign _T_31_r_bits_id = _T_239_bits_id;
  assign _T_31_r_bits_data = _T_239_bits_data;
  assign _T_31_r_bits_resp = _T_239_bits_resp;
  assign _T_31_r_bits_last = _T_239_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_207_valid;
  assign _T_89_aw_bits_id = _T_207_bits_id;
  assign _T_89_aw_bits_addr = _T_207_bits_addr;
  assign _T_89_aw_bits_len = _T_207_bits_len;
  assign _T_89_aw_bits_size = _T_207_bits_size;
  assign _T_89_aw_bits_burst = _T_207_bits_burst;
  assign _T_89_aw_bits_lock = _T_207_bits_lock;
  assign _T_89_aw_bits_cache = _T_207_bits_cache;
  assign _T_89_aw_bits_prot = _T_207_bits_prot;
  assign _T_89_aw_bits_qos = _T_207_bits_qos;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_215_valid;
  assign _T_89_w_bits_data = _T_215_bits_data;
  assign _T_89_w_bits_strb = _T_215_bits_strb;
  assign _T_89_w_bits_last = _T_215_bits_last;
  assign _T_89_b_ready = Queue_2_io_enq_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_231_valid;
  assign _T_89_ar_bits_id = _T_231_bits_id;
  assign _T_89_ar_bits_addr = _T_231_bits_addr;
  assign _T_89_ar_bits_len = _T_231_bits_len;
  assign _T_89_ar_bits_size = _T_231_bits_size;
  assign _T_89_ar_bits_burst = _T_231_bits_burst;
  assign _T_89_ar_bits_lock = _T_231_bits_lock;
  assign _T_89_ar_bits_cache = _T_231_bits_cache;
  assign _T_89_ar_bits_prot = _T_231_bits_prot;
  assign _T_89_ar_bits_qos = _T_231_bits_qos;
  assign _T_89_r_ready = Queue_4_io_enq_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_31_aw_valid;
  assign Queue_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_io_enq_bits_len = _T_31_aw_bits_len;
  assign Queue_io_enq_bits_size = _T_31_aw_bits_size;
  assign Queue_io_enq_bits_burst = _T_31_aw_bits_burst;
  assign Queue_io_enq_bits_lock = _T_31_aw_bits_lock;
  assign Queue_io_enq_bits_cache = _T_31_aw_bits_cache;
  assign Queue_io_enq_bits_prot = _T_31_aw_bits_prot;
  assign Queue_io_enq_bits_qos = _T_31_aw_bits_qos;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_89_aw_ready;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_len = Queue_io_deq_bits_len;
  assign _T_207_bits_size = Queue_io_deq_bits_size;
  assign _T_207_bits_burst = Queue_io_deq_bits_burst;
  assign _T_207_bits_lock = Queue_io_deq_bits_lock;
  assign _T_207_bits_cache = Queue_io_deq_bits_cache;
  assign _T_207_bits_prot = Queue_io_deq_bits_prot;
  assign _T_207_bits_qos = Queue_io_deq_bits_qos;
  assign Queue_1_io_enq_valid = _T_31_w_valid;
  assign Queue_1_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_1_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_1_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_1_io_deq_ready = _T_215_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_215_ready = _T_89_w_ready;
  assign _T_215_valid = Queue_1_io_deq_valid;
  assign _T_215_bits_data = Queue_1_io_deq_bits_data;
  assign _T_215_bits_strb = Queue_1_io_deq_bits_strb;
  assign _T_215_bits_last = Queue_1_io_deq_bits_last;
  assign Queue_2_io_enq_valid = _T_89_b_valid;
  assign Queue_2_io_enq_bits_id = _T_89_b_bits_id;
  assign Queue_2_io_enq_bits_resp = _T_89_b_bits_resp;
  assign Queue_2_io_deq_ready = _T_223_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_223_ready = _T_31_b_ready;
  assign _T_223_valid = Queue_2_io_deq_valid;
  assign _T_223_bits_id = Queue_2_io_deq_bits_id;
  assign _T_223_bits_resp = Queue_2_io_deq_bits_resp;
  assign Queue_3_io_enq_valid = _T_31_ar_valid;
  assign Queue_3_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_3_io_enq_bits_len = _T_31_ar_bits_len;
  assign Queue_3_io_enq_bits_size = _T_31_ar_bits_size;
  assign Queue_3_io_enq_bits_burst = _T_31_ar_bits_burst;
  assign Queue_3_io_enq_bits_lock = _T_31_ar_bits_lock;
  assign Queue_3_io_enq_bits_cache = _T_31_ar_bits_cache;
  assign Queue_3_io_enq_bits_prot = _T_31_ar_bits_prot;
  assign Queue_3_io_enq_bits_qos = _T_31_ar_bits_qos;
  assign Queue_3_io_deq_ready = _T_231_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign _T_231_ready = _T_89_ar_ready;
  assign _T_231_valid = Queue_3_io_deq_valid;
  assign _T_231_bits_id = Queue_3_io_deq_bits_id;
  assign _T_231_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_231_bits_len = Queue_3_io_deq_bits_len;
  assign _T_231_bits_size = Queue_3_io_deq_bits_size;
  assign _T_231_bits_burst = Queue_3_io_deq_bits_burst;
  assign _T_231_bits_lock = Queue_3_io_deq_bits_lock;
  assign _T_231_bits_cache = Queue_3_io_deq_bits_cache;
  assign _T_231_bits_prot = Queue_3_io_deq_bits_prot;
  assign _T_231_bits_qos = Queue_3_io_deq_bits_qos;
  assign Queue_4_io_enq_valid = _T_89_r_valid;
  assign Queue_4_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_4_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_4_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_4_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_4_io_deq_ready = _T_239_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign _T_239_ready = _T_31_r_ready;
  assign _T_239_valid = Queue_4_io_deq_valid;
  assign _T_239_bits_id = Queue_4_io_deq_bits_id;
  assign _T_239_bits_data = Queue_4_io_deq_bits_data;
  assign _T_239_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_239_bits_last = Queue_4_io_deq_bits_last;
endmodule
module Queue_76(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [8:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [8:0] io_deq_bits
);
  reg [8:0] ram [0:0];
  reg [31:0] _RAND_0;
  wire [8:0] ram__T_42_data;
  wire  ram__T_42_addr;
  wire [8:0] ram__T_33_data;
  wire  ram__T_33_addr;
  wire  ram__T_33_mask;
  wire  ram__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_1;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_4;
  wire  _T_38;
  assign ram__T_42_addr = 1'h0;
  assign ram__T_42_data = ram[ram__T_42_addr];
  assign ram__T_33_data = io_enq_bits;
  assign ram__T_33_addr = 1'h0;
  assign ram__T_33_mask = do_enq;
  assign ram__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_4 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign io_enq_ready = empty;
  assign io_deq_valid = _T_38;
  assign io_deq_bits = ram__T_42_data;
  assign do_enq = _T_28;
  assign do_deq = _T_30;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[8:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  maybe_full = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_33_en & ram__T_33_mask) begin
      ram[ram__T_33_addr] <= ram__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_77(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [8:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [8:0] io_deq_bits
);
  reg [8:0] ram [0:7];
  reg [31:0] _RAND_0;
  wire [8:0] ram__T_50_data;
  wire [2:0] ram__T_50_addr;
  wire [8:0] ram__T_36_data;
  wire [2:0] ram__T_36_addr;
  wire  ram__T_36_mask;
  wire  ram__T_36_en;
  reg [2:0] value;
  reg [31:0] _RAND_1;
  reg [2:0] value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [3:0] _T_39;
  wire [2:0] _T_40;
  wire [2:0] _GEN_4;
  wire [3:0] _T_43;
  wire [2:0] _T_44;
  wire [2:0] _GEN_5;
  wire  _T_45;
  wire  _GEN_6;
  wire  _T_47;
  wire  _T_49;
  assign ram__T_50_addr = value_1;
  assign ram__T_50_data = ram[ram__T_50_addr];
  assign ram__T_36_data = io_enq_bits;
  assign ram__T_36_addr = value;
  assign ram__T_36_mask = do_enq;
  assign ram__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 3'h1;
  assign _T_40 = _T_39[2:0];
  assign _GEN_4 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 3'h1;
  assign _T_44 = _T_43[2:0];
  assign _GEN_5 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_6 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits = ram__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[8:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_36_en & ram__T_36_mask) begin
      ram[ram__T_36_addr] <= ram__T_36_data;
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4UserYanker(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [30:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [8:0]  auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [8:0]  auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [30:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [8:0]  auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [8:0]  auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [30:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire [8:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [8:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [30:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire [8:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [8:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [30:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [30:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [8:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [8:0] Queue_io_deq_bits;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [8:0] Queue_1_io_enq_bits;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [8:0] Queue_1_io_deq_bits;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [8:0] Queue_2_io_enq_bits;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [8:0] Queue_2_io_deq_bits;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [8:0] Queue_3_io_enq_bits;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [8:0] Queue_3_io_deq_bits;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [8:0] Queue_4_io_enq_bits;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [8:0] Queue_4_io_deq_bits;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [8:0] Queue_5_io_enq_bits;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [8:0] Queue_5_io_deq_bits;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [8:0] Queue_6_io_enq_bits;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [8:0] Queue_6_io_deq_bits;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [8:0] Queue_7_io_enq_bits;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [8:0] Queue_7_io_deq_bits;
  wire  Queue_8_clock;
  wire  Queue_8_reset;
  wire  Queue_8_io_enq_ready;
  wire  Queue_8_io_enq_valid;
  wire [8:0] Queue_8_io_enq_bits;
  wire  Queue_8_io_deq_ready;
  wire  Queue_8_io_deq_valid;
  wire [8:0] Queue_8_io_deq_bits;
  wire  Queue_9_clock;
  wire  Queue_9_reset;
  wire  Queue_9_io_enq_ready;
  wire  Queue_9_io_enq_valid;
  wire [8:0] Queue_9_io_enq_bits;
  wire  Queue_9_io_deq_ready;
  wire  Queue_9_io_deq_valid;
  wire [8:0] Queue_9_io_deq_bits;
  wire  Queue_10_clock;
  wire  Queue_10_reset;
  wire  Queue_10_io_enq_ready;
  wire  Queue_10_io_enq_valid;
  wire [8:0] Queue_10_io_enq_bits;
  wire  Queue_10_io_deq_ready;
  wire  Queue_10_io_deq_valid;
  wire [8:0] Queue_10_io_deq_bits;
  wire  Queue_11_clock;
  wire  Queue_11_reset;
  wire  Queue_11_io_enq_ready;
  wire  Queue_11_io_enq_valid;
  wire [8:0] Queue_11_io_enq_bits;
  wire  Queue_11_io_deq_ready;
  wire  Queue_11_io_deq_valid;
  wire [8:0] Queue_11_io_deq_bits;
  wire  Queue_12_clock;
  wire  Queue_12_reset;
  wire  Queue_12_io_enq_ready;
  wire  Queue_12_io_enq_valid;
  wire [8:0] Queue_12_io_enq_bits;
  wire  Queue_12_io_deq_ready;
  wire  Queue_12_io_deq_valid;
  wire [8:0] Queue_12_io_deq_bits;
  wire  Queue_13_clock;
  wire  Queue_13_reset;
  wire  Queue_13_io_enq_ready;
  wire  Queue_13_io_enq_valid;
  wire [8:0] Queue_13_io_enq_bits;
  wire  Queue_13_io_deq_ready;
  wire  Queue_13_io_deq_valid;
  wire [8:0] Queue_13_io_deq_bits;
  wire  Queue_14_clock;
  wire  Queue_14_reset;
  wire  Queue_14_io_enq_ready;
  wire  Queue_14_io_enq_valid;
  wire [8:0] Queue_14_io_enq_bits;
  wire  Queue_14_io_deq_ready;
  wire  Queue_14_io_deq_valid;
  wire [8:0] Queue_14_io_deq_bits;
  wire  Queue_15_clock;
  wire  Queue_15_reset;
  wire  Queue_15_io_enq_ready;
  wire  Queue_15_io_enq_valid;
  wire [8:0] Queue_15_io_enq_bits;
  wire  Queue_15_io_deq_ready;
  wire  Queue_15_io_deq_valid;
  wire [8:0] Queue_15_io_deq_bits;
  wire  _T_861_0;
  wire  _T_861_1;
  wire  _T_861_2;
  wire  _T_861_3;
  wire  _T_861_4;
  wire  _T_861_5;
  wire  _T_861_6;
  wire  _T_861_7;
  wire  _GEN_0;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _T_881;
  wire  _GEN_1;
  wire  _T_882;
  wire  _T_885_0;
  wire  _T_885_1;
  wire  _T_885_2;
  wire  _T_885_3;
  wire  _T_885_4;
  wire  _T_885_5;
  wire  _T_885_6;
  wire  _T_885_7;
  wire [8:0] _T_907_0;
  wire [8:0] _T_907_1;
  wire [8:0] _T_907_2;
  wire [8:0] _T_907_3;
  wire [8:0] _T_907_4;
  wire [8:0] _T_907_5;
  wire [8:0] _T_907_6;
  wire [8:0] _T_907_7;
  wire  _T_928;
  wire  _GEN_2;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _T_929;
  wire  _T_931;
  wire  _T_933;
  wire [8:0] _GEN_3;
  wire [8:0] _GEN_38;
  wire [8:0] _GEN_39;
  wire [8:0] _GEN_40;
  wire [8:0] _GEN_41;
  wire [8:0] _GEN_42;
  wire [8:0] _GEN_43;
  wire [8:0] _GEN_44;
  wire [8:0] _GEN_45;
  wire [8:0] _GEN_46;
  wire [8:0] _GEN_47;
  wire [8:0] _GEN_48;
  wire [8:0] _GEN_49;
  wire [8:0] _GEN_50;
  wire [8:0] _GEN_51;
  wire [8:0] _GEN_52;
  wire [15:0] _T_936;
  wire  _T_938;
  wire  _T_939;
  wire  _T_940;
  wire  _T_941;
  wire  _T_942;
  wire  _T_943;
  wire  _T_944;
  wire  _T_945;
  wire [15:0] _T_956;
  wire  _T_958;
  wire  _T_959;
  wire  _T_960;
  wire  _T_961;
  wire  _T_962;
  wire  _T_963;
  wire  _T_964;
  wire  _T_965;
  wire  _T_974;
  wire  _T_975;
  wire  _T_976;
  wire  _T_977;
  wire  _T_978;
  wire  _T_980;
  wire  _T_981;
  wire  _T_983;
  wire  _T_985;
  wire  _T_986;
  wire  _T_988;
  wire  _T_990;
  wire  _T_991;
  wire  _T_993;
  wire  _T_995;
  wire  _T_996;
  wire  _T_998;
  wire  _T_1000;
  wire  _T_1001;
  wire  _T_1003;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1008;
  wire  _T_1010;
  wire  _T_1011;
  wire  _T_1013;
  wire  _T_1056_0;
  wire  _T_1056_1;
  wire  _T_1056_2;
  wire  _T_1056_3;
  wire  _T_1056_4;
  wire  _T_1056_5;
  wire  _T_1056_6;
  wire  _T_1056_7;
  wire  _GEN_4;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _T_1076;
  wire  _GEN_5;
  wire  _T_1077;
  wire  _T_1080_0;
  wire  _T_1080_1;
  wire  _T_1080_2;
  wire  _T_1080_3;
  wire  _T_1080_4;
  wire  _T_1080_5;
  wire  _T_1080_6;
  wire  _T_1080_7;
  wire [8:0] _T_1102_0;
  wire [8:0] _T_1102_1;
  wire [8:0] _T_1102_2;
  wire [8:0] _T_1102_3;
  wire [8:0] _T_1102_4;
  wire [8:0] _T_1102_5;
  wire [8:0] _T_1102_6;
  wire [8:0] _T_1102_7;
  wire  _T_1123;
  wire  _GEN_6;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _T_1124;
  wire  _T_1126;
  wire  _T_1128;
  wire [8:0] _GEN_7;
  wire [8:0] _GEN_83;
  wire [8:0] _GEN_84;
  wire [8:0] _GEN_85;
  wire [8:0] _GEN_86;
  wire [8:0] _GEN_87;
  wire [8:0] _GEN_88;
  wire [8:0] _GEN_89;
  wire [8:0] _GEN_90;
  wire [8:0] _GEN_91;
  wire [8:0] _GEN_92;
  wire [8:0] _GEN_93;
  wire [8:0] _GEN_94;
  wire [8:0] _GEN_95;
  wire [8:0] _GEN_96;
  wire [8:0] _GEN_97;
  wire [15:0] _T_1131;
  wire  _T_1133;
  wire  _T_1134;
  wire  _T_1135;
  wire  _T_1136;
  wire  _T_1137;
  wire  _T_1138;
  wire  _T_1139;
  wire  _T_1140;
  wire [15:0] _T_1151;
  wire  _T_1153;
  wire  _T_1154;
  wire  _T_1155;
  wire  _T_1156;
  wire  _T_1157;
  wire  _T_1158;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1169;
  wire  _T_1170;
  wire  _T_1171;
  wire  _T_1172;
  wire  _T_1174;
  wire  _T_1176;
  wire  _T_1178;
  wire  _T_1180;
  wire  _T_1182;
  wire  _T_1184;
  wire  _T_1186;
  wire  _T_1188;
  wire  _T_1190;
  wire  _T_1192;
  wire  _T_1194;
  wire  _T_1196;
  wire  _T_1198;
  wire  _T_1200;
  Queue_76 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_77 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_77 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_76 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  Queue_76 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_76 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  Queue_76 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  Queue_76 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  Queue_76 Queue_8 (
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits(Queue_8_io_enq_bits),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits(Queue_8_io_deq_bits)
  );
  Queue_77 Queue_9 (
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits(Queue_9_io_enq_bits),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits(Queue_9_io_deq_bits)
  );
  Queue_77 Queue_10 (
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  Queue_76 Queue_11 (
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits(Queue_11_io_enq_bits),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits(Queue_11_io_deq_bits)
  );
  Queue_76 Queue_12 (
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits(Queue_12_io_enq_bits),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits(Queue_12_io_deq_bits)
  );
  Queue_76 Queue_13 (
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits(Queue_13_io_enq_bits),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits(Queue_13_io_deq_bits)
  );
  Queue_76 Queue_14 (
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits(Queue_14_io_enq_bits),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits(Queue_14_io_deq_bits)
  );
  Queue_76 Queue_15 (
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits(Queue_15_io_enq_bits),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits(Queue_15_io_deq_bits)
  );
  assign _GEN_8 = 4'h1 == _T_31_ar_bits_id ? _T_861_1 : _T_861_0;
  assign _GEN_9 = 4'h2 == _T_31_ar_bits_id ? _T_861_2 : _GEN_8;
  assign _GEN_10 = 4'h3 == _T_31_ar_bits_id ? _T_861_3 : _GEN_9;
  assign _GEN_11 = 4'h4 == _T_31_ar_bits_id ? _T_861_4 : _GEN_10;
  assign _GEN_12 = 4'h5 == _T_31_ar_bits_id ? _T_861_5 : _GEN_11;
  assign _GEN_13 = 4'h6 == _T_31_ar_bits_id ? _T_861_6 : _GEN_12;
  assign _GEN_14 = 4'h7 == _T_31_ar_bits_id ? _T_861_7 : _GEN_13;
  assign _GEN_15 = 4'h8 == _T_31_ar_bits_id ? 1'h0 : _GEN_14;
  assign _GEN_16 = 4'h9 == _T_31_ar_bits_id ? 1'h0 : _GEN_15;
  assign _GEN_17 = 4'ha == _T_31_ar_bits_id ? 1'h0 : _GEN_16;
  assign _GEN_18 = 4'hb == _T_31_ar_bits_id ? 1'h0 : _GEN_17;
  assign _GEN_19 = 4'hc == _T_31_ar_bits_id ? 1'h0 : _GEN_18;
  assign _GEN_20 = 4'hd == _T_31_ar_bits_id ? 1'h0 : _GEN_19;
  assign _GEN_21 = 4'he == _T_31_ar_bits_id ? 1'h0 : _GEN_20;
  assign _GEN_22 = 4'hf == _T_31_ar_bits_id ? 1'h0 : _GEN_21;
  assign _T_881 = _T_89_ar_ready & _GEN_0;
  assign _T_882 = _T_31_ar_valid & _GEN_1;
  assign _T_928 = _T_89_r_valid == 1'h0;
  assign _GEN_23 = 4'h1 == _T_89_r_bits_id ? _T_885_1 : _T_885_0;
  assign _GEN_24 = 4'h2 == _T_89_r_bits_id ? _T_885_2 : _GEN_23;
  assign _GEN_25 = 4'h3 == _T_89_r_bits_id ? _T_885_3 : _GEN_24;
  assign _GEN_26 = 4'h4 == _T_89_r_bits_id ? _T_885_4 : _GEN_25;
  assign _GEN_27 = 4'h5 == _T_89_r_bits_id ? _T_885_5 : _GEN_26;
  assign _GEN_28 = 4'h6 == _T_89_r_bits_id ? _T_885_6 : _GEN_27;
  assign _GEN_29 = 4'h7 == _T_89_r_bits_id ? _T_885_7 : _GEN_28;
  assign _GEN_30 = 4'h8 == _T_89_r_bits_id ? 1'h0 : _GEN_29;
  assign _GEN_31 = 4'h9 == _T_89_r_bits_id ? 1'h0 : _GEN_30;
  assign _GEN_32 = 4'ha == _T_89_r_bits_id ? 1'h0 : _GEN_31;
  assign _GEN_33 = 4'hb == _T_89_r_bits_id ? 1'h0 : _GEN_32;
  assign _GEN_34 = 4'hc == _T_89_r_bits_id ? 1'h0 : _GEN_33;
  assign _GEN_35 = 4'hd == _T_89_r_bits_id ? 1'h0 : _GEN_34;
  assign _GEN_36 = 4'he == _T_89_r_bits_id ? 1'h0 : _GEN_35;
  assign _GEN_37 = 4'hf == _T_89_r_bits_id ? 1'h0 : _GEN_36;
  assign _T_929 = _T_928 | _GEN_2;
  assign _T_931 = _T_929 | reset;
  assign _T_933 = _T_931 == 1'h0;
  assign _GEN_38 = 4'h1 == _T_89_r_bits_id ? _T_907_1 : _T_907_0;
  assign _GEN_39 = 4'h2 == _T_89_r_bits_id ? _T_907_2 : _GEN_38;
  assign _GEN_40 = 4'h3 == _T_89_r_bits_id ? _T_907_3 : _GEN_39;
  assign _GEN_41 = 4'h4 == _T_89_r_bits_id ? _T_907_4 : _GEN_40;
  assign _GEN_42 = 4'h5 == _T_89_r_bits_id ? _T_907_5 : _GEN_41;
  assign _GEN_43 = 4'h6 == _T_89_r_bits_id ? _T_907_6 : _GEN_42;
  assign _GEN_44 = 4'h7 == _T_89_r_bits_id ? _T_907_7 : _GEN_43;
  assign _GEN_45 = 4'h8 == _T_89_r_bits_id ? 9'h0 : _GEN_44;
  assign _GEN_46 = 4'h9 == _T_89_r_bits_id ? 9'h0 : _GEN_45;
  assign _GEN_47 = 4'ha == _T_89_r_bits_id ? 9'h0 : _GEN_46;
  assign _GEN_48 = 4'hb == _T_89_r_bits_id ? 9'h0 : _GEN_47;
  assign _GEN_49 = 4'hc == _T_89_r_bits_id ? 9'h0 : _GEN_48;
  assign _GEN_50 = 4'hd == _T_89_r_bits_id ? 9'h0 : _GEN_49;
  assign _GEN_51 = 4'he == _T_89_r_bits_id ? 9'h0 : _GEN_50;
  assign _GEN_52 = 4'hf == _T_89_r_bits_id ? 9'h0 : _GEN_51;
  assign _T_936 = 16'h1 << _T_31_ar_bits_id;
  assign _T_938 = _T_936[0];
  assign _T_939 = _T_936[1];
  assign _T_940 = _T_936[2];
  assign _T_941 = _T_936[3];
  assign _T_942 = _T_936[4];
  assign _T_943 = _T_936[5];
  assign _T_944 = _T_936[6];
  assign _T_945 = _T_936[7];
  assign _T_956 = 16'h1 << _T_89_r_bits_id;
  assign _T_958 = _T_956[0];
  assign _T_959 = _T_956[1];
  assign _T_960 = _T_956[2];
  assign _T_961 = _T_956[3];
  assign _T_962 = _T_956[4];
  assign _T_963 = _T_956[5];
  assign _T_964 = _T_956[6];
  assign _T_965 = _T_956[7];
  assign _T_974 = _T_89_r_valid & _T_31_r_ready;
  assign _T_975 = _T_974 & _T_958;
  assign _T_976 = _T_975 & _T_89_r_bits_last;
  assign _T_977 = _T_31_ar_valid & _T_89_ar_ready;
  assign _T_978 = _T_977 & _T_938;
  assign _T_980 = _T_974 & _T_959;
  assign _T_981 = _T_980 & _T_89_r_bits_last;
  assign _T_983 = _T_977 & _T_939;
  assign _T_985 = _T_974 & _T_960;
  assign _T_986 = _T_985 & _T_89_r_bits_last;
  assign _T_988 = _T_977 & _T_940;
  assign _T_990 = _T_974 & _T_961;
  assign _T_991 = _T_990 & _T_89_r_bits_last;
  assign _T_993 = _T_977 & _T_941;
  assign _T_995 = _T_974 & _T_962;
  assign _T_996 = _T_995 & _T_89_r_bits_last;
  assign _T_998 = _T_977 & _T_942;
  assign _T_1000 = _T_974 & _T_963;
  assign _T_1001 = _T_1000 & _T_89_r_bits_last;
  assign _T_1003 = _T_977 & _T_943;
  assign _T_1005 = _T_974 & _T_964;
  assign _T_1006 = _T_1005 & _T_89_r_bits_last;
  assign _T_1008 = _T_977 & _T_944;
  assign _T_1010 = _T_974 & _T_965;
  assign _T_1011 = _T_1010 & _T_89_r_bits_last;
  assign _T_1013 = _T_977 & _T_945;
  assign _GEN_53 = 4'h1 == _T_31_aw_bits_id ? _T_1056_1 : _T_1056_0;
  assign _GEN_54 = 4'h2 == _T_31_aw_bits_id ? _T_1056_2 : _GEN_53;
  assign _GEN_55 = 4'h3 == _T_31_aw_bits_id ? _T_1056_3 : _GEN_54;
  assign _GEN_56 = 4'h4 == _T_31_aw_bits_id ? _T_1056_4 : _GEN_55;
  assign _GEN_57 = 4'h5 == _T_31_aw_bits_id ? _T_1056_5 : _GEN_56;
  assign _GEN_58 = 4'h6 == _T_31_aw_bits_id ? _T_1056_6 : _GEN_57;
  assign _GEN_59 = 4'h7 == _T_31_aw_bits_id ? _T_1056_7 : _GEN_58;
  assign _GEN_60 = 4'h8 == _T_31_aw_bits_id ? 1'h0 : _GEN_59;
  assign _GEN_61 = 4'h9 == _T_31_aw_bits_id ? 1'h0 : _GEN_60;
  assign _GEN_62 = 4'ha == _T_31_aw_bits_id ? 1'h0 : _GEN_61;
  assign _GEN_63 = 4'hb == _T_31_aw_bits_id ? 1'h0 : _GEN_62;
  assign _GEN_64 = 4'hc == _T_31_aw_bits_id ? 1'h0 : _GEN_63;
  assign _GEN_65 = 4'hd == _T_31_aw_bits_id ? 1'h0 : _GEN_64;
  assign _GEN_66 = 4'he == _T_31_aw_bits_id ? 1'h0 : _GEN_65;
  assign _GEN_67 = 4'hf == _T_31_aw_bits_id ? 1'h0 : _GEN_66;
  assign _T_1076 = _T_89_aw_ready & _GEN_4;
  assign _T_1077 = _T_31_aw_valid & _GEN_5;
  assign _T_1123 = _T_89_b_valid == 1'h0;
  assign _GEN_68 = 4'h1 == _T_89_b_bits_id ? _T_1080_1 : _T_1080_0;
  assign _GEN_69 = 4'h2 == _T_89_b_bits_id ? _T_1080_2 : _GEN_68;
  assign _GEN_70 = 4'h3 == _T_89_b_bits_id ? _T_1080_3 : _GEN_69;
  assign _GEN_71 = 4'h4 == _T_89_b_bits_id ? _T_1080_4 : _GEN_70;
  assign _GEN_72 = 4'h5 == _T_89_b_bits_id ? _T_1080_5 : _GEN_71;
  assign _GEN_73 = 4'h6 == _T_89_b_bits_id ? _T_1080_6 : _GEN_72;
  assign _GEN_74 = 4'h7 == _T_89_b_bits_id ? _T_1080_7 : _GEN_73;
  assign _GEN_75 = 4'h8 == _T_89_b_bits_id ? 1'h0 : _GEN_74;
  assign _GEN_76 = 4'h9 == _T_89_b_bits_id ? 1'h0 : _GEN_75;
  assign _GEN_77 = 4'ha == _T_89_b_bits_id ? 1'h0 : _GEN_76;
  assign _GEN_78 = 4'hb == _T_89_b_bits_id ? 1'h0 : _GEN_77;
  assign _GEN_79 = 4'hc == _T_89_b_bits_id ? 1'h0 : _GEN_78;
  assign _GEN_80 = 4'hd == _T_89_b_bits_id ? 1'h0 : _GEN_79;
  assign _GEN_81 = 4'he == _T_89_b_bits_id ? 1'h0 : _GEN_80;
  assign _GEN_82 = 4'hf == _T_89_b_bits_id ? 1'h0 : _GEN_81;
  assign _T_1124 = _T_1123 | _GEN_6;
  assign _T_1126 = _T_1124 | reset;
  assign _T_1128 = _T_1126 == 1'h0;
  assign _GEN_83 = 4'h1 == _T_89_b_bits_id ? _T_1102_1 : _T_1102_0;
  assign _GEN_84 = 4'h2 == _T_89_b_bits_id ? _T_1102_2 : _GEN_83;
  assign _GEN_85 = 4'h3 == _T_89_b_bits_id ? _T_1102_3 : _GEN_84;
  assign _GEN_86 = 4'h4 == _T_89_b_bits_id ? _T_1102_4 : _GEN_85;
  assign _GEN_87 = 4'h5 == _T_89_b_bits_id ? _T_1102_5 : _GEN_86;
  assign _GEN_88 = 4'h6 == _T_89_b_bits_id ? _T_1102_6 : _GEN_87;
  assign _GEN_89 = 4'h7 == _T_89_b_bits_id ? _T_1102_7 : _GEN_88;
  assign _GEN_90 = 4'h8 == _T_89_b_bits_id ? 9'h0 : _GEN_89;
  assign _GEN_91 = 4'h9 == _T_89_b_bits_id ? 9'h0 : _GEN_90;
  assign _GEN_92 = 4'ha == _T_89_b_bits_id ? 9'h0 : _GEN_91;
  assign _GEN_93 = 4'hb == _T_89_b_bits_id ? 9'h0 : _GEN_92;
  assign _GEN_94 = 4'hc == _T_89_b_bits_id ? 9'h0 : _GEN_93;
  assign _GEN_95 = 4'hd == _T_89_b_bits_id ? 9'h0 : _GEN_94;
  assign _GEN_96 = 4'he == _T_89_b_bits_id ? 9'h0 : _GEN_95;
  assign _GEN_97 = 4'hf == _T_89_b_bits_id ? 9'h0 : _GEN_96;
  assign _T_1131 = 16'h1 << _T_31_aw_bits_id;
  assign _T_1133 = _T_1131[0];
  assign _T_1134 = _T_1131[1];
  assign _T_1135 = _T_1131[2];
  assign _T_1136 = _T_1131[3];
  assign _T_1137 = _T_1131[4];
  assign _T_1138 = _T_1131[5];
  assign _T_1139 = _T_1131[6];
  assign _T_1140 = _T_1131[7];
  assign _T_1151 = 16'h1 << _T_89_b_bits_id;
  assign _T_1153 = _T_1151[0];
  assign _T_1154 = _T_1151[1];
  assign _T_1155 = _T_1151[2];
  assign _T_1156 = _T_1151[3];
  assign _T_1157 = _T_1151[4];
  assign _T_1158 = _T_1151[5];
  assign _T_1159 = _T_1151[6];
  assign _T_1160 = _T_1151[7];
  assign _T_1169 = _T_89_b_valid & _T_31_b_ready;
  assign _T_1170 = _T_1169 & _T_1153;
  assign _T_1171 = _T_31_aw_valid & _T_89_aw_ready;
  assign _T_1172 = _T_1171 & _T_1133;
  assign _T_1174 = _T_1169 & _T_1154;
  assign _T_1176 = _T_1171 & _T_1134;
  assign _T_1178 = _T_1169 & _T_1155;
  assign _T_1180 = _T_1171 & _T_1135;
  assign _T_1182 = _T_1169 & _T_1156;
  assign _T_1184 = _T_1171 & _T_1136;
  assign _T_1186 = _T_1169 & _T_1157;
  assign _T_1188 = _T_1171 & _T_1137;
  assign _T_1190 = _T_1169 & _T_1158;
  assign _T_1192 = _T_1171 & _T_1138;
  assign _T_1194 = _T_1169 & _T_1159;
  assign _T_1196 = _T_1171 & _T_1139;
  assign _T_1198 = _T_1169 & _T_1160;
  assign _T_1200 = _T_1171 & _T_1140;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_1076;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _GEN_7;
  assign _T_31_ar_ready = _T_881;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _GEN_3;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_1077;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id;
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_lock = _T_31_aw_bits_lock;
  assign _T_89_aw_bits_cache = _T_31_aw_bits_cache;
  assign _T_89_aw_bits_prot = _T_31_aw_bits_prot;
  assign _T_89_aw_bits_qos = _T_31_aw_bits_qos;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_882;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id;
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_lock = _T_31_ar_bits_lock;
  assign _T_89_ar_bits_cache = _T_31_ar_bits_cache;
  assign _T_89_ar_bits_prot = _T_31_ar_bits_prot;
  assign _T_89_ar_bits_qos = _T_31_ar_bits_qos;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_978;
  assign Queue_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_io_deq_ready = _T_976;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_983;
  assign Queue_1_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_1_io_deq_ready = _T_981;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_2_io_enq_valid = _T_988;
  assign Queue_2_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_2_io_deq_ready = _T_986;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_3_io_enq_valid = _T_993;
  assign Queue_3_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_3_io_deq_ready = _T_991;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_4_io_enq_valid = _T_998;
  assign Queue_4_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_4_io_deq_ready = _T_996;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_5_io_enq_valid = _T_1003;
  assign Queue_5_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_5_io_deq_ready = _T_1001;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_6_io_enq_valid = _T_1008;
  assign Queue_6_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_6_io_deq_ready = _T_1006;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_7_io_enq_valid = _T_1013;
  assign Queue_7_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_7_io_deq_ready = _T_1011;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_8_io_enq_valid = _T_1172;
  assign Queue_8_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_8_io_deq_ready = _T_1170;
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_9_io_enq_valid = _T_1176;
  assign Queue_9_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_9_io_deq_ready = _T_1174;
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_10_io_enq_valid = _T_1180;
  assign Queue_10_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_10_io_deq_ready = _T_1178;
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_11_io_enq_valid = _T_1184;
  assign Queue_11_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_11_io_deq_ready = _T_1182;
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_12_io_enq_valid = _T_1188;
  assign Queue_12_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_12_io_deq_ready = _T_1186;
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_13_io_enq_valid = _T_1192;
  assign Queue_13_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_13_io_deq_ready = _T_1190;
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_14_io_enq_valid = _T_1196;
  assign Queue_14_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_14_io_deq_ready = _T_1194;
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_15_io_enq_valid = _T_1200;
  assign Queue_15_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_15_io_deq_ready = _T_1198;
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign _T_861_0 = Queue_io_enq_ready;
  assign _T_861_1 = Queue_1_io_enq_ready;
  assign _T_861_2 = Queue_2_io_enq_ready;
  assign _T_861_3 = Queue_3_io_enq_ready;
  assign _T_861_4 = Queue_4_io_enq_ready;
  assign _T_861_5 = Queue_5_io_enq_ready;
  assign _T_861_6 = Queue_6_io_enq_ready;
  assign _T_861_7 = Queue_7_io_enq_ready;
  assign _GEN_0 = _GEN_22;
  assign _GEN_1 = _GEN_22;
  assign _T_885_0 = Queue_io_deq_valid;
  assign _T_885_1 = Queue_1_io_deq_valid;
  assign _T_885_2 = Queue_2_io_deq_valid;
  assign _T_885_3 = Queue_3_io_deq_valid;
  assign _T_885_4 = Queue_4_io_deq_valid;
  assign _T_885_5 = Queue_5_io_deq_valid;
  assign _T_885_6 = Queue_6_io_deq_valid;
  assign _T_885_7 = Queue_7_io_deq_valid;
  assign _T_907_0 = Queue_io_deq_bits;
  assign _T_907_1 = Queue_1_io_deq_bits;
  assign _T_907_2 = Queue_2_io_deq_bits;
  assign _T_907_3 = Queue_3_io_deq_bits;
  assign _T_907_4 = Queue_4_io_deq_bits;
  assign _T_907_5 = Queue_5_io_deq_bits;
  assign _T_907_6 = Queue_6_io_deq_bits;
  assign _T_907_7 = Queue_7_io_deq_bits;
  assign _GEN_2 = _GEN_37;
  assign _GEN_3 = _GEN_52;
  assign _T_1056_0 = Queue_8_io_enq_ready;
  assign _T_1056_1 = Queue_9_io_enq_ready;
  assign _T_1056_2 = Queue_10_io_enq_ready;
  assign _T_1056_3 = Queue_11_io_enq_ready;
  assign _T_1056_4 = Queue_12_io_enq_ready;
  assign _T_1056_5 = Queue_13_io_enq_ready;
  assign _T_1056_6 = Queue_14_io_enq_ready;
  assign _T_1056_7 = Queue_15_io_enq_ready;
  assign _GEN_4 = _GEN_67;
  assign _GEN_5 = _GEN_67;
  assign _T_1080_0 = Queue_8_io_deq_valid;
  assign _T_1080_1 = Queue_9_io_deq_valid;
  assign _T_1080_2 = Queue_10_io_deq_valid;
  assign _T_1080_3 = Queue_11_io_deq_valid;
  assign _T_1080_4 = Queue_12_io_deq_valid;
  assign _T_1080_5 = Queue_13_io_deq_valid;
  assign _T_1080_6 = Queue_14_io_deq_valid;
  assign _T_1080_7 = Queue_15_io_deq_valid;
  assign _T_1102_0 = Queue_8_io_deq_bits;
  assign _T_1102_1 = Queue_9_io_deq_bits;
  assign _T_1102_2 = Queue_10_io_deq_bits;
  assign _T_1102_3 = Queue_11_io_deq_bits;
  assign _T_1102_4 = Queue_12_io_deq_bits;
  assign _T_1102_5 = Queue_13_io_deq_bits;
  assign _T_1102_6 = Queue_14_io_deq_bits;
  assign _T_1102_7 = Queue_15_io_deq_bits;
  assign _GEN_6 = _GEN_82;
  assign _GEN_7 = _GEN_97;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_933) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_933) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1128) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_92(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input  [8:0]  io_enq_bits_user,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output [8:0]  io_deq_bits_user,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:7];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire [2:0] ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire [2:0] ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [63:0] ram_data [0:7];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_50_data;
  wire [2:0] ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire [2:0] ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg [1:0] ram_resp [0:7];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_50_data;
  wire [2:0] ram_resp__T_50_addr;
  wire [1:0] ram_resp__T_36_data;
  wire [2:0] ram_resp__T_36_addr;
  wire  ram_resp__T_36_mask;
  wire  ram_resp__T_36_en;
  reg [8:0] ram_user [0:7];
  reg [31:0] _RAND_3;
  wire [8:0] ram_user__T_50_data;
  wire [2:0] ram_user__T_50_addr;
  wire [8:0] ram_user__T_36_data;
  wire [2:0] ram_user__T_36_addr;
  wire  ram_user__T_36_mask;
  wire  ram_user__T_36_en;
  reg  ram_last [0:7];
  reg [31:0] _RAND_4;
  wire  ram_last__T_50_data;
  wire [2:0] ram_last__T_50_addr;
  wire  ram_last__T_36_data;
  wire [2:0] ram_last__T_36_addr;
  wire  ram_last__T_36_mask;
  wire  ram_last__T_36_en;
  reg [2:0] value;
  reg [31:0] _RAND_5;
  reg [2:0] value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [3:0] _T_39;
  wire [2:0] _T_40;
  wire [2:0] _GEN_8;
  wire [3:0] _T_43;
  wire [2:0] _T_44;
  wire [2:0] _GEN_9;
  wire  _T_45;
  wire  _GEN_10;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign ram_resp__T_50_addr = value_1;
  assign ram_resp__T_50_data = ram_resp[ram_resp__T_50_addr];
  assign ram_resp__T_36_data = io_enq_bits_resp;
  assign ram_resp__T_36_addr = value;
  assign ram_resp__T_36_mask = do_enq;
  assign ram_resp__T_36_en = do_enq;
  assign ram_user__T_50_addr = value_1;
  assign ram_user__T_50_data = ram_user[ram_user__T_50_addr];
  assign ram_user__T_36_data = io_enq_bits_user;
  assign ram_user__T_36_addr = value;
  assign ram_user__T_36_mask = do_enq;
  assign ram_user__T_36_en = do_enq;
  assign ram_last__T_50_addr = value_1;
  assign ram_last__T_50_data = ram_last[ram_last__T_50_addr];
  assign ram_last__T_36_data = io_enq_bits_last;
  assign ram_last__T_36_addr = value;
  assign ram_last__T_36_mask = do_enq;
  assign ram_last__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 3'h1;
  assign _T_40 = _T_39[2:0];
  assign _GEN_8 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 3'h1;
  assign _T_44 = _T_43[2:0];
  assign _GEN_9 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_10 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign io_deq_bits_resp = ram_resp__T_50_data;
  assign io_deq_bits_user = ram_user__T_50_data;
  assign io_deq_bits_last = ram_last__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_user[initvar] = _RAND_3[8:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_last[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if(ram_resp__T_36_en & ram_resp__T_36_mask) begin
      ram_resp[ram_resp__T_36_addr] <= ram_resp__T_36_data;
    end
    if(ram_user__T_36_en & ram_user__T_36_mask) begin
      ram_user[ram_user__T_36_addr] <= ram_user__T_36_data;
    end
    if(ram_last__T_36_en & ram_last__T_36_mask) begin
      ram_last[ram_last__T_36_addr] <= ram_last__T_36_data;
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Deinterleaver(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [30:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [8:0]  auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [8:0]  auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [30:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [8:0]  auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [8:0]  auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [8:0]  auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [8:0]  auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [8:0]  auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [8:0]  auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [30:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire [8:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [8:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [30:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire [8:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [8:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [30:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire [8:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [8:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [30:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire [8:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [8:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [63:0] Queue_io_enq_bits_data;
  wire [1:0] Queue_io_enq_bits_resp;
  wire [8:0] Queue_io_enq_bits_user;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [63:0] Queue_io_deq_bits_data;
  wire [1:0] Queue_io_deq_bits_resp;
  wire [8:0] Queue_io_deq_bits_user;
  wire  Queue_io_deq_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_id;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [1:0] Queue_1_io_enq_bits_resp;
  wire [8:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_id;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [1:0] Queue_1_io_deq_bits_resp;
  wire [8:0] Queue_1_io_deq_bits_user;
  wire  Queue_1_io_deq_bits_last;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire [8:0] Queue_2_io_enq_bits_user;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire [8:0] Queue_2_io_deq_bits_user;
  wire  Queue_2_io_deq_bits_last;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [63:0] Queue_3_io_enq_bits_data;
  wire [1:0] Queue_3_io_enq_bits_resp;
  wire [8:0] Queue_3_io_enq_bits_user;
  wire  Queue_3_io_enq_bits_last;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [63:0] Queue_3_io_deq_bits_data;
  wire [1:0] Queue_3_io_deq_bits_resp;
  wire [8:0] Queue_3_io_deq_bits_user;
  wire  Queue_3_io_deq_bits_last;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire [8:0] Queue_4_io_enq_bits_user;
  wire  Queue_4_io_enq_bits_last;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire [8:0] Queue_4_io_deq_bits_user;
  wire  Queue_4_io_deq_bits_last;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [3:0] Queue_5_io_enq_bits_id;
  wire [63:0] Queue_5_io_enq_bits_data;
  wire [1:0] Queue_5_io_enq_bits_resp;
  wire [8:0] Queue_5_io_enq_bits_user;
  wire  Queue_5_io_enq_bits_last;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [3:0] Queue_5_io_deq_bits_id;
  wire [63:0] Queue_5_io_deq_bits_data;
  wire [1:0] Queue_5_io_deq_bits_resp;
  wire [8:0] Queue_5_io_deq_bits_user;
  wire  Queue_5_io_deq_bits_last;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [3:0] Queue_6_io_enq_bits_id;
  wire [63:0] Queue_6_io_enq_bits_data;
  wire [1:0] Queue_6_io_enq_bits_resp;
  wire [8:0] Queue_6_io_enq_bits_user;
  wire  Queue_6_io_enq_bits_last;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [3:0] Queue_6_io_deq_bits_id;
  wire [63:0] Queue_6_io_deq_bits_data;
  wire [1:0] Queue_6_io_deq_bits_resp;
  wire [8:0] Queue_6_io_deq_bits_user;
  wire  Queue_6_io_deq_bits_last;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [3:0] Queue_7_io_enq_bits_id;
  wire [63:0] Queue_7_io_enq_bits_data;
  wire [1:0] Queue_7_io_enq_bits_resp;
  wire [8:0] Queue_7_io_enq_bits_user;
  wire  Queue_7_io_enq_bits_last;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [3:0] Queue_7_io_deq_bits_id;
  wire [63:0] Queue_7_io_deq_bits_data;
  wire [1:0] Queue_7_io_deq_bits_resp;
  wire [8:0] Queue_7_io_deq_bits_user;
  wire  Queue_7_io_deq_bits_last;
  reg  _T_533;
  reg [31:0] _RAND_0;
  reg [3:0] _T_535;
  reg [31:0] _RAND_1;
  wire [15:0] _T_538;
  wire [15:0] _T_542;
  reg [3:0] _T_546;
  reg [31:0] _RAND_2;
  wire [3:0] _T_547;
  wire  _T_548;
  wire  _T_549;
  wire  _T_550;
  wire  _T_551;
  wire  _T_552;
  wire  _T_553;
  wire  _T_554;
  wire  _T_555;
  wire [3:0] _GEN_0;
  wire [4:0] _T_556;
  wire [3:0] _T_557;
  wire [3:0] _GEN_1;
  wire [4:0] _T_558;
  wire [4:0] _T_559;
  wire [3:0] _T_560;
  wire  _T_562;
  wire  _T_564;
  wire  _T_565;
  wire  _T_567;
  wire  _T_569;
  wire  _T_571;
  wire  _T_573;
  wire  _T_574;
  wire  _T_576;
  wire  _T_578;
  wire  _T_580;
  reg [3:0] _T_583;
  reg [31:0] _RAND_3;
  wire [3:0] _T_584;
  wire  _T_585;
  wire  _T_587;
  wire  _T_588;
  wire  _T_589;
  wire  _T_591;
  wire  _T_592;
  wire [3:0] _GEN_2;
  wire [4:0] _T_593;
  wire [3:0] _T_594;
  wire [3:0] _GEN_3;
  wire [4:0] _T_595;
  wire [4:0] _T_596;
  wire [3:0] _T_597;
  wire  _T_599;
  wire  _T_601;
  wire  _T_602;
  wire  _T_604;
  wire  _T_606;
  wire  _T_608;
  wire  _T_610;
  wire  _T_611;
  wire  _T_613;
  wire  _T_615;
  wire  _T_617;
  reg [3:0] _T_620;
  reg [31:0] _RAND_4;
  wire [3:0] _T_621;
  wire  _T_622;
  wire  _T_624;
  wire  _T_625;
  wire  _T_626;
  wire  _T_628;
  wire  _T_629;
  wire [3:0] _GEN_4;
  wire [4:0] _T_630;
  wire [3:0] _T_631;
  wire [3:0] _GEN_98;
  wire [4:0] _T_632;
  wire [4:0] _T_633;
  wire [3:0] _T_634;
  wire  _T_636;
  wire  _T_638;
  wire  _T_639;
  wire  _T_641;
  wire  _T_643;
  wire  _T_645;
  wire  _T_647;
  wire  _T_648;
  wire  _T_650;
  wire  _T_652;
  wire  _T_654;
  reg [3:0] _T_657;
  reg [31:0] _RAND_5;
  wire [3:0] _T_658;
  wire  _T_659;
  wire  _T_661;
  wire  _T_662;
  wire  _T_663;
  wire  _T_665;
  wire  _T_666;
  wire [3:0] _GEN_99;
  wire [4:0] _T_667;
  wire [3:0] _T_668;
  wire [3:0] _GEN_100;
  wire [4:0] _T_669;
  wire [4:0] _T_670;
  wire [3:0] _T_671;
  wire  _T_673;
  wire  _T_675;
  wire  _T_676;
  wire  _T_678;
  wire  _T_680;
  wire  _T_682;
  wire  _T_684;
  wire  _T_685;
  wire  _T_687;
  wire  _T_689;
  wire  _T_691;
  reg [3:0] _T_694;
  reg [31:0] _RAND_6;
  wire [3:0] _T_695;
  wire  _T_696;
  wire  _T_698;
  wire  _T_699;
  wire  _T_700;
  wire  _T_702;
  wire  _T_703;
  wire [3:0] _GEN_101;
  wire [4:0] _T_704;
  wire [3:0] _T_705;
  wire [3:0] _GEN_102;
  wire [4:0] _T_706;
  wire [4:0] _T_707;
  wire [3:0] _T_708;
  wire  _T_710;
  wire  _T_712;
  wire  _T_713;
  wire  _T_715;
  wire  _T_717;
  wire  _T_719;
  wire  _T_721;
  wire  _T_722;
  wire  _T_724;
  wire  _T_726;
  wire  _T_728;
  reg [3:0] _T_731;
  reg [31:0] _RAND_7;
  wire [3:0] _T_732;
  wire  _T_733;
  wire  _T_735;
  wire  _T_736;
  wire  _T_737;
  wire  _T_739;
  wire  _T_740;
  wire [3:0] _GEN_103;
  wire [4:0] _T_741;
  wire [3:0] _T_742;
  wire [3:0] _GEN_104;
  wire [4:0] _T_743;
  wire [4:0] _T_744;
  wire [3:0] _T_745;
  wire  _T_747;
  wire  _T_749;
  wire  _T_750;
  wire  _T_752;
  wire  _T_754;
  wire  _T_756;
  wire  _T_758;
  wire  _T_759;
  wire  _T_761;
  wire  _T_763;
  wire  _T_765;
  reg [3:0] _T_768;
  reg [31:0] _RAND_8;
  wire [3:0] _T_769;
  wire  _T_770;
  wire  _T_772;
  wire  _T_773;
  wire  _T_774;
  wire  _T_776;
  wire  _T_777;
  wire [3:0] _GEN_105;
  wire [4:0] _T_778;
  wire [3:0] _T_779;
  wire [3:0] _GEN_106;
  wire [4:0] _T_780;
  wire [4:0] _T_781;
  wire [3:0] _T_782;
  wire  _T_784;
  wire  _T_786;
  wire  _T_787;
  wire  _T_789;
  wire  _T_791;
  wire  _T_793;
  wire  _T_795;
  wire  _T_796;
  wire  _T_798;
  wire  _T_800;
  wire  _T_802;
  reg [3:0] _T_805;
  reg [31:0] _RAND_9;
  wire [3:0] _T_806;
  wire  _T_807;
  wire  _T_809;
  wire  _T_810;
  wire  _T_811;
  wire  _T_813;
  wire  _T_814;
  wire [3:0] _GEN_107;
  wire [4:0] _T_815;
  wire [3:0] _T_816;
  wire [3:0] _GEN_108;
  wire [4:0] _T_817;
  wire [4:0] _T_818;
  wire [3:0] _T_819;
  wire  _T_821;
  wire  _T_823;
  wire  _T_824;
  wire  _T_826;
  wire  _T_828;
  wire  _T_830;
  wire  _T_832;
  wire  _T_833;
  wire  _T_835;
  wire  _T_837;
  wire  _T_839;
  wire [1:0] _T_848;
  wire [1:0] _T_849;
  wire [3:0] _T_850;
  wire [1:0] _T_851;
  wire [1:0] _T_852;
  wire [3:0] _T_853;
  wire [7:0] _T_854;
  wire [15:0] _T_862;
  wire [16:0] _GEN_109;
  wire [16:0] _T_863;
  wire [15:0] _T_864;
  wire [15:0] _T_865;
  wire [17:0] _GEN_110;
  wire [17:0] _T_866;
  wire [15:0] _T_867;
  wire [15:0] _T_868;
  wire [19:0] _GEN_111;
  wire [19:0] _T_869;
  wire [15:0] _T_870;
  wire [15:0] _T_871;
  wire [23:0] _GEN_112;
  wire [23:0] _T_872;
  wire [15:0] _T_873;
  wire [15:0] _T_874;
  wire [16:0] _GEN_113;
  wire [16:0] _T_876;
  wire [16:0] _T_877;
  wire [16:0] _T_878;
  wire  _T_880;
  wire  _T_882;
  wire  _T_883;
  wire  _T_885;
  wire  _T_886;
  wire [15:0] _T_887;
  wire [15:0] _GEN_115;
  wire [15:0] _T_890;
  wire [7:0] _T_891;
  wire [7:0] _T_892;
  wire  _T_894;
  wire [7:0] _T_895;
  wire [3:0] _T_896;
  wire [3:0] _T_897;
  wire  _T_899;
  wire [3:0] _T_900;
  wire [1:0] _T_901;
  wire [1:0] _T_902;
  wire  _T_904;
  wire [1:0] _T_905;
  wire  _T_906;
  wire [1:0] _T_907;
  wire [2:0] _T_908;
  wire [3:0] _T_909;
  wire [4:0] _T_910;
  wire  _GEN_6;
  wire [4:0] _GEN_7;
  wire [3:0] _T_913_0_id;
  wire [63:0] _T_913_0_data;
  wire [1:0] _T_913_0_resp;
  wire [8:0] _T_913_0_user;
  wire  _T_913_0_last;
  wire [3:0] _T_913_1_id;
  wire [63:0] _T_913_1_data;
  wire [1:0] _T_913_1_resp;
  wire [8:0] _T_913_1_user;
  wire  _T_913_1_last;
  wire [3:0] _T_913_2_id;
  wire [63:0] _T_913_2_data;
  wire [1:0] _T_913_2_resp;
  wire [8:0] _T_913_2_user;
  wire  _T_913_2_last;
  wire [3:0] _T_913_3_id;
  wire [63:0] _T_913_3_data;
  wire [1:0] _T_913_3_resp;
  wire [8:0] _T_913_3_user;
  wire  _T_913_3_last;
  wire [3:0] _T_913_4_id;
  wire [63:0] _T_913_4_data;
  wire [1:0] _T_913_4_resp;
  wire [8:0] _T_913_4_user;
  wire  _T_913_4_last;
  wire [3:0] _T_913_5_id;
  wire [63:0] _T_913_5_data;
  wire [1:0] _T_913_5_resp;
  wire [8:0] _T_913_5_user;
  wire  _T_913_5_last;
  wire [3:0] _T_913_6_id;
  wire [63:0] _T_913_6_data;
  wire [1:0] _T_913_6_resp;
  wire [8:0] _T_913_6_user;
  wire  _T_913_6_last;
  wire [3:0] _T_913_7_id;
  wire [63:0] _T_913_7_data;
  wire [1:0] _T_913_7_resp;
  wire [8:0] _T_913_7_user;
  wire  _T_913_7_last;
  wire [3:0] _GEN_0_id;
  wire [3:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [1:0] _GEN_10;
  wire [8:0] _GEN_11;
  wire  _GEN_12;
  wire [3:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [8:0] _GEN_16;
  wire  _GEN_17;
  wire [3:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [8:0] _GEN_21;
  wire  _GEN_22;
  wire [3:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [8:0] _GEN_26;
  wire  _GEN_27;
  wire [3:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [1:0] _GEN_30;
  wire [8:0] _GEN_31;
  wire  _GEN_32;
  wire [3:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [1:0] _GEN_35;
  wire [8:0] _GEN_36;
  wire  _GEN_37;
  wire [3:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [1:0] _GEN_40;
  wire [8:0] _GEN_41;
  wire  _GEN_42;
  wire [3:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [1:0] _GEN_45;
  wire [8:0] _GEN_46;
  wire  _GEN_47;
  wire [3:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [1:0] _GEN_50;
  wire [8:0] _GEN_51;
  wire  _GEN_52;
  wire [3:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [1:0] _GEN_55;
  wire [8:0] _GEN_56;
  wire  _GEN_57;
  wire [3:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [1:0] _GEN_60;
  wire [8:0] _GEN_61;
  wire  _GEN_62;
  wire [3:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [1:0] _GEN_65;
  wire [8:0] _GEN_66;
  wire  _GEN_67;
  wire [3:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [1:0] _GEN_70;
  wire [8:0] _GEN_71;
  wire  _GEN_72;
  wire [3:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [1:0] _GEN_75;
  wire [8:0] _GEN_76;
  wire  _GEN_77;
  wire [3:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [1:0] _GEN_80;
  wire [8:0] _GEN_81;
  wire  _GEN_82;
  wire [63:0] _GEN_1_data;
  wire [1:0] _GEN_2_resp;
  wire [8:0] _GEN_3_user;
  wire  _GEN_4_last;
  wire  _T_983_0;
  wire  _T_983_1;
  wire  _T_983_2;
  wire  _T_983_3;
  wire  _T_983_4;
  wire  _T_983_5;
  wire  _T_983_6;
  wire  _T_983_7;
  wire  _GEN_5;
  wire  _GEN_83;
  wire  _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1021;
  wire  _T_1022;
  wire  _T_1023;
  wire  _T_1024;
  wire  _T_1025;
  wire  _T_1026;
  Queue_92 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_user(Queue_io_deq_bits_user),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_92 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_92 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  Queue_92 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_enq_bits_resp(Queue_3_io_enq_bits_resp),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_enq_bits_last(Queue_3_io_enq_bits_last),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_resp(Queue_3_io_deq_bits_resp),
    .io_deq_bits_user(Queue_3_io_deq_bits_user),
    .io_deq_bits_last(Queue_3_io_deq_bits_last)
  );
  Queue_92 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_user(Queue_4_io_enq_bits_user),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_user(Queue_4_io_deq_bits_user),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  Queue_92 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_id(Queue_5_io_enq_bits_id),
    .io_enq_bits_data(Queue_5_io_enq_bits_data),
    .io_enq_bits_resp(Queue_5_io_enq_bits_resp),
    .io_enq_bits_user(Queue_5_io_enq_bits_user),
    .io_enq_bits_last(Queue_5_io_enq_bits_last),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_id(Queue_5_io_deq_bits_id),
    .io_deq_bits_data(Queue_5_io_deq_bits_data),
    .io_deq_bits_resp(Queue_5_io_deq_bits_resp),
    .io_deq_bits_user(Queue_5_io_deq_bits_user),
    .io_deq_bits_last(Queue_5_io_deq_bits_last)
  );
  Queue_92 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_id(Queue_6_io_enq_bits_id),
    .io_enq_bits_data(Queue_6_io_enq_bits_data),
    .io_enq_bits_resp(Queue_6_io_enq_bits_resp),
    .io_enq_bits_user(Queue_6_io_enq_bits_user),
    .io_enq_bits_last(Queue_6_io_enq_bits_last),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_id(Queue_6_io_deq_bits_id),
    .io_deq_bits_data(Queue_6_io_deq_bits_data),
    .io_deq_bits_resp(Queue_6_io_deq_bits_resp),
    .io_deq_bits_user(Queue_6_io_deq_bits_user),
    .io_deq_bits_last(Queue_6_io_deq_bits_last)
  );
  Queue_92 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_id(Queue_7_io_enq_bits_id),
    .io_enq_bits_data(Queue_7_io_enq_bits_data),
    .io_enq_bits_resp(Queue_7_io_enq_bits_resp),
    .io_enq_bits_user(Queue_7_io_enq_bits_user),
    .io_enq_bits_last(Queue_7_io_enq_bits_last),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_id(Queue_7_io_deq_bits_id),
    .io_deq_bits_data(Queue_7_io_deq_bits_data),
    .io_deq_bits_resp(Queue_7_io_deq_bits_resp),
    .io_deq_bits_user(Queue_7_io_deq_bits_user),
    .io_deq_bits_last(Queue_7_io_deq_bits_last)
  );
  assign _T_538 = 16'h1 << _T_535;
  assign _T_542 = 16'h1 << _T_89_r_bits_id;
  assign _T_548 = _T_542[0];
  assign _T_549 = _T_89_r_ready & _T_89_r_valid;
  assign _T_550 = _T_548 & _T_549;
  assign _T_551 = _T_550 & _T_89_r_bits_last;
  assign _T_552 = _T_538[0];
  assign _T_553 = _T_31_r_ready & _T_31_r_valid;
  assign _T_554 = _T_552 & _T_553;
  assign _T_555 = _T_554 & _T_31_r_bits_last;
  assign _GEN_0 = {{3'd0}, _T_551};
  assign _T_556 = _T_546 + _GEN_0;
  assign _T_557 = _T_556[3:0];
  assign _GEN_1 = {{3'd0}, _T_555};
  assign _T_558 = _T_557 - _GEN_1;
  assign _T_559 = $unsigned(_T_558);
  assign _T_560 = _T_559[3:0];
  assign _T_562 = _T_555 == 1'h0;
  assign _T_564 = _T_546 != 4'h0;
  assign _T_565 = _T_562 | _T_564;
  assign _T_567 = _T_565 | reset;
  assign _T_569 = _T_567 == 1'h0;
  assign _T_571 = _T_551 == 1'h0;
  assign _T_573 = _T_546 != 4'h8;
  assign _T_574 = _T_571 | _T_573;
  assign _T_576 = _T_574 | reset;
  assign _T_578 = _T_576 == 1'h0;
  assign _T_580 = _T_547 != 4'h0;
  assign _T_585 = _T_542[1];
  assign _T_587 = _T_585 & _T_549;
  assign _T_588 = _T_587 & _T_89_r_bits_last;
  assign _T_589 = _T_538[1];
  assign _T_591 = _T_589 & _T_553;
  assign _T_592 = _T_591 & _T_31_r_bits_last;
  assign _GEN_2 = {{3'd0}, _T_588};
  assign _T_593 = _T_583 + _GEN_2;
  assign _T_594 = _T_593[3:0];
  assign _GEN_3 = {{3'd0}, _T_592};
  assign _T_595 = _T_594 - _GEN_3;
  assign _T_596 = $unsigned(_T_595);
  assign _T_597 = _T_596[3:0];
  assign _T_599 = _T_592 == 1'h0;
  assign _T_601 = _T_583 != 4'h0;
  assign _T_602 = _T_599 | _T_601;
  assign _T_604 = _T_602 | reset;
  assign _T_606 = _T_604 == 1'h0;
  assign _T_608 = _T_588 == 1'h0;
  assign _T_610 = _T_583 != 4'h8;
  assign _T_611 = _T_608 | _T_610;
  assign _T_613 = _T_611 | reset;
  assign _T_615 = _T_613 == 1'h0;
  assign _T_617 = _T_584 != 4'h0;
  assign _T_622 = _T_542[2];
  assign _T_624 = _T_622 & _T_549;
  assign _T_625 = _T_624 & _T_89_r_bits_last;
  assign _T_626 = _T_538[2];
  assign _T_628 = _T_626 & _T_553;
  assign _T_629 = _T_628 & _T_31_r_bits_last;
  assign _GEN_4 = {{3'd0}, _T_625};
  assign _T_630 = _T_620 + _GEN_4;
  assign _T_631 = _T_630[3:0];
  assign _GEN_98 = {{3'd0}, _T_629};
  assign _T_632 = _T_631 - _GEN_98;
  assign _T_633 = $unsigned(_T_632);
  assign _T_634 = _T_633[3:0];
  assign _T_636 = _T_629 == 1'h0;
  assign _T_638 = _T_620 != 4'h0;
  assign _T_639 = _T_636 | _T_638;
  assign _T_641 = _T_639 | reset;
  assign _T_643 = _T_641 == 1'h0;
  assign _T_645 = _T_625 == 1'h0;
  assign _T_647 = _T_620 != 4'h8;
  assign _T_648 = _T_645 | _T_647;
  assign _T_650 = _T_648 | reset;
  assign _T_652 = _T_650 == 1'h0;
  assign _T_654 = _T_621 != 4'h0;
  assign _T_659 = _T_542[3];
  assign _T_661 = _T_659 & _T_549;
  assign _T_662 = _T_661 & _T_89_r_bits_last;
  assign _T_663 = _T_538[3];
  assign _T_665 = _T_663 & _T_553;
  assign _T_666 = _T_665 & _T_31_r_bits_last;
  assign _GEN_99 = {{3'd0}, _T_662};
  assign _T_667 = _T_657 + _GEN_99;
  assign _T_668 = _T_667[3:0];
  assign _GEN_100 = {{3'd0}, _T_666};
  assign _T_669 = _T_668 - _GEN_100;
  assign _T_670 = $unsigned(_T_669);
  assign _T_671 = _T_670[3:0];
  assign _T_673 = _T_666 == 1'h0;
  assign _T_675 = _T_657 != 4'h0;
  assign _T_676 = _T_673 | _T_675;
  assign _T_678 = _T_676 | reset;
  assign _T_680 = _T_678 == 1'h0;
  assign _T_682 = _T_662 == 1'h0;
  assign _T_684 = _T_657 != 4'h8;
  assign _T_685 = _T_682 | _T_684;
  assign _T_687 = _T_685 | reset;
  assign _T_689 = _T_687 == 1'h0;
  assign _T_691 = _T_658 != 4'h0;
  assign _T_696 = _T_542[4];
  assign _T_698 = _T_696 & _T_549;
  assign _T_699 = _T_698 & _T_89_r_bits_last;
  assign _T_700 = _T_538[4];
  assign _T_702 = _T_700 & _T_553;
  assign _T_703 = _T_702 & _T_31_r_bits_last;
  assign _GEN_101 = {{3'd0}, _T_699};
  assign _T_704 = _T_694 + _GEN_101;
  assign _T_705 = _T_704[3:0];
  assign _GEN_102 = {{3'd0}, _T_703};
  assign _T_706 = _T_705 - _GEN_102;
  assign _T_707 = $unsigned(_T_706);
  assign _T_708 = _T_707[3:0];
  assign _T_710 = _T_703 == 1'h0;
  assign _T_712 = _T_694 != 4'h0;
  assign _T_713 = _T_710 | _T_712;
  assign _T_715 = _T_713 | reset;
  assign _T_717 = _T_715 == 1'h0;
  assign _T_719 = _T_699 == 1'h0;
  assign _T_721 = _T_694 != 4'h8;
  assign _T_722 = _T_719 | _T_721;
  assign _T_724 = _T_722 | reset;
  assign _T_726 = _T_724 == 1'h0;
  assign _T_728 = _T_695 != 4'h0;
  assign _T_733 = _T_542[5];
  assign _T_735 = _T_733 & _T_549;
  assign _T_736 = _T_735 & _T_89_r_bits_last;
  assign _T_737 = _T_538[5];
  assign _T_739 = _T_737 & _T_553;
  assign _T_740 = _T_739 & _T_31_r_bits_last;
  assign _GEN_103 = {{3'd0}, _T_736};
  assign _T_741 = _T_731 + _GEN_103;
  assign _T_742 = _T_741[3:0];
  assign _GEN_104 = {{3'd0}, _T_740};
  assign _T_743 = _T_742 - _GEN_104;
  assign _T_744 = $unsigned(_T_743);
  assign _T_745 = _T_744[3:0];
  assign _T_747 = _T_740 == 1'h0;
  assign _T_749 = _T_731 != 4'h0;
  assign _T_750 = _T_747 | _T_749;
  assign _T_752 = _T_750 | reset;
  assign _T_754 = _T_752 == 1'h0;
  assign _T_756 = _T_736 == 1'h0;
  assign _T_758 = _T_731 != 4'h8;
  assign _T_759 = _T_756 | _T_758;
  assign _T_761 = _T_759 | reset;
  assign _T_763 = _T_761 == 1'h0;
  assign _T_765 = _T_732 != 4'h0;
  assign _T_770 = _T_542[6];
  assign _T_772 = _T_770 & _T_549;
  assign _T_773 = _T_772 & _T_89_r_bits_last;
  assign _T_774 = _T_538[6];
  assign _T_776 = _T_774 & _T_553;
  assign _T_777 = _T_776 & _T_31_r_bits_last;
  assign _GEN_105 = {{3'd0}, _T_773};
  assign _T_778 = _T_768 + _GEN_105;
  assign _T_779 = _T_778[3:0];
  assign _GEN_106 = {{3'd0}, _T_777};
  assign _T_780 = _T_779 - _GEN_106;
  assign _T_781 = $unsigned(_T_780);
  assign _T_782 = _T_781[3:0];
  assign _T_784 = _T_777 == 1'h0;
  assign _T_786 = _T_768 != 4'h0;
  assign _T_787 = _T_784 | _T_786;
  assign _T_789 = _T_787 | reset;
  assign _T_791 = _T_789 == 1'h0;
  assign _T_793 = _T_773 == 1'h0;
  assign _T_795 = _T_768 != 4'h8;
  assign _T_796 = _T_793 | _T_795;
  assign _T_798 = _T_796 | reset;
  assign _T_800 = _T_798 == 1'h0;
  assign _T_802 = _T_769 != 4'h0;
  assign _T_807 = _T_542[7];
  assign _T_809 = _T_807 & _T_549;
  assign _T_810 = _T_809 & _T_89_r_bits_last;
  assign _T_811 = _T_538[7];
  assign _T_813 = _T_811 & _T_553;
  assign _T_814 = _T_813 & _T_31_r_bits_last;
  assign _GEN_107 = {{3'd0}, _T_810};
  assign _T_815 = _T_805 + _GEN_107;
  assign _T_816 = _T_815[3:0];
  assign _GEN_108 = {{3'd0}, _T_814};
  assign _T_817 = _T_816 - _GEN_108;
  assign _T_818 = $unsigned(_T_817);
  assign _T_819 = _T_818[3:0];
  assign _T_821 = _T_814 == 1'h0;
  assign _T_823 = _T_805 != 4'h0;
  assign _T_824 = _T_821 | _T_823;
  assign _T_826 = _T_824 | reset;
  assign _T_828 = _T_826 == 1'h0;
  assign _T_830 = _T_810 == 1'h0;
  assign _T_832 = _T_805 != 4'h8;
  assign _T_833 = _T_830 | _T_832;
  assign _T_835 = _T_833 | reset;
  assign _T_837 = _T_835 == 1'h0;
  assign _T_839 = _T_806 != 4'h0;
  assign _T_848 = {_T_617,_T_580};
  assign _T_849 = {_T_691,_T_654};
  assign _T_850 = {_T_849,_T_848};
  assign _T_851 = {_T_765,_T_728};
  assign _T_852 = {_T_839,_T_802};
  assign _T_853 = {_T_852,_T_851};
  assign _T_854 = {_T_853,_T_850};
  assign _T_862 = {8'h0,_T_854};
  assign _GEN_109 = {{1'd0}, _T_862};
  assign _T_863 = _GEN_109 << 1;
  assign _T_864 = _T_863[15:0];
  assign _T_865 = _T_862 | _T_864;
  assign _GEN_110 = {{2'd0}, _T_865};
  assign _T_866 = _GEN_110 << 2;
  assign _T_867 = _T_866[15:0];
  assign _T_868 = _T_865 | _T_867;
  assign _GEN_111 = {{4'd0}, _T_868};
  assign _T_869 = _GEN_111 << 4;
  assign _T_870 = _T_869[15:0];
  assign _T_871 = _T_868 | _T_870;
  assign _GEN_112 = {{8'd0}, _T_871};
  assign _T_872 = _GEN_112 << 8;
  assign _T_873 = _T_872[15:0];
  assign _T_874 = _T_871 | _T_873;
  assign _GEN_113 = {{1'd0}, _T_874};
  assign _T_876 = _GEN_113 << 1;
  assign _T_877 = ~ _T_876;
  assign _T_878 = _GEN_109 & _T_877;
  assign _T_880 = _T_533 == 1'h0;
  assign _T_882 = _T_553 & _T_31_r_bits_last;
  assign _T_883 = _T_880 | _T_882;
  assign _T_885 = _T_862 != 16'h0;
  assign _T_886 = _T_878[16];
  assign _T_887 = _T_878[15:0];
  assign _GEN_115 = {{15'd0}, _T_886};
  assign _T_890 = _GEN_115 | _T_887;
  assign _T_891 = _T_890[15:8];
  assign _T_892 = _T_890[7:0];
  assign _T_894 = _T_891 != 8'h0;
  assign _T_895 = _T_891 | _T_892;
  assign _T_896 = _T_895[7:4];
  assign _T_897 = _T_895[3:0];
  assign _T_899 = _T_896 != 4'h0;
  assign _T_900 = _T_896 | _T_897;
  assign _T_901 = _T_900[3:2];
  assign _T_902 = _T_900[1:0];
  assign _T_904 = _T_901 != 2'h0;
  assign _T_905 = _T_901 | _T_902;
  assign _T_906 = _T_905[1];
  assign _T_907 = {_T_904,_T_906};
  assign _T_908 = {_T_899,_T_907};
  assign _T_909 = {_T_894,_T_908};
  assign _T_910 = {_T_886,_T_909};
  assign _GEN_6 = _T_883 ? _T_885 : _T_533;
  assign _GEN_7 = _T_883 ? _T_910 : {{1'd0}, _T_535};
  assign _GEN_8 = 4'h1 == _T_535 ? _T_913_1_id : _T_913_0_id;
  assign _GEN_9 = 4'h1 == _T_535 ? _T_913_1_data : _T_913_0_data;
  assign _GEN_10 = 4'h1 == _T_535 ? _T_913_1_resp : _T_913_0_resp;
  assign _GEN_11 = 4'h1 == _T_535 ? _T_913_1_user : _T_913_0_user;
  assign _GEN_12 = 4'h1 == _T_535 ? _T_913_1_last : _T_913_0_last;
  assign _GEN_13 = 4'h2 == _T_535 ? _T_913_2_id : _GEN_8;
  assign _GEN_14 = 4'h2 == _T_535 ? _T_913_2_data : _GEN_9;
  assign _GEN_15 = 4'h2 == _T_535 ? _T_913_2_resp : _GEN_10;
  assign _GEN_16 = 4'h2 == _T_535 ? _T_913_2_user : _GEN_11;
  assign _GEN_17 = 4'h2 == _T_535 ? _T_913_2_last : _GEN_12;
  assign _GEN_18 = 4'h3 == _T_535 ? _T_913_3_id : _GEN_13;
  assign _GEN_19 = 4'h3 == _T_535 ? _T_913_3_data : _GEN_14;
  assign _GEN_20 = 4'h3 == _T_535 ? _T_913_3_resp : _GEN_15;
  assign _GEN_21 = 4'h3 == _T_535 ? _T_913_3_user : _GEN_16;
  assign _GEN_22 = 4'h3 == _T_535 ? _T_913_3_last : _GEN_17;
  assign _GEN_23 = 4'h4 == _T_535 ? _T_913_4_id : _GEN_18;
  assign _GEN_24 = 4'h4 == _T_535 ? _T_913_4_data : _GEN_19;
  assign _GEN_25 = 4'h4 == _T_535 ? _T_913_4_resp : _GEN_20;
  assign _GEN_26 = 4'h4 == _T_535 ? _T_913_4_user : _GEN_21;
  assign _GEN_27 = 4'h4 == _T_535 ? _T_913_4_last : _GEN_22;
  assign _GEN_28 = 4'h5 == _T_535 ? _T_913_5_id : _GEN_23;
  assign _GEN_29 = 4'h5 == _T_535 ? _T_913_5_data : _GEN_24;
  assign _GEN_30 = 4'h5 == _T_535 ? _T_913_5_resp : _GEN_25;
  assign _GEN_31 = 4'h5 == _T_535 ? _T_913_5_user : _GEN_26;
  assign _GEN_32 = 4'h5 == _T_535 ? _T_913_5_last : _GEN_27;
  assign _GEN_33 = 4'h6 == _T_535 ? _T_913_6_id : _GEN_28;
  assign _GEN_34 = 4'h6 == _T_535 ? _T_913_6_data : _GEN_29;
  assign _GEN_35 = 4'h6 == _T_535 ? _T_913_6_resp : _GEN_30;
  assign _GEN_36 = 4'h6 == _T_535 ? _T_913_6_user : _GEN_31;
  assign _GEN_37 = 4'h6 == _T_535 ? _T_913_6_last : _GEN_32;
  assign _GEN_38 = 4'h7 == _T_535 ? _T_913_7_id : _GEN_33;
  assign _GEN_39 = 4'h7 == _T_535 ? _T_913_7_data : _GEN_34;
  assign _GEN_40 = 4'h7 == _T_535 ? _T_913_7_resp : _GEN_35;
  assign _GEN_41 = 4'h7 == _T_535 ? _T_913_7_user : _GEN_36;
  assign _GEN_42 = 4'h7 == _T_535 ? _T_913_7_last : _GEN_37;
  assign _GEN_43 = 4'h8 == _T_535 ? 4'h0 : _GEN_38;
  assign _GEN_44 = 4'h8 == _T_535 ? 64'h0 : _GEN_39;
  assign _GEN_45 = 4'h8 == _T_535 ? 2'h0 : _GEN_40;
  assign _GEN_46 = 4'h8 == _T_535 ? 9'h0 : _GEN_41;
  assign _GEN_47 = 4'h8 == _T_535 ? 1'h0 : _GEN_42;
  assign _GEN_48 = 4'h9 == _T_535 ? 4'h0 : _GEN_43;
  assign _GEN_49 = 4'h9 == _T_535 ? 64'h0 : _GEN_44;
  assign _GEN_50 = 4'h9 == _T_535 ? 2'h0 : _GEN_45;
  assign _GEN_51 = 4'h9 == _T_535 ? 9'h0 : _GEN_46;
  assign _GEN_52 = 4'h9 == _T_535 ? 1'h0 : _GEN_47;
  assign _GEN_53 = 4'ha == _T_535 ? 4'h0 : _GEN_48;
  assign _GEN_54 = 4'ha == _T_535 ? 64'h0 : _GEN_49;
  assign _GEN_55 = 4'ha == _T_535 ? 2'h0 : _GEN_50;
  assign _GEN_56 = 4'ha == _T_535 ? 9'h0 : _GEN_51;
  assign _GEN_57 = 4'ha == _T_535 ? 1'h0 : _GEN_52;
  assign _GEN_58 = 4'hb == _T_535 ? 4'h0 : _GEN_53;
  assign _GEN_59 = 4'hb == _T_535 ? 64'h0 : _GEN_54;
  assign _GEN_60 = 4'hb == _T_535 ? 2'h0 : _GEN_55;
  assign _GEN_61 = 4'hb == _T_535 ? 9'h0 : _GEN_56;
  assign _GEN_62 = 4'hb == _T_535 ? 1'h0 : _GEN_57;
  assign _GEN_63 = 4'hc == _T_535 ? 4'h0 : _GEN_58;
  assign _GEN_64 = 4'hc == _T_535 ? 64'h0 : _GEN_59;
  assign _GEN_65 = 4'hc == _T_535 ? 2'h0 : _GEN_60;
  assign _GEN_66 = 4'hc == _T_535 ? 9'h0 : _GEN_61;
  assign _GEN_67 = 4'hc == _T_535 ? 1'h0 : _GEN_62;
  assign _GEN_68 = 4'hd == _T_535 ? 4'h0 : _GEN_63;
  assign _GEN_69 = 4'hd == _T_535 ? 64'h0 : _GEN_64;
  assign _GEN_70 = 4'hd == _T_535 ? 2'h0 : _GEN_65;
  assign _GEN_71 = 4'hd == _T_535 ? 9'h0 : _GEN_66;
  assign _GEN_72 = 4'hd == _T_535 ? 1'h0 : _GEN_67;
  assign _GEN_73 = 4'he == _T_535 ? 4'h0 : _GEN_68;
  assign _GEN_74 = 4'he == _T_535 ? 64'h0 : _GEN_69;
  assign _GEN_75 = 4'he == _T_535 ? 2'h0 : _GEN_70;
  assign _GEN_76 = 4'he == _T_535 ? 9'h0 : _GEN_71;
  assign _GEN_77 = 4'he == _T_535 ? 1'h0 : _GEN_72;
  assign _GEN_78 = 4'hf == _T_535 ? 4'h0 : _GEN_73;
  assign _GEN_79 = 4'hf == _T_535 ? 64'h0 : _GEN_74;
  assign _GEN_80 = 4'hf == _T_535 ? 2'h0 : _GEN_75;
  assign _GEN_81 = 4'hf == _T_535 ? 9'h0 : _GEN_76;
  assign _GEN_82 = 4'hf == _T_535 ? 1'h0 : _GEN_77;
  assign _GEN_83 = 4'h1 == _T_89_r_bits_id ? _T_983_1 : _T_983_0;
  assign _GEN_84 = 4'h2 == _T_89_r_bits_id ? _T_983_2 : _GEN_83;
  assign _GEN_85 = 4'h3 == _T_89_r_bits_id ? _T_983_3 : _GEN_84;
  assign _GEN_86 = 4'h4 == _T_89_r_bits_id ? _T_983_4 : _GEN_85;
  assign _GEN_87 = 4'h5 == _T_89_r_bits_id ? _T_983_5 : _GEN_86;
  assign _GEN_88 = 4'h6 == _T_89_r_bits_id ? _T_983_6 : _GEN_87;
  assign _GEN_89 = 4'h7 == _T_89_r_bits_id ? _T_983_7 : _GEN_88;
  assign _GEN_90 = 4'h8 == _T_89_r_bits_id ? 1'h0 : _GEN_89;
  assign _GEN_91 = 4'h9 == _T_89_r_bits_id ? 1'h0 : _GEN_90;
  assign _GEN_92 = 4'ha == _T_89_r_bits_id ? 1'h0 : _GEN_91;
  assign _GEN_93 = 4'hb == _T_89_r_bits_id ? 1'h0 : _GEN_92;
  assign _GEN_94 = 4'hc == _T_89_r_bits_id ? 1'h0 : _GEN_93;
  assign _GEN_95 = 4'hd == _T_89_r_bits_id ? 1'h0 : _GEN_94;
  assign _GEN_96 = 4'he == _T_89_r_bits_id ? 1'h0 : _GEN_95;
  assign _GEN_97 = 4'hf == _T_89_r_bits_id ? 1'h0 : _GEN_96;
  assign _T_1019 = _T_548 & _T_89_r_valid;
  assign _T_1020 = _T_585 & _T_89_r_valid;
  assign _T_1021 = _T_622 & _T_89_r_valid;
  assign _T_1022 = _T_659 & _T_89_r_valid;
  assign _T_1023 = _T_696 & _T_89_r_valid;
  assign _T_1024 = _T_733 & _T_89_r_valid;
  assign _T_1025 = _T_770 & _T_89_r_valid;
  assign _T_1026 = _T_807 & _T_89_r_valid;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_89_aw_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _T_89_b_bits_user;
  assign _T_31_ar_ready = _T_89_ar_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_533;
  assign _T_31_r_bits_id = _GEN_0_id;
  assign _T_31_r_bits_data = _GEN_1_data;
  assign _T_31_r_bits_resp = _GEN_2_resp;
  assign _T_31_r_bits_user = _GEN_3_user;
  assign _T_31_r_bits_last = _GEN_4_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_31_aw_valid;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id;
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_lock = _T_31_aw_bits_lock;
  assign _T_89_aw_bits_cache = _T_31_aw_bits_cache;
  assign _T_89_aw_bits_prot = _T_31_aw_bits_prot;
  assign _T_89_aw_bits_qos = _T_31_aw_bits_qos;
  assign _T_89_aw_bits_user = _T_31_aw_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_31_ar_valid;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id;
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_lock = _T_31_ar_bits_lock;
  assign _T_89_ar_bits_cache = _T_31_ar_bits_cache;
  assign _T_89_ar_bits_prot = _T_31_ar_bits_prot;
  assign _T_89_ar_bits_qos = _T_31_ar_bits_qos;
  assign _T_89_ar_bits_user = _T_31_ar_bits_user;
  assign _T_89_r_ready = _GEN_5;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_1019;
  assign Queue_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_io_deq_ready = _T_554;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_1020;
  assign Queue_1_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_1_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_1_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_1_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_1_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_1_io_deq_ready = _T_591;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_2_io_enq_valid = _T_1021;
  assign Queue_2_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_2_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_2_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_2_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_2_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_2_io_deq_ready = _T_628;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_3_io_enq_valid = _T_1022;
  assign Queue_3_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_3_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_3_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_3_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_3_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_3_io_deq_ready = _T_665;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_4_io_enq_valid = _T_1023;
  assign Queue_4_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_4_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_4_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_4_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_4_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_4_io_deq_ready = _T_702;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_5_io_enq_valid = _T_1024;
  assign Queue_5_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_5_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_5_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_5_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_5_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_5_io_deq_ready = _T_739;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_6_io_enq_valid = _T_1025;
  assign Queue_6_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_6_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_6_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_6_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_6_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_6_io_deq_ready = _T_776;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_7_io_enq_valid = _T_1026;
  assign Queue_7_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_7_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_7_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_7_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_7_io_enq_bits_last = _T_89_r_bits_last;
  assign Queue_7_io_deq_ready = _T_813;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign _T_547 = _T_560;
  assign _T_584 = _T_597;
  assign _T_621 = _T_634;
  assign _T_658 = _T_671;
  assign _T_695 = _T_708;
  assign _T_732 = _T_745;
  assign _T_769 = _T_782;
  assign _T_806 = _T_819;
  assign _T_913_0_id = Queue_io_deq_bits_id;
  assign _T_913_0_data = Queue_io_deq_bits_data;
  assign _T_913_0_resp = Queue_io_deq_bits_resp;
  assign _T_913_0_user = Queue_io_deq_bits_user;
  assign _T_913_0_last = Queue_io_deq_bits_last;
  assign _T_913_1_id = Queue_1_io_deq_bits_id;
  assign _T_913_1_data = Queue_1_io_deq_bits_data;
  assign _T_913_1_resp = Queue_1_io_deq_bits_resp;
  assign _T_913_1_user = Queue_1_io_deq_bits_user;
  assign _T_913_1_last = Queue_1_io_deq_bits_last;
  assign _T_913_2_id = Queue_2_io_deq_bits_id;
  assign _T_913_2_data = Queue_2_io_deq_bits_data;
  assign _T_913_2_resp = Queue_2_io_deq_bits_resp;
  assign _T_913_2_user = Queue_2_io_deq_bits_user;
  assign _T_913_2_last = Queue_2_io_deq_bits_last;
  assign _T_913_3_id = Queue_3_io_deq_bits_id;
  assign _T_913_3_data = Queue_3_io_deq_bits_data;
  assign _T_913_3_resp = Queue_3_io_deq_bits_resp;
  assign _T_913_3_user = Queue_3_io_deq_bits_user;
  assign _T_913_3_last = Queue_3_io_deq_bits_last;
  assign _T_913_4_id = Queue_4_io_deq_bits_id;
  assign _T_913_4_data = Queue_4_io_deq_bits_data;
  assign _T_913_4_resp = Queue_4_io_deq_bits_resp;
  assign _T_913_4_user = Queue_4_io_deq_bits_user;
  assign _T_913_4_last = Queue_4_io_deq_bits_last;
  assign _T_913_5_id = Queue_5_io_deq_bits_id;
  assign _T_913_5_data = Queue_5_io_deq_bits_data;
  assign _T_913_5_resp = Queue_5_io_deq_bits_resp;
  assign _T_913_5_user = Queue_5_io_deq_bits_user;
  assign _T_913_5_last = Queue_5_io_deq_bits_last;
  assign _T_913_6_id = Queue_6_io_deq_bits_id;
  assign _T_913_6_data = Queue_6_io_deq_bits_data;
  assign _T_913_6_resp = Queue_6_io_deq_bits_resp;
  assign _T_913_6_user = Queue_6_io_deq_bits_user;
  assign _T_913_6_last = Queue_6_io_deq_bits_last;
  assign _T_913_7_id = Queue_7_io_deq_bits_id;
  assign _T_913_7_data = Queue_7_io_deq_bits_data;
  assign _T_913_7_resp = Queue_7_io_deq_bits_resp;
  assign _T_913_7_user = Queue_7_io_deq_bits_user;
  assign _T_913_7_last = Queue_7_io_deq_bits_last;
  assign _GEN_0_id = _GEN_78;
  assign _GEN_1_data = _GEN_79;
  assign _GEN_2_resp = _GEN_80;
  assign _GEN_3_user = _GEN_81;
  assign _GEN_4_last = _GEN_82;
  assign _T_983_0 = Queue_io_enq_ready;
  assign _T_983_1 = Queue_1_io_enq_ready;
  assign _T_983_2 = Queue_2_io_enq_ready;
  assign _T_983_3 = Queue_3_io_enq_ready;
  assign _T_983_4 = Queue_4_io_enq_ready;
  assign _T_983_5 = Queue_5_io_enq_ready;
  assign _T_983_6 = Queue_6_io_enq_ready;
  assign _T_983_7 = Queue_7_io_enq_ready;
  assign _GEN_5 = _GEN_97;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_533 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_535 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_546 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_583 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_620 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_657 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_694 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_731 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_768 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_805 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_533 <= 1'h0;
    end else begin
      if (_T_883) begin
        _T_533 <= _T_885;
      end
    end
    _T_535 <= _GEN_7[3:0];
    if (reset) begin
      _T_546 <= 4'h0;
    end else begin
      _T_546 <= _T_547;
    end
    if (reset) begin
      _T_583 <= 4'h0;
    end else begin
      _T_583 <= _T_584;
    end
    if (reset) begin
      _T_620 <= 4'h0;
    end else begin
      _T_620 <= _T_621;
    end
    if (reset) begin
      _T_657 <= 4'h0;
    end else begin
      _T_657 <= _T_658;
    end
    if (reset) begin
      _T_694 <= 4'h0;
    end else begin
      _T_694 <= _T_695;
    end
    if (reset) begin
      _T_731 <= 4'h0;
    end else begin
      _T_731 <= _T_732;
    end
    if (reset) begin
      _T_768 <= 4'h0;
    end else begin
      _T_768 <= _T_769;
    end
    if (reset) begin
      _T_805 <= 4'h0;
    end else begin
      _T_805 <= _T_806;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_569) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_569) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_578) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_578) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_606) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_615) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_615) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_643) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_643) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_680) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_680) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_689) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_689) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_726) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_726) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_754) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_754) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_763) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_763) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_791) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_791) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_800) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_800) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_828) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_828) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_837) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_837) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [2:0]  auto_in_aw_bits_id,
  input  [30:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [8:0]  auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [2:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [8:0]  auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [2:0]  auto_in_ar_bits_id,
  input  [30:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [8:0]  auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [2:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [8:0]  auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [8:0]  auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [8:0]  auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [8:0]  auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [8:0]  auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [2:0] _T_31_aw_bits_id;
  wire [30:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_aw_bits_lock;
  wire [3:0] _T_31_aw_bits_cache;
  wire [2:0] _T_31_aw_bits_prot;
  wire [3:0] _T_31_aw_bits_qos;
  wire [8:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [2:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [8:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [2:0] _T_31_ar_bits_id;
  wire [30:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_ar_bits_lock;
  wire [3:0] _T_31_ar_bits_cache;
  wire [2:0] _T_31_ar_bits_prot;
  wire [3:0] _T_31_ar_bits_qos;
  wire [8:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [2:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [8:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [30:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire [8:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [8:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [30:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire [8:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [8:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_89_aw_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_lock = auto_in_aw_bits_lock;
  assign _T_31_aw_bits_cache = auto_in_aw_bits_cache;
  assign _T_31_aw_bits_prot = auto_in_aw_bits_prot;
  assign _T_31_aw_bits_qos = auto_in_aw_bits_qos;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_89_b_bits_id[2:0];
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _T_89_b_bits_user;
  assign _T_31_ar_ready = _T_89_ar_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_lock = auto_in_ar_bits_lock;
  assign _T_31_ar_bits_cache = auto_in_ar_bits_cache;
  assign _T_31_ar_bits_prot = auto_in_ar_bits_prot;
  assign _T_31_ar_bits_qos = auto_in_ar_bits_qos;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id[2:0];
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _T_89_r_bits_user;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_31_aw_valid;
  assign _T_89_aw_bits_id = {{1'd0}, _T_31_aw_bits_id};
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_lock = _T_31_aw_bits_lock;
  assign _T_89_aw_bits_cache = _T_31_aw_bits_cache;
  assign _T_89_aw_bits_prot = _T_31_aw_bits_prot;
  assign _T_89_aw_bits_qos = _T_31_aw_bits_qos;
  assign _T_89_aw_bits_user = _T_31_aw_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_31_ar_valid;
  assign _T_89_ar_bits_id = {{1'd0}, _T_31_ar_bits_id};
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_lock = _T_31_ar_bits_lock;
  assign _T_89_ar_bits_cache = _T_31_ar_bits_cache;
  assign _T_89_ar_bits_prot = _T_31_ar_bits_prot;
  assign _T_89_ar_bits_qos = _T_31_ar_bits_qos;
  assign _T_89_ar_bits_user = _T_31_ar_bits_user;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
endmodule
module Queue_101(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_id,
  input  [30:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [8:0]  io_enq_bits_user,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [8:0]  io_deq_bits_user,
  output        io_deq_bits_wen
);
  reg [2:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire [2:0] ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [30:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [30:0] ram_addr__T_42_data;
  wire  ram_addr__T_42_addr;
  wire [30:0] ram_addr__T_33_data;
  wire  ram_addr__T_33_addr;
  wire  ram_addr__T_33_mask;
  wire  ram_addr__T_33_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_42_data;
  wire  ram_len__T_42_addr;
  wire [7:0] ram_len__T_33_data;
  wire  ram_len__T_33_addr;
  wire  ram_len__T_33_mask;
  wire  ram_len__T_33_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [2:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_42_data;
  wire  ram_burst__T_42_addr;
  wire [1:0] ram_burst__T_33_data;
  wire  ram_burst__T_33_addr;
  wire  ram_burst__T_33_mask;
  wire  ram_burst__T_33_en;
  reg  ram_lock [0:0];
  reg [31:0] _RAND_5;
  wire  ram_lock__T_42_data;
  wire  ram_lock__T_42_addr;
  wire  ram_lock__T_33_data;
  wire  ram_lock__T_33_addr;
  wire  ram_lock__T_33_mask;
  wire  ram_lock__T_33_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] _RAND_6;
  wire [3:0] ram_cache__T_42_data;
  wire  ram_cache__T_42_addr;
  wire [3:0] ram_cache__T_33_data;
  wire  ram_cache__T_33_addr;
  wire  ram_cache__T_33_mask;
  wire  ram_cache__T_33_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] _RAND_7;
  wire [2:0] ram_prot__T_42_data;
  wire  ram_prot__T_42_addr;
  wire [2:0] ram_prot__T_33_data;
  wire  ram_prot__T_33_addr;
  wire  ram_prot__T_33_mask;
  wire  ram_prot__T_33_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] _RAND_8;
  wire [3:0] ram_qos__T_42_data;
  wire  ram_qos__T_42_addr;
  wire [3:0] ram_qos__T_33_data;
  wire  ram_qos__T_33_addr;
  wire  ram_qos__T_33_mask;
  wire  ram_qos__T_33_en;
  reg [8:0] ram_user [0:0];
  reg [31:0] _RAND_9;
  wire [8:0] ram_user__T_42_data;
  wire  ram_user__T_42_addr;
  wire [8:0] ram_user__T_33_data;
  wire  ram_user__T_33_addr;
  wire  ram_user__T_33_mask;
  wire  ram_user__T_33_en;
  reg  ram_wen [0:0];
  reg [31:0] _RAND_10;
  wire  ram_wen__T_42_data;
  wire  ram_wen__T_42_addr;
  wire  ram_wen__T_33_data;
  wire  ram_wen__T_33_addr;
  wire  ram_wen__T_33_mask;
  wire  ram_wen__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_11;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_14;
  wire  _T_38;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire [8:0] _GEN_18;
  wire [3:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [3:0] _GEN_21;
  wire  _GEN_22;
  wire [1:0] _GEN_23;
  wire [2:0] _GEN_24;
  wire [7:0] _GEN_25;
  wire [30:0] _GEN_26;
  wire [2:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_addr__T_42_addr = 1'h0;
  assign ram_addr__T_42_data = ram_addr[ram_addr__T_42_addr];
  assign ram_addr__T_33_data = io_enq_bits_addr;
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_mask = do_enq;
  assign ram_addr__T_33_en = do_enq;
  assign ram_len__T_42_addr = 1'h0;
  assign ram_len__T_42_data = ram_len[ram_len__T_42_addr];
  assign ram_len__T_33_data = io_enq_bits_len;
  assign ram_len__T_33_addr = 1'h0;
  assign ram_len__T_33_mask = do_enq;
  assign ram_len__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_burst__T_42_addr = 1'h0;
  assign ram_burst__T_42_data = ram_burst[ram_burst__T_42_addr];
  assign ram_burst__T_33_data = 2'h1;
  assign ram_burst__T_33_addr = 1'h0;
  assign ram_burst__T_33_mask = do_enq;
  assign ram_burst__T_33_en = do_enq;
  assign ram_lock__T_42_addr = 1'h0;
  assign ram_lock__T_42_data = ram_lock[ram_lock__T_42_addr];
  assign ram_lock__T_33_data = 1'h0;
  assign ram_lock__T_33_addr = 1'h0;
  assign ram_lock__T_33_mask = do_enq;
  assign ram_lock__T_33_en = do_enq;
  assign ram_cache__T_42_addr = 1'h0;
  assign ram_cache__T_42_data = ram_cache[ram_cache__T_42_addr];
  assign ram_cache__T_33_data = 4'h0;
  assign ram_cache__T_33_addr = 1'h0;
  assign ram_cache__T_33_mask = do_enq;
  assign ram_cache__T_33_en = do_enq;
  assign ram_prot__T_42_addr = 1'h0;
  assign ram_prot__T_42_data = ram_prot[ram_prot__T_42_addr];
  assign ram_prot__T_33_data = 3'h1;
  assign ram_prot__T_33_addr = 1'h0;
  assign ram_prot__T_33_mask = do_enq;
  assign ram_prot__T_33_en = do_enq;
  assign ram_qos__T_42_addr = 1'h0;
  assign ram_qos__T_42_data = ram_qos[ram_qos__T_42_addr];
  assign ram_qos__T_33_data = 4'h0;
  assign ram_qos__T_33_addr = 1'h0;
  assign ram_qos__T_33_mask = do_enq;
  assign ram_qos__T_33_en = do_enq;
  assign ram_user__T_42_addr = 1'h0;
  assign ram_user__T_42_data = ram_user[ram_user__T_42_addr];
  assign ram_user__T_33_data = io_enq_bits_user;
  assign ram_user__T_33_addr = 1'h0;
  assign ram_user__T_33_mask = do_enq;
  assign ram_user__T_33_en = do_enq;
  assign ram_wen__T_42_addr = 1'h0;
  assign ram_wen__T_42_data = ram_wen[ram_wen__T_42_addr];
  assign ram_wen__T_33_data = io_enq_bits_wen;
  assign ram_wen__T_33_addr = 1'h0;
  assign ram_wen__T_33_mask = do_enq;
  assign ram_wen__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_14 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_15 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_16 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_17 = empty ? io_enq_bits_wen : ram_wen__T_42_data;
  assign _GEN_18 = empty ? io_enq_bits_user : ram_user__T_42_data;
  assign _GEN_19 = empty ? 4'h0 : ram_qos__T_42_data;
  assign _GEN_20 = empty ? 3'h1 : ram_prot__T_42_data;
  assign _GEN_21 = empty ? 4'h0 : ram_cache__T_42_data;
  assign _GEN_22 = empty ? 1'h0 : ram_lock__T_42_data;
  assign _GEN_23 = empty ? 2'h1 : ram_burst__T_42_data;
  assign _GEN_24 = empty ? io_enq_bits_size : ram_size__T_42_data;
  assign _GEN_25 = empty ? io_enq_bits_len : ram_len__T_42_data;
  assign _GEN_26 = empty ? io_enq_bits_addr : ram_addr__T_42_data;
  assign _GEN_27 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_28 = empty ? 1'h0 : _T_30;
  assign _GEN_29 = empty ? _GEN_16 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_15;
  assign io_deq_bits_id = _GEN_27;
  assign io_deq_bits_addr = _GEN_26;
  assign io_deq_bits_len = _GEN_25;
  assign io_deq_bits_size = _GEN_24;
  assign io_deq_bits_burst = _GEN_23;
  assign io_deq_bits_lock = _GEN_22;
  assign io_deq_bits_cache = _GEN_21;
  assign io_deq_bits_prot = _GEN_20;
  assign io_deq_bits_qos = _GEN_19;
  assign io_deq_bits_user = _GEN_18;
  assign io_deq_bits_wen = _GEN_17;
  assign do_enq = _GEN_29;
  assign do_deq = _GEN_28;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = _RAND_9[8:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  maybe_full = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_addr__T_33_en & ram_addr__T_33_mask) begin
      ram_addr[ram_addr__T_33_addr] <= ram_addr__T_33_data;
    end
    if(ram_len__T_33_en & ram_len__T_33_mask) begin
      ram_len[ram_len__T_33_addr] <= ram_len__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_burst__T_33_en & ram_burst__T_33_mask) begin
      ram_burst[ram_burst__T_33_addr] <= ram_burst__T_33_data;
    end
    if(ram_lock__T_33_en & ram_lock__T_33_mask) begin
      ram_lock[ram_lock__T_33_addr] <= ram_lock__T_33_data;
    end
    if(ram_cache__T_33_en & ram_cache__T_33_mask) begin
      ram_cache[ram_cache__T_33_addr] <= ram_cache__T_33_data;
    end
    if(ram_prot__T_33_en & ram_prot__T_33_mask) begin
      ram_prot[ram_prot__T_33_addr] <= ram_prot__T_33_data;
    end
    if(ram_qos__T_33_en & ram_qos__T_33_mask) begin
      ram_qos[ram_qos__T_33_addr] <= ram_qos__T_33_data;
    end
    if(ram_user__T_33_en & ram_user__T_33_mask) begin
      ram_user[ram_user__T_33_addr] <= ram_user__T_33_data;
    end
    if(ram_wen__T_33_en & ram_wen__T_33_mask) begin
      ram_wen[ram_wen__T_33_addr] <= ram_wen__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TLToAXI4(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [4:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [4:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [2:0]  auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [8:0]  auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [8:0]  auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [2:0]  auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [8:0]  auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [2:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [8:0]  auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [3:0] _T_31_a_bits_size;
  wire [4:0] _T_31_a_bits_source;
  wire [30:0] _T_31_a_bits_address;
  wire [7:0] _T_31_a_bits_mask;
  wire [63:0] _T_31_a_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [3:0] _T_31_d_bits_size;
  wire [4:0] _T_31_d_bits_source;
  wire [63:0] _T_31_d_bits_data;
  wire  _T_31_d_bits_error;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [2:0] _T_89_aw_bits_id;
  wire [30:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire  _T_89_aw_bits_lock;
  wire [3:0] _T_89_aw_bits_cache;
  wire [2:0] _T_89_aw_bits_prot;
  wire [3:0] _T_89_aw_bits_qos;
  wire [8:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [2:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [8:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [2:0] _T_89_ar_bits_id;
  wire [30:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire  _T_89_ar_bits_lock;
  wire [3:0] _T_89_ar_bits_cache;
  wire [2:0] _T_89_ar_bits_prot;
  wire [3:0] _T_89_ar_bits_qos;
  wire [8:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [2:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [8:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  _T_206_0;
  wire  _T_206_1;
  wire  _T_206_2;
  wire  _T_206_3;
  wire  _T_206_4;
  wire  _T_206_8;
  wire  _T_206_16;
  wire  _T_206_17;
  wire  _T_206_18;
  wire  _T_206_19;
  wire  _T_206_20;
  wire  _T_206_21;
  wire  _T_206_22;
  wire  _T_206_23;
  wire  _T_206_24;
  wire  _T_206_25;
  wire  _T_206_26;
  wire  _T_206_27;
  wire  _T_206_28;
  wire  _T_206_29;
  wire  _T_206_30;
  wire  _T_206_31;
  wire  _T_319_0;
  wire  _T_319_1;
  wire  _T_319_2;
  wire  _T_319_3;
  wire  _T_319_4;
  wire  _T_319_5;
  wire  _T_319_6;
  wire  _T_319_7;
  wire  _T_370;
  wire  _T_372;
  wire  _T_373;
  wire [22:0] _T_376;
  wire [7:0] _T_377;
  wire [7:0] _T_378;
  wire [4:0] _T_379;
  wire [4:0] _T_384;
  reg [4:0] _T_387;
  reg [31:0] _RAND_0;
  wire [5:0] _T_389;
  wire [5:0] _T_390;
  wire [4:0] _T_391;
  wire  _T_393;
  wire  _T_395;
  wire  _T_397;
  wire  _T_398;
  wire [4:0] _T_402;
  wire [4:0] _GEN_2;
  wire [8:0] _GEN_76;
  wire [8:0] _T_416;
  wire [8:0] _GEN_77;
  wire [8:0] _T_417;
  wire [4:0] _T_418;
  wire [3:0] _T_419;
  wire [4:0] _T_420;
  wire [3:0] _T_421;
  wire  _T_427_ready;
  wire  _T_427_valid;
  wire [2:0] _T_427_bits_id;
  wire [30:0] _T_427_bits_addr;
  wire [7:0] _T_427_bits_len;
  wire [2:0] _T_427_bits_size;
  wire [8:0] _T_427_bits_user;
  wire  _T_427_bits_wen;
  wire  _T_431_ready;
  wire  _T_431_valid;
  wire [63:0] _T_431_bits_data;
  wire [7:0] _T_431_bits_strb;
  wire  _T_431_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [63:0] Queue_io_enq_bits_data;
  wire [7:0] Queue_io_enq_bits_strb;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [63:0] Queue_io_deq_bits_data;
  wire [7:0] Queue_io_deq_bits_strb;
  wire  Queue_io_deq_bits_last;
  wire  _T_439_ready;
  wire  _T_439_valid;
  wire [63:0] _T_439_bits_data;
  wire [7:0] _T_439_bits_strb;
  wire  _T_439_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_id;
  wire [30:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [8:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_enq_bits_wen;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_id;
  wire [30:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire  Queue_1_io_deq_bits_lock;
  wire [3:0] Queue_1_io_deq_bits_cache;
  wire [2:0] Queue_1_io_deq_bits_prot;
  wire [3:0] Queue_1_io_deq_bits_qos;
  wire [8:0] Queue_1_io_deq_bits_user;
  wire  Queue_1_io_deq_bits_wen;
  wire  _T_447_ready;
  wire  _T_447_valid;
  wire [2:0] _T_447_bits_id;
  wire [30:0] _T_447_bits_addr;
  wire [7:0] _T_447_bits_len;
  wire [2:0] _T_447_bits_size;
  wire [1:0] _T_447_bits_burst;
  wire  _T_447_bits_lock;
  wire [3:0] _T_447_bits_cache;
  wire [2:0] _T_447_bits_prot;
  wire [3:0] _T_447_bits_qos;
  wire [8:0] _T_447_bits_user;
  wire  _T_447_bits_wen;
  wire  _T_452;
  wire  _T_453;
  wire  _T_454;
  wire  _T_455;
  reg  _T_459;
  reg [31:0] _RAND_1;
  wire  _T_462;
  wire  _GEN_3;
  wire [2:0] _GEN_0;
  wire [2:0] _GEN_4;
  wire [2:0] _GEN_5;
  wire [2:0] _GEN_6;
  wire [2:0] _GEN_7;
  wire [2:0] _GEN_8;
  wire [2:0] _GEN_9;
  wire [2:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire [2:0] _GEN_12;
  wire [2:0] _GEN_13;
  wire [2:0] _GEN_14;
  wire [2:0] _GEN_15;
  wire [2:0] _GEN_16;
  wire [2:0] _GEN_17;
  wire [2:0] _GEN_18;
  wire [2:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [2:0] _GEN_21;
  wire [2:0] _GEN_22;
  wire [2:0] _GEN_23;
  wire [2:0] _GEN_24;
  wire [2:0] _GEN_25;
  wire [2:0] _GEN_26;
  wire [2:0] _GEN_27;
  wire [2:0] _GEN_28;
  wire [2:0] _GEN_29;
  wire [2:0] _GEN_30;
  wire [2:0] _GEN_31;
  wire [2:0] _GEN_32;
  wire [2:0] _GEN_33;
  wire [2:0] _GEN_34;
  wire [25:0] _T_466;
  wire [10:0] _T_467;
  wire [10:0] _T_468;
  wire [7:0] _T_469;
  wire  _T_470;
  wire [3:0] _T_471;
  wire  _GEN_1;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _T_478;
  wire  _T_480;
  wire  _T_481;
  wire  _T_482;
  wire  _T_483;
  wire  _T_484;
  wire  _T_487;
  wire  _T_489;
  wire  _T_490;
  wire  _T_492;
  wire  _T_493;
  wire  _T_497;
  wire  _T_499;
  reg  _T_502;
  reg [31:0] _RAND_2;
  wire  _T_503;
  wire  _T_505;
  wire  _GEN_66;
  wire  _T_506;
  wire  _T_508;
  wire  _T_509;
  wire  _T_510;
  wire  _T_512;
  wire  _T_514;
  reg  _T_517;
  reg [31:0] _RAND_3;
  wire  _T_521;
  wire  _T_522;
  wire  _GEN_67;
  wire [3:0] _T_526_size;
  wire [4:0] _T_526_source;
  wire  _T_526_error;
  wire [3:0] _T_531_size;
  wire [4:0] _T_531_source;
  wire  _T_531_error;
  wire [2:0] _T_536_opcode;
  wire [3:0] _T_536_size;
  wire [4:0] _T_536_source;
  wire  _T_536_error;
  wire [7:0] _T_539;
  wire  _T_541;
  wire  _T_542;
  wire  _T_543;
  wire  _T_544;
  wire  _T_545;
  wire  _T_546;
  wire  _T_547;
  wire  _T_548;
  wire [2:0] _T_549;
  wire [7:0] _T_552;
  wire  _T_554;
  wire  _T_555;
  wire  _T_556;
  wire  _T_557;
  wire  _T_558;
  wire  _T_559;
  wire  _T_560;
  wire  _T_561;
  wire  _T_563;
  reg  _T_566;
  reg [31:0] _RAND_4;
  wire  _T_571;
  wire  _T_572;
  wire  _T_573;
  wire  _T_574;
  wire  _T_575;
  wire [1:0] _T_576;
  wire  _T_577;
  wire [1:0] _T_578;
  wire [1:0] _T_579;
  wire  _T_580;
  wire  _T_582;
  wire  _T_585;
  wire  _T_587;
  wire  _T_589;
  wire  _T_591;
  wire  _T_593;
  wire  _T_594;
  wire  _T_596;
  wire  _T_598;
  reg [3:0] _T_608;
  reg [31:0] _RAND_5;
  reg  _T_610;
  reg [31:0] _RAND_6;
  wire  _T_612;
  wire  _T_614;
  wire  _T_615;
  wire  _T_617;
  wire [3:0] _GEN_78;
  wire [4:0] _T_618;
  wire [3:0] _T_619;
  wire [3:0] _GEN_79;
  wire [4:0] _T_620;
  wire [4:0] _T_621;
  wire [3:0] _T_622;
  wire  _T_624;
  wire  _T_626;
  wire  _T_627;
  wire  _T_629;
  wire  _T_631;
  wire  _T_633;
  wire  _T_635;
  wire  _T_636;
  wire  _T_638;
  wire  _T_640;
  wire  _GEN_69;
  wire  _T_641;
  wire  _T_643;
  wire  _T_644;
  wire  _T_646;
  wire  _T_647;
  reg [3:0] _T_650;
  reg [31:0] _RAND_7;
  reg  _T_652;
  reg [31:0] _RAND_8;
  wire  _T_654;
  wire  _T_656;
  wire  _T_657;
  wire  _T_659;
  wire [3:0] _GEN_80;
  wire [4:0] _T_660;
  wire [3:0] _T_661;
  wire [3:0] _GEN_81;
  wire [4:0] _T_662;
  wire [4:0] _T_663;
  wire [3:0] _T_664;
  wire  _T_666;
  wire  _T_668;
  wire  _T_669;
  wire  _T_671;
  wire  _T_673;
  wire  _T_675;
  wire  _T_677;
  wire  _T_678;
  wire  _T_680;
  wire  _T_682;
  wire  _GEN_70;
  wire  _T_683;
  wire  _T_685;
  wire  _T_686;
  wire  _T_688;
  wire  _T_689;
  reg  _T_692;
  reg [31:0] _RAND_9;
  wire  _T_698;
  wire  _T_699;
  wire  _T_701;
  wire [1:0] _T_702;
  wire  _T_703;
  wire [1:0] _T_704;
  wire [1:0] _T_705;
  wire  _T_706;
  wire  _T_708;
  wire  _T_711;
  wire  _T_713;
  wire  _T_715;
  wire  _T_717;
  wire  _T_719;
  wire  _T_720;
  wire  _T_722;
  wire  _T_724;
  reg  _T_734;
  reg [31:0] _RAND_10;
  wire  _T_740;
  wire  _T_741;
  wire  _T_743;
  wire [1:0] _T_744;
  wire  _T_745;
  wire [1:0] _T_746;
  wire [1:0] _T_747;
  wire  _T_748;
  wire  _T_750;
  wire  _T_753;
  wire  _T_755;
  wire  _T_757;
  wire  _T_759;
  wire  _T_761;
  wire  _T_762;
  wire  _T_764;
  wire  _T_766;
  reg  _T_776;
  reg [31:0] _RAND_11;
  wire  _T_782;
  wire  _T_783;
  wire  _T_785;
  wire [1:0] _T_786;
  wire  _T_787;
  wire [1:0] _T_788;
  wire [1:0] _T_789;
  wire  _T_790;
  wire  _T_792;
  wire  _T_795;
  wire  _T_797;
  wire  _T_799;
  wire  _T_801;
  wire  _T_803;
  wire  _T_804;
  wire  _T_806;
  wire  _T_808;
  reg  _T_818;
  reg [31:0] _RAND_12;
  wire  _T_824;
  wire  _T_825;
  wire  _T_827;
  wire [1:0] _T_828;
  wire  _T_829;
  wire [1:0] _T_830;
  wire [1:0] _T_831;
  wire  _T_832;
  wire  _T_834;
  wire  _T_837;
  wire  _T_839;
  wire  _T_841;
  wire  _T_843;
  wire  _T_845;
  wire  _T_846;
  wire  _T_848;
  wire  _T_850;
  reg  _T_860;
  reg [31:0] _RAND_13;
  wire  _T_866;
  wire  _T_867;
  wire  _T_869;
  wire [1:0] _T_870;
  wire  _T_871;
  wire [1:0] _T_872;
  wire [1:0] _T_873;
  wire  _T_874;
  wire  _T_876;
  wire  _T_879;
  wire  _T_881;
  wire  _T_883;
  wire  _T_885;
  wire  _T_887;
  wire  _T_888;
  wire  _T_890;
  wire  _T_892;
  Queue_32 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_101 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_370 = _T_31_a_bits_opcode[2];
  assign _T_372 = _T_370 == 1'h0;
  assign _T_373 = _T_31_a_ready & _T_31_a_valid;
  assign _T_376 = 23'hff << _T_31_a_bits_size;
  assign _T_377 = _T_376[7:0];
  assign _T_378 = ~ _T_377;
  assign _T_379 = _T_378[7:3];
  assign _T_384 = _T_372 ? _T_379 : 5'h0;
  assign _T_389 = _T_387 - 5'h1;
  assign _T_390 = $unsigned(_T_389);
  assign _T_391 = _T_390[4:0];
  assign _T_393 = _T_387 == 5'h0;
  assign _T_395 = _T_387 == 5'h1;
  assign _T_397 = _T_384 == 5'h0;
  assign _T_398 = _T_395 | _T_397;
  assign _T_402 = _T_393 ? _T_384 : _T_391;
  assign _GEN_2 = _T_373 ? _T_402 : _T_387;
  assign _GEN_76 = {{5'd0}, _T_31_a_bits_size};
  assign _T_416 = _GEN_76 << 5;
  assign _GEN_77 = {{4'd0}, _T_31_a_bits_source};
  assign _T_417 = _GEN_77 | _T_416;
  assign _T_418 = _T_89_r_bits_user[4:0];
  assign _T_419 = _T_89_r_bits_user[8:5];
  assign _T_420 = _T_89_b_bits_user[4:0];
  assign _T_421 = _T_89_b_bits_user[8:5];
  assign _T_452 = _T_447_bits_wen == 1'h0;
  assign _T_453 = _T_447_valid & _T_452;
  assign _T_454 = _T_447_valid & _T_447_bits_wen;
  assign _T_455 = _T_447_bits_wen ? _T_89_aw_ready : _T_89_ar_ready;
  assign _T_462 = _T_398 == 1'h0;
  assign _GEN_3 = _T_373 ? _T_462 : _T_459;
  assign _GEN_4 = 5'h1 == _T_31_a_bits_source ? 3'h5 : 3'h4;
  assign _GEN_5 = 5'h2 == _T_31_a_bits_source ? 3'h6 : _GEN_4;
  assign _GEN_6 = 5'h3 == _T_31_a_bits_source ? 3'h7 : _GEN_5;
  assign _GEN_7 = 5'h4 == _T_31_a_bits_source ? 3'h3 : _GEN_6;
  assign _GEN_8 = 5'h5 == _T_31_a_bits_source ? 3'h0 : _GEN_7;
  assign _GEN_9 = 5'h6 == _T_31_a_bits_source ? 3'h0 : _GEN_8;
  assign _GEN_10 = 5'h7 == _T_31_a_bits_source ? 3'h0 : _GEN_9;
  assign _GEN_11 = 5'h8 == _T_31_a_bits_source ? 3'h0 : _GEN_10;
  assign _GEN_12 = 5'h9 == _T_31_a_bits_source ? 3'h0 : _GEN_11;
  assign _GEN_13 = 5'ha == _T_31_a_bits_source ? 3'h0 : _GEN_12;
  assign _GEN_14 = 5'hb == _T_31_a_bits_source ? 3'h0 : _GEN_13;
  assign _GEN_15 = 5'hc == _T_31_a_bits_source ? 3'h0 : _GEN_14;
  assign _GEN_16 = 5'hd == _T_31_a_bits_source ? 3'h0 : _GEN_15;
  assign _GEN_17 = 5'he == _T_31_a_bits_source ? 3'h0 : _GEN_16;
  assign _GEN_18 = 5'hf == _T_31_a_bits_source ? 3'h0 : _GEN_17;
  assign _GEN_19 = 5'h10 == _T_31_a_bits_source ? 3'h1 : _GEN_18;
  assign _GEN_20 = 5'h11 == _T_31_a_bits_source ? 3'h1 : _GEN_19;
  assign _GEN_21 = 5'h12 == _T_31_a_bits_source ? 3'h1 : _GEN_20;
  assign _GEN_22 = 5'h13 == _T_31_a_bits_source ? 3'h1 : _GEN_21;
  assign _GEN_23 = 5'h14 == _T_31_a_bits_source ? 3'h1 : _GEN_22;
  assign _GEN_24 = 5'h15 == _T_31_a_bits_source ? 3'h1 : _GEN_23;
  assign _GEN_25 = 5'h16 == _T_31_a_bits_source ? 3'h1 : _GEN_24;
  assign _GEN_26 = 5'h17 == _T_31_a_bits_source ? 3'h1 : _GEN_25;
  assign _GEN_27 = 5'h18 == _T_31_a_bits_source ? 3'h2 : _GEN_26;
  assign _GEN_28 = 5'h19 == _T_31_a_bits_source ? 3'h2 : _GEN_27;
  assign _GEN_29 = 5'h1a == _T_31_a_bits_source ? 3'h2 : _GEN_28;
  assign _GEN_30 = 5'h1b == _T_31_a_bits_source ? 3'h2 : _GEN_29;
  assign _GEN_31 = 5'h1c == _T_31_a_bits_source ? 3'h2 : _GEN_30;
  assign _GEN_32 = 5'h1d == _T_31_a_bits_source ? 3'h2 : _GEN_31;
  assign _GEN_33 = 5'h1e == _T_31_a_bits_source ? 3'h2 : _GEN_32;
  assign _GEN_34 = 5'h1f == _T_31_a_bits_source ? 3'h2 : _GEN_33;
  assign _T_466 = 26'h7ff << _T_31_a_bits_size;
  assign _T_467 = _T_466[10:0];
  assign _T_468 = ~ _T_467;
  assign _T_469 = _T_468[10:3];
  assign _T_470 = _T_31_a_bits_size >= 4'h3;
  assign _T_471 = _T_470 ? 4'h3 : _T_31_a_bits_size;
  assign _GEN_35 = 5'h1 == _T_31_a_bits_source ? _T_206_1 : _T_206_0;
  assign _GEN_36 = 5'h2 == _T_31_a_bits_source ? _T_206_2 : _GEN_35;
  assign _GEN_37 = 5'h3 == _T_31_a_bits_source ? _T_206_3 : _GEN_36;
  assign _GEN_38 = 5'h4 == _T_31_a_bits_source ? _T_206_4 : _GEN_37;
  assign _GEN_39 = 5'h5 == _T_31_a_bits_source ? 1'h0 : _GEN_38;
  assign _GEN_40 = 5'h6 == _T_31_a_bits_source ? 1'h0 : _GEN_39;
  assign _GEN_41 = 5'h7 == _T_31_a_bits_source ? 1'h0 : _GEN_40;
  assign _GEN_42 = 5'h8 == _T_31_a_bits_source ? _T_206_8 : _GEN_41;
  assign _GEN_43 = 5'h9 == _T_31_a_bits_source ? 1'h0 : _GEN_42;
  assign _GEN_44 = 5'ha == _T_31_a_bits_source ? 1'h0 : _GEN_43;
  assign _GEN_45 = 5'hb == _T_31_a_bits_source ? 1'h0 : _GEN_44;
  assign _GEN_46 = 5'hc == _T_31_a_bits_source ? 1'h0 : _GEN_45;
  assign _GEN_47 = 5'hd == _T_31_a_bits_source ? 1'h0 : _GEN_46;
  assign _GEN_48 = 5'he == _T_31_a_bits_source ? 1'h0 : _GEN_47;
  assign _GEN_49 = 5'hf == _T_31_a_bits_source ? 1'h0 : _GEN_48;
  assign _GEN_50 = 5'h10 == _T_31_a_bits_source ? _T_206_16 : _GEN_49;
  assign _GEN_51 = 5'h11 == _T_31_a_bits_source ? _T_206_17 : _GEN_50;
  assign _GEN_52 = 5'h12 == _T_31_a_bits_source ? _T_206_18 : _GEN_51;
  assign _GEN_53 = 5'h13 == _T_31_a_bits_source ? _T_206_19 : _GEN_52;
  assign _GEN_54 = 5'h14 == _T_31_a_bits_source ? _T_206_20 : _GEN_53;
  assign _GEN_55 = 5'h15 == _T_31_a_bits_source ? _T_206_21 : _GEN_54;
  assign _GEN_56 = 5'h16 == _T_31_a_bits_source ? _T_206_22 : _GEN_55;
  assign _GEN_57 = 5'h17 == _T_31_a_bits_source ? _T_206_23 : _GEN_56;
  assign _GEN_58 = 5'h18 == _T_31_a_bits_source ? _T_206_24 : _GEN_57;
  assign _GEN_59 = 5'h19 == _T_31_a_bits_source ? _T_206_25 : _GEN_58;
  assign _GEN_60 = 5'h1a == _T_31_a_bits_source ? _T_206_26 : _GEN_59;
  assign _GEN_61 = 5'h1b == _T_31_a_bits_source ? _T_206_27 : _GEN_60;
  assign _GEN_62 = 5'h1c == _T_31_a_bits_source ? _T_206_28 : _GEN_61;
  assign _GEN_63 = 5'h1d == _T_31_a_bits_source ? _T_206_29 : _GEN_62;
  assign _GEN_64 = 5'h1e == _T_31_a_bits_source ? _T_206_30 : _GEN_63;
  assign _GEN_65 = 5'h1f == _T_31_a_bits_source ? _T_206_31 : _GEN_64;
  assign _T_478 = _GEN_1 & _T_393;
  assign _T_480 = _T_478 == 1'h0;
  assign _T_481 = _T_459 | _T_427_ready;
  assign _T_482 = _T_481 & _T_431_ready;
  assign _T_483 = _T_372 ? _T_482 : _T_427_ready;
  assign _T_484 = _T_480 & _T_483;
  assign _T_487 = _T_480 & _T_31_a_valid;
  assign _T_489 = _T_459 == 1'h0;
  assign _T_490 = _T_489 & _T_431_ready;
  assign _T_492 = _T_372 ? _T_490 : 1'h1;
  assign _T_493 = _T_487 & _T_492;
  assign _T_497 = _T_487 & _T_372;
  assign _T_499 = _T_497 & _T_481;
  assign _T_503 = _T_89_r_ready & _T_89_r_valid;
  assign _T_505 = _T_89_r_bits_last == 1'h0;
  assign _GEN_66 = _T_503 ? _T_505 : _T_502;
  assign _T_506 = _T_89_r_valid | _T_502;
  assign _T_508 = _T_506 == 1'h0;
  assign _T_509 = _T_31_d_ready & _T_508;
  assign _T_510 = _T_506 ? _T_89_r_valid : _T_89_b_valid;
  assign _T_512 = _T_89_r_bits_resp != 2'h0;
  assign _T_514 = _T_89_b_bits_resp != 2'h0;
  assign _T_521 = _T_517 | _T_512;
  assign _T_522 = _T_505 & _T_521;
  assign _GEN_67 = _T_503 ? _T_522 : _T_517;
  assign _T_536_opcode = _T_506 ? 3'h1 : 3'h0;
  assign _T_536_size = _T_506 ? _T_526_size : _T_531_size;
  assign _T_536_source = _T_506 ? _T_526_source : _T_531_source;
  assign _T_536_error = _T_506 ? _T_526_error : _T_531_error;
  assign _T_539 = 8'h1 << _T_427_bits_id;
  assign _T_541 = _T_539[0];
  assign _T_542 = _T_539[1];
  assign _T_543 = _T_539[2];
  assign _T_544 = _T_539[3];
  assign _T_545 = _T_539[4];
  assign _T_546 = _T_539[5];
  assign _T_547 = _T_539[6];
  assign _T_548 = _T_539[7];
  assign _T_549 = _T_506 ? _T_89_r_bits_id : _T_89_b_bits_id;
  assign _T_552 = 8'h1 << _T_549;
  assign _T_554 = _T_552[0];
  assign _T_555 = _T_552[1];
  assign _T_556 = _T_552[2];
  assign _T_557 = _T_552[3];
  assign _T_558 = _T_552[4];
  assign _T_559 = _T_552[5];
  assign _T_560 = _T_552[6];
  assign _T_561 = _T_552[7];
  assign _T_563 = _T_506 ? _T_89_r_bits_last : 1'h1;
  assign _T_571 = _T_427_ready & _T_427_valid;
  assign _T_572 = _T_541 & _T_571;
  assign _T_573 = _T_554 & _T_563;
  assign _T_574 = _T_31_d_ready & _T_31_d_valid;
  assign _T_575 = _T_573 & _T_574;
  assign _T_576 = _T_566 + _T_572;
  assign _T_577 = _T_576[0:0];
  assign _T_578 = _T_577 - _T_575;
  assign _T_579 = $unsigned(_T_578);
  assign _T_580 = _T_579[0:0];
  assign _T_582 = _T_575 == 1'h0;
  assign _T_585 = _T_582 | _T_566;
  assign _T_587 = _T_585 | reset;
  assign _T_589 = _T_587 == 1'h0;
  assign _T_591 = _T_572 == 1'h0;
  assign _T_593 = _T_566 != 1'h1;
  assign _T_594 = _T_591 | _T_593;
  assign _T_596 = _T_594 | reset;
  assign _T_598 = _T_596 == 1'h0;
  assign _T_612 = _T_608 == 4'h0;
  assign _T_614 = _T_542 & _T_571;
  assign _T_615 = _T_555 & _T_563;
  assign _T_617 = _T_615 & _T_574;
  assign _GEN_78 = {{3'd0}, _T_614};
  assign _T_618 = _T_608 + _GEN_78;
  assign _T_619 = _T_618[3:0];
  assign _GEN_79 = {{3'd0}, _T_617};
  assign _T_620 = _T_619 - _GEN_79;
  assign _T_621 = $unsigned(_T_620);
  assign _T_622 = _T_621[3:0];
  assign _T_624 = _T_617 == 1'h0;
  assign _T_626 = _T_608 != 4'h0;
  assign _T_627 = _T_624 | _T_626;
  assign _T_629 = _T_627 | reset;
  assign _T_631 = _T_629 == 1'h0;
  assign _T_633 = _T_614 == 1'h0;
  assign _T_635 = _T_608 != 4'h8;
  assign _T_636 = _T_633 | _T_635;
  assign _T_638 = _T_636 | reset;
  assign _T_640 = _T_638 == 1'h0;
  assign _GEN_69 = _T_614 ? _T_427_bits_wen : _T_610;
  assign _T_641 = _T_610 != _T_427_bits_wen;
  assign _T_643 = _T_612 == 1'h0;
  assign _T_644 = _T_643 & _T_641;
  assign _T_646 = _T_608 == 4'h8;
  assign _T_647 = _T_644 | _T_646;
  assign _T_654 = _T_650 == 4'h0;
  assign _T_656 = _T_543 & _T_571;
  assign _T_657 = _T_556 & _T_563;
  assign _T_659 = _T_657 & _T_574;
  assign _GEN_80 = {{3'd0}, _T_656};
  assign _T_660 = _T_650 + _GEN_80;
  assign _T_661 = _T_660[3:0];
  assign _GEN_81 = {{3'd0}, _T_659};
  assign _T_662 = _T_661 - _GEN_81;
  assign _T_663 = $unsigned(_T_662);
  assign _T_664 = _T_663[3:0];
  assign _T_666 = _T_659 == 1'h0;
  assign _T_668 = _T_650 != 4'h0;
  assign _T_669 = _T_666 | _T_668;
  assign _T_671 = _T_669 | reset;
  assign _T_673 = _T_671 == 1'h0;
  assign _T_675 = _T_656 == 1'h0;
  assign _T_677 = _T_650 != 4'h8;
  assign _T_678 = _T_675 | _T_677;
  assign _T_680 = _T_678 | reset;
  assign _T_682 = _T_680 == 1'h0;
  assign _GEN_70 = _T_656 ? _T_427_bits_wen : _T_652;
  assign _T_683 = _T_652 != _T_427_bits_wen;
  assign _T_685 = _T_654 == 1'h0;
  assign _T_686 = _T_685 & _T_683;
  assign _T_688 = _T_650 == 4'h8;
  assign _T_689 = _T_686 | _T_688;
  assign _T_698 = _T_544 & _T_571;
  assign _T_699 = _T_557 & _T_563;
  assign _T_701 = _T_699 & _T_574;
  assign _T_702 = _T_692 + _T_698;
  assign _T_703 = _T_702[0:0];
  assign _T_704 = _T_703 - _T_701;
  assign _T_705 = $unsigned(_T_704);
  assign _T_706 = _T_705[0:0];
  assign _T_708 = _T_701 == 1'h0;
  assign _T_711 = _T_708 | _T_692;
  assign _T_713 = _T_711 | reset;
  assign _T_715 = _T_713 == 1'h0;
  assign _T_717 = _T_698 == 1'h0;
  assign _T_719 = _T_692 != 1'h1;
  assign _T_720 = _T_717 | _T_719;
  assign _T_722 = _T_720 | reset;
  assign _T_724 = _T_722 == 1'h0;
  assign _T_740 = _T_545 & _T_571;
  assign _T_741 = _T_558 & _T_563;
  assign _T_743 = _T_741 & _T_574;
  assign _T_744 = _T_734 + _T_740;
  assign _T_745 = _T_744[0:0];
  assign _T_746 = _T_745 - _T_743;
  assign _T_747 = $unsigned(_T_746);
  assign _T_748 = _T_747[0:0];
  assign _T_750 = _T_743 == 1'h0;
  assign _T_753 = _T_750 | _T_734;
  assign _T_755 = _T_753 | reset;
  assign _T_757 = _T_755 == 1'h0;
  assign _T_759 = _T_740 == 1'h0;
  assign _T_761 = _T_734 != 1'h1;
  assign _T_762 = _T_759 | _T_761;
  assign _T_764 = _T_762 | reset;
  assign _T_766 = _T_764 == 1'h0;
  assign _T_782 = _T_546 & _T_571;
  assign _T_783 = _T_559 & _T_563;
  assign _T_785 = _T_783 & _T_574;
  assign _T_786 = _T_776 + _T_782;
  assign _T_787 = _T_786[0:0];
  assign _T_788 = _T_787 - _T_785;
  assign _T_789 = $unsigned(_T_788);
  assign _T_790 = _T_789[0:0];
  assign _T_792 = _T_785 == 1'h0;
  assign _T_795 = _T_792 | _T_776;
  assign _T_797 = _T_795 | reset;
  assign _T_799 = _T_797 == 1'h0;
  assign _T_801 = _T_782 == 1'h0;
  assign _T_803 = _T_776 != 1'h1;
  assign _T_804 = _T_801 | _T_803;
  assign _T_806 = _T_804 | reset;
  assign _T_808 = _T_806 == 1'h0;
  assign _T_824 = _T_547 & _T_571;
  assign _T_825 = _T_560 & _T_563;
  assign _T_827 = _T_825 & _T_574;
  assign _T_828 = _T_818 + _T_824;
  assign _T_829 = _T_828[0:0];
  assign _T_830 = _T_829 - _T_827;
  assign _T_831 = $unsigned(_T_830);
  assign _T_832 = _T_831[0:0];
  assign _T_834 = _T_827 == 1'h0;
  assign _T_837 = _T_834 | _T_818;
  assign _T_839 = _T_837 | reset;
  assign _T_841 = _T_839 == 1'h0;
  assign _T_843 = _T_824 == 1'h0;
  assign _T_845 = _T_818 != 1'h1;
  assign _T_846 = _T_843 | _T_845;
  assign _T_848 = _T_846 | reset;
  assign _T_850 = _T_848 == 1'h0;
  assign _T_866 = _T_548 & _T_571;
  assign _T_867 = _T_561 & _T_563;
  assign _T_869 = _T_867 & _T_574;
  assign _T_870 = _T_860 + _T_866;
  assign _T_871 = _T_870[0:0];
  assign _T_872 = _T_871 - _T_869;
  assign _T_873 = $unsigned(_T_872);
  assign _T_874 = _T_873[0:0];
  assign _T_876 = _T_869 == 1'h0;
  assign _T_879 = _T_876 | _T_860;
  assign _T_881 = _T_879 | reset;
  assign _T_883 = _T_881 == 1'h0;
  assign _T_885 = _T_866 == 1'h0;
  assign _T_887 = _T_860 != 1'h1;
  assign _T_888 = _T_885 | _T_887;
  assign _T_890 = _T_888 | reset;
  assign _T_892 = _T_890 == 1'h0;
  assign auto_in_a_ready = _T_31_a_ready;
  assign auto_in_d_valid = _T_31_d_valid;
  assign auto_in_d_bits_opcode = _T_31_d_bits_opcode;
  assign auto_in_d_bits_size = _T_31_d_bits_size;
  assign auto_in_d_bits_source = _T_31_d_bits_source;
  assign auto_in_d_bits_data = _T_31_d_bits_data;
  assign auto_in_d_bits_error = _T_31_d_bits_error;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_lock = _T_89_aw_bits_lock;
  assign auto_out_aw_bits_cache = _T_89_aw_bits_cache;
  assign auto_out_aw_bits_prot = _T_89_aw_bits_prot;
  assign auto_out_aw_bits_qos = _T_89_aw_bits_qos;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_lock = _T_89_ar_bits_lock;
  assign auto_out_ar_bits_cache = _T_89_ar_bits_cache;
  assign auto_out_ar_bits_prot = _T_89_ar_bits_prot;
  assign auto_out_ar_bits_qos = _T_89_ar_bits_qos;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_a_ready = _T_484;
  assign _T_31_a_valid = auto_in_a_valid;
  assign _T_31_a_bits_opcode = auto_in_a_bits_opcode;
  assign _T_31_a_bits_size = auto_in_a_bits_size;
  assign _T_31_a_bits_source = auto_in_a_bits_source;
  assign _T_31_a_bits_address = auto_in_a_bits_address;
  assign _T_31_a_bits_mask = auto_in_a_bits_mask;
  assign _T_31_a_bits_data = auto_in_a_bits_data;
  assign _T_31_d_ready = auto_in_d_ready;
  assign _T_31_d_valid = _T_510;
  assign _T_31_d_bits_opcode = _T_536_opcode;
  assign _T_31_d_bits_size = _T_536_size;
  assign _T_31_d_bits_source = _T_536_source;
  assign _T_31_d_bits_data = _T_89_r_bits_data;
  assign _T_31_d_bits_error = _T_536_error;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_454;
  assign _T_89_aw_bits_id = _T_447_bits_id;
  assign _T_89_aw_bits_addr = _T_447_bits_addr;
  assign _T_89_aw_bits_len = _T_447_bits_len;
  assign _T_89_aw_bits_size = _T_447_bits_size;
  assign _T_89_aw_bits_burst = _T_447_bits_burst;
  assign _T_89_aw_bits_lock = _T_447_bits_lock;
  assign _T_89_aw_bits_cache = _T_447_bits_cache;
  assign _T_89_aw_bits_prot = _T_447_bits_prot;
  assign _T_89_aw_bits_qos = _T_447_bits_qos;
  assign _T_89_aw_bits_user = _T_447_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_439_valid;
  assign _T_89_w_bits_data = _T_439_bits_data;
  assign _T_89_w_bits_strb = _T_439_bits_strb;
  assign _T_89_w_bits_last = _T_439_bits_last;
  assign _T_89_b_ready = _T_509;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_453;
  assign _T_89_ar_bits_id = _T_447_bits_id;
  assign _T_89_ar_bits_addr = _T_447_bits_addr;
  assign _T_89_ar_bits_len = _T_447_bits_len;
  assign _T_89_ar_bits_size = _T_447_bits_size;
  assign _T_89_ar_bits_burst = _T_447_bits_burst;
  assign _T_89_ar_bits_lock = _T_447_bits_lock;
  assign _T_89_ar_bits_cache = _T_447_bits_cache;
  assign _T_89_ar_bits_prot = _T_447_bits_prot;
  assign _T_89_ar_bits_qos = _T_447_bits_qos;
  assign _T_89_ar_bits_user = _T_447_bits_user;
  assign _T_89_r_ready = _T_31_d_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign _T_206_0 = _T_319_4;
  assign _T_206_1 = _T_319_5;
  assign _T_206_2 = _T_319_6;
  assign _T_206_3 = _T_319_7;
  assign _T_206_4 = _T_319_3;
  assign _T_206_8 = _T_319_0;
  assign _T_206_16 = _T_319_1;
  assign _T_206_17 = _T_319_1;
  assign _T_206_18 = _T_319_1;
  assign _T_206_19 = _T_319_1;
  assign _T_206_20 = _T_319_1;
  assign _T_206_21 = _T_319_1;
  assign _T_206_22 = _T_319_1;
  assign _T_206_23 = _T_319_1;
  assign _T_206_24 = _T_319_2;
  assign _T_206_25 = _T_319_2;
  assign _T_206_26 = _T_319_2;
  assign _T_206_27 = _T_319_2;
  assign _T_206_28 = _T_319_2;
  assign _T_206_29 = _T_319_2;
  assign _T_206_30 = _T_319_2;
  assign _T_206_31 = _T_319_2;
  assign _T_319_0 = _T_566;
  assign _T_319_1 = _T_647;
  assign _T_319_2 = _T_689;
  assign _T_319_3 = _T_692;
  assign _T_319_4 = _T_734;
  assign _T_319_5 = _T_776;
  assign _T_319_6 = _T_818;
  assign _T_319_7 = _T_860;
  assign _T_427_ready = Queue_1_io_enq_ready;
  assign _T_427_valid = _T_493;
  assign _T_427_bits_id = _GEN_0;
  assign _T_427_bits_addr = _T_31_a_bits_address;
  assign _T_427_bits_len = _T_469;
  assign _T_427_bits_size = _T_471[2:0];
  assign _T_427_bits_user = _T_417;
  assign _T_427_bits_wen = _T_372;
  assign _T_431_ready = Queue_io_enq_ready;
  assign _T_431_valid = _T_499;
  assign _T_431_bits_data = _T_31_a_bits_data;
  assign _T_431_bits_strb = _T_31_a_bits_mask;
  assign _T_431_bits_last = _T_398;
  assign Queue_io_enq_valid = _T_431_valid;
  assign Queue_io_enq_bits_data = _T_431_bits_data;
  assign Queue_io_enq_bits_strb = _T_431_bits_strb;
  assign Queue_io_enq_bits_last = _T_431_bits_last;
  assign Queue_io_deq_ready = _T_439_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_439_ready = _T_89_w_ready;
  assign _T_439_valid = Queue_io_deq_valid;
  assign _T_439_bits_data = Queue_io_deq_bits_data;
  assign _T_439_bits_strb = Queue_io_deq_bits_strb;
  assign _T_439_bits_last = Queue_io_deq_bits_last;
  assign Queue_1_io_enq_valid = _T_427_valid;
  assign Queue_1_io_enq_bits_id = _T_427_bits_id;
  assign Queue_1_io_enq_bits_addr = _T_427_bits_addr;
  assign Queue_1_io_enq_bits_len = _T_427_bits_len;
  assign Queue_1_io_enq_bits_size = _T_427_bits_size;
  assign Queue_1_io_enq_bits_user = _T_427_bits_user;
  assign Queue_1_io_enq_bits_wen = _T_427_bits_wen;
  assign Queue_1_io_deq_ready = _T_447_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_447_ready = _T_455;
  assign _T_447_valid = Queue_1_io_deq_valid;
  assign _T_447_bits_id = Queue_1_io_deq_bits_id;
  assign _T_447_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_447_bits_len = Queue_1_io_deq_bits_len;
  assign _T_447_bits_size = Queue_1_io_deq_bits_size;
  assign _T_447_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_447_bits_lock = Queue_1_io_deq_bits_lock;
  assign _T_447_bits_cache = Queue_1_io_deq_bits_cache;
  assign _T_447_bits_prot = Queue_1_io_deq_bits_prot;
  assign _T_447_bits_qos = Queue_1_io_deq_bits_qos;
  assign _T_447_bits_user = Queue_1_io_deq_bits_user;
  assign _T_447_bits_wen = Queue_1_io_deq_bits_wen;
  assign _GEN_0 = _GEN_34;
  assign _GEN_1 = _GEN_65;
  assign _T_526_size = _T_419;
  assign _T_526_source = _T_418;
  assign _T_526_error = _T_521;
  assign _T_531_size = _T_421;
  assign _T_531_source = _T_420;
  assign _T_531_error = _T_514;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_387 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_459 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_502 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_517 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_566 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_608 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_610 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_650 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_652 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_692 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_734 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_776 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_818 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_860 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_387 <= 5'h0;
    end else begin
      if (_T_373) begin
        if (_T_393) begin
          if (_T_372) begin
            _T_387 <= _T_379;
          end else begin
            _T_387 <= 5'h0;
          end
        end else begin
          _T_387 <= _T_391;
        end
      end
    end
    if (reset) begin
      _T_459 <= 1'h0;
    end else begin
      if (_T_373) begin
        _T_459 <= _T_462;
      end
    end
    if (reset) begin
      _T_502 <= 1'h0;
    end else begin
      if (_T_503) begin
        _T_502 <= _T_505;
      end
    end
    if (reset) begin
      _T_517 <= 1'h0;
    end else begin
      if (_T_503) begin
        _T_517 <= _T_522;
      end
    end
    if (reset) begin
      _T_566 <= 1'h0;
    end else begin
      _T_566 <= _T_580;
    end
    if (reset) begin
      _T_608 <= 4'h0;
    end else begin
      _T_608 <= _T_622;
    end
    if (_T_614) begin
      _T_610 <= _T_427_bits_wen;
    end
    if (reset) begin
      _T_650 <= 4'h0;
    end else begin
      _T_650 <= _T_664;
    end
    if (_T_656) begin
      _T_652 <= _T_427_bits_wen;
    end
    if (reset) begin
      _T_692 <= 1'h0;
    end else begin
      _T_692 <= _T_706;
    end
    if (reset) begin
      _T_734 <= 1'h0;
    end else begin
      _T_734 <= _T_748;
    end
    if (reset) begin
      _T_776 <= 1'h0;
    end else begin
      _T_776 <= _T_790;
    end
    if (reset) begin
      _T_818 <= 1'h0;
    end else begin
      _T_818 <= _T_832;
    end
    if (reset) begin
      _T_860 <= 1'h0;
    end else begin
      _T_860 <= _T_874;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:106 assert (a_source  < UInt(BigInt(1) << sourceBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:107 assert (a_size    < UInt(BigInt(1) << sizeBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_589) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_589) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_598) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_598) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_631) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_631) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_640) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_640) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_682) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_682) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_715) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_715) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_724) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_724) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_757) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_757) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_766) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_766) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_799) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_799) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_808) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_808) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_841) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_841) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_850) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_850) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_883) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:210 assert (!dec || count =/= UInt(0))        // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_883) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_892) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:211 assert (!inc || count =/= UInt(maxCount)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_892) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module TLBuffer_SystemBus_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [2:0]  auto_out_d_bits_sink,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_error
);
  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [2:0] _T_31_a_bits_param;
  wire [3:0] _T_31_a_bits_size;
  wire [3:0] _T_31_a_bits_source;
  wire [31:0] _T_31_a_bits_address;
  wire [7:0] _T_31_a_bits_mask;
  wire [63:0] _T_31_a_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [3:0] _T_31_d_bits_size;
  wire [3:0] _T_31_d_bits_source;
  wire [63:0] _T_31_d_bits_data;
  wire  _T_31_d_bits_error;
  wire  _T_89_a_ready;
  wire  _T_89_a_valid;
  wire [2:0] _T_89_a_bits_opcode;
  wire [2:0] _T_89_a_bits_param;
  wire [3:0] _T_89_a_bits_size;
  wire [3:0] _T_89_a_bits_source;
  wire [31:0] _T_89_a_bits_address;
  wire [7:0] _T_89_a_bits_mask;
  wire [63:0] _T_89_a_bits_data;
  wire  _T_89_d_ready;
  wire  _T_89_d_valid;
  wire [2:0] _T_89_d_bits_opcode;
  wire [1:0] _T_89_d_bits_param;
  wire [3:0] _T_89_d_bits_size;
  wire [3:0] _T_89_d_bits_source;
  wire [2:0] _T_89_d_bits_sink;
  wire [63:0] _T_89_d_bits_data;
  wire  _T_89_d_bits_error;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [3:0] Queue_io_enq_bits_size;
  wire [3:0] Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [7:0] Queue_io_enq_bits_mask;
  wire [63:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [3:0] Queue_io_deq_bits_size;
  wire [3:0] Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [7:0] Queue_io_deq_bits_mask;
  wire [63:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [1:0] Queue_1_io_enq_bits_param;
  wire [3:0] Queue_1_io_enq_bits_size;
  wire [3:0] Queue_1_io_enq_bits_source;
  wire [2:0] Queue_1_io_enq_bits_sink;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [1:0] Queue_1_io_deq_bits_param;
  wire [3:0] Queue_1_io_deq_bits_size;
  wire [3:0] Queue_1_io_deq_bits_source;
  wire [2:0] Queue_1_io_deq_bits_sink;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  Queue_27 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_28 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  assign auto_in_a_ready = _T_31_a_ready;
  assign auto_in_d_valid = _T_31_d_valid;
  assign auto_in_d_bits_opcode = _T_31_d_bits_opcode;
  assign auto_in_d_bits_size = _T_31_d_bits_size;
  assign auto_in_d_bits_source = _T_31_d_bits_source;
  assign auto_in_d_bits_data = _T_31_d_bits_data;
  assign auto_in_d_bits_error = _T_31_d_bits_error;
  assign auto_out_a_valid = _T_89_a_valid;
  assign auto_out_a_bits_opcode = _T_89_a_bits_opcode;
  assign auto_out_a_bits_param = _T_89_a_bits_param;
  assign auto_out_a_bits_size = _T_89_a_bits_size;
  assign auto_out_a_bits_source = _T_89_a_bits_source;
  assign auto_out_a_bits_address = _T_89_a_bits_address;
  assign auto_out_a_bits_mask = _T_89_a_bits_mask;
  assign auto_out_a_bits_data = _T_89_a_bits_data;
  assign auto_out_d_ready = _T_89_d_ready;
  assign _T_31_a_ready = Queue_io_enq_ready;
  assign _T_31_a_valid = auto_in_a_valid;
  assign _T_31_a_bits_opcode = auto_in_a_bits_opcode;
  assign _T_31_a_bits_param = auto_in_a_bits_param;
  assign _T_31_a_bits_size = auto_in_a_bits_size;
  assign _T_31_a_bits_source = auto_in_a_bits_source;
  assign _T_31_a_bits_address = auto_in_a_bits_address;
  assign _T_31_a_bits_mask = auto_in_a_bits_mask;
  assign _T_31_a_bits_data = auto_in_a_bits_data;
  assign _T_31_d_ready = auto_in_d_ready;
  assign _T_31_d_valid = Queue_1_io_deq_valid;
  assign _T_31_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign _T_31_d_bits_size = Queue_1_io_deq_bits_size;
  assign _T_31_d_bits_source = Queue_1_io_deq_bits_source;
  assign _T_31_d_bits_data = Queue_1_io_deq_bits_data;
  assign _T_31_d_bits_error = Queue_1_io_deq_bits_error;
  assign _T_89_a_ready = auto_out_a_ready;
  assign _T_89_a_valid = Queue_io_deq_valid;
  assign _T_89_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign _T_89_a_bits_param = Queue_io_deq_bits_param;
  assign _T_89_a_bits_size = Queue_io_deq_bits_size;
  assign _T_89_a_bits_source = Queue_io_deq_bits_source;
  assign _T_89_a_bits_address = Queue_io_deq_bits_address;
  assign _T_89_a_bits_mask = Queue_io_deq_bits_mask;
  assign _T_89_a_bits_data = Queue_io_deq_bits_data;
  assign _T_89_d_ready = Queue_1_io_enq_ready;
  assign _T_89_d_valid = auto_out_d_valid;
  assign _T_89_d_bits_opcode = auto_out_d_bits_opcode;
  assign _T_89_d_bits_param = auto_out_d_bits_param;
  assign _T_89_d_bits_size = auto_out_d_bits_size;
  assign _T_89_d_bits_source = auto_out_d_bits_source;
  assign _T_89_d_bits_sink = auto_out_d_bits_sink;
  assign _T_89_d_bits_data = auto_out_d_bits_data;
  assign _T_89_d_bits_error = auto_out_d_bits_error;
  assign Queue_io_enq_valid = _T_31_a_valid;
  assign Queue_io_enq_bits_opcode = _T_31_a_bits_opcode;
  assign Queue_io_enq_bits_param = _T_31_a_bits_param;
  assign Queue_io_enq_bits_size = _T_31_a_bits_size;
  assign Queue_io_enq_bits_source = _T_31_a_bits_source;
  assign Queue_io_enq_bits_address = _T_31_a_bits_address;
  assign Queue_io_enq_bits_mask = _T_31_a_bits_mask;
  assign Queue_io_enq_bits_data = _T_31_a_bits_data;
  assign Queue_io_deq_ready = _T_89_a_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_89_d_valid;
  assign Queue_1_io_enq_bits_opcode = _T_89_d_bits_opcode;
  assign Queue_1_io_enq_bits_param = _T_89_d_bits_param;
  assign Queue_1_io_enq_bits_size = _T_89_d_bits_size;
  assign Queue_1_io_enq_bits_source = _T_89_d_bits_source;
  assign Queue_1_io_enq_bits_sink = _T_89_d_bits_sink;
  assign Queue_1_io_enq_bits_data = _T_89_d_bits_data;
  assign Queue_1_io_enq_bits_error = _T_89_d_bits_error;
  assign Queue_1_io_deq_ready = _T_31_d_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
endmodule
module TLWidthWidget_SystemBus(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_error
);
  wire  _T_31_a_ready;
  wire  _T_31_a_valid;
  wire [2:0] _T_31_a_bits_opcode;
  wire [2:0] _T_31_a_bits_param;
  wire [3:0] _T_31_a_bits_size;
  wire [3:0] _T_31_a_bits_source;
  wire [31:0] _T_31_a_bits_address;
  wire [7:0] _T_31_a_bits_mask;
  wire [63:0] _T_31_a_bits_data;
  wire  _T_31_d_ready;
  wire  _T_31_d_valid;
  wire [2:0] _T_31_d_bits_opcode;
  wire [3:0] _T_31_d_bits_size;
  wire [3:0] _T_31_d_bits_source;
  wire [63:0] _T_31_d_bits_data;
  wire  _T_31_d_bits_error;
  wire  _T_89_a_ready;
  wire  _T_89_a_valid;
  wire [2:0] _T_89_a_bits_opcode;
  wire [2:0] _T_89_a_bits_param;
  wire [3:0] _T_89_a_bits_size;
  wire [3:0] _T_89_a_bits_source;
  wire [31:0] _T_89_a_bits_address;
  wire [7:0] _T_89_a_bits_mask;
  wire [63:0] _T_89_a_bits_data;
  wire  _T_89_d_ready;
  wire  _T_89_d_valid;
  wire [2:0] _T_89_d_bits_opcode;
  wire [3:0] _T_89_d_bits_size;
  wire [3:0] _T_89_d_bits_source;
  wire [63:0] _T_89_d_bits_data;
  wire  _T_89_d_bits_error;
  assign auto_in_a_ready = _T_31_a_ready;
  assign auto_in_d_valid = _T_31_d_valid;
  assign auto_in_d_bits_opcode = _T_31_d_bits_opcode;
  assign auto_in_d_bits_size = _T_31_d_bits_size;
  assign auto_in_d_bits_source = _T_31_d_bits_source;
  assign auto_in_d_bits_data = _T_31_d_bits_data;
  assign auto_in_d_bits_error = _T_31_d_bits_error;
  assign auto_out_a_valid = _T_89_a_valid;
  assign auto_out_a_bits_opcode = _T_89_a_bits_opcode;
  assign auto_out_a_bits_param = _T_89_a_bits_param;
  assign auto_out_a_bits_size = _T_89_a_bits_size;
  assign auto_out_a_bits_source = _T_89_a_bits_source;
  assign auto_out_a_bits_address = _T_89_a_bits_address;
  assign auto_out_a_bits_mask = _T_89_a_bits_mask;
  assign auto_out_a_bits_data = _T_89_a_bits_data;
  assign auto_out_d_ready = _T_89_d_ready;
  assign _T_31_a_ready = _T_89_a_ready;
  assign _T_31_a_valid = auto_in_a_valid;
  assign _T_31_a_bits_opcode = auto_in_a_bits_opcode;
  assign _T_31_a_bits_param = auto_in_a_bits_param;
  assign _T_31_a_bits_size = auto_in_a_bits_size;
  assign _T_31_a_bits_source = auto_in_a_bits_source;
  assign _T_31_a_bits_address = auto_in_a_bits_address;
  assign _T_31_a_bits_mask = auto_in_a_bits_mask;
  assign _T_31_a_bits_data = auto_in_a_bits_data;
  assign _T_31_d_ready = auto_in_d_ready;
  assign _T_31_d_valid = _T_89_d_valid;
  assign _T_31_d_bits_opcode = _T_89_d_bits_opcode;
  assign _T_31_d_bits_size = _T_89_d_bits_size;
  assign _T_31_d_bits_source = _T_89_d_bits_source;
  assign _T_31_d_bits_data = _T_89_d_bits_data;
  assign _T_31_d_bits_error = _T_89_d_bits_error;
  assign _T_89_a_ready = auto_out_a_ready;
  assign _T_89_a_valid = _T_31_a_valid;
  assign _T_89_a_bits_opcode = _T_31_a_bits_opcode;
  assign _T_89_a_bits_param = _T_31_a_bits_param;
  assign _T_89_a_bits_size = _T_31_a_bits_size;
  assign _T_89_a_bits_source = _T_31_a_bits_source;
  assign _T_89_a_bits_address = _T_31_a_bits_address;
  assign _T_89_a_bits_mask = _T_31_a_bits_mask;
  assign _T_89_a_bits_data = _T_31_a_bits_data;
  assign _T_89_d_ready = _T_31_d_ready;
  assign _T_89_d_valid = auto_out_d_valid;
  assign _T_89_d_bits_opcode = auto_out_d_bits_opcode;
  assign _T_89_d_bits_size = auto_out_d_bits_size;
  assign _T_89_d_bits_source = auto_out_d_bits_source;
  assign _T_89_d_bits_data = auto_out_d_bits_data;
  assign _T_89_d_bits_error = auto_out_d_bits_error;
endmodule
module Queue_104(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire  ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_42_data;
  wire  ram_data__T_42_addr;
  wire [63:0] ram_data__T_33_data;
  wire  ram_data__T_33_addr;
  wire  ram_data__T_33_mask;
  wire  ram_data__T_33_en;
  reg [1:0] ram_resp [0:0];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_42_data;
  wire  ram_resp__T_42_addr;
  wire [1:0] ram_resp__T_33_data;
  wire  ram_resp__T_33_addr;
  wire  ram_resp__T_33_mask;
  wire  ram_resp__T_33_en;
  reg  ram_last [0:0];
  reg [31:0] _RAND_3;
  wire  ram_last__T_42_data;
  wire  ram_last__T_42_addr;
  wire  ram_last__T_33_data;
  wire  ram_last__T_33_addr;
  wire  ram_last__T_33_mask;
  wire  ram_last__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_4;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_7;
  wire  _T_38;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire [1:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_data__T_42_addr = 1'h0;
  assign ram_data__T_42_data = ram_data[ram_data__T_42_addr];
  assign ram_data__T_33_data = io_enq_bits_data;
  assign ram_data__T_33_addr = 1'h0;
  assign ram_data__T_33_mask = do_enq;
  assign ram_data__T_33_en = do_enq;
  assign ram_resp__T_42_addr = 1'h0;
  assign ram_resp__T_42_data = ram_resp[ram_resp__T_42_addr];
  assign ram_resp__T_33_data = io_enq_bits_resp;
  assign ram_resp__T_33_addr = 1'h0;
  assign ram_resp__T_33_mask = do_enq;
  assign ram_resp__T_33_en = do_enq;
  assign ram_last__T_42_addr = 1'h0;
  assign ram_last__T_42_data = ram_last[ram_last__T_42_addr];
  assign ram_last__T_33_data = io_enq_bits_last;
  assign ram_last__T_33_addr = 1'h0;
  assign ram_last__T_33_mask = do_enq;
  assign ram_last__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_7 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_8 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_10 = empty ? io_enq_bits_last : ram_last__T_42_data;
  assign _GEN_11 = empty ? io_enq_bits_resp : ram_resp__T_42_data;
  assign _GEN_12 = empty ? io_enq_bits_data : ram_data__T_42_data;
  assign _GEN_13 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_14 = empty ? 1'h0 : _T_30;
  assign _GEN_15 = empty ? _GEN_9 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_8;
  assign io_deq_bits_id = _GEN_13;
  assign io_deq_bits_data = _GEN_12;
  assign io_deq_bits_resp = _GEN_11;
  assign io_deq_bits_last = _GEN_10;
  assign do_enq = _GEN_15;
  assign do_deq = _GEN_14;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  maybe_full = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_data__T_33_en & ram_data__T_33_mask) begin
      ram_data[ram_data__T_33_addr] <= ram_data__T_33_data;
    end
    if(ram_resp__T_33_en & ram_resp__T_33_mask) begin
      ram_resp[ram_resp__T_33_addr] <= ram_resp__T_33_data;
    end
    if(ram_last__T_33_en & ram_last__T_33_mask) begin
      ram_last[ram_last__T_33_addr] <= ram_last__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_105(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire  ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [1:0] ram_resp [0:0];
  reg [31:0] _RAND_1;
  wire [1:0] ram_resp__T_42_data;
  wire  ram_resp__T_42_addr;
  wire [1:0] ram_resp__T_33_data;
  wire  ram_resp__T_33_addr;
  wire  ram_resp__T_33_mask;
  wire  ram_resp__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_2;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_5;
  wire  _T_38;
  wire  _GEN_6;
  wire  _GEN_7;
  wire [1:0] _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_resp__T_42_addr = 1'h0;
  assign ram_resp__T_42_data = ram_resp[ram_resp__T_42_addr];
  assign ram_resp__T_33_data = io_enq_bits_resp;
  assign ram_resp__T_33_addr = 1'h0;
  assign ram_resp__T_33_mask = do_enq;
  assign ram_resp__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_5 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_6 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_7 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_8 = empty ? io_enq_bits_resp : ram_resp__T_42_data;
  assign _GEN_9 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_10 = empty ? 1'h0 : _T_30;
  assign _GEN_11 = empty ? _GEN_7 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_6;
  assign io_deq_bits_id = _GEN_9;
  assign io_deq_bits_resp = _GEN_8;
  assign do_enq = _GEN_11;
  assign do_deq = _GEN_10;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  maybe_full = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_resp__T_33_en & ram_resp__T_33_mask) begin
      ram_resp[ram_resp__T_33_addr] <= ram_resp__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4ToTL(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_error
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire  _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire  _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire  _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire  _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_a_ready;
  wire  _T_89_a_valid;
  wire [2:0] _T_89_a_bits_opcode;
  wire [2:0] _T_89_a_bits_param;
  wire [3:0] _T_89_a_bits_size;
  wire [3:0] _T_89_a_bits_source;
  wire [31:0] _T_89_a_bits_address;
  wire [7:0] _T_89_a_bits_mask;
  wire [63:0] _T_89_a_bits_data;
  wire  _T_89_d_ready;
  wire  _T_89_d_valid;
  wire [2:0] _T_89_d_bits_opcode;
  wire [3:0] _T_89_d_bits_size;
  wire [3:0] _T_89_d_bits_source;
  wire [63:0] _T_89_d_bits_data;
  wire  _T_89_d_bits_error;
  wire  _T_203_ready;
  wire  _T_203_valid;
  wire [3:0] _T_203_bits_size;
  wire [3:0] _T_203_bits_source;
  wire [31:0] _T_203_bits_address;
  wire [7:0] _T_203_bits_mask;
  wire [15:0] _T_208;
  wire [22:0] _GEN_16;
  wire [22:0] _T_209;
  wire [14:0] _T_210;
  wire [15:0] _GEN_17;
  wire [15:0] _T_211;
  wire [15:0] _T_213;
  wire [15:0] _T_215;
  wire [15:0] _T_216;
  wire [15:0] _T_217;
  wire [7:0] _T_218;
  wire [7:0] _T_219;
  wire  _T_221;
  wire [7:0] _T_222;
  wire [3:0] _T_223;
  wire [3:0] _T_224;
  wire  _T_226;
  wire [3:0] _T_227;
  wire [1:0] _T_228;
  wire [1:0] _T_229;
  wire  _T_231;
  wire [1:0] _T_232;
  wire  _T_233;
  wire [1:0] _T_234;
  wire [2:0] _T_235;
  wire [3:0] _T_236;
  wire  _T_241;
  wire [31:0] _T_245;
  wire [32:0] _T_246;
  wire [32:0] _T_248;
  wire [32:0] _T_249;
  wire  _T_251;
  wire  _T_252;
  wire  _T_257;
  wire [31:0] _T_261;
  wire [32:0] _T_262;
  wire [32:0] _T_264;
  wire [32:0] _T_265;
  wire  _T_267;
  wire [31:0] _T_269;
  wire [32:0] _T_270;
  wire [32:0] _T_272;
  wire [32:0] _T_273;
  wire  _T_275;
  wire [32:0] _T_278;
  wire [32:0] _T_280;
  wire [32:0] _T_281;
  wire  _T_283;
  wire [31:0] _T_285;
  wire [32:0] _T_286;
  wire [32:0] _T_288;
  wire [32:0] _T_289;
  wire  _T_291;
  wire [31:0] _T_293;
  wire [32:0] _T_294;
  wire [32:0] _T_296;
  wire [32:0] _T_297;
  wire  _T_299;
  wire [31:0] _T_301;
  wire [32:0] _T_302;
  wire [32:0] _T_304;
  wire [32:0] _T_305;
  wire  _T_307;
  wire  _T_308;
  wire  _T_309;
  wire  _T_310;
  wire  _T_311;
  wire  _T_312;
  wire  _T_313;
  wire  _T_316;
  wire [2:0] _T_318;
  wire [13:0] _GEN_18;
  wire [13:0] _T_319;
  wire [31:0] _T_320;
  reg [2:0] _T_338_0;
  reg [31:0] _RAND_0;
  reg [2:0] _T_338_1;
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_0;
  wire [2:0] _GEN_4;
  wire [1:0] _T_352;
  wire [2:0] _T_354;
  wire [3:0] _T_355;
  wire  _T_357;
  wire [29:0] _T_360;
  wire [14:0] _T_361;
  wire [14:0] _T_362;
  wire  _T_363;
  wire  _T_364;
  wire  _T_366;
  wire  _T_368;
  wire [3:0] _T_450_size;
  wire [3:0] _T_450_source;
  wire [31:0] _T_450_address;
  wire [7:0] _T_450_mask;
  wire [1:0] _T_453;
  wire [3:0] _T_455;
  wire [2:0] _T_456;
  wire [2:0] _T_458;
  wire  _T_460;
  wire  _T_462;
  wire  _T_463;
  wire  _T_465;
  wire  _T_467;
  wire  _T_468;
  wire  _T_470;
  wire  _T_471;
  wire  _T_472;
  wire  _T_473;
  wire  _T_475;
  wire  _T_476;
  wire  _T_477;
  wire  _T_478;
  wire  _T_479;
  wire  _T_480;
  wire  _T_481;
  wire  _T_482;
  wire  _T_483;
  wire  _T_484;
  wire  _T_485;
  wire  _T_486;
  wire  _T_487;
  wire  _T_488;
  wire  _T_489;
  wire  _T_491;
  wire  _T_492;
  wire  _T_493;
  wire  _T_494;
  wire  _T_495;
  wire  _T_496;
  wire  _T_497;
  wire  _T_498;
  wire  _T_499;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire  _T_507;
  wire  _T_508;
  wire  _T_509;
  wire  _T_510;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_515;
  wire [1:0] _T_516;
  wire [1:0] _T_517;
  wire [3:0] _T_518;
  wire [1:0] _T_519;
  wire [1:0] _T_520;
  wire [3:0] _T_521;
  wire [7:0] _T_522;
  wire [1:0] _T_526;
  wire  _T_528;
  wire  _T_529;
  wire  _T_530;
  wire  _T_531;
  wire [3:0] _T_533;
  wire [2:0] _T_534;
  wire [2:0] _GEN_5;
  wire  _T_536;
  wire [3:0] _T_538;
  wire [2:0] _T_539;
  wire [2:0] _GEN_6;
  wire  _T_540_ready;
  wire  _T_540_valid;
  wire [3:0] _T_540_bits_size;
  wire [3:0] _T_540_bits_source;
  wire [31:0] _T_540_bits_address;
  wire [7:0] _T_540_bits_mask;
  wire [63:0] _T_540_bits_data;
  wire [15:0] _T_545;
  wire [22:0] _GEN_19;
  wire [22:0] _T_546;
  wire [14:0] _T_547;
  wire [15:0] _GEN_20;
  wire [15:0] _T_548;
  wire [15:0] _T_550;
  wire [15:0] _T_552;
  wire [15:0] _T_553;
  wire [15:0] _T_554;
  wire [7:0] _T_555;
  wire [7:0] _T_556;
  wire  _T_558;
  wire [7:0] _T_559;
  wire [3:0] _T_560;
  wire [3:0] _T_561;
  wire  _T_563;
  wire [3:0] _T_564;
  wire [1:0] _T_565;
  wire [1:0] _T_566;
  wire  _T_568;
  wire [1:0] _T_569;
  wire  _T_570;
  wire [1:0] _T_571;
  wire [2:0] _T_572;
  wire [3:0] _T_573;
  wire  _T_578;
  wire [31:0] _T_582;
  wire [32:0] _T_583;
  wire [32:0] _T_585;
  wire [32:0] _T_586;
  wire  _T_588;
  wire  _T_589;
  wire  _T_594;
  wire [31:0] _T_598;
  wire [32:0] _T_599;
  wire [32:0] _T_601;
  wire [32:0] _T_602;
  wire  _T_604;
  wire [31:0] _T_606;
  wire [32:0] _T_607;
  wire [32:0] _T_609;
  wire [32:0] _T_610;
  wire  _T_612;
  wire [32:0] _T_615;
  wire [32:0] _T_617;
  wire [32:0] _T_618;
  wire  _T_620;
  wire [31:0] _T_622;
  wire [32:0] _T_623;
  wire [32:0] _T_625;
  wire [32:0] _T_626;
  wire  _T_628;
  wire  _T_629;
  wire  _T_630;
  wire  _T_631;
  wire  _T_632;
  wire  _T_637;
  wire [31:0] _T_641;
  wire [32:0] _T_642;
  wire [32:0] _T_644;
  wire [32:0] _T_645;
  wire  _T_647;
  wire  _T_648;
  wire  _T_663;
  wire  _T_664;
  wire [2:0] _T_667;
  wire [13:0] _GEN_21;
  wire [13:0] _T_668;
  wire [31:0] _T_669;
  reg [2:0] _T_687_0;
  reg [31:0] _RAND_2;
  reg [2:0] _T_687_1;
  reg [31:0] _RAND_3;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_7;
  wire [1:0] _T_701;
  wire [2:0] _T_703;
  wire [3:0] _T_704;
  wire  _T_706;
  wire [29:0] _T_709;
  wire [14:0] _T_710;
  wire [14:0] _T_711;
  wire  _T_712;
  wire  _T_713;
  wire  _T_715;
  wire  _T_717;
  wire  _T_721;
  wire  _T_722;
  wire  _T_724;
  wire  _T_725;
  wire  _T_727;
  wire  _T_729;
  wire  _T_730;
  wire  _T_731;
  wire  _T_732;
  wire  _T_733;
  wire [3:0] _T_827_size;
  wire [3:0] _T_827_source;
  wire [31:0] _T_827_address;
  wire [7:0] _T_827_mask;
  wire [63:0] _T_827_data;
  wire [1:0] _T_832;
  wire  _T_834;
  wire  _T_835;
  wire  _T_836;
  wire  _T_837;
  wire [3:0] _T_839;
  wire [2:0] _T_840;
  wire [2:0] _GEN_8;
  wire  _T_842;
  wire [3:0] _T_844;
  wire [2:0] _T_845;
  wire [2:0] _GEN_9;
  reg [7:0] _T_849;
  reg [31:0] _RAND_4;
  wire  _T_851;
  wire  _T_852;
  wire [1:0] _T_853;
  wire  _T_855;
  wire  _T_857;
  wire  _T_859;
  reg [1:0] _T_863;
  reg [31:0] _RAND_5;
  wire [1:0] _T_864;
  wire [1:0] _T_865;
  wire [3:0] _T_866;
  wire [2:0] _T_867;
  wire [3:0] _GEN_22;
  wire [3:0] _T_868;
  wire [2:0] _T_870;
  wire [3:0] _GEN_23;
  wire [3:0] _T_871;
  wire [3:0] _GEN_24;
  wire [3:0] _T_872;
  wire [1:0] _T_873;
  wire [1:0] _T_874;
  wire [1:0] _T_875;
  wire [1:0] _T_876;
  wire  _T_878;
  wire  _T_879;
  wire [1:0] _T_880;
  wire [2:0] _GEN_25;
  wire [2:0] _T_881;
  wire [1:0] _T_882;
  wire [1:0] _T_883;
  wire [1:0] _GEN_10;
  wire  _T_886;
  wire  _T_887;
  wire  _T_890_0;
  wire  _T_890_1;
  wire  _T_895;
  wire  _T_896;
  wire  _T_899_0;
  wire  _T_899_1;
  wire  _T_906;
  wire  _T_910;
  wire  _T_915;
  wire  _T_916;
  wire  _T_919;
  wire  _T_921;
  wire  _T_922;
  wire  _T_924;
  wire  _T_926;
  wire  _T_928;
  wire  _T_930;
  wire [7:0] _T_934;
  wire  _T_936;
  wire [7:0] _GEN_26;
  wire [8:0] _T_937;
  wire [8:0] _T_938;
  wire [7:0] _T_939;
  wire [7:0] _T_940;
  reg  _T_958_0;
  reg [31:0] _RAND_6;
  reg  _T_958_1;
  reg [31:0] _RAND_7;
  wire  _T_969_0;
  wire  _T_969_1;
  wire  _T_977_0;
  wire  _T_977_1;
  wire  _T_985;
  wire  _T_986;
  wire  _T_990;
  wire  _T_992;
  wire  _T_993;
  wire  _T_995;
  wire  _T_996;
  wire [39:0] _T_998;
  wire [103:0] _T_999;
  wire [7:0] _T_1000;
  wire [13:0] _T_1002;
  wire [117:0] _T_1003;
  wire [117:0] _T_1005;
  wire [39:0] _T_1006;
  wire [103:0] _T_1007;
  wire [7:0] _T_1008;
  wire [13:0] _T_1010;
  wire [117:0] _T_1011;
  wire [117:0] _T_1013;
  wire [117:0] _T_1014;
  wire [2:0] _T_1016_opcode;
  wire [2:0] _T_1016_param;
  wire [3:0] _T_1016_size;
  wire [3:0] _T_1016_source;
  wire [31:0] _T_1016_address;
  wire [7:0] _T_1016_mask;
  wire [63:0] _T_1016_data;
  wire [117:0] _T_1018;
  wire [63:0] _T_1019;
  wire [7:0] _T_1020;
  wire [31:0] _T_1021;
  wire [3:0] _T_1022;
  wire [3:0] _T_1023;
  wire [2:0] _T_1024;
  wire [2:0] _T_1025;
  wire  _T_1026_ready;
  wire  _T_1026_valid;
  wire  _T_1026_bits_id;
  wire [1:0] _T_1026_bits_resp;
  wire  _T_1030_ready;
  wire  _T_1030_valid;
  wire  _T_1030_bits_id;
  wire [63:0] _T_1030_bits_data;
  wire [1:0] _T_1030_bits_resp;
  wire  _T_1030_bits_last;
  wire [1:0] _T_1036;
  wire  _T_1037;
  wire  _T_1038;
  wire [26:0] _T_1041;
  wire [11:0] _T_1042;
  wire [11:0] _T_1043;
  wire [8:0] _T_1044;
  wire [8:0] _T_1047;
  reg [8:0] _T_1050;
  reg [31:0] _RAND_8;
  wire [9:0] _T_1052;
  wire [9:0] _T_1053;
  wire [8:0] _T_1054;
  wire  _T_1056;
  wire  _T_1058;
  wire  _T_1060;
  wire  _T_1061;
  wire [8:0] _T_1065;
  wire [8:0] _GEN_11;
  wire  _T_1066;
  wire  _T_1067;
  wire  _T_1069;
  wire  _T_1070;
  wire  _T_1071;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits_id;
  wire [63:0] Queue_io_enq_bits_data;
  wire [1:0] Queue_io_enq_bits_resp;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits_id;
  wire [63:0] Queue_io_deq_bits_data;
  wire [1:0] Queue_io_deq_bits_resp;
  wire  Queue_io_deq_bits_last;
  wire  _T_1076_ready;
  wire  _T_1076_valid;
  wire  _T_1076_bits_id;
  wire [63:0] _T_1076_bits_data;
  wire [1:0] _T_1076_bits_resp;
  wire  _T_1076_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_id;
  wire [1:0] Queue_1_io_enq_bits_resp;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_id;
  wire [1:0] Queue_1_io_deq_bits_resp;
  wire  _T_1085_ready;
  wire  _T_1085_valid;
  wire  _T_1085_bits_id;
  wire [1:0] _T_1085_bits_resp;
  reg [2:0] _T_1106_0;
  reg [31:0] _RAND_9;
  reg [2:0] _T_1106_1;
  reg [31:0] _RAND_10;
  wire [2:0] _GEN_2;
  wire [2:0] _GEN_12;
  wire [2:0] _GEN_3;
  wire [2:0] _GEN_13;
  wire  _T_1123;
  wire [1:0] _T_1126;
  wire  _T_1128;
  wire  _T_1129;
  wire  _T_1130;
  wire  _T_1131;
  wire [3:0] _T_1133;
  wire [2:0] _T_1134;
  wire [2:0] _GEN_14;
  wire  _T_1136;
  wire [3:0] _T_1138;
  wire [2:0] _T_1139;
  wire [2:0] _GEN_15;
  wire  _T_1140;
  wire  _T_1141;
  Queue_104 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_105 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp)
  );
  assign _T_208 = {_T_31_ar_bits_len,8'hff};
  assign _GEN_16 = {{7'd0}, _T_208};
  assign _T_209 = _GEN_16 << _T_31_ar_bits_size;
  assign _T_210 = _T_209[22:8];
  assign _GEN_17 = {{1'd0}, _T_210};
  assign _T_211 = _GEN_17 << 1;
  assign _T_213 = _T_211 | 16'h1;
  assign _T_215 = {1'h0,_T_210};
  assign _T_216 = ~ _T_215;
  assign _T_217 = _T_213 & _T_216;
  assign _T_218 = _T_217[15:8];
  assign _T_219 = _T_217[7:0];
  assign _T_221 = _T_218 != 8'h0;
  assign _T_222 = _T_218 | _T_219;
  assign _T_223 = _T_222[7:4];
  assign _T_224 = _T_222[3:0];
  assign _T_226 = _T_223 != 4'h0;
  assign _T_227 = _T_223 | _T_224;
  assign _T_228 = _T_227[3:2];
  assign _T_229 = _T_227[1:0];
  assign _T_231 = _T_228 != 2'h0;
  assign _T_232 = _T_228 | _T_229;
  assign _T_233 = _T_232[1];
  assign _T_234 = {_T_231,_T_233};
  assign _T_235 = {_T_226,_T_234};
  assign _T_236 = {_T_221,_T_235};
  assign _T_241 = _T_236 <= 4'hc;
  assign _T_245 = _T_31_ar_bits_addr ^ 32'h3000;
  assign _T_246 = {1'b0,$signed(_T_245)};
  assign _T_248 = $signed(_T_246) & $signed(-33'sh1000);
  assign _T_249 = $signed(_T_248);
  assign _T_251 = $signed(_T_249) == $signed(33'sh0);
  assign _T_252 = _T_241 & _T_251;
  assign _T_257 = _T_236 <= 4'h6;
  assign _T_261 = _T_31_ar_bits_addr ^ 32'hc000000;
  assign _T_262 = {1'b0,$signed(_T_261)};
  assign _T_264 = $signed(_T_262) & $signed(-33'sh4000000);
  assign _T_265 = $signed(_T_264);
  assign _T_267 = $signed(_T_265) == $signed(33'sh0);
  assign _T_269 = _T_31_ar_bits_addr ^ 32'h2000000;
  assign _T_270 = {1'b0,$signed(_T_269)};
  assign _T_272 = $signed(_T_270) & $signed(-33'sh10000);
  assign _T_273 = $signed(_T_272);
  assign _T_275 = $signed(_T_273) == $signed(33'sh0);
  assign _T_278 = {1'b0,$signed(_T_31_ar_bits_addr)};
  assign _T_280 = $signed(_T_278) & $signed(-33'sh1000);
  assign _T_281 = $signed(_T_280);
  assign _T_283 = $signed(_T_281) == $signed(33'sh0);
  assign _T_285 = _T_31_ar_bits_addr ^ 32'h10000;
  assign _T_286 = {1'b0,$signed(_T_285)};
  assign _T_288 = $signed(_T_286) & $signed(-33'sh10000);
  assign _T_289 = $signed(_T_288);
  assign _T_291 = $signed(_T_289) == $signed(33'sh0);
  assign _T_293 = _T_31_ar_bits_addr ^ 32'h60000000;
  assign _T_294 = {1'b0,$signed(_T_293)};
  assign _T_296 = $signed(_T_294) & $signed(-33'sh20000000);
  assign _T_297 = $signed(_T_296);
  assign _T_299 = $signed(_T_297) == $signed(33'sh0);
  assign _T_301 = _T_31_ar_bits_addr ^ 32'h80000000;
  assign _T_302 = {1'b0,$signed(_T_301)};
  assign _T_304 = $signed(_T_302) & $signed(-33'sh10000000);
  assign _T_305 = $signed(_T_304);
  assign _T_307 = $signed(_T_305) == $signed(33'sh0);
  assign _T_308 = _T_267 | _T_275;
  assign _T_309 = _T_308 | _T_283;
  assign _T_310 = _T_309 | _T_291;
  assign _T_311 = _T_310 | _T_299;
  assign _T_312 = _T_311 | _T_307;
  assign _T_313 = _T_257 & _T_312;
  assign _T_316 = _T_252 | _T_313;
  assign _T_318 = _T_31_ar_bits_addr[2:0];
  assign _GEN_18 = {{11'd0}, _T_318};
  assign _T_319 = 14'h3000 | _GEN_18;
  assign _T_320 = _T_316 ? _T_31_ar_bits_addr : {{18'd0}, _T_319};
  assign _GEN_4 = _T_31_ar_bits_id ? _T_338_1 : _T_338_0;
  assign _T_352 = _GEN_0[1:0];
  assign _T_354 = {_T_31_ar_bits_id,_T_352};
  assign _T_355 = {_T_354,1'h0};
  assign _T_357 = _T_31_ar_valid == 1'h0;
  assign _T_360 = 30'h7fff << _T_236;
  assign _T_361 = _T_360[14:0];
  assign _T_362 = ~ _T_361;
  assign _T_363 = _T_210 == _T_362;
  assign _T_364 = _T_357 | _T_363;
  assign _T_366 = _T_364 | reset;
  assign _T_368 = _T_366 == 1'h0;
  assign _T_453 = _T_236[1:0];
  assign _T_455 = 4'h1 << _T_453;
  assign _T_456 = _T_455[2:0];
  assign _T_458 = _T_456 | 3'h1;
  assign _T_460 = _T_236 >= 4'h3;
  assign _T_462 = _T_458[2];
  assign _T_463 = _T_320[2];
  assign _T_465 = _T_463 == 1'h0;
  assign _T_467 = _T_462 & _T_465;
  assign _T_468 = _T_460 | _T_467;
  assign _T_470 = _T_462 & _T_463;
  assign _T_471 = _T_460 | _T_470;
  assign _T_472 = _T_458[1];
  assign _T_473 = _T_320[1];
  assign _T_475 = _T_473 == 1'h0;
  assign _T_476 = _T_465 & _T_475;
  assign _T_477 = _T_472 & _T_476;
  assign _T_478 = _T_468 | _T_477;
  assign _T_479 = _T_465 & _T_473;
  assign _T_480 = _T_472 & _T_479;
  assign _T_481 = _T_468 | _T_480;
  assign _T_482 = _T_463 & _T_475;
  assign _T_483 = _T_472 & _T_482;
  assign _T_484 = _T_471 | _T_483;
  assign _T_485 = _T_463 & _T_473;
  assign _T_486 = _T_472 & _T_485;
  assign _T_487 = _T_471 | _T_486;
  assign _T_488 = _T_458[0];
  assign _T_489 = _T_320[0];
  assign _T_491 = _T_489 == 1'h0;
  assign _T_492 = _T_476 & _T_491;
  assign _T_493 = _T_488 & _T_492;
  assign _T_494 = _T_478 | _T_493;
  assign _T_495 = _T_476 & _T_489;
  assign _T_496 = _T_488 & _T_495;
  assign _T_497 = _T_478 | _T_496;
  assign _T_498 = _T_479 & _T_491;
  assign _T_499 = _T_488 & _T_498;
  assign _T_500 = _T_481 | _T_499;
  assign _T_501 = _T_479 & _T_489;
  assign _T_502 = _T_488 & _T_501;
  assign _T_503 = _T_481 | _T_502;
  assign _T_504 = _T_482 & _T_491;
  assign _T_505 = _T_488 & _T_504;
  assign _T_506 = _T_484 | _T_505;
  assign _T_507 = _T_482 & _T_489;
  assign _T_508 = _T_488 & _T_507;
  assign _T_509 = _T_484 | _T_508;
  assign _T_510 = _T_485 & _T_491;
  assign _T_511 = _T_488 & _T_510;
  assign _T_512 = _T_487 | _T_511;
  assign _T_513 = _T_485 & _T_489;
  assign _T_514 = _T_488 & _T_513;
  assign _T_515 = _T_487 | _T_514;
  assign _T_516 = {_T_497,_T_494};
  assign _T_517 = {_T_503,_T_500};
  assign _T_518 = {_T_517,_T_516};
  assign _T_519 = {_T_509,_T_506};
  assign _T_520 = {_T_515,_T_512};
  assign _T_521 = {_T_520,_T_519};
  assign _T_522 = {_T_521,_T_518};
  assign _T_526 = 2'h1 << _T_31_ar_bits_id;
  assign _T_528 = _T_526[0];
  assign _T_529 = _T_526[1];
  assign _T_530 = _T_31_ar_ready & _T_31_ar_valid;
  assign _T_531 = _T_530 & _T_528;
  assign _T_533 = _T_338_0 + 3'h1;
  assign _T_534 = _T_533[2:0];
  assign _GEN_5 = _T_531 ? _T_534 : _T_338_0;
  assign _T_536 = _T_530 & _T_529;
  assign _T_538 = _T_338_1 + 3'h1;
  assign _T_539 = _T_538[2:0];
  assign _GEN_6 = _T_536 ? _T_539 : _T_338_1;
  assign _T_545 = {_T_31_aw_bits_len,8'hff};
  assign _GEN_19 = {{7'd0}, _T_545};
  assign _T_546 = _GEN_19 << _T_31_aw_bits_size;
  assign _T_547 = _T_546[22:8];
  assign _GEN_20 = {{1'd0}, _T_547};
  assign _T_548 = _GEN_20 << 1;
  assign _T_550 = _T_548 | 16'h1;
  assign _T_552 = {1'h0,_T_547};
  assign _T_553 = ~ _T_552;
  assign _T_554 = _T_550 & _T_553;
  assign _T_555 = _T_554[15:8];
  assign _T_556 = _T_554[7:0];
  assign _T_558 = _T_555 != 8'h0;
  assign _T_559 = _T_555 | _T_556;
  assign _T_560 = _T_559[7:4];
  assign _T_561 = _T_559[3:0];
  assign _T_563 = _T_560 != 4'h0;
  assign _T_564 = _T_560 | _T_561;
  assign _T_565 = _T_564[3:2];
  assign _T_566 = _T_564[1:0];
  assign _T_568 = _T_565 != 2'h0;
  assign _T_569 = _T_565 | _T_566;
  assign _T_570 = _T_569[1];
  assign _T_571 = {_T_568,_T_570};
  assign _T_572 = {_T_563,_T_571};
  assign _T_573 = {_T_558,_T_572};
  assign _T_578 = _T_573 <= 4'hc;
  assign _T_582 = _T_31_aw_bits_addr ^ 32'h3000;
  assign _T_583 = {1'b0,$signed(_T_582)};
  assign _T_585 = $signed(_T_583) & $signed(-33'sh1000);
  assign _T_586 = $signed(_T_585);
  assign _T_588 = $signed(_T_586) == $signed(33'sh0);
  assign _T_589 = _T_578 & _T_588;
  assign _T_594 = _T_573 <= 4'h6;
  assign _T_598 = _T_31_aw_bits_addr ^ 32'hc000000;
  assign _T_599 = {1'b0,$signed(_T_598)};
  assign _T_601 = $signed(_T_599) & $signed(-33'sh4000000);
  assign _T_602 = $signed(_T_601);
  assign _T_604 = $signed(_T_602) == $signed(33'sh0);
  assign _T_606 = _T_31_aw_bits_addr ^ 32'h2000000;
  assign _T_607 = {1'b0,$signed(_T_606)};
  assign _T_609 = $signed(_T_607) & $signed(-33'sh10000);
  assign _T_610 = $signed(_T_609);
  assign _T_612 = $signed(_T_610) == $signed(33'sh0);
  assign _T_615 = {1'b0,$signed(_T_31_aw_bits_addr)};
  assign _T_617 = $signed(_T_615) & $signed(-33'sh1000);
  assign _T_618 = $signed(_T_617);
  assign _T_620 = $signed(_T_618) == $signed(33'sh0);
  assign _T_622 = _T_31_aw_bits_addr ^ 32'h80000000;
  assign _T_623 = {1'b0,$signed(_T_622)};
  assign _T_625 = $signed(_T_623) & $signed(-33'sh10000000);
  assign _T_626 = $signed(_T_625);
  assign _T_628 = $signed(_T_626) == $signed(33'sh0);
  assign _T_629 = _T_604 | _T_612;
  assign _T_630 = _T_629 | _T_620;
  assign _T_631 = _T_630 | _T_628;
  assign _T_632 = _T_594 & _T_631;
  assign _T_637 = _T_573 <= 4'h8;
  assign _T_641 = _T_31_aw_bits_addr ^ 32'h60000000;
  assign _T_642 = {1'b0,$signed(_T_641)};
  assign _T_644 = $signed(_T_642) & $signed(-33'sh20000000);
  assign _T_645 = $signed(_T_644);
  assign _T_647 = $signed(_T_645) == $signed(33'sh0);
  assign _T_648 = _T_637 & _T_647;
  assign _T_663 = _T_589 | _T_632;
  assign _T_664 = _T_663 | _T_648;
  assign _T_667 = _T_31_aw_bits_addr[2:0];
  assign _GEN_21 = {{11'd0}, _T_667};
  assign _T_668 = 14'h3000 | _GEN_21;
  assign _T_669 = _T_664 ? _T_31_aw_bits_addr : {{18'd0}, _T_668};
  assign _GEN_7 = _T_31_aw_bits_id ? _T_687_1 : _T_687_0;
  assign _T_701 = _GEN_1[1:0];
  assign _T_703 = {_T_31_aw_bits_id,_T_701};
  assign _T_704 = {_T_703,1'h1};
  assign _T_706 = _T_31_aw_valid == 1'h0;
  assign _T_709 = 30'h7fff << _T_573;
  assign _T_710 = _T_709[14:0];
  assign _T_711 = ~ _T_710;
  assign _T_712 = _T_547 == _T_711;
  assign _T_713 = _T_706 | _T_712;
  assign _T_715 = _T_713 | reset;
  assign _T_717 = _T_715 == 1'h0;
  assign _T_721 = _T_31_aw_bits_len == 8'h0;
  assign _T_722 = _T_706 | _T_721;
  assign _T_724 = _T_31_aw_bits_size == 3'h3;
  assign _T_725 = _T_722 | _T_724;
  assign _T_727 = _T_725 | reset;
  assign _T_729 = _T_727 == 1'h0;
  assign _T_730 = _T_540_ready & _T_31_w_valid;
  assign _T_731 = _T_730 & _T_31_w_bits_last;
  assign _T_732 = _T_540_ready & _T_31_aw_valid;
  assign _T_733 = _T_31_aw_valid & _T_31_w_valid;
  assign _T_832 = 2'h1 << _T_31_aw_bits_id;
  assign _T_834 = _T_832[0];
  assign _T_835 = _T_832[1];
  assign _T_836 = _T_31_aw_ready & _T_31_aw_valid;
  assign _T_837 = _T_836 & _T_834;
  assign _T_839 = _T_687_0 + 3'h1;
  assign _T_840 = _T_839[2:0];
  assign _GEN_8 = _T_837 ? _T_840 : _T_687_0;
  assign _T_842 = _T_836 & _T_835;
  assign _T_844 = _T_687_1 + 3'h1;
  assign _T_845 = _T_844[2:0];
  assign _GEN_9 = _T_842 ? _T_845 : _T_687_1;
  assign _T_851 = _T_849 == 8'h0;
  assign _T_852 = _T_851 & _T_89_a_ready;
  assign _T_853 = {_T_540_valid,_T_203_valid};
  assign _T_855 = _T_853 == _T_853;
  assign _T_857 = _T_855 | reset;
  assign _T_859 = _T_857 == 1'h0;
  assign _T_864 = ~ _T_863;
  assign _T_865 = _T_853 & _T_864;
  assign _T_866 = {_T_865,_T_853};
  assign _T_867 = _T_866[3:1];
  assign _GEN_22 = {{1'd0}, _T_867};
  assign _T_868 = _T_866 | _GEN_22;
  assign _T_870 = _T_868[3:1];
  assign _GEN_23 = {{2'd0}, _T_863};
  assign _T_871 = _GEN_23 << 2;
  assign _GEN_24 = {{1'd0}, _T_870};
  assign _T_872 = _GEN_24 | _T_871;
  assign _T_873 = _T_872[3:2];
  assign _T_874 = _T_872[1:0];
  assign _T_875 = _T_873 & _T_874;
  assign _T_876 = ~ _T_875;
  assign _T_878 = _T_853 != 2'h0;
  assign _T_879 = _T_852 & _T_878;
  assign _T_880 = _T_876 & _T_853;
  assign _GEN_25 = {{1'd0}, _T_880};
  assign _T_881 = _GEN_25 << 1;
  assign _T_882 = _T_881[1:0];
  assign _T_883 = _T_880 | _T_882;
  assign _GEN_10 = _T_879 ? _T_883 : _T_863;
  assign _T_886 = _T_876[0];
  assign _T_887 = _T_876[1];
  assign _T_895 = _T_890_0 & _T_203_valid;
  assign _T_896 = _T_890_1 & _T_540_valid;
  assign _T_906 = _T_899_0 | _T_899_1;
  assign _T_910 = _T_899_0 == 1'h0;
  assign _T_915 = _T_899_1 == 1'h0;
  assign _T_916 = _T_910 | _T_915;
  assign _T_919 = _T_916 | reset;
  assign _T_921 = _T_919 == 1'h0;
  assign _T_922 = _T_203_valid | _T_540_valid;
  assign _T_924 = _T_922 == 1'h0;
  assign _T_926 = _T_924 | _T_906;
  assign _T_928 = _T_926 | reset;
  assign _T_930 = _T_928 == 1'h0;
  assign _T_934 = _T_899_1 ? _T_31_aw_bits_len : 8'h0;
  assign _T_936 = _T_89_a_ready & _T_89_a_valid;
  assign _GEN_26 = {{7'd0}, _T_936};
  assign _T_937 = _T_849 - _GEN_26;
  assign _T_938 = $unsigned(_T_937);
  assign _T_939 = _T_938[7:0];
  assign _T_940 = _T_852 ? _T_934 : _T_939;
  assign _T_969_0 = _T_851 ? _T_899_0 : _T_958_0;
  assign _T_969_1 = _T_851 ? _T_899_1 : _T_958_1;
  assign _T_977_0 = _T_851 ? _T_890_0 : _T_958_0;
  assign _T_977_1 = _T_851 ? _T_890_1 : _T_958_1;
  assign _T_985 = _T_89_a_ready & _T_977_0;
  assign _T_986 = _T_89_a_ready & _T_977_1;
  assign _T_990 = _T_958_0 ? _T_203_valid : 1'h0;
  assign _T_992 = _T_958_1 ? _T_540_valid : 1'h0;
  assign _T_993 = _T_990 | _T_992;
  assign _T_996 = _T_851 ? _T_922 : _T_995;
  assign _T_998 = {_T_203_bits_address,_T_203_bits_mask};
  assign _T_999 = {_T_998,64'h0};
  assign _T_1000 = {_T_203_bits_size,_T_203_bits_source};
  assign _T_1002 = {6'h20,_T_1000};
  assign _T_1003 = {_T_1002,_T_999};
  assign _T_1005 = _T_969_0 ? _T_1003 : 118'h0;
  assign _T_1006 = {_T_540_bits_address,_T_540_bits_mask};
  assign _T_1007 = {_T_1006,_T_540_bits_data};
  assign _T_1008 = {_T_540_bits_size,_T_540_bits_source};
  assign _T_1010 = {6'h8,_T_1008};
  assign _T_1011 = {_T_1010,_T_1007};
  assign _T_1013 = _T_969_1 ? _T_1011 : 118'h0;
  assign _T_1014 = _T_1005 | _T_1013;
  assign _T_1019 = _T_1018[63:0];
  assign _T_1020 = _T_1018[71:64];
  assign _T_1021 = _T_1018[103:72];
  assign _T_1022 = _T_1018[107:104];
  assign _T_1023 = _T_1018[111:108];
  assign _T_1024 = _T_1018[114:112];
  assign _T_1025 = _T_1018[117:115];
  assign _T_1036 = _T_89_d_bits_error ? 2'h2 : 2'h0;
  assign _T_1037 = _T_89_d_bits_opcode[0];
  assign _T_1038 = _T_89_d_ready & _T_89_d_valid;
  assign _T_1041 = 27'hfff << _T_89_d_bits_size;
  assign _T_1042 = _T_1041[11:0];
  assign _T_1043 = ~ _T_1042;
  assign _T_1044 = _T_1043[11:3];
  assign _T_1047 = _T_1037 ? _T_1044 : 9'h0;
  assign _T_1052 = _T_1050 - 9'h1;
  assign _T_1053 = $unsigned(_T_1052);
  assign _T_1054 = _T_1053[8:0];
  assign _T_1056 = _T_1050 == 9'h0;
  assign _T_1058 = _T_1050 == 9'h1;
  assign _T_1060 = _T_1047 == 9'h0;
  assign _T_1061 = _T_1058 | _T_1060;
  assign _T_1065 = _T_1056 ? _T_1047 : _T_1054;
  assign _GEN_11 = _T_1038 ? _T_1065 : _T_1050;
  assign _T_1066 = _T_1037 ? _T_1030_ready : _T_1026_ready;
  assign _T_1067 = _T_89_d_valid & _T_1037;
  assign _T_1069 = _T_1037 == 1'h0;
  assign _T_1070 = _T_89_d_valid & _T_1069;
  assign _T_1071 = _T_89_d_bits_source[3:3];
  assign _GEN_12 = _T_31_b_bits_id ? _T_1106_1 : _T_1106_0;
  assign _GEN_13 = _T_31_b_bits_id ? _T_687_1 : _T_687_0;
  assign _T_1123 = _GEN_2 != _GEN_3;
  assign _T_1126 = 2'h1 << _T_31_b_bits_id;
  assign _T_1128 = _T_1126[0];
  assign _T_1129 = _T_1126[1];
  assign _T_1130 = _T_31_b_ready & _T_31_b_valid;
  assign _T_1131 = _T_1130 & _T_1128;
  assign _T_1133 = _T_1106_0 + 3'h1;
  assign _T_1134 = _T_1133[2:0];
  assign _GEN_14 = _T_1131 ? _T_1134 : _T_1106_0;
  assign _T_1136 = _T_1130 & _T_1129;
  assign _T_1138 = _T_1106_1 + 3'h1;
  assign _T_1139 = _T_1138[2:0];
  assign _GEN_15 = _T_1136 ? _T_1139 : _T_1106_1;
  assign _T_1140 = _T_1085_valid & _T_1123;
  assign _T_1141 = _T_31_b_ready & _T_1123;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_a_valid = _T_89_a_valid;
  assign auto_out_a_bits_opcode = _T_89_a_bits_opcode;
  assign auto_out_a_bits_param = _T_89_a_bits_param;
  assign auto_out_a_bits_size = _T_89_a_bits_size;
  assign auto_out_a_bits_source = _T_89_a_bits_source;
  assign auto_out_a_bits_address = _T_89_a_bits_address;
  assign auto_out_a_bits_mask = _T_89_a_bits_mask;
  assign auto_out_a_bits_data = _T_89_a_bits_data;
  assign auto_out_d_ready = _T_89_d_ready;
  assign _T_31_aw_ready = _T_731;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_w_ready = _T_732;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_1140;
  assign _T_31_b_bits_id = _T_1085_bits_id;
  assign _T_31_b_bits_resp = _T_1085_bits_resp;
  assign _T_31_ar_ready = _T_203_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_1076_valid;
  assign _T_31_r_bits_id = _T_1076_bits_id;
  assign _T_31_r_bits_data = _T_1076_bits_data;
  assign _T_31_r_bits_resp = _T_1076_bits_resp;
  assign _T_31_r_bits_last = _T_1076_bits_last;
  assign _T_89_a_ready = auto_out_a_ready;
  assign _T_89_a_valid = _T_996;
  assign _T_89_a_bits_opcode = _T_1016_opcode;
  assign _T_89_a_bits_param = _T_1016_param;
  assign _T_89_a_bits_size = _T_1016_size;
  assign _T_89_a_bits_source = _T_1016_source;
  assign _T_89_a_bits_address = _T_1016_address;
  assign _T_89_a_bits_mask = _T_1016_mask;
  assign _T_89_a_bits_data = _T_1016_data;
  assign _T_89_d_ready = _T_1066;
  assign _T_89_d_valid = auto_out_d_valid;
  assign _T_89_d_bits_opcode = auto_out_d_bits_opcode;
  assign _T_89_d_bits_size = auto_out_d_bits_size;
  assign _T_89_d_bits_source = auto_out_d_bits_source;
  assign _T_89_d_bits_data = auto_out_d_bits_data;
  assign _T_89_d_bits_error = auto_out_d_bits_error;
  assign _T_203_ready = _T_985;
  assign _T_203_valid = _T_31_ar_valid;
  assign _T_203_bits_size = _T_450_size;
  assign _T_203_bits_source = _T_450_source;
  assign _T_203_bits_address = _T_450_address;
  assign _T_203_bits_mask = _T_450_mask;
  assign _GEN_0 = _GEN_4;
  assign _T_450_size = _T_236;
  assign _T_450_source = _T_355;
  assign _T_450_address = _T_320;
  assign _T_450_mask = _T_522;
  assign _T_540_ready = _T_986;
  assign _T_540_valid = _T_733;
  assign _T_540_bits_size = _T_827_size;
  assign _T_540_bits_source = _T_827_source;
  assign _T_540_bits_address = _T_827_address;
  assign _T_540_bits_mask = _T_827_mask;
  assign _T_540_bits_data = _T_827_data;
  assign _GEN_1 = _GEN_7;
  assign _T_827_size = _T_573;
  assign _T_827_source = _T_704;
  assign _T_827_address = _T_669;
  assign _T_827_mask = _T_31_w_bits_strb;
  assign _T_827_data = _T_31_w_bits_data;
  assign _T_890_0 = _T_886;
  assign _T_890_1 = _T_887;
  assign _T_899_0 = _T_895;
  assign _T_899_1 = _T_896;
  assign _T_995 = _T_993;
  assign _T_1016_opcode = _T_1025;
  assign _T_1016_param = _T_1024;
  assign _T_1016_size = _T_1023;
  assign _T_1016_source = _T_1022;
  assign _T_1016_address = _T_1021;
  assign _T_1016_mask = _T_1020;
  assign _T_1016_data = _T_1019;
  assign _T_1018 = _T_1014;
  assign _T_1026_ready = Queue_1_io_enq_ready;
  assign _T_1026_valid = _T_1070;
  assign _T_1026_bits_id = _T_1071;
  assign _T_1026_bits_resp = _T_1036;
  assign _T_1030_ready = Queue_io_enq_ready;
  assign _T_1030_valid = _T_1067;
  assign _T_1030_bits_id = _T_1071;
  assign _T_1030_bits_data = _T_89_d_bits_data;
  assign _T_1030_bits_resp = _T_1036;
  assign _T_1030_bits_last = _T_1061;
  assign Queue_io_enq_valid = _T_1030_valid;
  assign Queue_io_enq_bits_id = _T_1030_bits_id;
  assign Queue_io_enq_bits_data = _T_1030_bits_data;
  assign Queue_io_enq_bits_resp = _T_1030_bits_resp;
  assign Queue_io_enq_bits_last = _T_1030_bits_last;
  assign Queue_io_deq_ready = _T_1076_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_1076_ready = _T_31_r_ready;
  assign _T_1076_valid = Queue_io_deq_valid;
  assign _T_1076_bits_id = Queue_io_deq_bits_id;
  assign _T_1076_bits_data = Queue_io_deq_bits_data;
  assign _T_1076_bits_resp = Queue_io_deq_bits_resp;
  assign _T_1076_bits_last = Queue_io_deq_bits_last;
  assign Queue_1_io_enq_valid = _T_1026_valid;
  assign Queue_1_io_enq_bits_id = _T_1026_bits_id;
  assign Queue_1_io_enq_bits_resp = _T_1026_bits_resp;
  assign Queue_1_io_deq_ready = _T_1085_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_1085_ready = _T_1141;
  assign _T_1085_valid = Queue_1_io_deq_valid;
  assign _T_1085_bits_id = Queue_1_io_deq_bits_id;
  assign _T_1085_bits_resp = Queue_1_io_deq_bits_resp;
  assign _GEN_2 = _GEN_12;
  assign _GEN_3 = _GEN_13;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_338_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_338_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_687_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_687_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_849 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_863 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_958_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_958_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_1050 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_1106_0 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_1106_1 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_338_0 <= 3'h0;
    end else begin
      if (_T_531) begin
        _T_338_0 <= _T_534;
      end
    end
    if (reset) begin
      _T_338_1 <= 3'h0;
    end else begin
      if (_T_536) begin
        _T_338_1 <= _T_539;
      end
    end
    if (reset) begin
      _T_687_0 <= 3'h0;
    end else begin
      if (_T_837) begin
        _T_687_0 <= _T_840;
      end
    end
    if (reset) begin
      _T_687_1 <= 3'h0;
    end else begin
      if (_T_842) begin
        _T_687_1 <= _T_845;
      end
    end
    if (reset) begin
      _T_849 <= 8'h0;
    end else begin
      if (_T_852) begin
        if (_T_899_1) begin
          _T_849 <= _T_31_aw_bits_len;
        end else begin
          _T_849 <= 8'h0;
        end
      end else begin
        _T_849 <= _T_939;
      end
    end
    if (reset) begin
      _T_863 <= 2'h3;
    end else begin
      if (_T_879) begin
        _T_863 <= _T_883;
      end
    end
    if (reset) begin
      _T_958_0 <= 1'h0;
    end else begin
      if (_T_851) begin
        _T_958_0 <= _T_899_0;
      end
    end
    if (reset) begin
      _T_958_1 <= 1'h0;
    end else begin
      if (_T_851) begin
        _T_958_1 <= _T_899_1;
      end
    end
    if (reset) begin
      _T_1050 <= 9'h0;
    end else begin
      if (_T_1038) begin
        if (_T_1056) begin
          if (_T_1037) begin
            _T_1050 <= _T_1044;
          end else begin
            _T_1050 <= 9'h0;
          end
        end else begin
          _T_1050 <= _T_1054;
        end
      end
    end
    if (reset) begin
      _T_1106_0 <= 3'h0;
    end else begin
      if (_T_1131) begin
        _T_1106_0 <= _T_1134;
      end
    end
    if (reset) begin
      _T_1106_1 <= 3'h0;
    end else begin
      if (_T_1136) begin
        _T_1106_1 <= _T_1139;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_368) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:76 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_368) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:94 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_729) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:95 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_729) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_859) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_859) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_921) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_921) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_930) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_930) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_106(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  reg [7:0] ram [0:3];
  reg [31:0] _RAND_0;
  wire [7:0] ram__T_50_data;
  wire [1:0] ram__T_50_addr;
  wire [7:0] ram__T_36_data;
  wire [1:0] ram__T_36_addr;
  wire  ram__T_36_mask;
  wire  ram__T_36_en;
  reg [1:0] value;
  reg [31:0] _RAND_1;
  reg [1:0] value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [2:0] _T_39;
  wire [1:0] _T_40;
  wire [1:0] _GEN_4;
  wire [2:0] _T_43;
  wire [1:0] _T_44;
  wire [1:0] _GEN_5;
  wire  _T_45;
  wire  _GEN_6;
  wire  _T_47;
  wire  _T_49;
  assign ram__T_50_addr = value_1;
  assign ram__T_50_data = ram[ram__T_50_addr];
  assign ram__T_36_data = io_enq_bits;
  assign ram__T_36_addr = value;
  assign ram__T_36_mask = do_enq;
  assign ram__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 2'h1;
  assign _T_40 = _T_39[1:0];
  assign _GEN_4 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 2'h1;
  assign _T_44 = _T_43[1:0];
  assign _GEN_5 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_6 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits = ram__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_36_en & ram__T_36_mask) begin
      ram[ram__T_36_addr] <= ram__T_36_data;
    end
    if (reset) begin
      value <= 2'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4UserYanker_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [7:0]  auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [7:0]  auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [7:0]  auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [7:0]  auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire  _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [7:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire  _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [7:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire  _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [7:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire  _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [7:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire  _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire  _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire  _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire  _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [7:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [7:0] Queue_io_deq_bits;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [7:0] Queue_1_io_enq_bits;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [7:0] Queue_1_io_deq_bits;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [7:0] Queue_2_io_enq_bits;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [7:0] Queue_2_io_deq_bits;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [7:0] Queue_3_io_enq_bits;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [7:0] Queue_3_io_deq_bits;
  wire  _T_205_0;
  wire  _T_205_1;
  wire  _GEN_0;
  wire  _GEN_8;
  wire  _T_211;
  wire  _GEN_1;
  wire  _T_212;
  wire  _T_215_0;
  wire  _T_215_1;
  wire [7:0] _T_223_0;
  wire [7:0] _T_223_1;
  wire  _T_230;
  wire  _GEN_2;
  wire  _GEN_9;
  wire  _T_231;
  wire  _T_233;
  wire  _T_235;
  wire [7:0] _GEN_3;
  wire [7:0] _GEN_10;
  wire [1:0] _T_238;
  wire  _T_240;
  wire  _T_241;
  wire [1:0] _T_244;
  wire  _T_246;
  wire  _T_247;
  wire  _T_248;
  wire  _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_252;
  wire  _T_254;
  wire  _T_255;
  wire  _T_257;
  wire  _T_260_0;
  wire  _T_260_1;
  wire  _GEN_4;
  wire  _GEN_11;
  wire  _T_266;
  wire  _GEN_5;
  wire  _T_267;
  wire  _T_270_0;
  wire  _T_270_1;
  wire [7:0] _T_278_0;
  wire [7:0] _T_278_1;
  wire  _T_285;
  wire  _GEN_6;
  wire  _GEN_12;
  wire  _T_286;
  wire  _T_288;
  wire  _T_290;
  wire [7:0] _GEN_7;
  wire [7:0] _GEN_13;
  wire [1:0] _T_293;
  wire  _T_295;
  wire  _T_296;
  wire [1:0] _T_299;
  wire  _T_301;
  wire  _T_302;
  wire  _T_303;
  wire  _T_304;
  wire  _T_305;
  wire  _T_306;
  wire  _T_308;
  wire  _T_310;
  Queue_106 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_106 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_106 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_106 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  assign _GEN_8 = _T_31_ar_bits_id ? _T_205_1 : _T_205_0;
  assign _T_211 = _T_89_ar_ready & _GEN_0;
  assign _T_212 = _T_31_ar_valid & _GEN_1;
  assign _T_230 = _T_89_r_valid == 1'h0;
  assign _GEN_9 = _T_89_r_bits_id ? _T_215_1 : _T_215_0;
  assign _T_231 = _T_230 | _GEN_2;
  assign _T_233 = _T_231 | reset;
  assign _T_235 = _T_233 == 1'h0;
  assign _GEN_10 = _T_89_r_bits_id ? _T_223_1 : _T_223_0;
  assign _T_238 = 2'h1 << _T_31_ar_bits_id;
  assign _T_240 = _T_238[0];
  assign _T_241 = _T_238[1];
  assign _T_244 = 2'h1 << _T_89_r_bits_id;
  assign _T_246 = _T_244[0];
  assign _T_247 = _T_244[1];
  assign _T_248 = _T_89_r_valid & _T_31_r_ready;
  assign _T_249 = _T_248 & _T_246;
  assign _T_250 = _T_249 & _T_89_r_bits_last;
  assign _T_251 = _T_31_ar_valid & _T_89_ar_ready;
  assign _T_252 = _T_251 & _T_240;
  assign _T_254 = _T_248 & _T_247;
  assign _T_255 = _T_254 & _T_89_r_bits_last;
  assign _T_257 = _T_251 & _T_241;
  assign _GEN_11 = _T_31_aw_bits_id ? _T_260_1 : _T_260_0;
  assign _T_266 = _T_89_aw_ready & _GEN_4;
  assign _T_267 = _T_31_aw_valid & _GEN_5;
  assign _T_285 = _T_89_b_valid == 1'h0;
  assign _GEN_12 = _T_89_b_bits_id ? _T_270_1 : _T_270_0;
  assign _T_286 = _T_285 | _GEN_6;
  assign _T_288 = _T_286 | reset;
  assign _T_290 = _T_288 == 1'h0;
  assign _GEN_13 = _T_89_b_bits_id ? _T_278_1 : _T_278_0;
  assign _T_293 = 2'h1 << _T_31_aw_bits_id;
  assign _T_295 = _T_293[0];
  assign _T_296 = _T_293[1];
  assign _T_299 = 2'h1 << _T_89_b_bits_id;
  assign _T_301 = _T_299[0];
  assign _T_302 = _T_299[1];
  assign _T_303 = _T_89_b_valid & _T_31_b_ready;
  assign _T_304 = _T_303 & _T_301;
  assign _T_305 = _T_31_aw_valid & _T_89_aw_ready;
  assign _T_306 = _T_305 & _T_295;
  assign _T_308 = _T_303 & _T_302;
  assign _T_310 = _T_305 & _T_296;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_266;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_b_bits_user = _GEN_7;
  assign _T_31_ar_ready = _T_211;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _GEN_3;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_267;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id;
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_212;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id;
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_252;
  assign Queue_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_io_deq_ready = _T_250;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_1_io_enq_valid = _T_257;
  assign Queue_1_io_enq_bits = _T_31_ar_bits_user;
  assign Queue_1_io_deq_ready = _T_255;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_2_io_enq_valid = _T_306;
  assign Queue_2_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_2_io_deq_ready = _T_304;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_3_io_enq_valid = _T_310;
  assign Queue_3_io_enq_bits = _T_31_aw_bits_user;
  assign Queue_3_io_deq_ready = _T_308;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign _T_205_0 = Queue_io_enq_ready;
  assign _T_205_1 = Queue_1_io_enq_ready;
  assign _GEN_0 = _GEN_8;
  assign _GEN_1 = _GEN_8;
  assign _T_215_0 = Queue_io_deq_valid;
  assign _T_215_1 = Queue_1_io_deq_valid;
  assign _T_223_0 = Queue_io_deq_bits;
  assign _T_223_1 = Queue_1_io_deq_bits;
  assign _GEN_2 = _GEN_9;
  assign _GEN_3 = _GEN_10;
  assign _T_260_0 = Queue_2_io_enq_ready;
  assign _T_260_1 = Queue_3_io_enq_ready;
  assign _GEN_4 = _GEN_11;
  assign _GEN_5 = _GEN_11;
  assign _T_270_0 = Queue_2_io_deq_valid;
  assign _T_270_1 = Queue_3_io_deq_valid;
  assign _T_278_0 = Queue_2_io_deq_bits;
  assign _T_278_1 = Queue_3_io_deq_bits;
  assign _GEN_6 = _GEN_12;
  assign _GEN_7 = _GEN_13;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_235) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_290) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_110(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [6:0]  io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [6:0]  io_deq_bits_user
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire  ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [31:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [31:0] ram_addr__T_42_data;
  wire  ram_addr__T_42_addr;
  wire [31:0] ram_addr__T_33_data;
  wire  ram_addr__T_33_addr;
  wire  ram_addr__T_33_mask;
  wire  ram_addr__T_33_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_42_data;
  wire  ram_len__T_42_addr;
  wire [7:0] ram_len__T_33_data;
  wire  ram_len__T_33_addr;
  wire  ram_len__T_33_mask;
  wire  ram_len__T_33_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [2:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_42_data;
  wire  ram_burst__T_42_addr;
  wire [1:0] ram_burst__T_33_data;
  wire  ram_burst__T_33_addr;
  wire  ram_burst__T_33_mask;
  wire  ram_burst__T_33_en;
  reg [6:0] ram_user [0:0];
  reg [31:0] _RAND_5;
  wire [6:0] ram_user__T_42_data;
  wire  ram_user__T_42_addr;
  wire [6:0] ram_user__T_33_data;
  wire  ram_user__T_33_addr;
  wire  ram_user__T_33_mask;
  wire  ram_user__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_13;
  wire  _T_38;
  wire  _GEN_14;
  wire  _GEN_15;
  wire [6:0] _GEN_16;
  wire [1:0] _GEN_21;
  wire [2:0] _GEN_22;
  wire [7:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_addr__T_42_addr = 1'h0;
  assign ram_addr__T_42_data = ram_addr[ram_addr__T_42_addr];
  assign ram_addr__T_33_data = io_enq_bits_addr;
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_mask = do_enq;
  assign ram_addr__T_33_en = do_enq;
  assign ram_len__T_42_addr = 1'h0;
  assign ram_len__T_42_data = ram_len[ram_len__T_42_addr];
  assign ram_len__T_33_data = io_enq_bits_len;
  assign ram_len__T_33_addr = 1'h0;
  assign ram_len__T_33_mask = do_enq;
  assign ram_len__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_burst__T_42_addr = 1'h0;
  assign ram_burst__T_42_data = ram_burst[ram_burst__T_42_addr];
  assign ram_burst__T_33_data = io_enq_bits_burst;
  assign ram_burst__T_33_addr = 1'h0;
  assign ram_burst__T_33_mask = do_enq;
  assign ram_burst__T_33_en = do_enq;
  assign ram_user__T_42_addr = 1'h0;
  assign ram_user__T_42_data = ram_user[ram_user__T_42_addr];
  assign ram_user__T_33_data = io_enq_bits_user;
  assign ram_user__T_33_addr = 1'h0;
  assign ram_user__T_33_mask = do_enq;
  assign ram_user__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_13 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_14 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_15 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_16 = empty ? io_enq_bits_user : ram_user__T_42_data;
  assign _GEN_21 = empty ? io_enq_bits_burst : ram_burst__T_42_data;
  assign _GEN_22 = empty ? io_enq_bits_size : ram_size__T_42_data;
  assign _GEN_23 = empty ? io_enq_bits_len : ram_len__T_42_data;
  assign _GEN_24 = empty ? io_enq_bits_addr : ram_addr__T_42_data;
  assign _GEN_25 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_26 = empty ? 1'h0 : _T_30;
  assign _GEN_27 = empty ? _GEN_15 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_14;
  assign io_deq_bits_id = _GEN_25;
  assign io_deq_bits_addr = _GEN_24;
  assign io_deq_bits_len = _GEN_23;
  assign io_deq_bits_size = _GEN_22;
  assign io_deq_bits_burst = _GEN_21;
  assign io_deq_bits_user = _GEN_16;
  assign do_enq = _GEN_27;
  assign do_deq = _GEN_26;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = _RAND_5[6:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_addr__T_33_en & ram_addr__T_33_mask) begin
      ram_addr[ram_addr__T_33_addr] <= ram_addr__T_33_data;
    end
    if(ram_len__T_33_en & ram_len__T_33_mask) begin
      ram_len[ram_len__T_33_addr] <= ram_len__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_burst__T_33_en & ram_burst__T_33_mask) begin
      ram_burst[ram_burst__T_33_addr] <= ram_burst__T_33_data;
    end
    if(ram_user__T_33_en & ram_user__T_33_mask) begin
      ram_user[ram_user__T_33_addr] <= ram_user__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input  [6:0]  auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [6:0]  auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input  [6:0]  auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [6:0]  auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [7:0]  auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [7:0]  auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [7:0]  auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [7:0]  auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire  _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire [6:0] _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire  _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire [6:0] _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire  _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire [6:0] _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire  _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire [6:0] _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire  _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [7:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire  _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [7:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire  _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [7:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire  _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [7:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits_id;
  wire [31:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire [6:0] Queue_io_enq_bits_user;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits_id;
  wire [31:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire [6:0] Queue_io_deq_bits_user;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire  _T_207_bits_id;
  wire [31:0] _T_207_bits_addr;
  wire [7:0] _T_207_bits_len;
  wire [2:0] _T_207_bits_size;
  wire [1:0] _T_207_bits_burst;
  wire [6:0] _T_207_bits_user;
  wire  _T_211_ready;
  wire  _T_211_valid;
  wire  _T_211_bits_id;
  wire [31:0] _T_211_bits_addr;
  wire [7:0] _T_211_bits_len;
  wire [2:0] _T_211_bits_size;
  wire [6:0] _T_211_bits_user;
  reg  _T_217;
  reg [31:0] _RAND_0;
  reg [31:0] _T_219;
  reg [31:0] _RAND_1;
  reg [7:0] _T_221;
  reg [31:0] _RAND_2;
  wire [7:0] _T_222;
  wire [31:0] _T_223;
  wire [28:0] _T_225;
  wire [7:0] _T_226;
  wire [31:0] _T_228;
  wire [32:0] _T_229;
  wire [32:0] _T_231;
  wire [32:0] _T_232;
  wire  _T_234;
  wire [31:0] _T_236;
  wire [32:0] _T_237;
  wire [32:0] _T_239;
  wire [32:0] _T_240;
  wire  _T_242;
  wire [32:0] _T_245;
  wire [32:0] _T_247;
  wire [32:0] _T_248;
  wire  _T_250;
  wire [31:0] _T_252;
  wire [32:0] _T_253;
  wire [32:0] _T_255;
  wire [32:0] _T_256;
  wire  _T_258;
  wire [31:0] _T_260;
  wire [32:0] _T_261;
  wire [32:0] _T_263;
  wire [32:0] _T_264;
  wire  _T_266;
  wire [31:0] _T_268;
  wire [32:0] _T_269;
  wire [32:0] _T_271;
  wire [32:0] _T_272;
  wire  _T_274;
  wire  _T_275;
  wire  _T_276;
  wire  _T_277;
  wire  _T_278;
  wire  _T_279;
  wire [31:0] _T_282;
  wire [32:0] _T_283;
  wire [32:0] _T_285;
  wire [32:0] _T_286;
  wire  _T_288;
  wire [2:0] _T_292;
  wire [7:0] _T_294;
  wire [7:0] _GEN_16;
  wire [7:0] _T_295;
  wire [7:0] _T_297;
  wire [6:0] _T_298;
  wire [7:0] _GEN_17;
  wire [7:0] _T_299;
  wire [5:0] _T_300;
  wire [7:0] _GEN_18;
  wire [7:0] _T_301;
  wire [3:0] _T_302;
  wire [7:0] _GEN_19;
  wire [7:0] _T_303;
  wire [6:0] _T_305;
  wire [7:0] _T_306;
  wire [8:0] _GEN_20;
  wire [8:0] _T_307;
  wire [7:0] _T_308;
  wire [7:0] _T_309;
  wire [9:0] _GEN_21;
  wire [9:0] _T_310;
  wire [7:0] _T_311;
  wire [7:0] _T_312;
  wire [11:0] _GEN_22;
  wire [11:0] _T_313;
  wire [7:0] _T_314;
  wire [7:0] _T_315;
  wire [7:0] _T_317;
  wire [7:0] _GEN_23;
  wire [7:0] _T_318;
  wire [8:0] _GEN_24;
  wire [8:0] _T_319;
  wire [7:0] _T_320;
  wire [7:0] _T_321;
  wire [9:0] _GEN_25;
  wire [9:0] _T_322;
  wire [7:0] _T_323;
  wire [7:0] _T_324;
  wire [11:0] _GEN_26;
  wire [11:0] _T_325;
  wire [7:0] _T_326;
  wire [7:0] _T_327;
  wire [7:0] _T_329;
  wire [7:0] _T_330;
  wire [7:0] _T_331;
  wire  _T_333;
  wire  _T_335;
  wire  _T_336;
  wire [7:0] _T_338;
  wire [8:0] _GEN_27;
  wire [8:0] _T_339;
  wire [8:0] _T_341;
  wire [8:0] _T_343;
  wire [8:0] _T_344;
  wire [8:0] _T_345;
  wire [15:0] _GEN_28;
  wire [15:0] _T_346;
  wire [31:0] _GEN_29;
  wire [32:0] _T_347;
  wire [31:0] _T_348;
  wire [15:0] _T_350;
  wire [22:0] _GEN_30;
  wire [22:0] _T_351;
  wire [14:0] _T_352;
  wire [31:0] _T_354;
  wire  _T_356;
  wire [31:0] _GEN_31;
  wire [31:0] _T_357;
  wire [31:0] _T_358;
  wire [31:0] _T_359;
  wire [31:0] _T_360;
  wire [31:0] _T_361;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire  _T_364;
  wire  _T_365;
  wire [31:0] _T_366;
  wire [9:0] _T_369;
  wire [2:0] _T_370;
  wire [2:0] _T_371;
  wire [31:0] _GEN_33;
  wire [31:0] _T_372;
  wire [31:0] _T_373;
  wire  _T_374;
  wire  _T_376;
  wire [8:0] _GEN_34;
  wire [9:0] _T_377;
  wire [9:0] _T_378;
  wire [8:0] _T_379;
  wire  _GEN_3;
  wire [31:0] _GEN_4;
  wire [8:0] _GEN_5;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_id;
  wire [31:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire [6:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_id;
  wire [31:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire [6:0] Queue_1_io_deq_bits_user;
  wire  _T_384_ready;
  wire  _T_384_valid;
  wire  _T_384_bits_id;
  wire [31:0] _T_384_bits_addr;
  wire [7:0] _T_384_bits_len;
  wire [2:0] _T_384_bits_size;
  wire [1:0] _T_384_bits_burst;
  wire [6:0] _T_384_bits_user;
  wire  _T_388_ready;
  wire  _T_388_valid;
  wire  _T_388_bits_id;
  wire [31:0] _T_388_bits_addr;
  wire [7:0] _T_388_bits_len;
  wire [2:0] _T_388_bits_size;
  wire [6:0] _T_388_bits_user;
  reg  _T_394;
  reg [31:0] _RAND_3;
  reg [31:0] _T_396;
  reg [31:0] _RAND_4;
  reg [7:0] _T_398;
  reg [31:0] _RAND_5;
  wire [7:0] _T_399;
  wire [31:0] _T_400;
  wire [28:0] _T_402;
  wire [7:0] _T_403;
  wire [31:0] _T_405;
  wire [32:0] _T_406;
  wire [32:0] _T_408;
  wire [32:0] _T_409;
  wire  _T_411;
  wire [31:0] _T_414;
  wire [32:0] _T_415;
  wire [32:0] _T_417;
  wire [32:0] _T_418;
  wire  _T_420;
  wire [31:0] _T_422;
  wire [32:0] _T_423;
  wire [32:0] _T_425;
  wire [32:0] _T_426;
  wire  _T_428;
  wire [32:0] _T_431;
  wire [32:0] _T_433;
  wire [32:0] _T_434;
  wire  _T_436;
  wire [31:0] _T_438;
  wire [32:0] _T_439;
  wire [32:0] _T_441;
  wire [32:0] _T_442;
  wire  _T_444;
  wire  _T_445;
  wire  _T_446;
  wire  _T_447;
  wire [31:0] _T_450;
  wire [32:0] _T_451;
  wire [32:0] _T_453;
  wire [32:0] _T_454;
  wire  _T_456;
  wire [4:0] _T_460;
  wire [2:0] _T_462;
  wire [7:0] _T_464;
  wire [4:0] _GEN_35;
  wire [4:0] _T_465;
  wire [7:0] _GEN_36;
  wire [7:0] _T_466;
  wire [7:0] _T_468;
  wire [6:0] _T_469;
  wire [7:0] _GEN_37;
  wire [7:0] _T_470;
  wire [5:0] _T_471;
  wire [7:0] _GEN_38;
  wire [7:0] _T_472;
  wire [3:0] _T_473;
  wire [7:0] _GEN_39;
  wire [7:0] _T_474;
  wire [6:0] _T_476;
  wire [7:0] _T_477;
  wire [8:0] _GEN_40;
  wire [8:0] _T_478;
  wire [7:0] _T_479;
  wire [7:0] _T_480;
  wire [9:0] _GEN_41;
  wire [9:0] _T_481;
  wire [7:0] _T_482;
  wire [7:0] _T_483;
  wire [11:0] _GEN_42;
  wire [11:0] _T_484;
  wire [7:0] _T_485;
  wire [7:0] _T_486;
  wire [7:0] _T_488;
  wire [7:0] _GEN_43;
  wire [7:0] _T_489;
  wire [8:0] _GEN_44;
  wire [8:0] _T_490;
  wire [7:0] _T_491;
  wire [7:0] _T_492;
  wire [9:0] _GEN_45;
  wire [9:0] _T_493;
  wire [7:0] _T_494;
  wire [7:0] _T_495;
  wire [11:0] _GEN_46;
  wire [11:0] _T_496;
  wire [7:0] _T_497;
  wire [7:0] _T_498;
  wire [7:0] _T_500;
  wire [7:0] _T_501;
  wire [7:0] _T_502;
  wire  _T_504;
  wire  _T_506;
  wire  _T_507;
  wire [7:0] _T_509;
  wire [8:0] _GEN_47;
  wire [8:0] _T_510;
  wire [8:0] _T_512;
  wire [8:0] _T_514;
  wire [8:0] _T_515;
  wire [8:0] _T_516;
  wire [15:0] _GEN_48;
  wire [15:0] _T_517;
  wire [31:0] _GEN_49;
  wire [32:0] _T_518;
  wire [31:0] _T_519;
  wire [15:0] _T_521;
  wire [22:0] _GEN_50;
  wire [22:0] _T_522;
  wire [14:0] _T_523;
  wire [31:0] _T_525;
  wire  _T_527;
  wire [31:0] _GEN_51;
  wire [31:0] _T_528;
  wire [31:0] _T_529;
  wire [31:0] _T_530;
  wire [31:0] _T_531;
  wire [31:0] _T_532;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_535;
  wire  _T_536;
  wire [31:0] _T_537;
  wire [9:0] _T_540;
  wire [2:0] _T_541;
  wire [2:0] _T_542;
  wire [31:0] _GEN_53;
  wire [31:0] _T_543;
  wire [31:0] _T_544;
  wire  _T_545;
  wire  _T_547;
  wire [8:0] _GEN_54;
  wire [9:0] _T_548;
  wire [9:0] _T_549;
  wire [8:0] _T_550;
  wire  _GEN_8;
  wire [31:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [7:0] Queue_2_io_enq_bits_strb;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [7:0] Queue_2_io_deq_bits_strb;
  wire  Queue_2_io_deq_bits_last;
  wire  _T_555_ready;
  wire  _T_555_valid;
  wire [63:0] _T_555_bits_data;
  wire [7:0] _T_555_bits_strb;
  wire  _T_555_bits_last;
  wire [7:0] _T_559;
  reg  _T_562;
  reg [31:0] _RAND_6;
  wire  _T_564;
  wire  _T_566;
  wire  _T_567;
  wire  _GEN_11;
  wire  _T_569;
  wire  _GEN_12;
  wire  _T_571;
  wire  _T_572;
  wire  _T_574;
  wire  _T_576;
  wire  _T_577;
  wire [7:0] _T_578;
  reg [8:0] _T_581;
  reg [31:0] _RAND_7;
  wire  _T_583;
  wire [8:0] _T_585;
  wire [8:0] _T_586;
  wire  _T_588;
  wire  _T_589;
  wire [8:0] _GEN_55;
  wire [9:0] _T_590;
  wire [9:0] _T_591;
  wire [8:0] _T_592;
  wire  _T_595;
  wire  _T_597;
  wire  _T_598;
  wire  _T_600;
  wire  _T_602;
  wire  _T_604;
  wire  _T_605;
  wire  _T_606;
  wire  _T_610;
  wire  _T_612;
  wire  _T_614;
  wire  _T_615;
  wire  _T_616;
  wire  _T_618;
  wire  _T_620;
  wire  _T_621;
  wire  _T_622;
  wire [6:0] _T_623;
  wire  _T_624;
  wire  _T_625;
  wire  _T_627;
  wire  _T_628;
  wire [6:0] _T_629;
  reg [1:0] _T_647_0;
  reg [31:0] _RAND_8;
  reg [1:0] _T_647_1;
  reg [31:0] _RAND_9;
  wire [1:0] _GEN_0;
  wire [1:0] _GEN_13;
  wire [1:0] _T_661;
  wire [1:0] _T_664;
  wire  _T_666;
  wire  _T_667;
  wire  _T_668;
  wire  _T_669;
  wire [1:0] _T_671;
  wire [1:0] _T_672;
  wire [1:0] _GEN_14;
  wire  _T_674;
  wire [1:0] _T_676;
  wire [1:0] _T_677;
  wire [1:0] _GEN_15;
  Queue_110 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  Queue_110 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_user(Queue_1_io_deq_bits_user)
  );
  Queue_32 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign _T_222 = _T_217 ? _T_221 : _T_207_bits_len;
  assign _T_223 = _T_217 ? _T_219 : _T_207_bits_addr;
  assign _T_225 = _T_223[31:3];
  assign _T_226 = _T_225[7:0];
  assign _T_228 = _T_223 ^ 32'h8000000;
  assign _T_229 = {1'b0,$signed(_T_228)};
  assign _T_231 = $signed(_T_229) & $signed(33'shc8000000);
  assign _T_232 = $signed(_T_231);
  assign _T_234 = $signed(_T_232) == $signed(33'sh0);
  assign _T_236 = _T_223 ^ 32'h2000000;
  assign _T_237 = {1'b0,$signed(_T_236)};
  assign _T_239 = $signed(_T_237) & $signed(33'shca010000);
  assign _T_240 = $signed(_T_239);
  assign _T_242 = $signed(_T_240) == $signed(33'sh0);
  assign _T_245 = {1'b0,$signed(_T_223)};
  assign _T_247 = $signed(_T_245) & $signed(33'shca012000);
  assign _T_248 = $signed(_T_247);
  assign _T_250 = $signed(_T_248) == $signed(33'sh0);
  assign _T_252 = _T_223 ^ 32'h10000;
  assign _T_253 = {1'b0,$signed(_T_252)};
  assign _T_255 = $signed(_T_253) & $signed(33'shca010000);
  assign _T_256 = $signed(_T_255);
  assign _T_258 = $signed(_T_256) == $signed(33'sh0);
  assign _T_260 = _T_223 ^ 32'h40000000;
  assign _T_261 = {1'b0,$signed(_T_260)};
  assign _T_263 = $signed(_T_261) & $signed(33'shc0000000);
  assign _T_264 = $signed(_T_263);
  assign _T_266 = $signed(_T_264) == $signed(33'sh0);
  assign _T_268 = _T_223 ^ 32'h80000000;
  assign _T_269 = {1'b0,$signed(_T_268)};
  assign _T_271 = $signed(_T_269) & $signed(33'shc0000000);
  assign _T_272 = $signed(_T_271);
  assign _T_274 = $signed(_T_272) == $signed(33'sh0);
  assign _T_275 = _T_234 | _T_242;
  assign _T_276 = _T_275 | _T_250;
  assign _T_277 = _T_276 | _T_258;
  assign _T_278 = _T_277 | _T_266;
  assign _T_279 = _T_278 | _T_274;
  assign _T_282 = _T_223 ^ 32'h2000;
  assign _T_283 = {1'b0,$signed(_T_282)};
  assign _T_285 = $signed(_T_283) & $signed(33'shca012000);
  assign _T_286 = $signed(_T_285);
  assign _T_288 = $signed(_T_286) == $signed(33'sh0);
  assign _T_292 = _T_279 ? 3'h7 : 3'h0;
  assign _T_294 = _T_288 ? 8'hff : 8'h0;
  assign _GEN_16 = {{5'd0}, _T_292};
  assign _T_295 = _GEN_16 | _T_294;
  assign _T_298 = _T_222[7:1];
  assign _GEN_17 = {{1'd0}, _T_298};
  assign _T_299 = _T_222 | _GEN_17;
  assign _T_300 = _T_299[7:2];
  assign _GEN_18 = {{2'd0}, _T_300};
  assign _T_301 = _T_299 | _GEN_18;
  assign _T_302 = _T_301[7:4];
  assign _GEN_19 = {{4'd0}, _T_302};
  assign _T_303 = _T_301 | _GEN_19;
  assign _T_305 = _T_303[7:1];
  assign _T_306 = ~ _T_222;
  assign _GEN_20 = {{1'd0}, _T_306};
  assign _T_307 = _GEN_20 << 1;
  assign _T_308 = _T_307[7:0];
  assign _T_309 = _T_306 | _T_308;
  assign _GEN_21 = {{2'd0}, _T_309};
  assign _T_310 = _GEN_21 << 2;
  assign _T_311 = _T_310[7:0];
  assign _T_312 = _T_309 | _T_311;
  assign _GEN_22 = {{4'd0}, _T_312};
  assign _T_313 = _GEN_22 << 4;
  assign _T_314 = _T_313[7:0];
  assign _T_315 = _T_312 | _T_314;
  assign _T_317 = ~ _T_315;
  assign _GEN_23 = {{1'd0}, _T_305};
  assign _T_318 = _GEN_23 | _T_317;
  assign _GEN_24 = {{1'd0}, _T_226};
  assign _T_319 = _GEN_24 << 1;
  assign _T_320 = _T_319[7:0];
  assign _T_321 = _T_226 | _T_320;
  assign _GEN_25 = {{2'd0}, _T_321};
  assign _T_322 = _GEN_25 << 2;
  assign _T_323 = _T_322[7:0];
  assign _T_324 = _T_321 | _T_323;
  assign _GEN_26 = {{4'd0}, _T_324};
  assign _T_325 = _GEN_26 << 4;
  assign _T_326 = _T_325[7:0];
  assign _T_327 = _T_324 | _T_326;
  assign _T_329 = ~ _T_327;
  assign _T_330 = _T_318 & _T_329;
  assign _T_331 = _T_330 & _T_297;
  assign _T_333 = _T_207_bits_burst == 2'h0;
  assign _T_335 = _T_207_bits_size != 3'h3;
  assign _T_336 = _T_333 | _T_335;
  assign _T_338 = _T_336 ? 8'h0 : _T_331;
  assign _GEN_27 = {{1'd0}, _T_338};
  assign _T_339 = _GEN_27 << 1;
  assign _T_341 = _T_339 | 9'h1;
  assign _T_343 = {1'h0,_T_338};
  assign _T_344 = ~ _T_343;
  assign _T_345 = _T_341 & _T_344;
  assign _GEN_28 = {{7'd0}, _T_345};
  assign _T_346 = _GEN_28 << _T_207_bits_size;
  assign _GEN_29 = {{16'd0}, _T_346};
  assign _T_347 = _T_223 + _GEN_29;
  assign _T_348 = _T_347[31:0];
  assign _T_350 = {_T_207_bits_len,8'hff};
  assign _GEN_30 = {{7'd0}, _T_350};
  assign _T_351 = _GEN_30 << _T_207_bits_size;
  assign _T_352 = _T_351[22:8];
  assign _T_356 = _T_207_bits_burst == 2'h2;
  assign _GEN_31 = {{17'd0}, _T_352};
  assign _T_357 = _T_348 & _GEN_31;
  assign _T_358 = ~ _T_207_bits_addr;
  assign _T_359 = _T_358 | _GEN_31;
  assign _T_360 = ~ _T_359;
  assign _T_361 = _T_357 | _T_360;
  assign _GEN_1 = _T_356 ? _T_361 : _T_348;
  assign _GEN_2 = _T_333 ? _T_207_bits_addr : _GEN_1;
  assign _T_364 = _T_338 == _T_222;
  assign _T_365 = _T_211_ready & _T_364;
  assign _T_366 = ~ _T_223;
  assign _T_369 = 10'h7 << _T_207_bits_size;
  assign _T_370 = _T_369[2:0];
  assign _T_371 = ~ _T_370;
  assign _GEN_33 = {{29'd0}, _T_371};
  assign _T_372 = _T_366 | _GEN_33;
  assign _T_373 = ~ _T_372;
  assign _T_374 = _T_211_ready & _T_211_valid;
  assign _T_376 = _T_364 == 1'h0;
  assign _GEN_34 = {{1'd0}, _T_222};
  assign _T_377 = _GEN_34 - _T_345;
  assign _T_378 = $unsigned(_T_377);
  assign _T_379 = _T_378[8:0];
  assign _GEN_3 = _T_374 ? _T_376 : _T_217;
  assign _GEN_4 = _T_374 ? _T_354 : _T_219;
  assign _GEN_5 = _T_374 ? _T_379 : {{1'd0}, _T_221};
  assign _T_399 = _T_394 ? _T_398 : _T_384_bits_len;
  assign _T_400 = _T_394 ? _T_396 : _T_384_bits_addr;
  assign _T_402 = _T_400[31:3];
  assign _T_403 = _T_402[7:0];
  assign _T_405 = _T_400 ^ 32'h40000000;
  assign _T_406 = {1'b0,$signed(_T_405)};
  assign _T_408 = $signed(_T_406) & $signed(33'shc0000000);
  assign _T_409 = $signed(_T_408);
  assign _T_411 = $signed(_T_409) == $signed(33'sh0);
  assign _T_414 = _T_400 ^ 32'h8000000;
  assign _T_415 = {1'b0,$signed(_T_414)};
  assign _T_417 = $signed(_T_415) & $signed(33'shc8000000);
  assign _T_418 = $signed(_T_417);
  assign _T_420 = $signed(_T_418) == $signed(33'sh0);
  assign _T_422 = _T_400 ^ 32'h2000000;
  assign _T_423 = {1'b0,$signed(_T_422)};
  assign _T_425 = $signed(_T_423) & $signed(33'shca000000);
  assign _T_426 = $signed(_T_425);
  assign _T_428 = $signed(_T_426) == $signed(33'sh0);
  assign _T_431 = {1'b0,$signed(_T_400)};
  assign _T_433 = $signed(_T_431) & $signed(33'shca002000);
  assign _T_434 = $signed(_T_433);
  assign _T_436 = $signed(_T_434) == $signed(33'sh0);
  assign _T_438 = _T_400 ^ 32'h80000000;
  assign _T_439 = {1'b0,$signed(_T_438)};
  assign _T_441 = $signed(_T_439) & $signed(33'shc0000000);
  assign _T_442 = $signed(_T_441);
  assign _T_444 = $signed(_T_442) == $signed(33'sh0);
  assign _T_445 = _T_420 | _T_428;
  assign _T_446 = _T_445 | _T_436;
  assign _T_447 = _T_446 | _T_444;
  assign _T_450 = _T_400 ^ 32'h2000;
  assign _T_451 = {1'b0,$signed(_T_450)};
  assign _T_453 = $signed(_T_451) & $signed(33'shca002000);
  assign _T_454 = $signed(_T_453);
  assign _T_456 = $signed(_T_454) == $signed(33'sh0);
  assign _T_460 = _T_411 ? 5'h1f : 5'h0;
  assign _T_462 = _T_447 ? 3'h7 : 3'h0;
  assign _T_464 = _T_456 ? 8'hff : 8'h0;
  assign _GEN_35 = {{2'd0}, _T_462};
  assign _T_465 = _T_460 | _GEN_35;
  assign _GEN_36 = {{3'd0}, _T_465};
  assign _T_466 = _GEN_36 | _T_464;
  assign _T_469 = _T_399[7:1];
  assign _GEN_37 = {{1'd0}, _T_469};
  assign _T_470 = _T_399 | _GEN_37;
  assign _T_471 = _T_470[7:2];
  assign _GEN_38 = {{2'd0}, _T_471};
  assign _T_472 = _T_470 | _GEN_38;
  assign _T_473 = _T_472[7:4];
  assign _GEN_39 = {{4'd0}, _T_473};
  assign _T_474 = _T_472 | _GEN_39;
  assign _T_476 = _T_474[7:1];
  assign _T_477 = ~ _T_399;
  assign _GEN_40 = {{1'd0}, _T_477};
  assign _T_478 = _GEN_40 << 1;
  assign _T_479 = _T_478[7:0];
  assign _T_480 = _T_477 | _T_479;
  assign _GEN_41 = {{2'd0}, _T_480};
  assign _T_481 = _GEN_41 << 2;
  assign _T_482 = _T_481[7:0];
  assign _T_483 = _T_480 | _T_482;
  assign _GEN_42 = {{4'd0}, _T_483};
  assign _T_484 = _GEN_42 << 4;
  assign _T_485 = _T_484[7:0];
  assign _T_486 = _T_483 | _T_485;
  assign _T_488 = ~ _T_486;
  assign _GEN_43 = {{1'd0}, _T_476};
  assign _T_489 = _GEN_43 | _T_488;
  assign _GEN_44 = {{1'd0}, _T_403};
  assign _T_490 = _GEN_44 << 1;
  assign _T_491 = _T_490[7:0];
  assign _T_492 = _T_403 | _T_491;
  assign _GEN_45 = {{2'd0}, _T_492};
  assign _T_493 = _GEN_45 << 2;
  assign _T_494 = _T_493[7:0];
  assign _T_495 = _T_492 | _T_494;
  assign _GEN_46 = {{4'd0}, _T_495};
  assign _T_496 = _GEN_46 << 4;
  assign _T_497 = _T_496[7:0];
  assign _T_498 = _T_495 | _T_497;
  assign _T_500 = ~ _T_498;
  assign _T_501 = _T_489 & _T_500;
  assign _T_502 = _T_501 & _T_468;
  assign _T_504 = _T_384_bits_burst == 2'h0;
  assign _T_506 = _T_384_bits_size != 3'h3;
  assign _T_507 = _T_504 | _T_506;
  assign _T_509 = _T_507 ? 8'h0 : _T_502;
  assign _GEN_47 = {{1'd0}, _T_509};
  assign _T_510 = _GEN_47 << 1;
  assign _T_512 = _T_510 | 9'h1;
  assign _T_514 = {1'h0,_T_509};
  assign _T_515 = ~ _T_514;
  assign _T_516 = _T_512 & _T_515;
  assign _GEN_48 = {{7'd0}, _T_516};
  assign _T_517 = _GEN_48 << _T_384_bits_size;
  assign _GEN_49 = {{16'd0}, _T_517};
  assign _T_518 = _T_400 + _GEN_49;
  assign _T_519 = _T_518[31:0];
  assign _T_521 = {_T_384_bits_len,8'hff};
  assign _GEN_50 = {{7'd0}, _T_521};
  assign _T_522 = _GEN_50 << _T_384_bits_size;
  assign _T_523 = _T_522[22:8];
  assign _T_527 = _T_384_bits_burst == 2'h2;
  assign _GEN_51 = {{17'd0}, _T_523};
  assign _T_528 = _T_519 & _GEN_51;
  assign _T_529 = ~ _T_384_bits_addr;
  assign _T_530 = _T_529 | _GEN_51;
  assign _T_531 = ~ _T_530;
  assign _T_532 = _T_528 | _T_531;
  assign _GEN_6 = _T_527 ? _T_532 : _T_519;
  assign _GEN_7 = _T_504 ? _T_384_bits_addr : _GEN_6;
  assign _T_535 = _T_509 == _T_399;
  assign _T_536 = _T_388_ready & _T_535;
  assign _T_537 = ~ _T_400;
  assign _T_540 = 10'h7 << _T_384_bits_size;
  assign _T_541 = _T_540[2:0];
  assign _T_542 = ~ _T_541;
  assign _GEN_53 = {{29'd0}, _T_542};
  assign _T_543 = _T_537 | _GEN_53;
  assign _T_544 = ~ _T_543;
  assign _T_545 = _T_388_ready & _T_388_valid;
  assign _T_547 = _T_535 == 1'h0;
  assign _GEN_54 = {{1'd0}, _T_399};
  assign _T_548 = _GEN_54 - _T_516;
  assign _T_549 = $unsigned(_T_548);
  assign _T_550 = _T_549[8:0];
  assign _GEN_8 = _T_545 ? _T_547 : _T_394;
  assign _GEN_9 = _T_545 ? _T_525 : _T_396;
  assign _GEN_10 = _T_545 ? _T_550 : {{1'd0}, _T_398};
  assign _T_559 = {_T_211_bits_user,_T_364};
  assign _T_567 = _T_566 & _T_564;
  assign _GEN_11 = _T_567 ? 1'h1 : _T_562;
  assign _T_569 = _T_89_aw_ready & _T_89_aw_valid;
  assign _GEN_12 = _T_569 ? 1'h0 : _GEN_11;
  assign _T_571 = _T_564 | _T_562;
  assign _T_572 = _T_388_valid & _T_571;
  assign _T_574 = _T_89_aw_ready & _T_571;
  assign _T_576 = _T_562 == 1'h0;
  assign _T_577 = _T_388_valid & _T_576;
  assign _T_578 = {_T_388_bits_user,_T_535};
  assign _T_583 = _T_581 == 9'h0;
  assign _T_585 = _T_566 ? _T_516 : 9'h0;
  assign _T_586 = _T_583 ? _T_585 : _T_581;
  assign _T_588 = _T_586 == 9'h1;
  assign _T_589 = _T_89_w_ready & _T_89_w_valid;
  assign _GEN_55 = {{8'd0}, _T_589};
  assign _T_590 = _T_586 - _GEN_55;
  assign _T_591 = $unsigned(_T_590);
  assign _T_592 = _T_591[8:0];
  assign _T_595 = _T_589 == 1'h0;
  assign _T_597 = _T_586 != 9'h0;
  assign _T_598 = _T_595 | _T_597;
  assign _T_600 = _T_598 | reset;
  assign _T_602 = _T_600 == 1'h0;
  assign _T_604 = _T_564 == 1'h0;
  assign _T_605 = _T_604 | _T_566;
  assign _T_606 = _T_555_valid & _T_605;
  assign _T_610 = _T_89_w_ready & _T_605;
  assign _T_612 = _T_89_w_valid == 1'h0;
  assign _T_614 = _T_555_bits_last == 1'h0;
  assign _T_615 = _T_612 | _T_614;
  assign _T_616 = _T_615 | _T_588;
  assign _T_618 = _T_616 | reset;
  assign _T_620 = _T_618 == 1'h0;
  assign _T_621 = _T_89_r_bits_user[0];
  assign _T_622 = _T_89_r_bits_last & _T_621;
  assign _T_623 = _T_89_r_bits_user[7:1];
  assign _T_624 = _T_89_b_bits_user[0];
  assign _T_625 = _T_89_b_valid & _T_624;
  assign _T_627 = _T_624 == 1'h0;
  assign _T_628 = _T_31_b_ready | _T_627;
  assign _T_629 = _T_89_b_bits_user[7:1];
  assign _GEN_13 = _T_89_b_bits_id ? _T_647_1 : _T_647_0;
  assign _T_661 = _T_89_b_bits_resp | _GEN_0;
  assign _T_664 = 2'h1 << _T_89_b_bits_id;
  assign _T_666 = _T_664[0];
  assign _T_667 = _T_664[1];
  assign _T_668 = _T_89_b_ready & _T_89_b_valid;
  assign _T_669 = _T_666 & _T_668;
  assign _T_671 = _T_647_0 | _T_89_b_bits_resp;
  assign _T_672 = _T_624 ? 2'h0 : _T_671;
  assign _GEN_14 = _T_669 ? _T_672 : _T_647_0;
  assign _T_674 = _T_667 & _T_668;
  assign _T_676 = _T_647_1 | _T_89_b_bits_resp;
  assign _T_677 = _T_624 ? 2'h0 : _T_676;
  assign _GEN_15 = _T_674 ? _T_677 : _T_647_1;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_1_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = Queue_2_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_625;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_661;
  assign _T_31_b_bits_user = _T_629;
  assign _T_31_ar_ready = Queue_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_user = _T_623;
  assign _T_31_r_bits_last = _T_622;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_572;
  assign _T_89_aw_bits_id = _T_388_bits_id;
  assign _T_89_aw_bits_addr = _T_388_bits_addr;
  assign _T_89_aw_bits_len = _T_388_bits_len;
  assign _T_89_aw_bits_size = _T_388_bits_size;
  assign _T_89_aw_bits_user = _T_578;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_606;
  assign _T_89_w_bits_data = _T_555_bits_data;
  assign _T_89_w_bits_strb = _T_555_bits_strb;
  assign _T_89_w_bits_last = _T_588;
  assign _T_89_b_ready = _T_628;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_211_valid;
  assign _T_89_ar_bits_id = _T_211_bits_id;
  assign _T_89_ar_bits_addr = _T_211_bits_addr;
  assign _T_89_ar_bits_len = _T_211_bits_len;
  assign _T_89_ar_bits_size = _T_211_bits_size;
  assign _T_89_ar_bits_user = _T_559;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_31_ar_valid;
  assign Queue_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_io_enq_bits_len = _T_31_ar_bits_len;
  assign Queue_io_enq_bits_size = _T_31_ar_bits_size;
  assign Queue_io_enq_bits_burst = _T_31_ar_bits_burst;
  assign Queue_io_enq_bits_user = _T_31_ar_bits_user;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_365;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_len = Queue_io_deq_bits_len;
  assign _T_207_bits_size = Queue_io_deq_bits_size;
  assign _T_207_bits_burst = Queue_io_deq_bits_burst;
  assign _T_207_bits_user = Queue_io_deq_bits_user;
  assign _T_211_ready = _T_89_ar_ready;
  assign _T_211_valid = _T_207_valid;
  assign _T_211_bits_id = _T_207_bits_id;
  assign _T_211_bits_addr = _T_373;
  assign _T_211_bits_len = _T_338;
  assign _T_211_bits_size = _T_207_bits_size;
  assign _T_211_bits_user = _T_207_bits_user;
  assign _T_297 = _T_295;
  assign _T_354 = _GEN_2;
  assign Queue_1_io_enq_valid = _T_31_aw_valid;
  assign Queue_1_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_1_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_1_io_enq_bits_len = _T_31_aw_bits_len;
  assign Queue_1_io_enq_bits_size = _T_31_aw_bits_size;
  assign Queue_1_io_enq_bits_burst = _T_31_aw_bits_burst;
  assign Queue_1_io_enq_bits_user = _T_31_aw_bits_user;
  assign Queue_1_io_deq_ready = _T_384_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_384_ready = _T_536;
  assign _T_384_valid = Queue_1_io_deq_valid;
  assign _T_384_bits_id = Queue_1_io_deq_bits_id;
  assign _T_384_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_384_bits_len = Queue_1_io_deq_bits_len;
  assign _T_384_bits_size = Queue_1_io_deq_bits_size;
  assign _T_384_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_384_bits_user = Queue_1_io_deq_bits_user;
  assign _T_388_ready = _T_574;
  assign _T_388_valid = _T_384_valid;
  assign _T_388_bits_id = _T_384_bits_id;
  assign _T_388_bits_addr = _T_544;
  assign _T_388_bits_len = _T_509;
  assign _T_388_bits_size = _T_384_bits_size;
  assign _T_388_bits_user = _T_384_bits_user;
  assign _T_468 = _T_466;
  assign _T_525 = _GEN_7;
  assign Queue_2_io_enq_valid = _T_31_w_valid;
  assign Queue_2_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_2_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_2_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_2_io_deq_ready = _T_555_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_555_ready = _T_610;
  assign _T_555_valid = Queue_2_io_deq_valid;
  assign _T_555_bits_data = Queue_2_io_deq_bits_data;
  assign _T_555_bits_strb = Queue_2_io_deq_bits_strb;
  assign _T_555_bits_last = Queue_2_io_deq_bits_last;
  assign _T_564 = _T_583;
  assign _T_566 = _T_577;
  assign _GEN_0 = _GEN_13;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_217 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_219 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_221 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_394 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_396 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_398 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_562 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_581 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_647_0 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_647_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_217 <= 1'h0;
    end else begin
      if (_T_374) begin
        _T_217 <= _T_376;
      end
    end
    if (_T_374) begin
      _T_219 <= _T_354;
    end
    _T_221 <= _GEN_5[7:0];
    if (reset) begin
      _T_394 <= 1'h0;
    end else begin
      if (_T_545) begin
        _T_394 <= _T_547;
      end
    end
    if (_T_545) begin
      _T_396 <= _T_525;
    end
    _T_398 <= _GEN_10[7:0];
    if (reset) begin
      _T_562 <= 1'h0;
    end else begin
      if (_T_569) begin
        _T_562 <= 1'h0;
      end else begin
        if (_T_567) begin
          _T_562 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_581 <= 9'h0;
    end else begin
      _T_581 <= _T_592;
    end
    if (reset) begin
      _T_647_0 <= 2'h0;
    end else begin
      if (_T_669) begin
        if (_T_624) begin
          _T_647_0 <= 2'h0;
        end else begin
          _T_647_0 <= _T_671;
        end
      end
    end
    if (reset) begin
      _T_647_1 <= 2'h0;
    end else begin
      if (_T_674) begin
        if (_T_624) begin
          _T_647_1 <= 2'h0;
        end else begin
          _T_647_1 <= _T_676;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_602) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:166 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_602) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_620) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:175 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_620) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_1(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [7:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [7:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [7:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [7:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output [6:0]  auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [6:0]  auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output [6:0]  auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [6:0]  auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [7:0] _T_31_aw_bits_id;
  wire [31:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [7:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [7:0] _T_31_ar_bits_id;
  wire [31:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [7:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire  _T_89_aw_bits_id;
  wire [31:0] _T_89_aw_bits_addr;
  wire [7:0] _T_89_aw_bits_len;
  wire [2:0] _T_89_aw_bits_size;
  wire [1:0] _T_89_aw_bits_burst;
  wire [6:0] _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire  _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire [6:0] _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire  _T_89_ar_bits_id;
  wire [31:0] _T_89_ar_bits_addr;
  wire [7:0] _T_89_ar_bits_len;
  wire [2:0] _T_89_ar_bits_size;
  wire [1:0] _T_89_ar_bits_burst;
  wire [6:0] _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire  _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire [6:0] _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire [6:0] _T_203;
  wire [6:0] _T_204;
  wire [7:0] _T_205;
  wire [7:0] _T_206;
  assign _T_203 = _T_31_ar_bits_id[7:1];
  assign _T_204 = _T_31_aw_bits_id[7:1];
  assign _T_205 = {_T_89_r_bits_user,_T_89_r_bits_id};
  assign _T_206 = {_T_89_b_bits_user,_T_89_b_bits_id};
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_len = _T_89_aw_bits_len;
  assign auto_out_aw_bits_size = _T_89_aw_bits_size;
  assign auto_out_aw_bits_burst = _T_89_aw_bits_burst;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_len = _T_89_ar_bits_len;
  assign auto_out_ar_bits_size = _T_89_ar_bits_size;
  assign auto_out_ar_bits_burst = _T_89_ar_bits_burst;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = _T_89_aw_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_w_ready = _T_89_w_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_89_b_valid;
  assign _T_31_b_bits_id = _T_206;
  assign _T_31_b_bits_resp = _T_89_b_bits_resp;
  assign _T_31_ar_ready = _T_89_ar_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_205;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_last = _T_89_r_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_31_aw_valid;
  assign _T_89_aw_bits_id = _T_31_aw_bits_id[0];
  assign _T_89_aw_bits_addr = _T_31_aw_bits_addr;
  assign _T_89_aw_bits_len = _T_31_aw_bits_len;
  assign _T_89_aw_bits_size = _T_31_aw_bits_size;
  assign _T_89_aw_bits_burst = _T_31_aw_bits_burst;
  assign _T_89_aw_bits_user = _T_204;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_31_w_valid;
  assign _T_89_w_bits_data = _T_31_w_bits_data;
  assign _T_89_w_bits_strb = _T_31_w_bits_strb;
  assign _T_89_w_bits_last = _T_31_w_bits_last;
  assign _T_89_b_ready = _T_31_b_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_31_ar_valid;
  assign _T_89_ar_bits_id = _T_31_ar_bits_id[0];
  assign _T_89_ar_bits_addr = _T_31_ar_bits_addr;
  assign _T_89_ar_bits_len = _T_31_ar_bits_len;
  assign _T_89_ar_bits_size = _T_31_ar_bits_size;
  assign _T_89_ar_bits_burst = _T_31_ar_bits_burst;
  assign _T_89_ar_bits_user = _T_203;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
endmodule
module TLROM_bootrom(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [1:0]  auto_in_a_bits_size,
  input  [8:0]  auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [8:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data
);
  wire  in_a_ready;
  wire  in_a_valid;
  wire [1:0] in_a_bits_size;
  wire [8:0] in_a_bits_source;
  wire [16:0] in_a_bits_address;
  wire  in_d_ready;
  wire  in_d_valid;
  wire [1:0] in_d_bits_size;
  wire [8:0] in_d_bits_source;
  wire [63:0] in_d_bits_data;
  wire [8:0] index;
  wire [3:0] high;
  wire  _T_1145;
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire [63:0] _GEN_5;
  wire [63:0] _GEN_6;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire [63:0] _GEN_17;
  wire [63:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire [63:0] _GEN_26;
  wire [63:0] _GEN_27;
  wire [63:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire [63:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [63:0] _GEN_35;
  wire [63:0] _GEN_36;
  wire [63:0] _GEN_37;
  wire [63:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [63:0] _GEN_40;
  wire [63:0] _GEN_41;
  wire [63:0] _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [63:0] _GEN_45;
  wire [63:0] _GEN_46;
  wire [63:0] _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [63:0] _GEN_50;
  wire [63:0] _GEN_51;
  wire [63:0] _GEN_52;
  wire [63:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [63:0] _GEN_55;
  wire [63:0] _GEN_56;
  wire [63:0] _GEN_57;
  wire [63:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [63:0] _GEN_60;
  wire [63:0] _GEN_61;
  wire [63:0] _GEN_62;
  wire [63:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [63:0] _GEN_65;
  wire [63:0] _GEN_66;
  wire [63:0] _GEN_67;
  wire [63:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [63:0] _GEN_70;
  wire [63:0] _GEN_71;
  wire [63:0] _GEN_72;
  wire [63:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [63:0] _GEN_75;
  wire [63:0] _GEN_76;
  wire [63:0] _GEN_77;
  wire [63:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [63:0] _GEN_80;
  wire [63:0] _GEN_81;
  wire [63:0] _GEN_82;
  wire [63:0] _GEN_83;
  wire [63:0] _GEN_84;
  wire [63:0] _GEN_85;
  wire [63:0] _GEN_86;
  wire [63:0] _GEN_87;
  wire [63:0] _GEN_88;
  wire [63:0] _GEN_89;
  wire [63:0] _GEN_90;
  wire [63:0] _GEN_91;
  wire [63:0] _GEN_92;
  wire [63:0] _GEN_93;
  wire [63:0] _GEN_94;
  wire [63:0] _GEN_95;
  wire [63:0] _GEN_96;
  wire [63:0] _GEN_97;
  wire [63:0] _GEN_98;
  wire [63:0] _GEN_99;
  wire [63:0] _GEN_100;
  wire [63:0] _GEN_101;
  wire [63:0] _GEN_102;
  wire [63:0] _GEN_103;
  wire [63:0] _GEN_104;
  wire [63:0] _GEN_105;
  wire [63:0] _GEN_106;
  wire [63:0] _GEN_107;
  wire [63:0] _GEN_108;
  wire [63:0] _GEN_109;
  wire [63:0] _GEN_110;
  wire [63:0] _GEN_111;
  wire [63:0] _GEN_112;
  wire [63:0] _GEN_113;
  wire [63:0] _GEN_114;
  wire [63:0] _GEN_115;
  wire [63:0] _GEN_116;
  wire [63:0] _GEN_117;
  wire [63:0] _GEN_118;
  wire [63:0] _GEN_119;
  wire [63:0] _GEN_120;
  wire [63:0] _GEN_121;
  wire [63:0] _GEN_122;
  wire [63:0] _GEN_123;
  wire [63:0] _GEN_124;
  wire [63:0] _GEN_125;
  wire [63:0] _GEN_126;
  wire [63:0] _GEN_127;
  wire [63:0] _GEN_128;
  wire [63:0] _GEN_129;
  wire [63:0] _GEN_130;
  wire [63:0] _GEN_131;
  wire [63:0] _GEN_132;
  wire [63:0] _GEN_133;
  wire [63:0] _GEN_134;
  wire [63:0] _GEN_135;
  wire [63:0] _GEN_136;
  wire [63:0] _GEN_137;
  wire [63:0] _GEN_138;
  wire [63:0] _GEN_139;
  wire [63:0] _GEN_140;
  wire [63:0] _GEN_141;
  wire [63:0] _GEN_142;
  wire [63:0] _GEN_143;
  wire [63:0] _GEN_144;
  wire [63:0] _GEN_145;
  wire [63:0] _GEN_146;
  wire [63:0] _GEN_147;
  wire [63:0] _GEN_148;
  wire [63:0] _GEN_149;
  wire [63:0] _GEN_150;
  wire [63:0] _GEN_151;
  wire [63:0] _GEN_152;
  wire [63:0] _GEN_153;
  wire [63:0] _GEN_154;
  wire [63:0] _GEN_155;
  wire [63:0] _GEN_156;
  wire [63:0] _GEN_157;
  wire [63:0] _GEN_158;
  wire [63:0] _GEN_159;
  wire [63:0] _GEN_160;
  wire [63:0] _GEN_161;
  wire [63:0] _GEN_162;
  wire [63:0] _GEN_163;
  wire [63:0] _GEN_164;
  wire [63:0] _GEN_165;
  wire [63:0] _GEN_166;
  wire [63:0] _GEN_167;
  wire [63:0] _GEN_168;
  wire [63:0] _GEN_169;
  wire [63:0] _GEN_170;
  wire [63:0] _GEN_171;
  wire [63:0] _GEN_172;
  wire [63:0] _GEN_173;
  wire [63:0] _GEN_174;
  wire [63:0] _GEN_175;
  wire [63:0] _GEN_176;
  wire [63:0] _GEN_177;
  wire [63:0] _GEN_178;
  wire [63:0] _GEN_179;
  wire [63:0] _GEN_180;
  wire [63:0] _GEN_181;
  wire [63:0] _GEN_182;
  wire [63:0] _GEN_183;
  wire [63:0] _GEN_184;
  wire [63:0] _GEN_185;
  wire [63:0] _GEN_186;
  wire [63:0] _GEN_187;
  wire [63:0] _GEN_188;
  wire [63:0] _GEN_189;
  wire [63:0] _GEN_190;
  wire [63:0] _GEN_191;
  wire [63:0] _GEN_192;
  wire [63:0] _GEN_193;
  wire [63:0] _GEN_194;
  wire [63:0] _GEN_195;
  wire [63:0] _GEN_196;
  wire [63:0] _GEN_197;
  wire [63:0] _GEN_198;
  wire [63:0] _GEN_199;
  wire [63:0] _GEN_200;
  wire [63:0] _GEN_201;
  wire [63:0] _GEN_202;
  wire [63:0] _GEN_203;
  wire [63:0] _GEN_204;
  wire [63:0] _GEN_205;
  wire [63:0] _GEN_206;
  wire [63:0] _GEN_207;
  wire [63:0] _GEN_208;
  wire [63:0] _GEN_209;
  wire [63:0] _GEN_210;
  wire [63:0] _GEN_211;
  wire [63:0] _GEN_212;
  wire [63:0] _GEN_213;
  wire [63:0] _GEN_214;
  wire [63:0] _GEN_215;
  wire [63:0] _GEN_216;
  wire [63:0] _GEN_217;
  wire [63:0] _GEN_218;
  wire [63:0] _GEN_219;
  wire [63:0] _GEN_220;
  wire [63:0] _GEN_221;
  wire [63:0] _GEN_222;
  wire [63:0] _GEN_223;
  wire [63:0] _GEN_224;
  wire [63:0] _GEN_225;
  wire [63:0] _GEN_226;
  wire [63:0] _GEN_227;
  wire [63:0] _GEN_228;
  wire [63:0] _GEN_229;
  wire [63:0] _GEN_230;
  wire [63:0] _GEN_231;
  wire [63:0] _GEN_232;
  wire [63:0] _GEN_233;
  wire [63:0] _GEN_234;
  wire [63:0] _GEN_235;
  wire [63:0] _GEN_236;
  wire [63:0] _GEN_237;
  wire [63:0] _GEN_238;
  wire [63:0] _GEN_239;
  wire [63:0] _GEN_240;
  wire [63:0] _GEN_241;
  wire [63:0] _GEN_242;
  wire [63:0] _GEN_243;
  wire [63:0] _GEN_244;
  wire [63:0] _GEN_245;
  wire [63:0] _GEN_246;
  wire [63:0] _GEN_247;
  wire [63:0] _GEN_248;
  wire [63:0] _GEN_249;
  wire [63:0] _GEN_250;
  wire [63:0] _GEN_251;
  wire [63:0] _GEN_252;
  wire [63:0] _GEN_253;
  wire [63:0] _GEN_254;
  wire [63:0] _GEN_255;
  wire [63:0] _GEN_256;
  wire [63:0] _GEN_257;
  wire [63:0] _GEN_258;
  wire [63:0] _GEN_259;
  wire [63:0] _GEN_260;
  wire [63:0] _GEN_261;
  wire [63:0] _GEN_262;
  wire [63:0] _GEN_263;
  wire [63:0] _GEN_264;
  wire [63:0] _GEN_265;
  wire [63:0] _GEN_266;
  wire [63:0] _GEN_267;
  wire [63:0] _GEN_268;
  wire [63:0] _GEN_269;
  wire [63:0] _GEN_270;
  wire [63:0] _GEN_271;
  wire [63:0] _GEN_272;
  wire [63:0] _GEN_273;
  wire [63:0] _GEN_274;
  wire [63:0] _GEN_275;
  wire [63:0] _GEN_276;
  wire [63:0] _GEN_277;
  wire [63:0] _GEN_278;
  wire [63:0] _GEN_279;
  wire [63:0] _GEN_280;
  wire [63:0] _GEN_281;
  wire [63:0] _GEN_282;
  wire [63:0] _GEN_283;
  wire [63:0] _GEN_284;
  wire [63:0] _GEN_285;
  wire [63:0] _GEN_286;
  wire [63:0] _GEN_287;
  wire [63:0] _GEN_288;
  wire [63:0] _GEN_289;
  wire [63:0] _GEN_290;
  wire [63:0] _GEN_291;
  wire [63:0] _GEN_292;
  wire [63:0] _GEN_293;
  wire [63:0] _GEN_294;
  wire [63:0] _GEN_295;
  wire [63:0] _GEN_296;
  wire [63:0] _GEN_297;
  wire [63:0] _GEN_298;
  wire [63:0] _GEN_299;
  wire [63:0] _GEN_300;
  wire [63:0] _GEN_301;
  wire [63:0] _GEN_302;
  wire [63:0] _GEN_303;
  wire [63:0] _GEN_304;
  wire [63:0] _GEN_305;
  wire [63:0] _GEN_306;
  wire [63:0] _GEN_307;
  wire [63:0] _GEN_308;
  wire [63:0] _GEN_309;
  wire [63:0] _GEN_310;
  wire [63:0] _GEN_311;
  wire [63:0] _GEN_312;
  wire [63:0] _GEN_313;
  wire [63:0] _GEN_314;
  wire [63:0] _GEN_315;
  wire [63:0] _GEN_316;
  wire [63:0] _GEN_317;
  wire [63:0] _GEN_318;
  wire [63:0] _GEN_319;
  wire [63:0] _GEN_320;
  wire [63:0] _GEN_321;
  wire [63:0] _GEN_322;
  wire [63:0] _GEN_323;
  wire [63:0] _GEN_324;
  wire [63:0] _GEN_325;
  wire [63:0] _GEN_326;
  wire [63:0] _GEN_327;
  wire [63:0] _GEN_328;
  wire [63:0] _GEN_329;
  wire [63:0] _GEN_330;
  wire [63:0] _GEN_331;
  wire [63:0] _GEN_332;
  wire [63:0] _GEN_333;
  wire [63:0] _GEN_334;
  wire [63:0] _GEN_335;
  wire [63:0] _GEN_336;
  wire [63:0] _GEN_337;
  wire [63:0] _GEN_338;
  wire [63:0] _GEN_339;
  wire [63:0] _GEN_340;
  wire [63:0] _GEN_341;
  wire [63:0] _GEN_342;
  wire [63:0] _GEN_343;
  wire [63:0] _GEN_344;
  wire [63:0] _GEN_345;
  wire [63:0] _GEN_346;
  wire [63:0] _GEN_347;
  wire [63:0] _GEN_348;
  wire [63:0] _GEN_349;
  wire [63:0] _GEN_350;
  wire [63:0] _GEN_351;
  wire [63:0] _GEN_352;
  wire [63:0] _GEN_353;
  wire [63:0] _GEN_354;
  wire [63:0] _GEN_355;
  wire [63:0] _GEN_356;
  wire [63:0] _GEN_357;
  wire [63:0] _GEN_358;
  wire [63:0] _GEN_359;
  wire [63:0] _GEN_360;
  wire [63:0] _GEN_361;
  wire [63:0] _GEN_362;
  wire [63:0] _GEN_363;
  wire [63:0] _GEN_364;
  wire [63:0] _GEN_365;
  wire [63:0] _GEN_366;
  wire [63:0] _GEN_367;
  wire [63:0] _GEN_368;
  wire [63:0] _GEN_369;
  wire [63:0] _GEN_370;
  wire [63:0] _GEN_371;
  wire [63:0] _GEN_372;
  wire [63:0] _GEN_373;
  wire [63:0] _GEN_374;
  wire [63:0] _GEN_375;
  wire [63:0] _GEN_376;
  wire [63:0] _GEN_377;
  wire [63:0] _GEN_378;
  wire [63:0] _GEN_379;
  wire [63:0] _GEN_380;
  wire [63:0] _GEN_381;
  wire [63:0] _GEN_382;
  wire [63:0] _GEN_383;
  wire [63:0] _GEN_384;
  wire [63:0] _GEN_385;
  wire [63:0] _GEN_386;
  wire [63:0] _GEN_387;
  wire [63:0] _GEN_388;
  wire [63:0] _GEN_389;
  wire [63:0] _GEN_390;
  wire [63:0] _GEN_391;
  wire [63:0] _GEN_392;
  wire [63:0] _GEN_393;
  wire [63:0] _GEN_394;
  wire [63:0] _GEN_395;
  wire [63:0] _GEN_396;
  wire [63:0] _GEN_397;
  wire [63:0] _GEN_398;
  wire [63:0] _GEN_399;
  wire [63:0] _GEN_400;
  wire [63:0] _GEN_401;
  wire [63:0] _GEN_402;
  wire [63:0] _GEN_403;
  wire [63:0] _GEN_404;
  wire [63:0] _GEN_405;
  wire [63:0] _GEN_406;
  wire [63:0] _GEN_407;
  wire [63:0] _GEN_408;
  wire [63:0] _GEN_409;
  wire [63:0] _GEN_410;
  wire [63:0] _GEN_411;
  wire [63:0] _GEN_412;
  wire [63:0] _GEN_413;
  wire [63:0] _GEN_414;
  wire [63:0] _GEN_415;
  wire [63:0] _GEN_416;
  wire [63:0] _GEN_417;
  wire [63:0] _GEN_418;
  wire [63:0] _GEN_419;
  wire [63:0] _GEN_420;
  wire [63:0] _GEN_421;
  wire [63:0] _GEN_422;
  wire [63:0] _GEN_423;
  wire [63:0] _GEN_424;
  wire [63:0] _GEN_425;
  wire [63:0] _GEN_426;
  wire [63:0] _GEN_427;
  wire [63:0] _GEN_428;
  wire [63:0] _GEN_429;
  wire [63:0] _GEN_430;
  wire [63:0] _GEN_431;
  wire [63:0] _GEN_432;
  wire [63:0] _GEN_433;
  wire [63:0] _GEN_434;
  wire [63:0] _GEN_435;
  wire [63:0] _GEN_436;
  wire [63:0] _GEN_437;
  wire [63:0] _GEN_438;
  wire [63:0] _GEN_439;
  wire [63:0] _GEN_440;
  wire [63:0] _GEN_441;
  wire [63:0] _GEN_442;
  wire [63:0] _GEN_443;
  wire [63:0] _GEN_444;
  wire [63:0] _GEN_445;
  wire [63:0] _GEN_446;
  wire [63:0] _GEN_447;
  wire [63:0] _GEN_448;
  wire [63:0] _GEN_449;
  wire [63:0] _GEN_450;
  wire [63:0] _GEN_451;
  wire [63:0] _GEN_452;
  wire [63:0] _GEN_453;
  wire [63:0] _GEN_454;
  wire [63:0] _GEN_455;
  wire [63:0] _GEN_456;
  wire [63:0] _GEN_457;
  wire [63:0] _GEN_458;
  wire [63:0] _GEN_459;
  wire [63:0] _GEN_460;
  wire [63:0] _GEN_461;
  wire [63:0] _GEN_462;
  wire [63:0] _GEN_463;
  wire [63:0] _GEN_464;
  wire [63:0] _GEN_465;
  wire [63:0] _GEN_466;
  wire [63:0] _GEN_467;
  wire [63:0] _GEN_468;
  wire [63:0] _GEN_469;
  wire [63:0] _GEN_470;
  wire [63:0] _GEN_471;
  wire [63:0] _GEN_472;
  wire [63:0] _GEN_473;
  wire [63:0] _GEN_474;
  wire [63:0] _GEN_475;
  wire [63:0] _GEN_476;
  wire [63:0] _GEN_477;
  wire [63:0] _GEN_478;
  wire [63:0] _GEN_479;
  wire [63:0] _GEN_480;
  wire [63:0] _GEN_481;
  wire [63:0] _GEN_482;
  wire [63:0] _GEN_483;
  wire [63:0] _GEN_484;
  wire [63:0] _GEN_485;
  wire [63:0] _GEN_486;
  wire [63:0] _GEN_487;
  wire [63:0] _GEN_488;
  wire [63:0] _GEN_489;
  wire [63:0] _GEN_490;
  wire [63:0] _GEN_491;
  wire [63:0] _GEN_492;
  wire [63:0] _GEN_493;
  wire [63:0] _GEN_494;
  wire [63:0] _GEN_495;
  wire [63:0] _GEN_496;
  wire [63:0] _GEN_497;
  wire [63:0] _GEN_498;
  wire [63:0] _GEN_499;
  wire [63:0] _GEN_500;
  wire [63:0] _GEN_501;
  wire [63:0] _GEN_502;
  wire [63:0] _GEN_503;
  wire [63:0] _GEN_504;
  wire [63:0] _GEN_505;
  wire [63:0] _GEN_506;
  wire [63:0] _GEN_507;
  wire [63:0] _GEN_508;
  wire [63:0] _GEN_509;
  wire [63:0] _GEN_510;
  wire [63:0] _GEN_511;
  wire [63:0] _T_1148;
  wire [1:0] _T_1151_size;
  wire [8:0] _T_1151_source;
  wire [63:0] _T_1151_data;
  assign index = in_a_bits_address[11:3];
  assign high = in_a_bits_address[15:12];
  assign _T_1145 = high != 4'h0;
  assign _GEN_1 = 9'h1 == index ? 64'h597f1402573 : 64'h1f414130010041b;
  assign _GEN_2 = 9'h2 == index ? 64'h840207458593 : _GEN_1;
  assign _GEN_3 = 9'h3 == index ? 64'h0 : _GEN_2;
  assign _GEN_4 = 9'h4 == index ? 64'h0 : _GEN_3;
  assign _GEN_5 = 9'h5 == index ? 64'h0 : _GEN_4;
  assign _GEN_6 = 9'h6 == index ? 64'h0 : _GEN_5;
  assign _GEN_7 = 9'h7 == index ? 64'h0 : _GEN_6;
  assign _GEN_8 = 9'h8 == index ? 64'h597f1402573 : _GEN_7;
  assign _GEN_9 = 9'h9 == index ? 64'h1050007303c58593 : _GEN_8;
  assign _GEN_10 = 9'ha == index ? 64'hbff5 : _GEN_9;
  assign _GEN_11 = 9'hb == index ? 64'h0 : _GEN_10;
  assign _GEN_12 = 9'hc == index ? 64'h0 : _GEN_11;
  assign _GEN_13 = 9'hd == index ? 64'h0 : _GEN_12;
  assign _GEN_14 = 9'he == index ? 64'h0 : _GEN_13;
  assign _GEN_15 = 9'hf == index ? 64'h0 : _GEN_14;
  assign _GEN_16 = 9'h10 == index ? 64'h4c080000edfe0dd0 : _GEN_15;
  assign _GEN_17 = 9'h11 == index ? 64'hb806000038000000 : _GEN_16;
  assign _GEN_18 = 9'h12 == index ? 64'h1100000028000000 : _GEN_17;
  assign _GEN_19 = 9'h13 == index ? 64'h10000000 : _GEN_18;
  assign _GEN_20 = 9'h14 == index ? 64'h8006000094010000 : _GEN_19;
  assign _GEN_21 = 9'h15 == index ? 64'h0 : _GEN_20;
  assign _GEN_22 = 9'h16 == index ? 64'h0 : _GEN_21;
  assign _GEN_23 = 9'h17 == index ? 64'h1000000 : _GEN_22;
  assign _GEN_24 = 9'h18 == index ? 64'h400000003000000 : _GEN_23;
  assign _GEN_25 = 9'h19 == index ? 64'h100000000000000 : _GEN_24;
  assign _GEN_26 = 9'h1a == index ? 64'h400000003000000 : _GEN_25;
  assign _GEN_27 = 9'h1b == index ? 64'h10000000f000000 : _GEN_26;
  assign _GEN_28 = 9'h1c == index ? 64'h2100000003000000 : _GEN_27;
  assign _GEN_29 = 9'h1d == index ? 64'h656572661b000000 : _GEN_28;
  assign _GEN_30 = 9'h1e == index ? 64'h6f722c7370696863 : _GEN_29;
  assign _GEN_31 = 9'h1f == index ? 64'h7069686374656b63 : _GEN_30;
  assign _GEN_32 = 9'h20 == index ? 64'h6e776f6e6b6e752d : _GEN_31;
  assign _GEN_33 = 9'h21 == index ? 64'h7665642d : _GEN_32;
  assign _GEN_34 = 9'h22 == index ? 64'h1d00000003000000 : _GEN_33;
  assign _GEN_35 = 9'h23 == index ? 64'h6565726626000000 : _GEN_34;
  assign _GEN_36 = 9'h24 == index ? 64'h6f722c7370696863 : _GEN_35;
  assign _GEN_37 = 9'h25 == index ? 64'h7069686374656b63 : _GEN_36;
  assign _GEN_38 = 9'h26 == index ? 64'h6e776f6e6b6e752d : _GEN_37;
  assign _GEN_39 = 9'h27 == index ? 64'h100000000000000 : _GEN_38;
  assign _GEN_40 = 9'h28 == index ? 64'h73757063 : _GEN_39;
  assign _GEN_41 = 9'h29 == index ? 64'h400000003000000 : _GEN_40;
  assign _GEN_42 = 9'h2a == index ? 64'h100000000000000 : _GEN_41;
  assign _GEN_43 = 9'h2b == index ? 64'h400000003000000 : _GEN_42;
  assign _GEN_44 = 9'h2c == index ? 64'hf000000 : _GEN_43;
  assign _GEN_45 = 9'h2d == index ? 64'h4075706301000000 : _GEN_44;
  assign _GEN_46 = 9'h2e == index ? 64'h300000000000030 : _GEN_45;
  assign _GEN_47 = 9'h2f == index ? 64'h2c00000004000000 : _GEN_46;
  assign _GEN_48 = 9'h30 == index ? 64'h300000000000000 : _GEN_47;
  assign _GEN_49 = 9'h31 == index ? 64'h1b00000015000000 : _GEN_48;
  assign _GEN_50 = 9'h32 == index ? 64'h722c657669666973 : _GEN_49;
  assign _GEN_51 = 9'h33 == index ? 64'h72003074656b636f : _GEN_50;
  assign _GEN_52 = 9'h34 == index ? 64'h76637369 : _GEN_51;
  assign _GEN_53 = 9'h35 == index ? 64'h400000003000000 : _GEN_52;
  assign _GEN_54 = 9'h36 == index ? 64'h400000003c000000 : _GEN_53;
  assign _GEN_55 = 9'h37 == index ? 64'h400000003000000 : _GEN_54;
  assign _GEN_56 = 9'h38 == index ? 64'h400000004f000000 : _GEN_55;
  assign _GEN_57 = 9'h39 == index ? 64'h400000003000000 : _GEN_56;
  assign _GEN_58 = 9'h3a == index ? 64'h8000005c000000 : _GEN_57;
  assign _GEN_59 = 9'h3b == index ? 64'h400000003000000 : _GEN_58;
  assign _GEN_60 = 9'h3c == index ? 64'h100000069000000 : _GEN_59;
  assign _GEN_61 = 9'h3d == index ? 64'h400000003000000 : _GEN_60;
  assign _GEN_62 = 9'h3e == index ? 64'h1000000074000000 : _GEN_61;
  assign _GEN_63 = 9'h3f == index ? 64'h400000003000000 : _GEN_62;
  assign _GEN_64 = 9'h40 == index ? 64'h7570637f000000 : _GEN_63;
  assign _GEN_65 = 9'h41 == index ? 64'h400000003000000 : _GEN_64;
  assign _GEN_66 = 9'h42 == index ? 64'h400000008b000000 : _GEN_65;
  assign _GEN_67 = 9'h43 == index ? 64'h400000003000000 : _GEN_66;
  assign _GEN_68 = 9'h44 == index ? 64'h400000009e000000 : _GEN_67;
  assign _GEN_69 = 9'h45 == index ? 64'h400000003000000 : _GEN_68;
  assign _GEN_70 = 9'h46 == index ? 64'h800000ab000000 : _GEN_69;
  assign _GEN_71 = 9'h47 == index ? 64'h400000003000000 : _GEN_70;
  assign _GEN_72 = 9'h48 == index ? 64'h1000000b8000000 : _GEN_71;
  assign _GEN_73 = 9'h49 == index ? 64'h400000003000000 : _GEN_72;
  assign _GEN_74 = 9'h4a == index ? 64'h20000000c3000000 : _GEN_73;
  assign _GEN_75 = 9'h4b == index ? 64'hb00000003000000 : _GEN_74;
  assign _GEN_76 = 9'h4c == index ? 64'h63736972ce000000 : _GEN_75;
  assign _GEN_77 = 9'h4d == index ? 64'h393376732c76 : _GEN_76;
  assign _GEN_78 = 9'h4e == index ? 64'h800000003000000 : _GEN_77;
  assign _GEN_79 = 9'h4f == index ? 64'h1000000d7000000 : _GEN_78;
  assign _GEN_80 = 9'h50 == index ? 64'h300000002000000 : _GEN_79;
  assign _GEN_81 = 9'h51 == index ? 64'he800000004000000 : _GEN_80;
  assign _GEN_82 = 9'h52 == index ? 64'h300000000000000 : _GEN_81;
  assign _GEN_83 = 9'h53 == index ? 64'hec0000000a000000 : _GEN_82;
  assign _GEN_84 = 9'h54 == index ? 64'h66616d6934367672 : _GEN_83;
  assign _GEN_85 = 9'h55 == index ? 64'h300000000000064 : _GEN_84;
  assign _GEN_86 = 9'h56 == index ? 64'hf600000005000000 : _GEN_85;
  assign _GEN_87 = 9'h57 == index ? 64'h79616b6f : _GEN_86;
  assign _GEN_88 = 9'h58 == index ? 64'h3000000 : _GEN_87;
  assign _GEN_89 = 9'h59 == index ? 64'h1000000fd000000 : _GEN_88;
  assign _GEN_90 = 9'h5a == index ? 64'h7075727265746e69 : _GEN_89;
  assign _GEN_91 = 9'h5b == index ? 64'h6f72746e6f632d74 : _GEN_90;
  assign _GEN_92 = 9'h5c == index ? 64'h72656c6c : _GEN_91;
  assign _GEN_93 = 9'h5d == index ? 64'h400000003000000 : _GEN_92;
  assign _GEN_94 = 9'h5e == index ? 64'h100000007010000 : _GEN_93;
  assign _GEN_95 = 9'h5f == index ? 64'hf00000003000000 : _GEN_94;
  assign _GEN_96 = 9'h60 == index ? 64'h637369721b000000 : _GEN_95;
  assign _GEN_97 = 9'h61 == index ? 64'h6e692d7570632c76 : _GEN_96;
  assign _GEN_98 = 9'h62 == index ? 64'h300000000006374 : _GEN_97;
  assign _GEN_99 = 9'h63 == index ? 64'h1801000000000000 : _GEN_98;
  assign _GEN_100 = 9'h64 == index ? 64'h400000003000000 : _GEN_99;
  assign _GEN_101 = 9'h65 == index ? 64'h30000002d010000 : _GEN_100;
  assign _GEN_102 = 9'h66 == index ? 64'h200000002000000 : _GEN_101;
  assign _GEN_103 = 9'h67 == index ? 64'h100000002000000 : _GEN_102;
  assign _GEN_104 = 9'h68 == index ? 64'h384079726f6d656d : _GEN_103;
  assign _GEN_105 = 9'h69 == index ? 64'h30303030303030 : _GEN_104;
  assign _GEN_106 = 9'h6a == index ? 64'h700000003000000 : _GEN_105;
  assign _GEN_107 = 9'h6b == index ? 64'h6f6d656d7f000000 : _GEN_106;
  assign _GEN_108 = 9'h6c == index ? 64'h300000000007972 : _GEN_107;
  assign _GEN_109 = 9'h6d == index ? 64'he800000008000000 : _GEN_108;
  assign _GEN_110 = 9'h6e == index ? 64'h1000000080 : _GEN_109;
  assign _GEN_111 = 9'h6f == index ? 64'h400000003000000 : _GEN_110;
  assign _GEN_112 = 9'h70 == index ? 64'h20000002d010000 : _GEN_111;
  assign _GEN_113 = 9'h71 == index ? 64'h100000002000000 : _GEN_112;
  assign _GEN_114 = 9'h72 == index ? 64'h300000000636f73 : _GEN_113;
  assign _GEN_115 = 9'h73 == index ? 64'h4000000 : _GEN_114;
  assign _GEN_116 = 9'h74 == index ? 64'h300000001000000 : _GEN_115;
  assign _GEN_117 = 9'h75 == index ? 64'hf00000004000000 : _GEN_116;
  assign _GEN_118 = 9'h76 == index ? 64'h300000001000000 : _GEN_117;
  assign _GEN_119 = 9'h77 == index ? 64'h1b0000002c000000 : _GEN_118;
  assign _GEN_120 = 9'h78 == index ? 64'h7069686365657266 : _GEN_119;
  assign _GEN_121 = 9'h79 == index ? 64'h74656b636f722c73 : _GEN_120;
  assign _GEN_122 = 9'h7a == index ? 64'h6b6e752d70696863 : _GEN_121;
  assign _GEN_123 = 9'h7b == index ? 64'h636f732d6e776f6e : _GEN_122;
  assign _GEN_124 = 9'h7c == index ? 64'h2d656c706d697300 : _GEN_123;
  assign _GEN_125 = 9'h7d == index ? 64'h300000000737562 : _GEN_124;
  assign _GEN_126 = 9'h7e == index ? 64'h3501000000000000 : _GEN_125;
  assign _GEN_127 = 9'h7f == index ? 64'h6e696c6301000000 : _GEN_126;
  assign _GEN_128 = 9'h80 == index ? 64'h3030303030324074 : _GEN_127;
  assign _GEN_129 = 9'h81 == index ? 64'h300000000000030 : _GEN_128;
  assign _GEN_130 = 9'h82 == index ? 64'h1b0000000d000000 : _GEN_129;
  assign _GEN_131 = 9'h83 == index ? 64'h6c632c7663736972 : _GEN_130;
  assign _GEN_132 = 9'h84 == index ? 64'h30746e69 : _GEN_131;
  assign _GEN_133 = 9'h85 == index ? 64'h1000000003000000 : _GEN_132;
  assign _GEN_134 = 9'h86 == index ? 64'h30000003c010000 : _GEN_133;
  assign _GEN_135 = 9'h87 == index ? 64'h300000003000000 : _GEN_134;
  assign _GEN_136 = 9'h88 == index ? 64'h300000007000000 : _GEN_135;
  assign _GEN_137 = 9'h89 == index ? 64'he800000008000000 : _GEN_136;
  assign _GEN_138 = 9'h8a == index ? 64'h10000000002 : _GEN_137;
  assign _GEN_139 = 9'h8b == index ? 64'h800000003000000 : _GEN_138;
  assign _GEN_140 = 9'h8c == index ? 64'h746e6f6350010000 : _GEN_139;
  assign _GEN_141 = 9'h8d == index ? 64'h2000000006c6f72 : _GEN_140;
  assign _GEN_142 = 9'h8e == index ? 64'h7562656401000000 : _GEN_141;
  assign _GEN_143 = 9'h8f == index ? 64'h6f72746e6f632d67 : _GEN_142;
  assign _GEN_144 = 9'h90 == index ? 64'h304072656c6c : _GEN_143;
  assign _GEN_145 = 9'h91 == index ? 64'h2100000003000000 : _GEN_144;
  assign _GEN_146 = 9'h92 == index ? 64'h696669731b000000 : _GEN_145;
  assign _GEN_147 = 9'h93 == index ? 64'h67756265642c6576 : _GEN_146;
  assign _GEN_148 = 9'h94 == index ? 64'h736972003331302d : _GEN_147;
  assign _GEN_149 = 9'h95 == index ? 64'h67756265642c7663 : _GEN_148;
  assign _GEN_150 = 9'h96 == index ? 64'h3331302d : _GEN_149;
  assign _GEN_151 = 9'h97 == index ? 64'h800000003000000 : _GEN_150;
  assign _GEN_152 = 9'h98 == index ? 64'h30000003c010000 : _GEN_151;
  assign _GEN_153 = 9'h99 == index ? 64'h3000000ffff0000 : _GEN_152;
  assign _GEN_154 = 9'h9a == index ? 64'he800000008000000 : _GEN_153;
  assign _GEN_155 = 9'h9b == index ? 64'h10000000000000 : _GEN_154;
  assign _GEN_156 = 9'h9c == index ? 64'h800000003000000 : _GEN_155;
  assign _GEN_157 = 9'h9d == index ? 64'h746e6f6350010000 : _GEN_156;
  assign _GEN_158 = 9'h9e == index ? 64'h2000000006c6f72 : _GEN_157;
  assign _GEN_159 = 9'h9f == index ? 64'h6f72726501000000 : _GEN_158;
  assign _GEN_160 = 9'ha0 == index ? 64'h6563697665642d72 : _GEN_159;
  assign _GEN_161 = 9'ha1 == index ? 64'h3030303340 : _GEN_160;
  assign _GEN_162 = 9'ha2 == index ? 64'he00000003000000 : _GEN_161;
  assign _GEN_163 = 9'ha3 == index ? 64'h696669731b000000 : _GEN_162;
  assign _GEN_164 = 9'ha4 == index ? 64'h726f7272652c6576 : _GEN_163;
  assign _GEN_165 = 9'ha5 == index ? 64'h300000000000030 : _GEN_164;
  assign _GEN_166 = 9'ha6 == index ? 64'he800000008000000 : _GEN_165;
  assign _GEN_167 = 9'ha7 == index ? 64'h10000000300000 : _GEN_166;
  assign _GEN_168 = 9'ha8 == index ? 64'h400000003000000 : _GEN_167;
  assign _GEN_169 = 9'ha9 == index ? 64'h6d656d50010000 : _GEN_168;
  assign _GEN_170 = 9'haa == index ? 64'h400000003000000 : _GEN_169;
  assign _GEN_171 = 9'hab == index ? 64'h10000002d010000 : _GEN_170;
  assign _GEN_172 = 9'hac == index ? 64'h100000002000000 : _GEN_171;
  assign _GEN_173 = 9'had == index ? 64'h6c616e7265747865 : _GEN_172;
  assign _GEN_174 = 9'hae == index ? 64'h75727265746e692d : _GEN_173;
  assign _GEN_175 = 9'haf == index ? 64'h300000000737470 : _GEN_174;
  assign _GEN_176 = 9'hb0 == index ? 64'h5a01000004000000 : _GEN_175;
  assign _GEN_177 = 9'hb1 == index ? 64'h300000004000000 : _GEN_176;
  assign _GEN_178 = 9'hb2 == index ? 64'h6b01000008000000 : _GEN_177;
  assign _GEN_179 = 9'hb3 == index ? 64'h200000001000000 : _GEN_178;
  assign _GEN_180 = 9'hb4 == index ? 64'h100000002000000 : _GEN_179;
  assign _GEN_181 = 9'hb5 == index ? 64'h7075727265746e69 : _GEN_180;
  assign _GEN_182 = 9'hb6 == index ? 64'h6f72746e6f632d74 : _GEN_181;
  assign _GEN_183 = 9'hb7 == index ? 64'h3030634072656c6c : _GEN_182;
  assign _GEN_184 = 9'hb8 == index ? 64'h30303030 : _GEN_183;
  assign _GEN_185 = 9'hb9 == index ? 64'h400000003000000 : _GEN_184;
  assign _GEN_186 = 9'hba == index ? 64'h100000007010000 : _GEN_185;
  assign _GEN_187 = 9'hbb == index ? 64'hc00000003000000 : _GEN_186;
  assign _GEN_188 = 9'hbc == index ? 64'h637369721b000000 : _GEN_187;
  assign _GEN_189 = 9'hbd == index ? 64'h3063696c702c76 : _GEN_188;
  assign _GEN_190 = 9'hbe == index ? 64'h3000000 : _GEN_189;
  assign _GEN_191 = 9'hbf == index ? 64'h300000018010000 : _GEN_190;
  assign _GEN_192 = 9'hc0 == index ? 64'h3c01000010000000 : _GEN_191;
  assign _GEN_193 = 9'hc1 == index ? 64'hb00000003000000 : _GEN_192;
  assign _GEN_194 = 9'hc2 == index ? 64'h900000003000000 : _GEN_193;
  assign _GEN_195 = 9'hc3 == index ? 64'h800000003000000 : _GEN_194;
  assign _GEN_196 = 9'hc4 == index ? 64'hce8000000 : _GEN_195;
  assign _GEN_197 = 9'hc5 == index ? 64'h300000000000004 : _GEN_196;
  assign _GEN_198 = 9'hc6 == index ? 64'h5001000008000000 : _GEN_197;
  assign _GEN_199 = 9'hc7 == index ? 64'h6c6f72746e6f63 : _GEN_198;
  assign _GEN_200 = 9'hc8 == index ? 64'h400000003000000 : _GEN_199;
  assign _GEN_201 = 9'hc9 == index ? 64'h700000076010000 : _GEN_200;
  assign _GEN_202 = 9'hca == index ? 64'h400000003000000 : _GEN_201;
  assign _GEN_203 = 9'hcb == index ? 64'h200000089010000 : _GEN_202;
  assign _GEN_204 = 9'hcc == index ? 64'h400000003000000 : _GEN_203;
  assign _GEN_205 = 9'hcd == index ? 64'h40000002d010000 : _GEN_204;
  assign _GEN_206 = 9'hce == index ? 64'h100000002000000 : _GEN_205;
  assign _GEN_207 = 9'hcf == index ? 64'h303036406f696d6d : _GEN_206;
  assign _GEN_208 = 9'hd0 == index ? 64'h3030303030 : _GEN_207;
  assign _GEN_209 = 9'hd1 == index ? 64'h400000003000000 : _GEN_208;
  assign _GEN_210 = 9'hd2 == index ? 64'h100000000000000 : _GEN_209;
  assign _GEN_211 = 9'hd3 == index ? 64'h400000003000000 : _GEN_210;
  assign _GEN_212 = 9'hd4 == index ? 64'h10000000f000000 : _GEN_211;
  assign _GEN_213 = 9'hd5 == index ? 64'hb00000003000000 : _GEN_212;
  assign _GEN_214 = 9'hd6 == index ? 64'h706d69731b000000 : _GEN_213;
  assign _GEN_215 = 9'hd7 == index ? 64'h7375622d656c : _GEN_214;
  assign _GEN_216 = 9'hd8 == index ? 64'hc00000003000000 : _GEN_215;
  assign _GEN_217 = 9'hd9 == index ? 64'h6035010000 : _GEN_216;
  assign _GEN_218 = 9'hda == index ? 64'h2000000060 : _GEN_217;
  assign _GEN_219 = 9'hdb == index ? 64'h100000002000000 : _GEN_218;
  assign _GEN_220 = 9'hdc == index ? 64'h30303031406d6f72 : _GEN_219;
  assign _GEN_221 = 9'hdd == index ? 64'h300000000000030 : _GEN_220;
  assign _GEN_222 = 9'hde == index ? 64'h1b0000000c000000 : _GEN_221;
  assign _GEN_223 = 9'hdf == index ? 64'h722c657669666973 : _GEN_222;
  assign _GEN_224 = 9'he0 == index ? 64'h300000000306d6f : _GEN_223;
  assign _GEN_225 = 9'he1 == index ? 64'he800000008000000 : _GEN_224;
  assign _GEN_226 = 9'he2 == index ? 64'h10000000100 : _GEN_225;
  assign _GEN_227 = 9'he3 == index ? 64'h400000003000000 : _GEN_226;
  assign _GEN_228 = 9'he4 == index ? 64'h6d656d50010000 : _GEN_227;
  assign _GEN_229 = 9'he5 == index ? 64'h200000002000000 : _GEN_228;
  assign _GEN_230 = 9'he6 == index ? 64'h900000002000000 : _GEN_229;
  assign _GEN_231 = 9'he7 == index ? 64'h7373657264646123 : _GEN_230;
  assign _GEN_232 = 9'he8 == index ? 64'h2300736c6c65632d : _GEN_231;
  assign _GEN_233 = 9'he9 == index ? 64'h6c65632d657a6973 : _GEN_232;
  assign _GEN_234 = 9'hea == index ? 64'h61706d6f6300736c : _GEN_233;
  assign _GEN_235 = 9'heb == index ? 64'h6f6d00656c626974 : _GEN_234;
  assign _GEN_236 = 9'hec == index ? 64'h636f6c63006c6564 : _GEN_235;
  assign _GEN_237 = 9'hed == index ? 64'h6575716572662d6b : _GEN_236;
  assign _GEN_238 = 9'hee == index ? 64'h61632d640079636e : _GEN_237;
  assign _GEN_239 = 9'hef == index ? 64'h636f6c622d656863 : _GEN_238;
  assign _GEN_240 = 9'hf0 == index ? 64'h6400657a69732d6b : _GEN_239;
  assign _GEN_241 = 9'hf1 == index ? 64'h732d65686361632d : _GEN_240;
  assign _GEN_242 = 9'hf2 == index ? 64'h61632d6400737465 : _GEN_241;
  assign _GEN_243 = 9'hf3 == index ? 64'h657a69732d656863 : _GEN_242;
  assign _GEN_244 = 9'hf4 == index ? 64'h732d626c742d6400 : _GEN_243;
  assign _GEN_245 = 9'hf5 == index ? 64'h6c742d6400737465 : _GEN_244;
  assign _GEN_246 = 9'hf6 == index ? 64'h6400657a69732d62 : _GEN_245;
  assign _GEN_247 = 9'hf7 == index ? 64'h79745f6563697665 : _GEN_246;
  assign _GEN_248 = 9'hf8 == index ? 64'h6361632d69006570 : _GEN_247;
  assign _GEN_249 = 9'hf9 == index ? 64'h6b636f6c622d6568 : _GEN_248;
  assign _GEN_250 = 9'hfa == index ? 64'h2d6900657a69732d : _GEN_249;
  assign _GEN_251 = 9'hfb == index ? 64'h65732d6568636163 : _GEN_250;
  assign _GEN_252 = 9'hfc == index ? 64'h6361632d69007374 : _GEN_251;
  assign _GEN_253 = 9'hfd == index ? 64'h657a69732d6568 : _GEN_252;
  assign _GEN_254 = 9'hfe == index ? 64'h65732d626c742d69 : _GEN_253;
  assign _GEN_255 = 9'hff == index ? 64'h626c742d69007374 : _GEN_254;
  assign _GEN_256 = 9'h100 == index ? 64'h6d6d00657a69732d : _GEN_255;
  assign _GEN_257 = 9'h101 == index ? 64'h6e00657079742d75 : _GEN_256;
  assign _GEN_258 = 9'h102 == index ? 64'h6576656c2d747865 : _GEN_257;
  assign _GEN_259 = 9'h103 == index ? 64'h65686361632d6c : _GEN_258;
  assign _GEN_260 = 9'h104 == index ? 64'h6373697200676572 : _GEN_259;
  assign _GEN_261 = 9'h105 == index ? 64'h7473006173692c76 : _GEN_260;
  assign _GEN_262 = 9'h106 == index ? 64'h626c740073757461 : _GEN_261;
  assign _GEN_263 = 9'h107 == index ? 64'h230074696c70732d : _GEN_262;
  assign _GEN_264 = 9'h108 == index ? 64'h7075727265746e69 : _GEN_263;
  assign _GEN_265 = 9'h109 == index ? 64'h736c6c65632d74 : _GEN_264;
  assign _GEN_266 = 9'h10a == index ? 64'h7075727265746e69 : _GEN_265;
  assign _GEN_267 = 9'h10b == index ? 64'h6f72746e6f632d74 : _GEN_266;
  assign _GEN_268 = 9'h10c == index ? 64'h6168700072656c6c : _GEN_267;
  assign _GEN_269 = 9'h10d == index ? 64'h6e617200656c646e : _GEN_268;
  assign _GEN_270 = 9'h10e == index ? 64'h65746e6900736567 : _GEN_269;
  assign _GEN_271 = 9'h10f == index ? 64'h652d737470757272 : _GEN_270;
  assign _GEN_272 = 9'h110 == index ? 64'h6465646e657478 : _GEN_271;
  assign _GEN_273 = 9'h111 == index ? 64'h656d616e2d676572 : _GEN_272;
  assign _GEN_274 = 9'h112 == index ? 64'h727265746e690073 : _GEN_273;
  assign _GEN_275 = 9'h113 == index ? 64'h657261702d747075 : _GEN_274;
  assign _GEN_276 = 9'h114 == index ? 64'h7265746e6900746e : _GEN_275;
  assign _GEN_277 = 9'h115 == index ? 64'h6972007374707572 : _GEN_276;
  assign _GEN_278 = 9'h116 == index ? 64'h2d78616d2c766373 : _GEN_277;
  assign _GEN_279 = 9'h117 == index ? 64'h797469726f697270 : _GEN_278;
  assign _GEN_280 = 9'h118 == index ? 64'h6e2c766373697200 : _GEN_279;
  assign _GEN_281 = 9'h119 == index ? 64'h766564 : _GEN_280;
  assign _GEN_282 = 9'h11a == index ? 64'h0 : _GEN_281;
  assign _GEN_283 = 9'h11b == index ? 64'h0 : _GEN_282;
  assign _GEN_284 = 9'h11c == index ? 64'h0 : _GEN_283;
  assign _GEN_285 = 9'h11d == index ? 64'h0 : _GEN_284;
  assign _GEN_286 = 9'h11e == index ? 64'h0 : _GEN_285;
  assign _GEN_287 = 9'h11f == index ? 64'h0 : _GEN_286;
  assign _GEN_288 = 9'h120 == index ? 64'h0 : _GEN_287;
  assign _GEN_289 = 9'h121 == index ? 64'h0 : _GEN_288;
  assign _GEN_290 = 9'h122 == index ? 64'h0 : _GEN_289;
  assign _GEN_291 = 9'h123 == index ? 64'h0 : _GEN_290;
  assign _GEN_292 = 9'h124 == index ? 64'h0 : _GEN_291;
  assign _GEN_293 = 9'h125 == index ? 64'h0 : _GEN_292;
  assign _GEN_294 = 9'h126 == index ? 64'h0 : _GEN_293;
  assign _GEN_295 = 9'h127 == index ? 64'h0 : _GEN_294;
  assign _GEN_296 = 9'h128 == index ? 64'h0 : _GEN_295;
  assign _GEN_297 = 9'h129 == index ? 64'h0 : _GEN_296;
  assign _GEN_298 = 9'h12a == index ? 64'h0 : _GEN_297;
  assign _GEN_299 = 9'h12b == index ? 64'h0 : _GEN_298;
  assign _GEN_300 = 9'h12c == index ? 64'h0 : _GEN_299;
  assign _GEN_301 = 9'h12d == index ? 64'h0 : _GEN_300;
  assign _GEN_302 = 9'h12e == index ? 64'h0 : _GEN_301;
  assign _GEN_303 = 9'h12f == index ? 64'h0 : _GEN_302;
  assign _GEN_304 = 9'h130 == index ? 64'h0 : _GEN_303;
  assign _GEN_305 = 9'h131 == index ? 64'h0 : _GEN_304;
  assign _GEN_306 = 9'h132 == index ? 64'h0 : _GEN_305;
  assign _GEN_307 = 9'h133 == index ? 64'h0 : _GEN_306;
  assign _GEN_308 = 9'h134 == index ? 64'h0 : _GEN_307;
  assign _GEN_309 = 9'h135 == index ? 64'h0 : _GEN_308;
  assign _GEN_310 = 9'h136 == index ? 64'h0 : _GEN_309;
  assign _GEN_311 = 9'h137 == index ? 64'h0 : _GEN_310;
  assign _GEN_312 = 9'h138 == index ? 64'h0 : _GEN_311;
  assign _GEN_313 = 9'h139 == index ? 64'h0 : _GEN_312;
  assign _GEN_314 = 9'h13a == index ? 64'h0 : _GEN_313;
  assign _GEN_315 = 9'h13b == index ? 64'h0 : _GEN_314;
  assign _GEN_316 = 9'h13c == index ? 64'h0 : _GEN_315;
  assign _GEN_317 = 9'h13d == index ? 64'h0 : _GEN_316;
  assign _GEN_318 = 9'h13e == index ? 64'h0 : _GEN_317;
  assign _GEN_319 = 9'h13f == index ? 64'h0 : _GEN_318;
  assign _GEN_320 = 9'h140 == index ? 64'h0 : _GEN_319;
  assign _GEN_321 = 9'h141 == index ? 64'h0 : _GEN_320;
  assign _GEN_322 = 9'h142 == index ? 64'h0 : _GEN_321;
  assign _GEN_323 = 9'h143 == index ? 64'h0 : _GEN_322;
  assign _GEN_324 = 9'h144 == index ? 64'h0 : _GEN_323;
  assign _GEN_325 = 9'h145 == index ? 64'h0 : _GEN_324;
  assign _GEN_326 = 9'h146 == index ? 64'h0 : _GEN_325;
  assign _GEN_327 = 9'h147 == index ? 64'h0 : _GEN_326;
  assign _GEN_328 = 9'h148 == index ? 64'h0 : _GEN_327;
  assign _GEN_329 = 9'h149 == index ? 64'h0 : _GEN_328;
  assign _GEN_330 = 9'h14a == index ? 64'h0 : _GEN_329;
  assign _GEN_331 = 9'h14b == index ? 64'h0 : _GEN_330;
  assign _GEN_332 = 9'h14c == index ? 64'h0 : _GEN_331;
  assign _GEN_333 = 9'h14d == index ? 64'h0 : _GEN_332;
  assign _GEN_334 = 9'h14e == index ? 64'h0 : _GEN_333;
  assign _GEN_335 = 9'h14f == index ? 64'h0 : _GEN_334;
  assign _GEN_336 = 9'h150 == index ? 64'h0 : _GEN_335;
  assign _GEN_337 = 9'h151 == index ? 64'h0 : _GEN_336;
  assign _GEN_338 = 9'h152 == index ? 64'h0 : _GEN_337;
  assign _GEN_339 = 9'h153 == index ? 64'h0 : _GEN_338;
  assign _GEN_340 = 9'h154 == index ? 64'h0 : _GEN_339;
  assign _GEN_341 = 9'h155 == index ? 64'h0 : _GEN_340;
  assign _GEN_342 = 9'h156 == index ? 64'h0 : _GEN_341;
  assign _GEN_343 = 9'h157 == index ? 64'h0 : _GEN_342;
  assign _GEN_344 = 9'h158 == index ? 64'h0 : _GEN_343;
  assign _GEN_345 = 9'h159 == index ? 64'h0 : _GEN_344;
  assign _GEN_346 = 9'h15a == index ? 64'h0 : _GEN_345;
  assign _GEN_347 = 9'h15b == index ? 64'h0 : _GEN_346;
  assign _GEN_348 = 9'h15c == index ? 64'h0 : _GEN_347;
  assign _GEN_349 = 9'h15d == index ? 64'h0 : _GEN_348;
  assign _GEN_350 = 9'h15e == index ? 64'h0 : _GEN_349;
  assign _GEN_351 = 9'h15f == index ? 64'h0 : _GEN_350;
  assign _GEN_352 = 9'h160 == index ? 64'h0 : _GEN_351;
  assign _GEN_353 = 9'h161 == index ? 64'h0 : _GEN_352;
  assign _GEN_354 = 9'h162 == index ? 64'h0 : _GEN_353;
  assign _GEN_355 = 9'h163 == index ? 64'h0 : _GEN_354;
  assign _GEN_356 = 9'h164 == index ? 64'h0 : _GEN_355;
  assign _GEN_357 = 9'h165 == index ? 64'h0 : _GEN_356;
  assign _GEN_358 = 9'h166 == index ? 64'h0 : _GEN_357;
  assign _GEN_359 = 9'h167 == index ? 64'h0 : _GEN_358;
  assign _GEN_360 = 9'h168 == index ? 64'h0 : _GEN_359;
  assign _GEN_361 = 9'h169 == index ? 64'h0 : _GEN_360;
  assign _GEN_362 = 9'h16a == index ? 64'h0 : _GEN_361;
  assign _GEN_363 = 9'h16b == index ? 64'h0 : _GEN_362;
  assign _GEN_364 = 9'h16c == index ? 64'h0 : _GEN_363;
  assign _GEN_365 = 9'h16d == index ? 64'h0 : _GEN_364;
  assign _GEN_366 = 9'h16e == index ? 64'h0 : _GEN_365;
  assign _GEN_367 = 9'h16f == index ? 64'h0 : _GEN_366;
  assign _GEN_368 = 9'h170 == index ? 64'h0 : _GEN_367;
  assign _GEN_369 = 9'h171 == index ? 64'h0 : _GEN_368;
  assign _GEN_370 = 9'h172 == index ? 64'h0 : _GEN_369;
  assign _GEN_371 = 9'h173 == index ? 64'h0 : _GEN_370;
  assign _GEN_372 = 9'h174 == index ? 64'h0 : _GEN_371;
  assign _GEN_373 = 9'h175 == index ? 64'h0 : _GEN_372;
  assign _GEN_374 = 9'h176 == index ? 64'h0 : _GEN_373;
  assign _GEN_375 = 9'h177 == index ? 64'h0 : _GEN_374;
  assign _GEN_376 = 9'h178 == index ? 64'h0 : _GEN_375;
  assign _GEN_377 = 9'h179 == index ? 64'h0 : _GEN_376;
  assign _GEN_378 = 9'h17a == index ? 64'h0 : _GEN_377;
  assign _GEN_379 = 9'h17b == index ? 64'h0 : _GEN_378;
  assign _GEN_380 = 9'h17c == index ? 64'h0 : _GEN_379;
  assign _GEN_381 = 9'h17d == index ? 64'h0 : _GEN_380;
  assign _GEN_382 = 9'h17e == index ? 64'h0 : _GEN_381;
  assign _GEN_383 = 9'h17f == index ? 64'h0 : _GEN_382;
  assign _GEN_384 = 9'h180 == index ? 64'h0 : _GEN_383;
  assign _GEN_385 = 9'h181 == index ? 64'h0 : _GEN_384;
  assign _GEN_386 = 9'h182 == index ? 64'h0 : _GEN_385;
  assign _GEN_387 = 9'h183 == index ? 64'h0 : _GEN_386;
  assign _GEN_388 = 9'h184 == index ? 64'h0 : _GEN_387;
  assign _GEN_389 = 9'h185 == index ? 64'h0 : _GEN_388;
  assign _GEN_390 = 9'h186 == index ? 64'h0 : _GEN_389;
  assign _GEN_391 = 9'h187 == index ? 64'h0 : _GEN_390;
  assign _GEN_392 = 9'h188 == index ? 64'h0 : _GEN_391;
  assign _GEN_393 = 9'h189 == index ? 64'h0 : _GEN_392;
  assign _GEN_394 = 9'h18a == index ? 64'h0 : _GEN_393;
  assign _GEN_395 = 9'h18b == index ? 64'h0 : _GEN_394;
  assign _GEN_396 = 9'h18c == index ? 64'h0 : _GEN_395;
  assign _GEN_397 = 9'h18d == index ? 64'h0 : _GEN_396;
  assign _GEN_398 = 9'h18e == index ? 64'h0 : _GEN_397;
  assign _GEN_399 = 9'h18f == index ? 64'h0 : _GEN_398;
  assign _GEN_400 = 9'h190 == index ? 64'h0 : _GEN_399;
  assign _GEN_401 = 9'h191 == index ? 64'h0 : _GEN_400;
  assign _GEN_402 = 9'h192 == index ? 64'h0 : _GEN_401;
  assign _GEN_403 = 9'h193 == index ? 64'h0 : _GEN_402;
  assign _GEN_404 = 9'h194 == index ? 64'h0 : _GEN_403;
  assign _GEN_405 = 9'h195 == index ? 64'h0 : _GEN_404;
  assign _GEN_406 = 9'h196 == index ? 64'h0 : _GEN_405;
  assign _GEN_407 = 9'h197 == index ? 64'h0 : _GEN_406;
  assign _GEN_408 = 9'h198 == index ? 64'h0 : _GEN_407;
  assign _GEN_409 = 9'h199 == index ? 64'h0 : _GEN_408;
  assign _GEN_410 = 9'h19a == index ? 64'h0 : _GEN_409;
  assign _GEN_411 = 9'h19b == index ? 64'h0 : _GEN_410;
  assign _GEN_412 = 9'h19c == index ? 64'h0 : _GEN_411;
  assign _GEN_413 = 9'h19d == index ? 64'h0 : _GEN_412;
  assign _GEN_414 = 9'h19e == index ? 64'h0 : _GEN_413;
  assign _GEN_415 = 9'h19f == index ? 64'h0 : _GEN_414;
  assign _GEN_416 = 9'h1a0 == index ? 64'h0 : _GEN_415;
  assign _GEN_417 = 9'h1a1 == index ? 64'h0 : _GEN_416;
  assign _GEN_418 = 9'h1a2 == index ? 64'h0 : _GEN_417;
  assign _GEN_419 = 9'h1a3 == index ? 64'h0 : _GEN_418;
  assign _GEN_420 = 9'h1a4 == index ? 64'h0 : _GEN_419;
  assign _GEN_421 = 9'h1a5 == index ? 64'h0 : _GEN_420;
  assign _GEN_422 = 9'h1a6 == index ? 64'h0 : _GEN_421;
  assign _GEN_423 = 9'h1a7 == index ? 64'h0 : _GEN_422;
  assign _GEN_424 = 9'h1a8 == index ? 64'h0 : _GEN_423;
  assign _GEN_425 = 9'h1a9 == index ? 64'h0 : _GEN_424;
  assign _GEN_426 = 9'h1aa == index ? 64'h0 : _GEN_425;
  assign _GEN_427 = 9'h1ab == index ? 64'h0 : _GEN_426;
  assign _GEN_428 = 9'h1ac == index ? 64'h0 : _GEN_427;
  assign _GEN_429 = 9'h1ad == index ? 64'h0 : _GEN_428;
  assign _GEN_430 = 9'h1ae == index ? 64'h0 : _GEN_429;
  assign _GEN_431 = 9'h1af == index ? 64'h0 : _GEN_430;
  assign _GEN_432 = 9'h1b0 == index ? 64'h0 : _GEN_431;
  assign _GEN_433 = 9'h1b1 == index ? 64'h0 : _GEN_432;
  assign _GEN_434 = 9'h1b2 == index ? 64'h0 : _GEN_433;
  assign _GEN_435 = 9'h1b3 == index ? 64'h0 : _GEN_434;
  assign _GEN_436 = 9'h1b4 == index ? 64'h0 : _GEN_435;
  assign _GEN_437 = 9'h1b5 == index ? 64'h0 : _GEN_436;
  assign _GEN_438 = 9'h1b6 == index ? 64'h0 : _GEN_437;
  assign _GEN_439 = 9'h1b7 == index ? 64'h0 : _GEN_438;
  assign _GEN_440 = 9'h1b8 == index ? 64'h0 : _GEN_439;
  assign _GEN_441 = 9'h1b9 == index ? 64'h0 : _GEN_440;
  assign _GEN_442 = 9'h1ba == index ? 64'h0 : _GEN_441;
  assign _GEN_443 = 9'h1bb == index ? 64'h0 : _GEN_442;
  assign _GEN_444 = 9'h1bc == index ? 64'h0 : _GEN_443;
  assign _GEN_445 = 9'h1bd == index ? 64'h0 : _GEN_444;
  assign _GEN_446 = 9'h1be == index ? 64'h0 : _GEN_445;
  assign _GEN_447 = 9'h1bf == index ? 64'h0 : _GEN_446;
  assign _GEN_448 = 9'h1c0 == index ? 64'h0 : _GEN_447;
  assign _GEN_449 = 9'h1c1 == index ? 64'h0 : _GEN_448;
  assign _GEN_450 = 9'h1c2 == index ? 64'h0 : _GEN_449;
  assign _GEN_451 = 9'h1c3 == index ? 64'h0 : _GEN_450;
  assign _GEN_452 = 9'h1c4 == index ? 64'h0 : _GEN_451;
  assign _GEN_453 = 9'h1c5 == index ? 64'h0 : _GEN_452;
  assign _GEN_454 = 9'h1c6 == index ? 64'h0 : _GEN_453;
  assign _GEN_455 = 9'h1c7 == index ? 64'h0 : _GEN_454;
  assign _GEN_456 = 9'h1c8 == index ? 64'h0 : _GEN_455;
  assign _GEN_457 = 9'h1c9 == index ? 64'h0 : _GEN_456;
  assign _GEN_458 = 9'h1ca == index ? 64'h0 : _GEN_457;
  assign _GEN_459 = 9'h1cb == index ? 64'h0 : _GEN_458;
  assign _GEN_460 = 9'h1cc == index ? 64'h0 : _GEN_459;
  assign _GEN_461 = 9'h1cd == index ? 64'h0 : _GEN_460;
  assign _GEN_462 = 9'h1ce == index ? 64'h0 : _GEN_461;
  assign _GEN_463 = 9'h1cf == index ? 64'h0 : _GEN_462;
  assign _GEN_464 = 9'h1d0 == index ? 64'h0 : _GEN_463;
  assign _GEN_465 = 9'h1d1 == index ? 64'h0 : _GEN_464;
  assign _GEN_466 = 9'h1d2 == index ? 64'h0 : _GEN_465;
  assign _GEN_467 = 9'h1d3 == index ? 64'h0 : _GEN_466;
  assign _GEN_468 = 9'h1d4 == index ? 64'h0 : _GEN_467;
  assign _GEN_469 = 9'h1d5 == index ? 64'h0 : _GEN_468;
  assign _GEN_470 = 9'h1d6 == index ? 64'h0 : _GEN_469;
  assign _GEN_471 = 9'h1d7 == index ? 64'h0 : _GEN_470;
  assign _GEN_472 = 9'h1d8 == index ? 64'h0 : _GEN_471;
  assign _GEN_473 = 9'h1d9 == index ? 64'h0 : _GEN_472;
  assign _GEN_474 = 9'h1da == index ? 64'h0 : _GEN_473;
  assign _GEN_475 = 9'h1db == index ? 64'h0 : _GEN_474;
  assign _GEN_476 = 9'h1dc == index ? 64'h0 : _GEN_475;
  assign _GEN_477 = 9'h1dd == index ? 64'h0 : _GEN_476;
  assign _GEN_478 = 9'h1de == index ? 64'h0 : _GEN_477;
  assign _GEN_479 = 9'h1df == index ? 64'h0 : _GEN_478;
  assign _GEN_480 = 9'h1e0 == index ? 64'h0 : _GEN_479;
  assign _GEN_481 = 9'h1e1 == index ? 64'h0 : _GEN_480;
  assign _GEN_482 = 9'h1e2 == index ? 64'h0 : _GEN_481;
  assign _GEN_483 = 9'h1e3 == index ? 64'h0 : _GEN_482;
  assign _GEN_484 = 9'h1e4 == index ? 64'h0 : _GEN_483;
  assign _GEN_485 = 9'h1e5 == index ? 64'h0 : _GEN_484;
  assign _GEN_486 = 9'h1e6 == index ? 64'h0 : _GEN_485;
  assign _GEN_487 = 9'h1e7 == index ? 64'h0 : _GEN_486;
  assign _GEN_488 = 9'h1e8 == index ? 64'h0 : _GEN_487;
  assign _GEN_489 = 9'h1e9 == index ? 64'h0 : _GEN_488;
  assign _GEN_490 = 9'h1ea == index ? 64'h0 : _GEN_489;
  assign _GEN_491 = 9'h1eb == index ? 64'h0 : _GEN_490;
  assign _GEN_492 = 9'h1ec == index ? 64'h0 : _GEN_491;
  assign _GEN_493 = 9'h1ed == index ? 64'h0 : _GEN_492;
  assign _GEN_494 = 9'h1ee == index ? 64'h0 : _GEN_493;
  assign _GEN_495 = 9'h1ef == index ? 64'h0 : _GEN_494;
  assign _GEN_496 = 9'h1f0 == index ? 64'h0 : _GEN_495;
  assign _GEN_497 = 9'h1f1 == index ? 64'h0 : _GEN_496;
  assign _GEN_498 = 9'h1f2 == index ? 64'h0 : _GEN_497;
  assign _GEN_499 = 9'h1f3 == index ? 64'h0 : _GEN_498;
  assign _GEN_500 = 9'h1f4 == index ? 64'h0 : _GEN_499;
  assign _GEN_501 = 9'h1f5 == index ? 64'h0 : _GEN_500;
  assign _GEN_502 = 9'h1f6 == index ? 64'h0 : _GEN_501;
  assign _GEN_503 = 9'h1f7 == index ? 64'h0 : _GEN_502;
  assign _GEN_504 = 9'h1f8 == index ? 64'h0 : _GEN_503;
  assign _GEN_505 = 9'h1f9 == index ? 64'h0 : _GEN_504;
  assign _GEN_506 = 9'h1fa == index ? 64'h0 : _GEN_505;
  assign _GEN_507 = 9'h1fb == index ? 64'h0 : _GEN_506;
  assign _GEN_508 = 9'h1fc == index ? 64'h0 : _GEN_507;
  assign _GEN_509 = 9'h1fd == index ? 64'h0 : _GEN_508;
  assign _GEN_510 = 9'h1fe == index ? 64'h0 : _GEN_509;
  assign _GEN_511 = 9'h1ff == index ? 64'h0 : _GEN_510;
  assign _T_1148 = _T_1145 ? 64'h0 : _GEN_0;
  assign auto_in_a_ready = in_a_ready;
  assign auto_in_d_valid = in_d_valid;
  assign auto_in_d_bits_size = in_d_bits_size;
  assign auto_in_d_bits_source = in_d_bits_source;
  assign auto_in_d_bits_data = in_d_bits_data;
  assign in_a_ready = in_d_ready;
  assign in_a_valid = auto_in_a_valid;
  assign in_a_bits_size = auto_in_a_bits_size;
  assign in_a_bits_source = auto_in_a_bits_source;
  assign in_a_bits_address = auto_in_a_bits_address;
  assign in_d_ready = auto_in_d_ready;
  assign in_d_valid = in_a_valid;
  assign in_d_bits_size = _T_1151_size;
  assign in_d_bits_source = _T_1151_source;
  assign in_d_bits_data = _T_1151_data;
  assign _GEN_0 = _GEN_511;
  assign _T_1151_size = in_a_bits_size;
  assign _T_1151_source = in_a_bits_source;
  assign _T_1151_data = _T_1148;
endmodule
module Queue_113(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_42_data;
  wire  ram_opcode__T_42_addr;
  wire [2:0] ram_opcode__T_33_data;
  wire  ram_opcode__T_33_addr;
  wire  ram_opcode__T_33_mask;
  wire  ram_opcode__T_33_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [3:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_42_data;
  wire  ram_source__T_42_addr;
  wire [4:0] ram_source__T_33_data;
  wire  ram_source__T_33_addr;
  wire  ram_source__T_33_mask;
  wire  ram_source__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_10;
  wire  _T_38;
  assign ram_opcode__T_42_addr = 1'h0;
  assign ram_opcode__T_42_data = ram_opcode[ram_opcode__T_42_addr];
  assign ram_opcode__T_33_data = io_enq_bits_opcode;
  assign ram_opcode__T_33_addr = 1'h0;
  assign ram_opcode__T_33_mask = do_enq;
  assign ram_opcode__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_source__T_42_addr = 1'h0;
  assign ram_source__T_42_data = ram_source[ram_source__T_42_addr];
  assign ram_source__T_33_data = io_enq_bits_source;
  assign ram_source__T_33_addr = 1'h0;
  assign ram_source__T_33_mask = do_enq;
  assign ram_source__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_10 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign io_enq_ready = empty;
  assign io_deq_valid = _T_38;
  assign io_deq_bits_opcode = ram_opcode__T_42_data;
  assign io_deq_bits_size = ram_size__T_42_data;
  assign io_deq_bits_source = ram_source__T_42_data;
  assign do_enq = _T_28;
  assign do_deq = _T_30;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_33_en & ram_opcode__T_33_mask) begin
      ram_opcode[ram_opcode__T_33_addr] <= ram_opcode__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_source__T_33_en & ram_source__T_33_mask) begin
      ram_source[ram_source__T_33_addr] <= ram_source__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_114(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [2:0] io_enq_bits_param,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_42_data;
  wire  ram_opcode__T_42_addr;
  wire [2:0] ram_opcode__T_33_data;
  wire  ram_opcode__T_33_addr;
  wire  ram_opcode__T_33_mask;
  wire  ram_opcode__T_33_en;
  reg [2:0] ram_param [0:0];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_42_data;
  wire  ram_param__T_42_addr;
  wire [2:0] ram_param__T_33_data;
  wire  ram_param__T_33_addr;
  wire  ram_param__T_33_mask;
  wire  ram_param__T_33_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [3:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_42_data;
  wire  ram_source__T_42_addr;
  wire [4:0] ram_source__T_33_data;
  wire  ram_source__T_33_addr;
  wire  ram_source__T_33_mask;
  wire  ram_source__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_4;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_10;
  wire  _T_38;
  assign ram_opcode__T_42_addr = 1'h0;
  assign ram_opcode__T_42_data = ram_opcode[ram_opcode__T_42_addr];
  assign ram_opcode__T_33_data = io_enq_bits_opcode;
  assign ram_opcode__T_33_addr = 1'h0;
  assign ram_opcode__T_33_mask = do_enq;
  assign ram_opcode__T_33_en = do_enq;
  assign ram_param__T_42_addr = 1'h0;
  assign ram_param__T_42_data = ram_param[ram_param__T_42_addr];
  assign ram_param__T_33_data = io_enq_bits_param;
  assign ram_param__T_33_addr = 1'h0;
  assign ram_param__T_33_mask = do_enq;
  assign ram_param__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_source__T_42_addr = 1'h0;
  assign ram_source__T_42_data = ram_source[ram_source__T_42_addr];
  assign ram_source__T_33_data = io_enq_bits_source;
  assign ram_source__T_33_addr = 1'h0;
  assign ram_source__T_33_mask = do_enq;
  assign ram_source__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_10 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign io_enq_ready = empty;
  assign io_deq_valid = _T_38;
  assign io_deq_bits_opcode = ram_opcode__T_42_data;
  assign io_deq_bits_param = ram_param__T_42_data;
  assign io_deq_bits_size = ram_size__T_42_data;
  assign io_deq_bits_source = ram_source__T_42_data;
  assign do_enq = _T_28;
  assign do_deq = _T_30;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  maybe_full = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_33_en & ram_opcode__T_33_mask) begin
      ram_opcode[ram_opcode__T_33_addr] <= ram_opcode__T_33_data;
    end
    if(ram_param__T_33_en & ram_param__T_33_mask) begin
      ram_param[ram_param__T_33_addr] <= ram_param__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_source__T_33_en & ram_source__T_33_mask) begin
      ram_source[ram_source__T_33_addr] <= ram_source__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TLError_error(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [4:0]  auto_in_a_bits_source,
  output        auto_in_c_ready,
  input         auto_in_c_valid,
  input  [2:0]  auto_in_c_bits_opcode,
  input  [2:0]  auto_in_c_bits_param,
  input  [3:0]  auto_in_c_bits_size,
  input  [4:0]  auto_in_c_bits_source,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_param,
  output [3:0]  auto_in_d_bits_size,
  output [4:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_sink,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_error
);
  wire  in_a_ready;
  wire  in_a_valid;
  wire [2:0] in_a_bits_opcode;
  wire [3:0] in_a_bits_size;
  wire [4:0] in_a_bits_source;
  wire  in_c_ready;
  wire  in_c_valid;
  wire [2:0] in_c_bits_opcode;
  wire [2:0] in_c_bits_param;
  wire [3:0] in_c_bits_size;
  wire [4:0] in_c_bits_source;
  wire  in_d_ready;
  wire  in_d_valid;
  wire [2:0] in_d_bits_opcode;
  wire [1:0] in_d_bits_param;
  wire [3:0] in_d_bits_size;
  wire [4:0] in_d_bits_source;
  wire  in_d_bits_sink;
  wire [63:0] in_d_bits_data;
  wire  in_d_bits_error;
  wire  a_clock;
  wire  a_reset;
  wire  a_io_enq_ready;
  wire  a_io_enq_valid;
  wire [2:0] a_io_enq_bits_opcode;
  wire [3:0] a_io_enq_bits_size;
  wire [4:0] a_io_enq_bits_source;
  wire  a_io_deq_ready;
  wire  a_io_deq_valid;
  wire [2:0] a_io_deq_bits_opcode;
  wire [3:0] a_io_deq_bits_size;
  wire [4:0] a_io_deq_bits_source;
  wire  c_clock;
  wire  c_reset;
  wire  c_io_enq_ready;
  wire  c_io_enq_valid;
  wire [2:0] c_io_enq_bits_opcode;
  wire [2:0] c_io_enq_bits_param;
  wire [3:0] c_io_enq_bits_size;
  wire [4:0] c_io_enq_bits_source;
  wire  c_io_deq_ready;
  wire  c_io_deq_valid;
  wire [2:0] c_io_deq_bits_opcode;
  wire [2:0] c_io_deq_bits_param;
  wire [3:0] c_io_deq_bits_size;
  wire [4:0] c_io_deq_bits_source;
  wire  da_ready;
  wire  da_valid;
  wire [2:0] da_bits_opcode;
  wire [3:0] da_bits_size;
  wire [4:0] da_bits_source;
  wire  dc_ready;
  wire  dc_valid;
  wire [1:0] dc_bits_param;
  wire [3:0] dc_bits_size;
  wire [4:0] dc_bits_source;
  wire  _T_122;
  wire [26:0] _T_125;
  wire [11:0] _T_126;
  wire [11:0] _T_127;
  wire [8:0] _T_128;
  wire  _T_129;
  wire  _T_131;
  wire [8:0] _T_133;
  reg [8:0] _T_136;
  reg [31:0] _RAND_0;
  wire [9:0] _T_138;
  wire [9:0] _T_139;
  wire [8:0] _T_140;
  wire  _T_142;
  wire  _T_144;
  wire  _T_146;
  wire  a_last;
  wire [8:0] _T_150;
  wire [8:0] _GEN_2;
  wire  _T_151;
  wire [26:0] _T_154;
  wire [11:0] _T_155;
  wire [11:0] _T_156;
  wire [8:0] _T_157;
  wire  _T_158;
  wire [8:0] _T_160;
  reg [8:0] _T_163;
  reg [31:0] _RAND_1;
  wire [9:0] _T_165;
  wire [9:0] _T_166;
  wire [8:0] _T_167;
  wire  _T_169;
  wire  _T_171;
  wire  _T_173;
  wire  c_last;
  wire [8:0] _T_177;
  wire [8:0] _GEN_3;
  wire  _T_178;
  wire [26:0] _T_181;
  wire [11:0] _T_182;
  wire [11:0] _T_183;
  wire [8:0] _T_184;
  wire  _T_185;
  wire [8:0] _T_187;
  reg [8:0] _T_190;
  reg [31:0] _RAND_2;
  wire [9:0] _T_192;
  wire [9:0] _T_193;
  wire [8:0] _T_194;
  wire  _T_196;
  wire  _T_198;
  wire  _T_200;
  wire  da_last;
  wire [8:0] _T_204;
  wire [8:0] _GEN_4;
  wire  _T_232;
  wire  _T_234;
  wire  _T_235;
  wire  _T_236;
  wire [2:0] _GEN_0;
  wire [2:0] _GEN_7;
  wire [2:0] _GEN_8;
  wire [2:0] _GEN_9;
  wire [2:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire  _T_262;
  wire  _T_263;
  wire  _T_264;
  wire [1:0] _T_278;
  wire [1:0] _GEN_1;
  wire [1:0] _GEN_12;
  wire [1:0] _GEN_13;
  reg [8:0] _T_302;
  reg [31:0] _RAND_3;
  wire  _T_304;
  wire  _T_305;
  wire [1:0] _T_306;
  wire [2:0] _GEN_14;
  wire [2:0] _T_307;
  wire [1:0] _T_308;
  wire [1:0] _T_309;
  wire [2:0] _GEN_15;
  wire [2:0] _T_311;
  wire [1:0] _T_312;
  wire [1:0] _T_313;
  wire  _T_314;
  wire  _T_315;
  wire  _T_318_0;
  wire  _T_318_1;
  wire  _T_323;
  wire  _T_324;
  wire  _T_327_0;
  wire  _T_327_1;
  wire  _T_334;
  wire  _T_338;
  wire  _T_343;
  wire  _T_344;
  wire  _T_347;
  wire  _T_349;
  wire  _T_350;
  wire  _T_352;
  wire  _T_354;
  wire  _T_356;
  wire  _T_358;
  wire [8:0] _T_362;
  wire  _T_364;
  wire [8:0] _GEN_16;
  wire [9:0] _T_365;
  wire [9:0] _T_366;
  wire [8:0] _T_367;
  wire [8:0] _T_368;
  reg  _T_386_0;
  reg [31:0] _RAND_4;
  reg  _T_386_1;
  reg [31:0] _RAND_5;
  wire  _T_397_0;
  wire  _T_397_1;
  wire  _T_405_0;
  wire  _T_405_1;
  wire  _T_413;
  wire  _T_414;
  wire  _T_418;
  wire  _T_420;
  wire  _T_421;
  wire  _T_423;
  wire  _T_424;
  wire [8:0] _T_428;
  wire [4:0] _T_429;
  wire [13:0] _T_430;
  wire [79:0] _T_431;
  wire [79:0] _T_433;
  wire [8:0] _T_436;
  wire [4:0] _T_437;
  wire [13:0] _T_438;
  wire [79:0] _T_439;
  wire [79:0] _T_441;
  wire [79:0] _T_442;
  wire [2:0] _T_444_opcode;
  wire [1:0] _T_444_param;
  wire [3:0] _T_444_size;
  wire [4:0] _T_444_source;
  wire  _T_444_sink;
  wire [63:0] _T_444_data;
  wire  _T_444_error;
  wire [79:0] _T_446;
  wire  _T_447;
  wire [63:0] _T_448;
  wire  _T_449;
  wire [4:0] _T_450;
  wire [3:0] _T_451;
  wire [1:0] _T_452;
  wire [2:0] _T_453;
  Queue_113 a (
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  Queue_114 c (
    .clock(c_clock),
    .reset(c_reset),
    .io_enq_ready(c_io_enq_ready),
    .io_enq_valid(c_io_enq_valid),
    .io_enq_bits_opcode(c_io_enq_bits_opcode),
    .io_enq_bits_param(c_io_enq_bits_param),
    .io_enq_bits_size(c_io_enq_bits_size),
    .io_enq_bits_source(c_io_enq_bits_source),
    .io_deq_ready(c_io_deq_ready),
    .io_deq_valid(c_io_deq_valid),
    .io_deq_bits_opcode(c_io_deq_bits_opcode),
    .io_deq_bits_param(c_io_deq_bits_param),
    .io_deq_bits_size(c_io_deq_bits_size),
    .io_deq_bits_source(c_io_deq_bits_source)
  );
  assign _T_122 = a_io_deq_ready & a_io_deq_valid;
  assign _T_125 = 27'hfff << a_io_deq_bits_size;
  assign _T_126 = _T_125[11:0];
  assign _T_127 = ~ _T_126;
  assign _T_128 = _T_127[11:3];
  assign _T_129 = a_io_deq_bits_opcode[2];
  assign _T_131 = _T_129 == 1'h0;
  assign _T_133 = _T_131 ? _T_128 : 9'h0;
  assign _T_138 = _T_136 - 9'h1;
  assign _T_139 = $unsigned(_T_138);
  assign _T_140 = _T_139[8:0];
  assign _T_142 = _T_136 == 9'h0;
  assign _T_144 = _T_136 == 9'h1;
  assign _T_146 = _T_133 == 9'h0;
  assign a_last = _T_144 | _T_146;
  assign _T_150 = _T_142 ? _T_133 : _T_140;
  assign _GEN_2 = _T_122 ? _T_150 : _T_136;
  assign _T_151 = c_io_deq_ready & c_io_deq_valid;
  assign _T_154 = 27'hfff << c_io_deq_bits_size;
  assign _T_155 = _T_154[11:0];
  assign _T_156 = ~ _T_155;
  assign _T_157 = _T_156[11:3];
  assign _T_158 = c_io_deq_bits_opcode[0];
  assign _T_160 = _T_158 ? _T_157 : 9'h0;
  assign _T_165 = _T_163 - 9'h1;
  assign _T_166 = $unsigned(_T_165);
  assign _T_167 = _T_166[8:0];
  assign _T_169 = _T_163 == 9'h0;
  assign _T_171 = _T_163 == 9'h1;
  assign _T_173 = _T_160 == 9'h0;
  assign c_last = _T_171 | _T_173;
  assign _T_177 = _T_169 ? _T_160 : _T_167;
  assign _GEN_3 = _T_151 ? _T_177 : _T_163;
  assign _T_178 = da_ready & da_valid;
  assign _T_181 = 27'hfff << da_bits_size;
  assign _T_182 = _T_181[11:0];
  assign _T_183 = ~ _T_182;
  assign _T_184 = _T_183[11:3];
  assign _T_185 = da_bits_opcode[0];
  assign _T_187 = _T_185 ? _T_184 : 9'h0;
  assign _T_192 = _T_190 - 9'h1;
  assign _T_193 = $unsigned(_T_192);
  assign _T_194 = _T_193[8:0];
  assign _T_196 = _T_190 == 9'h0;
  assign _T_198 = _T_190 == 9'h1;
  assign _T_200 = _T_187 == 9'h0;
  assign da_last = _T_198 | _T_200;
  assign _T_204 = _T_196 ? _T_187 : _T_194;
  assign _GEN_4 = _T_178 ? _T_204 : _T_190;
  assign _T_232 = da_ready & da_last;
  assign _T_234 = a_last == 1'h0;
  assign _T_235 = _T_232 | _T_234;
  assign _T_236 = a_io_deq_valid & a_last;
  assign _GEN_7 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0;
  assign _GEN_8 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_7;
  assign _GEN_9 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_8;
  assign _GEN_10 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_9;
  assign _GEN_11 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_10;
  assign _T_262 = c_last == 1'h0;
  assign _T_263 = dc_ready | _T_262;
  assign _T_264 = c_io_deq_valid & c_last;
  assign _T_278 = c_io_deq_bits_param[1:0];
  assign _GEN_12 = 2'h1 == _T_278 ? 2'h2 : 2'h1;
  assign _GEN_13 = 2'h2 == _T_278 ? 2'h2 : _GEN_12;
  assign _T_304 = _T_302 == 9'h0;
  assign _T_305 = _T_304 & in_d_ready;
  assign _T_306 = {da_valid,dc_valid};
  assign _GEN_14 = {{1'd0}, _T_306};
  assign _T_307 = _GEN_14 << 1;
  assign _T_308 = _T_307[1:0];
  assign _T_309 = _T_306 | _T_308;
  assign _GEN_15 = {{1'd0}, _T_309};
  assign _T_311 = _GEN_15 << 1;
  assign _T_312 = _T_311[1:0];
  assign _T_313 = ~ _T_312;
  assign _T_314 = _T_313[0];
  assign _T_315 = _T_313[1];
  assign _T_323 = _T_318_0 & dc_valid;
  assign _T_324 = _T_318_1 & da_valid;
  assign _T_334 = _T_327_0 | _T_327_1;
  assign _T_338 = _T_327_0 == 1'h0;
  assign _T_343 = _T_327_1 == 1'h0;
  assign _T_344 = _T_338 | _T_343;
  assign _T_347 = _T_344 | reset;
  assign _T_349 = _T_347 == 1'h0;
  assign _T_350 = dc_valid | da_valid;
  assign _T_352 = _T_350 == 1'h0;
  assign _T_354 = _T_352 | _T_334;
  assign _T_356 = _T_354 | reset;
  assign _T_358 = _T_356 == 1'h0;
  assign _T_362 = _T_327_1 ? _T_187 : 9'h0;
  assign _T_364 = in_d_ready & in_d_valid;
  assign _GEN_16 = {{8'd0}, _T_364};
  assign _T_365 = _T_302 - _GEN_16;
  assign _T_366 = $unsigned(_T_365);
  assign _T_367 = _T_366[8:0];
  assign _T_368 = _T_305 ? _T_362 : _T_367;
  assign _T_397_0 = _T_304 ? _T_327_0 : _T_386_0;
  assign _T_397_1 = _T_304 ? _T_327_1 : _T_386_1;
  assign _T_405_0 = _T_304 ? _T_318_0 : _T_386_0;
  assign _T_405_1 = _T_304 ? _T_318_1 : _T_386_1;
  assign _T_413 = in_d_ready & _T_405_0;
  assign _T_414 = in_d_ready & _T_405_1;
  assign _T_418 = _T_386_0 ? dc_valid : 1'h0;
  assign _T_420 = _T_386_1 ? da_valid : 1'h0;
  assign _T_421 = _T_418 | _T_420;
  assign _T_424 = _T_304 ? _T_350 : _T_423;
  assign _T_428 = {dc_bits_size,dc_bits_source};
  assign _T_429 = {3'h6,dc_bits_param};
  assign _T_430 = {_T_429,_T_428};
  assign _T_431 = {_T_430,66'h1};
  assign _T_433 = _T_397_0 ? _T_431 : 80'h0;
  assign _T_436 = {da_bits_size,da_bits_source};
  assign _T_437 = {da_bits_opcode,2'h0};
  assign _T_438 = {_T_437,_T_436};
  assign _T_439 = {_T_438,66'h1};
  assign _T_441 = _T_397_1 ? _T_439 : 80'h0;
  assign _T_442 = _T_433 | _T_441;
  assign _T_447 = _T_446[0];
  assign _T_448 = _T_446[64:1];
  assign _T_449 = _T_446[65];
  assign _T_450 = _T_446[70:66];
  assign _T_451 = _T_446[74:71];
  assign _T_452 = _T_446[76:75];
  assign _T_453 = _T_446[79:77];
  assign auto_in_a_ready = in_a_ready;
  assign auto_in_c_ready = in_c_ready;
  assign auto_in_d_valid = in_d_valid;
  assign auto_in_d_bits_opcode = in_d_bits_opcode;
  assign auto_in_d_bits_param = in_d_bits_param;
  assign auto_in_d_bits_size = in_d_bits_size;
  assign auto_in_d_bits_source = in_d_bits_source;
  assign auto_in_d_bits_sink = in_d_bits_sink;
  assign auto_in_d_bits_data = in_d_bits_data;
  assign auto_in_d_bits_error = in_d_bits_error;
  assign in_a_ready = a_io_enq_ready;
  assign in_a_valid = auto_in_a_valid;
  assign in_a_bits_opcode = auto_in_a_bits_opcode;
  assign in_a_bits_size = auto_in_a_bits_size;
  assign in_a_bits_source = auto_in_a_bits_source;
  assign in_c_ready = c_io_enq_ready;
  assign in_c_valid = auto_in_c_valid;
  assign in_c_bits_opcode = auto_in_c_bits_opcode;
  assign in_c_bits_param = auto_in_c_bits_param;
  assign in_c_bits_size = auto_in_c_bits_size;
  assign in_c_bits_source = auto_in_c_bits_source;
  assign in_d_ready = auto_in_d_ready;
  assign in_d_valid = _T_424;
  assign in_d_bits_opcode = _T_444_opcode;
  assign in_d_bits_param = _T_444_param;
  assign in_d_bits_size = _T_444_size;
  assign in_d_bits_source = _T_444_source;
  assign in_d_bits_sink = _T_444_sink;
  assign in_d_bits_data = _T_444_data;
  assign in_d_bits_error = _T_444_error;
  assign a_io_enq_valid = in_a_valid;
  assign a_io_enq_bits_opcode = in_a_bits_opcode;
  assign a_io_enq_bits_size = in_a_bits_size;
  assign a_io_enq_bits_source = in_a_bits_source;
  assign a_io_deq_ready = _T_235;
  assign a_clock = clock;
  assign a_reset = reset;
  assign c_io_enq_valid = in_c_valid;
  assign c_io_enq_bits_opcode = in_c_bits_opcode;
  assign c_io_enq_bits_param = in_c_bits_param;
  assign c_io_enq_bits_size = in_c_bits_size;
  assign c_io_enq_bits_source = in_c_bits_source;
  assign c_io_deq_ready = _T_263;
  assign c_clock = clock;
  assign c_reset = reset;
  assign da_ready = _T_414;
  assign da_valid = _T_236;
  assign da_bits_opcode = _GEN_0;
  assign da_bits_size = a_io_deq_bits_size;
  assign da_bits_source = a_io_deq_bits_source;
  assign dc_ready = _T_413;
  assign dc_valid = _T_264;
  assign dc_bits_param = _GEN_1;
  assign dc_bits_size = c_io_deq_bits_size;
  assign dc_bits_source = c_io_deq_bits_source;
  assign _GEN_0 = _GEN_11;
  assign _GEN_1 = _GEN_13;
  assign _T_318_0 = _T_314;
  assign _T_318_1 = _T_315;
  assign _T_327_0 = _T_323;
  assign _T_327_1 = _T_324;
  assign _T_423 = _T_421;
  assign _T_444_opcode = _T_453;
  assign _T_444_param = _T_452;
  assign _T_444_size = _T_451;
  assign _T_444_source = _T_450;
  assign _T_444_sink = _T_449;
  assign _T_444_data = _T_448;
  assign _T_444_error = _T_447;
  assign _T_446 = _T_442;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_136 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_163 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_190 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_302 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_386_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_386_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_136 <= 9'h0;
    end else begin
      if (_T_122) begin
        if (_T_142) begin
          if (_T_131) begin
            _T_136 <= _T_128;
          end else begin
            _T_136 <= 9'h0;
          end
        end else begin
          _T_136 <= _T_140;
        end
      end
    end
    if (reset) begin
      _T_163 <= 9'h0;
    end else begin
      if (_T_151) begin
        if (_T_169) begin
          if (_T_158) begin
            _T_163 <= _T_157;
          end else begin
            _T_163 <= 9'h0;
          end
        end else begin
          _T_163 <= _T_167;
        end
      end
    end
    if (reset) begin
      _T_190 <= 9'h0;
    end else begin
      if (_T_178) begin
        if (_T_196) begin
          if (_T_185) begin
            _T_190 <= _T_184;
          end else begin
            _T_190 <= 9'h0;
          end
        end else begin
          _T_190 <= _T_194;
        end
      end
    end
    if (reset) begin
      _T_302 <= 9'h0;
    end else begin
      if (_T_305) begin
        if (_T_327_1) begin
          if (_T_185) begin
            _T_302 <= _T_184;
          end else begin
            _T_302 <= 9'h0;
          end
        end else begin
          _T_302 <= 9'h0;
        end
      end else begin
        _T_302 <= _T_367;
      end
    end
    if (reset) begin
      _T_386_0 <= 1'h0;
    end else begin
      if (_T_304) begin
        _T_386_0 <= _T_327_0;
      end
    end
    if (reset) begin
      _T_386_1 <= 1'h0;
    end else begin
      if (_T_304) begin
        _T_386_1 <= _T_327_1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_349) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_349) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_358) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_358) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ExampleBoomSystem(
  input         clock,
  input         reset,
  output        debug_clockeddmi_dmi_req_ready,
  input         debug_clockeddmi_dmi_req_valid,
  input  [6:0]  debug_clockeddmi_dmi_req_bits_addr,
  input  [31:0] debug_clockeddmi_dmi_req_bits_data,
  input  [1:0]  debug_clockeddmi_dmi_req_bits_op,
  input         debug_clockeddmi_dmi_resp_ready,
  output        debug_clockeddmi_dmi_resp_valid,
  output [31:0] debug_clockeddmi_dmi_resp_bits_data,
  output [1:0]  debug_clockeddmi_dmi_resp_bits_resp,
  input         debug_clockeddmi_dmiClock,
  input         debug_clockeddmi_dmiReset,
  output        debug_ndreset,
  output        debug_dmactive,
  input  [1:0]  interrupts,
  input         mem_axi4_0_aw_ready,
  output        mem_axi4_0_aw_valid,
  output [3:0]  mem_axi4_0_aw_bits_id,
  output [31:0] mem_axi4_0_aw_bits_addr,
  output [7:0]  mem_axi4_0_aw_bits_len,
  output [2:0]  mem_axi4_0_aw_bits_size,
  output [1:0]  mem_axi4_0_aw_bits_burst,
  output        mem_axi4_0_aw_bits_lock,
  output [3:0]  mem_axi4_0_aw_bits_cache,
  output [2:0]  mem_axi4_0_aw_bits_prot,
  output [3:0]  mem_axi4_0_aw_bits_qos,
  input         mem_axi4_0_w_ready,
  output        mem_axi4_0_w_valid,
  output [63:0] mem_axi4_0_w_bits_data,
  output [7:0]  mem_axi4_0_w_bits_strb,
  output        mem_axi4_0_w_bits_last,
  output        mem_axi4_0_b_ready,
  input         mem_axi4_0_b_valid,
  input  [3:0]  mem_axi4_0_b_bits_id,
  input  [1:0]  mem_axi4_0_b_bits_resp,
  input         mem_axi4_0_ar_ready,
  output        mem_axi4_0_ar_valid,
  output [3:0]  mem_axi4_0_ar_bits_id,
  output [31:0] mem_axi4_0_ar_bits_addr,
  output [7:0]  mem_axi4_0_ar_bits_len,
  output [2:0]  mem_axi4_0_ar_bits_size,
  output [1:0]  mem_axi4_0_ar_bits_burst,
  output        mem_axi4_0_ar_bits_lock,
  output [3:0]  mem_axi4_0_ar_bits_cache,
  output [2:0]  mem_axi4_0_ar_bits_prot,
  output [3:0]  mem_axi4_0_ar_bits_qos,
  output        mem_axi4_0_r_ready,
  input         mem_axi4_0_r_valid,
  input  [3:0]  mem_axi4_0_r_bits_id,
  input  [63:0] mem_axi4_0_r_bits_data,
  input  [1:0]  mem_axi4_0_r_bits_resp,
  input         mem_axi4_0_r_bits_last,
  input         mmio_axi4_0_aw_ready,
  output        mmio_axi4_0_aw_valid,
  output [3:0]  mmio_axi4_0_aw_bits_id,
  output [30:0] mmio_axi4_0_aw_bits_addr,
  output [7:0]  mmio_axi4_0_aw_bits_len,
  output [2:0]  mmio_axi4_0_aw_bits_size,
  output [1:0]  mmio_axi4_0_aw_bits_burst,
  output        mmio_axi4_0_aw_bits_lock,
  output [3:0]  mmio_axi4_0_aw_bits_cache,
  output [2:0]  mmio_axi4_0_aw_bits_prot,
  output [3:0]  mmio_axi4_0_aw_bits_qos,
  input         mmio_axi4_0_w_ready,
  output        mmio_axi4_0_w_valid,
  output [63:0] mmio_axi4_0_w_bits_data,
  output [7:0]  mmio_axi4_0_w_bits_strb,
  output        mmio_axi4_0_w_bits_last,
  output        mmio_axi4_0_b_ready,
  input         mmio_axi4_0_b_valid,
  input  [3:0]  mmio_axi4_0_b_bits_id,
  input  [1:0]  mmio_axi4_0_b_bits_resp,
  input         mmio_axi4_0_ar_ready,
  output        mmio_axi4_0_ar_valid,
  output [3:0]  mmio_axi4_0_ar_bits_id,
  output [30:0] mmio_axi4_0_ar_bits_addr,
  output [7:0]  mmio_axi4_0_ar_bits_len,
  output [2:0]  mmio_axi4_0_ar_bits_size,
  output [1:0]  mmio_axi4_0_ar_bits_burst,
  output        mmio_axi4_0_ar_bits_lock,
  output [3:0]  mmio_axi4_0_ar_bits_cache,
  output [2:0]  mmio_axi4_0_ar_bits_prot,
  output [3:0]  mmio_axi4_0_ar_bits_qos,
  output        mmio_axi4_0_r_ready,
  input         mmio_axi4_0_r_valid,
  input  [3:0]  mmio_axi4_0_r_bits_id,
  input  [63:0] mmio_axi4_0_r_bits_data,
  input  [1:0]  mmio_axi4_0_r_bits_resp,
  input         mmio_axi4_0_r_bits_last,
  output        l2_frontend_bus_axi4_0_aw_ready,
  input         l2_frontend_bus_axi4_0_aw_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_aw_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_aw_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_aw_bits_burst,
  input         l2_frontend_bus_axi4_0_aw_bits_lock,
  input  [3:0]  l2_frontend_bus_axi4_0_aw_bits_cache,
  input  [2:0]  l2_frontend_bus_axi4_0_aw_bits_prot,
  input  [3:0]  l2_frontend_bus_axi4_0_aw_bits_qos,
  output        l2_frontend_bus_axi4_0_w_ready,
  input         l2_frontend_bus_axi4_0_w_valid,
  input  [63:0] l2_frontend_bus_axi4_0_w_bits_data,
  input  [7:0]  l2_frontend_bus_axi4_0_w_bits_strb,
  input         l2_frontend_bus_axi4_0_w_bits_last,
  input         l2_frontend_bus_axi4_0_b_ready,
  output        l2_frontend_bus_axi4_0_b_valid,
  output [7:0]  l2_frontend_bus_axi4_0_b_bits_id,
  output [1:0]  l2_frontend_bus_axi4_0_b_bits_resp,
  output        l2_frontend_bus_axi4_0_ar_ready,
  input         l2_frontend_bus_axi4_0_ar_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_ar_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_ar_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_ar_bits_burst,
  input         l2_frontend_bus_axi4_0_ar_bits_lock,
  input  [3:0]  l2_frontend_bus_axi4_0_ar_bits_cache,
  input  [2:0]  l2_frontend_bus_axi4_0_ar_bits_prot,
  input  [3:0]  l2_frontend_bus_axi4_0_ar_bits_qos,
  input         l2_frontend_bus_axi4_0_r_ready,
  output        l2_frontend_bus_axi4_0_r_valid,
  output [7:0]  l2_frontend_bus_axi4_0_r_bits_id,
  output [63:0] l2_frontend_bus_axi4_0_r_bits_data,
  output [1:0]  l2_frontend_bus_axi4_0_r_bits_resp,
  output        l2_frontend_bus_axi4_0_r_bits_last
);
  wire  IntXbar_auto_int_in_0;
  wire  IntXbar_auto_int_in_1;
  wire  IntXbar_auto_int_out_0;
  wire  IntXbar_auto_int_out_1;
  wire  sbus_clock;
  wire  sbus_reset;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_a_ready;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_a_valid;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_opcode;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_param;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_size;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_source;
  wire [31:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_address;
  wire [7:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_mask;
  wire [63:0] sbus_auto_SystemBusFromTiletile_anon_in_a_bits_data;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_b_ready;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_b_valid;
  wire [1:0] sbus_auto_SystemBusFromTiletile_anon_in_b_bits_param;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_b_bits_size;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_b_bits_source;
  wire [31:0] sbus_auto_SystemBusFromTiletile_anon_in_b_bits_address;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_c_ready;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_c_valid;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_opcode;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_param;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_size;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_source;
  wire [31:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_address;
  wire [63:0] sbus_auto_SystemBusFromTiletile_anon_in_c_bits_data;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_d_ready;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_d_valid;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_opcode;
  wire [1:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_param;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_size;
  wire [3:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_source;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_sink;
  wire [63:0] sbus_auto_SystemBusFromTiletile_anon_in_d_bits_data;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_d_bits_error;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_e_ready;
  wire  sbus_auto_SystemBusFromTiletile_anon_in_e_valid;
  wire [2:0] sbus_auto_SystemBusFromTiletile_anon_in_e_bits_sink;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_ready;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_valid;
  wire [2:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_opcode;
  wire [2:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_param;
  wire [2:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_size;
  wire [4:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_source;
  wire [27:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_address;
  wire [7:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_mask;
  wire [63:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_data;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_ready;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_valid;
  wire [2:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_opcode;
  wire [1:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_param;
  wire [2:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_size;
  wire [4:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_source;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_sink;
  wire [63:0] sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_data;
  wire  sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_error;
  wire  sbus_auto_SystemBus_port_TLFIFOFixer_in_a_ready;
  wire  sbus_auto_SystemBus_port_TLFIFOFixer_in_a_valid;
  wire [2:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_opcode;
  wire [2:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_param;
  wire [3:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_size;
  wire [3:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_source;
  wire [31:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_address;
  wire [7:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_mask;
  wire [63:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_data;
  wire  sbus_auto_SystemBus_port_TLFIFOFixer_in_d_ready;
  wire  sbus_auto_SystemBus_port_TLFIFOFixer_in_d_valid;
  wire [2:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_opcode;
  wire [1:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_param;
  wire [3:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_size;
  wire [3:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_source;
  wire [2:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_sink;
  wire [63:0] sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_data;
  wire  sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_error;
  wire  sbus_auto_SystemBus_slave_TLWidthWidget_out_a_ready;
  wire  sbus_auto_SystemBus_slave_TLWidthWidget_out_a_valid;
  wire [2:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_opcode;
  wire [3:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_size;
  wire [4:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_source;
  wire [30:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_address;
  wire [7:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_mask;
  wire [63:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_data;
  wire  sbus_auto_SystemBus_slave_TLWidthWidget_out_d_ready;
  wire  sbus_auto_SystemBus_slave_TLWidthWidget_out_d_valid;
  wire [2:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_opcode;
  wire [3:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_size;
  wire [4:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_source;
  wire [63:0] sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_data;
  wire  sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_error;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_a_ready;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_a_valid;
  wire [2:0] sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_opcode;
  wire [3:0] sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_size;
  wire [4:0] sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_source;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_c_ready;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_c_valid;
  wire [2:0] sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_opcode;
  wire [2:0] sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_param;
  wire [3:0] sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_size;
  wire [4:0] sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_source;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_d_ready;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_d_valid;
  wire [2:0] sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_opcode;
  wire [1:0] sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_param;
  wire [3:0] sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_size;
  wire [4:0] sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_source;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_sink;
  wire [63:0] sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_data;
  wire  sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_error;
  wire  sbus_auto_SystemBus_out_a_ready;
  wire  sbus_auto_SystemBus_out_a_valid;
  wire [2:0] sbus_auto_SystemBus_out_a_bits_opcode;
  wire [2:0] sbus_auto_SystemBus_out_a_bits_param;
  wire [2:0] sbus_auto_SystemBus_out_a_bits_size;
  wire [4:0] sbus_auto_SystemBus_out_a_bits_source;
  wire [31:0] sbus_auto_SystemBus_out_a_bits_address;
  wire [7:0] sbus_auto_SystemBus_out_a_bits_mask;
  wire [63:0] sbus_auto_SystemBus_out_a_bits_data;
  wire  sbus_auto_SystemBus_out_b_ready;
  wire  sbus_auto_SystemBus_out_b_valid;
  wire [1:0] sbus_auto_SystemBus_out_b_bits_param;
  wire [31:0] sbus_auto_SystemBus_out_b_bits_address;
  wire  sbus_auto_SystemBus_out_c_ready;
  wire  sbus_auto_SystemBus_out_c_valid;
  wire [2:0] sbus_auto_SystemBus_out_c_bits_opcode;
  wire [2:0] sbus_auto_SystemBus_out_c_bits_size;
  wire [4:0] sbus_auto_SystemBus_out_c_bits_source;
  wire [31:0] sbus_auto_SystemBus_out_c_bits_address;
  wire [63:0] sbus_auto_SystemBus_out_c_bits_data;
  wire  sbus_auto_SystemBus_out_d_ready;
  wire  sbus_auto_SystemBus_out_d_valid;
  wire [2:0] sbus_auto_SystemBus_out_d_bits_opcode;
  wire [1:0] sbus_auto_SystemBus_out_d_bits_param;
  wire [2:0] sbus_auto_SystemBus_out_d_bits_size;
  wire [4:0] sbus_auto_SystemBus_out_d_bits_source;
  wire [1:0] sbus_auto_SystemBus_out_d_bits_sink;
  wire [63:0] sbus_auto_SystemBus_out_d_bits_data;
  wire  sbus_auto_SystemBus_out_d_bits_error;
  wire  sbus_auto_SystemBus_out_e_valid;
  wire [1:0] sbus_auto_SystemBus_out_e_bits_sink;
  wire  pbus_clock;
  wire  pbus_reset;
  wire  pbus_auto_anon_in_a_ready;
  wire  pbus_auto_anon_in_a_valid;
  wire [2:0] pbus_auto_anon_in_a_bits_opcode;
  wire [2:0] pbus_auto_anon_in_a_bits_param;
  wire [2:0] pbus_auto_anon_in_a_bits_size;
  wire [4:0] pbus_auto_anon_in_a_bits_source;
  wire [27:0] pbus_auto_anon_in_a_bits_address;
  wire [7:0] pbus_auto_anon_in_a_bits_mask;
  wire [63:0] pbus_auto_anon_in_a_bits_data;
  wire  pbus_auto_anon_in_d_ready;
  wire  pbus_auto_anon_in_d_valid;
  wire [2:0] pbus_auto_anon_in_d_bits_opcode;
  wire [1:0] pbus_auto_anon_in_d_bits_param;
  wire [2:0] pbus_auto_anon_in_d_bits_size;
  wire [4:0] pbus_auto_anon_in_d_bits_source;
  wire  pbus_auto_anon_in_d_bits_sink;
  wire [63:0] pbus_auto_anon_in_d_bits_data;
  wire  pbus_auto_anon_in_d_bits_error;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_valid;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_source;
  wire [16:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_address;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_valid;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_source;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_source;
  wire [11:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_address;
  wire [7:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_mask;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_source;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_source;
  wire [25:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_address;
  wire [7:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_mask;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_source;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_source;
  wire [27:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_address;
  wire [7:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_mask;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_data;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_ready;
  wire  pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_valid;
  wire [2:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_opcode;
  wire [1:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_size;
  wire [8:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_source;
  wire [63:0] pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_data;
  wire  TLBroadcast_clock;
  wire  TLBroadcast_reset;
  wire  TLBroadcast_auto_in_a_ready;
  wire  TLBroadcast_auto_in_a_valid;
  wire [2:0] TLBroadcast_auto_in_a_bits_opcode;
  wire [2:0] TLBroadcast_auto_in_a_bits_param;
  wire [2:0] TLBroadcast_auto_in_a_bits_size;
  wire [4:0] TLBroadcast_auto_in_a_bits_source;
  wire [31:0] TLBroadcast_auto_in_a_bits_address;
  wire [7:0] TLBroadcast_auto_in_a_bits_mask;
  wire [63:0] TLBroadcast_auto_in_a_bits_data;
  wire  TLBroadcast_auto_in_b_ready;
  wire  TLBroadcast_auto_in_b_valid;
  wire [1:0] TLBroadcast_auto_in_b_bits_param;
  wire [31:0] TLBroadcast_auto_in_b_bits_address;
  wire  TLBroadcast_auto_in_c_ready;
  wire  TLBroadcast_auto_in_c_valid;
  wire [2:0] TLBroadcast_auto_in_c_bits_opcode;
  wire [2:0] TLBroadcast_auto_in_c_bits_size;
  wire [4:0] TLBroadcast_auto_in_c_bits_source;
  wire [31:0] TLBroadcast_auto_in_c_bits_address;
  wire [63:0] TLBroadcast_auto_in_c_bits_data;
  wire  TLBroadcast_auto_in_d_ready;
  wire  TLBroadcast_auto_in_d_valid;
  wire [2:0] TLBroadcast_auto_in_d_bits_opcode;
  wire [1:0] TLBroadcast_auto_in_d_bits_param;
  wire [2:0] TLBroadcast_auto_in_d_bits_size;
  wire [4:0] TLBroadcast_auto_in_d_bits_source;
  wire [1:0] TLBroadcast_auto_in_d_bits_sink;
  wire [63:0] TLBroadcast_auto_in_d_bits_data;
  wire  TLBroadcast_auto_in_d_bits_error;
  wire  TLBroadcast_auto_in_e_valid;
  wire [1:0] TLBroadcast_auto_in_e_bits_sink;
  wire  TLBroadcast_auto_out_a_ready;
  wire  TLBroadcast_auto_out_a_valid;
  wire [2:0] TLBroadcast_auto_out_a_bits_opcode;
  wire [2:0] TLBroadcast_auto_out_a_bits_size;
  wire [6:0] TLBroadcast_auto_out_a_bits_source;
  wire [31:0] TLBroadcast_auto_out_a_bits_address;
  wire [7:0] TLBroadcast_auto_out_a_bits_mask;
  wire [63:0] TLBroadcast_auto_out_a_bits_data;
  wire  TLBroadcast_auto_out_d_ready;
  wire  TLBroadcast_auto_out_d_valid;
  wire [2:0] TLBroadcast_auto_out_d_bits_opcode;
  wire [1:0] TLBroadcast_auto_out_d_bits_param;
  wire [2:0] TLBroadcast_auto_out_d_bits_size;
  wire [6:0] TLBroadcast_auto_out_d_bits_source;
  wire [63:0] TLBroadcast_auto_out_d_bits_data;
  wire  TLBroadcast_auto_out_d_bits_error;
  wire  TLWidthWidget_auto_in_a_ready;
  wire  TLWidthWidget_auto_in_a_valid;
  wire [2:0] TLWidthWidget_auto_in_a_bits_opcode;
  wire [2:0] TLWidthWidget_auto_in_a_bits_size;
  wire [6:0] TLWidthWidget_auto_in_a_bits_source;
  wire [31:0] TLWidthWidget_auto_in_a_bits_address;
  wire [7:0] TLWidthWidget_auto_in_a_bits_mask;
  wire [63:0] TLWidthWidget_auto_in_a_bits_data;
  wire  TLWidthWidget_auto_in_d_ready;
  wire  TLWidthWidget_auto_in_d_valid;
  wire [2:0] TLWidthWidget_auto_in_d_bits_opcode;
  wire [1:0] TLWidthWidget_auto_in_d_bits_param;
  wire [2:0] TLWidthWidget_auto_in_d_bits_size;
  wire [6:0] TLWidthWidget_auto_in_d_bits_source;
  wire [63:0] TLWidthWidget_auto_in_d_bits_data;
  wire  TLWidthWidget_auto_in_d_bits_error;
  wire  TLWidthWidget_auto_out_a_ready;
  wire  TLWidthWidget_auto_out_a_valid;
  wire [2:0] TLWidthWidget_auto_out_a_bits_opcode;
  wire [2:0] TLWidthWidget_auto_out_a_bits_size;
  wire [6:0] TLWidthWidget_auto_out_a_bits_source;
  wire [31:0] TLWidthWidget_auto_out_a_bits_address;
  wire [7:0] TLWidthWidget_auto_out_a_bits_mask;
  wire [63:0] TLWidthWidget_auto_out_a_bits_data;
  wire  TLWidthWidget_auto_out_d_ready;
  wire  TLWidthWidget_auto_out_d_valid;
  wire [2:0] TLWidthWidget_auto_out_d_bits_opcode;
  wire [1:0] TLWidthWidget_auto_out_d_bits_param;
  wire [2:0] TLWidthWidget_auto_out_d_bits_size;
  wire [6:0] TLWidthWidget_auto_out_d_bits_source;
  wire [63:0] TLWidthWidget_auto_out_d_bits_data;
  wire  TLWidthWidget_auto_out_d_bits_error;
  wire  memBuses_0_clock;
  wire  memBuses_0_reset;
  wire  memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_ready;
  wire  memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_valid;
  wire [2:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_opcode;
  wire [2:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_size;
  wire [6:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_source;
  wire [31:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_address;
  wire [7:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_mask;
  wire [63:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_data;
  wire  memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_ready;
  wire  memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_valid;
  wire [2:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_opcode;
  wire [2:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_size;
  wire [6:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_source;
  wire [63:0] memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_data;
  wire  memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_error;
  wire  memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_ready;
  wire  memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_valid;
  wire [2:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_opcode;
  wire [2:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_size;
  wire [6:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_source;
  wire [31:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_address;
  wire [7:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_mask;
  wire [63:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_data;
  wire  memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_ready;
  wire  memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_valid;
  wire [2:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_opcode;
  wire [1:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_param;
  wire [2:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_size;
  wire [6:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_source;
  wire [63:0] memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_data;
  wire  memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_error;
  wire  TLFilter_auto_in_a_ready;
  wire  TLFilter_auto_in_a_valid;
  wire [2:0] TLFilter_auto_in_a_bits_opcode;
  wire [2:0] TLFilter_auto_in_a_bits_size;
  wire [6:0] TLFilter_auto_in_a_bits_source;
  wire [31:0] TLFilter_auto_in_a_bits_address;
  wire [7:0] TLFilter_auto_in_a_bits_mask;
  wire [63:0] TLFilter_auto_in_a_bits_data;
  wire  TLFilter_auto_in_d_ready;
  wire  TLFilter_auto_in_d_valid;
  wire [2:0] TLFilter_auto_in_d_bits_opcode;
  wire [1:0] TLFilter_auto_in_d_bits_param;
  wire [2:0] TLFilter_auto_in_d_bits_size;
  wire [6:0] TLFilter_auto_in_d_bits_source;
  wire [63:0] TLFilter_auto_in_d_bits_data;
  wire  TLFilter_auto_in_d_bits_error;
  wire  TLFilter_auto_out_a_ready;
  wire  TLFilter_auto_out_a_valid;
  wire [2:0] TLFilter_auto_out_a_bits_opcode;
  wire [2:0] TLFilter_auto_out_a_bits_size;
  wire [6:0] TLFilter_auto_out_a_bits_source;
  wire [31:0] TLFilter_auto_out_a_bits_address;
  wire [7:0] TLFilter_auto_out_a_bits_mask;
  wire [63:0] TLFilter_auto_out_a_bits_data;
  wire  TLFilter_auto_out_d_ready;
  wire  TLFilter_auto_out_d_valid;
  wire [2:0] TLFilter_auto_out_d_bits_opcode;
  wire [1:0] TLFilter_auto_out_d_bits_param;
  wire [2:0] TLFilter_auto_out_d_bits_size;
  wire [6:0] TLFilter_auto_out_d_bits_source;
  wire [63:0] TLFilter_auto_out_d_bits_data;
  wire  TLFilter_auto_out_d_bits_error;
  wire  plic_clock;
  wire  plic_reset;
  wire  plic_auto_int_in_0;
  wire  plic_auto_int_in_1;
  wire  plic_auto_int_out_1_0;
  wire  plic_auto_int_out_0_0;
  wire  plic_auto_in_a_ready;
  wire  plic_auto_in_a_valid;
  wire [2:0] plic_auto_in_a_bits_opcode;
  wire [1:0] plic_auto_in_a_bits_size;
  wire [8:0] plic_auto_in_a_bits_source;
  wire [27:0] plic_auto_in_a_bits_address;
  wire [7:0] plic_auto_in_a_bits_mask;
  wire [63:0] plic_auto_in_a_bits_data;
  wire  plic_auto_in_d_ready;
  wire  plic_auto_in_d_valid;
  wire [2:0] plic_auto_in_d_bits_opcode;
  wire [1:0] plic_auto_in_d_bits_size;
  wire [8:0] plic_auto_in_d_bits_source;
  wire [63:0] plic_auto_in_d_bits_data;
  wire  clint_clock;
  wire  clint_reset;
  wire  clint_auto_int_out_0;
  wire  clint_auto_int_out_1;
  wire  clint_auto_in_a_ready;
  wire  clint_auto_in_a_valid;
  wire [2:0] clint_auto_in_a_bits_opcode;
  wire [1:0] clint_auto_in_a_bits_size;
  wire [8:0] clint_auto_in_a_bits_source;
  wire [25:0] clint_auto_in_a_bits_address;
  wire [7:0] clint_auto_in_a_bits_mask;
  wire [63:0] clint_auto_in_a_bits_data;
  wire  clint_auto_in_d_ready;
  wire  clint_auto_in_d_valid;
  wire [2:0] clint_auto_in_d_bits_opcode;
  wire [1:0] clint_auto_in_d_bits_size;
  wire [8:0] clint_auto_in_d_bits_source;
  wire [63:0] clint_auto_in_d_bits_data;
  wire  clint_io_rtcTick;
  wire  debug_1_clock;
  wire  debug_1_reset;
  wire  debug_1_auto_dmInner_dmInner_tl_in_a_ready;
  wire  debug_1_auto_dmInner_dmInner_tl_in_a_valid;
  wire [2:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode;
  wire [1:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_size;
  wire [8:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_source;
  wire [11:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_address;
  wire [7:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask;
  wire [63:0] debug_1_auto_dmInner_dmInner_tl_in_a_bits_data;
  wire  debug_1_auto_dmInner_dmInner_tl_in_d_ready;
  wire  debug_1_auto_dmInner_dmInner_tl_in_d_valid;
  wire [2:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode;
  wire [1:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_size;
  wire [8:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_source;
  wire [63:0] debug_1_auto_dmInner_dmInner_tl_in_d_bits_data;
  wire  debug_1_auto_dmOuter_anon_out_sync_0;
  wire  debug_1_io_ctrl_ndreset;
  wire  debug_1_io_ctrl_dmactive;
  wire  debug_1_io_dmi_dmi_req_ready;
  wire  debug_1_io_dmi_dmi_req_valid;
  wire [6:0] debug_1_io_dmi_dmi_req_bits_addr;
  wire [31:0] debug_1_io_dmi_dmi_req_bits_data;
  wire [1:0] debug_1_io_dmi_dmi_req_bits_op;
  wire  debug_1_io_dmi_dmi_resp_ready;
  wire  debug_1_io_dmi_dmi_resp_valid;
  wire [31:0] debug_1_io_dmi_dmi_resp_bits_data;
  wire [1:0] debug_1_io_dmi_dmi_resp_bits_resp;
  wire  debug_1_io_dmi_dmiClock;
  wire  debug_1_io_dmi_dmiReset;
  wire  tile_clock;
  wire  tile_reset;
  wire  tile_auto_anon_in_3_sync_0;
  wire  tile_auto_anon_in_2_sync_0;
  wire  tile_auto_anon_in_1_sync_0;
  wire  tile_auto_anon_in_1_sync_1;
  wire  tile_auto_anon_in_0_sync_0;
  wire  tile_auto_anon_out_a_ready;
  wire  tile_auto_anon_out_a_valid;
  wire [2:0] tile_auto_anon_out_a_bits_opcode;
  wire [2:0] tile_auto_anon_out_a_bits_param;
  wire [3:0] tile_auto_anon_out_a_bits_size;
  wire [3:0] tile_auto_anon_out_a_bits_source;
  wire [31:0] tile_auto_anon_out_a_bits_address;
  wire [7:0] tile_auto_anon_out_a_bits_mask;
  wire [63:0] tile_auto_anon_out_a_bits_data;
  wire  tile_auto_anon_out_b_ready;
  wire  tile_auto_anon_out_b_valid;
  wire [1:0] tile_auto_anon_out_b_bits_param;
  wire [3:0] tile_auto_anon_out_b_bits_size;
  wire [3:0] tile_auto_anon_out_b_bits_source;
  wire [31:0] tile_auto_anon_out_b_bits_address;
  wire  tile_auto_anon_out_c_ready;
  wire  tile_auto_anon_out_c_valid;
  wire [2:0] tile_auto_anon_out_c_bits_opcode;
  wire [2:0] tile_auto_anon_out_c_bits_param;
  wire [3:0] tile_auto_anon_out_c_bits_size;
  wire [3:0] tile_auto_anon_out_c_bits_source;
  wire [31:0] tile_auto_anon_out_c_bits_address;
  wire [63:0] tile_auto_anon_out_c_bits_data;
  wire  tile_auto_anon_out_d_ready;
  wire  tile_auto_anon_out_d_valid;
  wire [2:0] tile_auto_anon_out_d_bits_opcode;
  wire [1:0] tile_auto_anon_out_d_bits_param;
  wire [3:0] tile_auto_anon_out_d_bits_size;
  wire [3:0] tile_auto_anon_out_d_bits_source;
  wire [2:0] tile_auto_anon_out_d_bits_sink;
  wire [63:0] tile_auto_anon_out_d_bits_data;
  wire  tile_auto_anon_out_d_bits_error;
  wire  tile_auto_anon_out_e_ready;
  wire  tile_auto_anon_out_e_valid;
  wire [2:0] tile_auto_anon_out_e_bits_sink;
  wire  IntSyncCrossingSource_clock;
  wire  IntSyncCrossingSource_reset;
  wire  IntSyncCrossingSource_auto_in_2_0;
  wire  IntSyncCrossingSource_auto_in_1_0;
  wire  IntSyncCrossingSource_auto_in_0_0;
  wire  IntSyncCrossingSource_auto_in_0_1;
  wire  IntSyncCrossingSource_auto_out_2_sync_0;
  wire  IntSyncCrossingSource_auto_out_1_sync_0;
  wire  IntSyncCrossingSource_auto_out_0_sync_0;
  wire  IntSyncCrossingSource_auto_out_0_sync_1;
  wire  IntXing_clock;
  wire  IntXing_auto_int_in_0;
  wire  IntXing_auto_int_in_1;
  wire  IntXing_auto_int_out_0;
  wire  IntXing_auto_int_out_1;
  wire  converter_clock;
  wire  converter_reset;
  wire  converter_auto_in_a_ready;
  wire  converter_auto_in_a_valid;
  wire [2:0] converter_auto_in_a_bits_opcode;
  wire [2:0] converter_auto_in_a_bits_size;
  wire [6:0] converter_auto_in_a_bits_source;
  wire [31:0] converter_auto_in_a_bits_address;
  wire [7:0] converter_auto_in_a_bits_mask;
  wire [63:0] converter_auto_in_a_bits_data;
  wire  converter_auto_in_d_ready;
  wire  converter_auto_in_d_valid;
  wire [2:0] converter_auto_in_d_bits_opcode;
  wire [2:0] converter_auto_in_d_bits_size;
  wire [6:0] converter_auto_in_d_bits_source;
  wire [63:0] converter_auto_in_d_bits_data;
  wire  converter_auto_in_d_bits_error;
  wire  converter_auto_out_aw_ready;
  wire  converter_auto_out_aw_valid;
  wire [6:0] converter_auto_out_aw_bits_id;
  wire [31:0] converter_auto_out_aw_bits_addr;
  wire [7:0] converter_auto_out_aw_bits_len;
  wire [2:0] converter_auto_out_aw_bits_size;
  wire [1:0] converter_auto_out_aw_bits_burst;
  wire  converter_auto_out_aw_bits_lock;
  wire [3:0] converter_auto_out_aw_bits_cache;
  wire [2:0] converter_auto_out_aw_bits_prot;
  wire [3:0] converter_auto_out_aw_bits_qos;
  wire [10:0] converter_auto_out_aw_bits_user;
  wire  converter_auto_out_w_ready;
  wire  converter_auto_out_w_valid;
  wire [63:0] converter_auto_out_w_bits_data;
  wire [7:0] converter_auto_out_w_bits_strb;
  wire  converter_auto_out_w_bits_last;
  wire  converter_auto_out_b_ready;
  wire  converter_auto_out_b_valid;
  wire [6:0] converter_auto_out_b_bits_id;
  wire [1:0] converter_auto_out_b_bits_resp;
  wire [10:0] converter_auto_out_b_bits_user;
  wire  converter_auto_out_ar_ready;
  wire  converter_auto_out_ar_valid;
  wire [6:0] converter_auto_out_ar_bits_id;
  wire [31:0] converter_auto_out_ar_bits_addr;
  wire [7:0] converter_auto_out_ar_bits_len;
  wire [2:0] converter_auto_out_ar_bits_size;
  wire [1:0] converter_auto_out_ar_bits_burst;
  wire  converter_auto_out_ar_bits_lock;
  wire [3:0] converter_auto_out_ar_bits_cache;
  wire [2:0] converter_auto_out_ar_bits_prot;
  wire [3:0] converter_auto_out_ar_bits_qos;
  wire [10:0] converter_auto_out_ar_bits_user;
  wire  converter_auto_out_r_ready;
  wire  converter_auto_out_r_valid;
  wire [6:0] converter_auto_out_r_bits_id;
  wire [63:0] converter_auto_out_r_bits_data;
  wire [1:0] converter_auto_out_r_bits_resp;
  wire [10:0] converter_auto_out_r_bits_user;
  wire  converter_auto_out_r_bits_last;
  wire  trim_auto_in_aw_ready;
  wire  trim_auto_in_aw_valid;
  wire [6:0] trim_auto_in_aw_bits_id;
  wire [31:0] trim_auto_in_aw_bits_addr;
  wire [7:0] trim_auto_in_aw_bits_len;
  wire [2:0] trim_auto_in_aw_bits_size;
  wire [1:0] trim_auto_in_aw_bits_burst;
  wire  trim_auto_in_aw_bits_lock;
  wire [3:0] trim_auto_in_aw_bits_cache;
  wire [2:0] trim_auto_in_aw_bits_prot;
  wire [3:0] trim_auto_in_aw_bits_qos;
  wire [10:0] trim_auto_in_aw_bits_user;
  wire  trim_auto_in_w_ready;
  wire  trim_auto_in_w_valid;
  wire [63:0] trim_auto_in_w_bits_data;
  wire [7:0] trim_auto_in_w_bits_strb;
  wire  trim_auto_in_w_bits_last;
  wire  trim_auto_in_b_ready;
  wire  trim_auto_in_b_valid;
  wire [6:0] trim_auto_in_b_bits_id;
  wire [1:0] trim_auto_in_b_bits_resp;
  wire [10:0] trim_auto_in_b_bits_user;
  wire  trim_auto_in_ar_ready;
  wire  trim_auto_in_ar_valid;
  wire [6:0] trim_auto_in_ar_bits_id;
  wire [31:0] trim_auto_in_ar_bits_addr;
  wire [7:0] trim_auto_in_ar_bits_len;
  wire [2:0] trim_auto_in_ar_bits_size;
  wire [1:0] trim_auto_in_ar_bits_burst;
  wire  trim_auto_in_ar_bits_lock;
  wire [3:0] trim_auto_in_ar_bits_cache;
  wire [2:0] trim_auto_in_ar_bits_prot;
  wire [3:0] trim_auto_in_ar_bits_qos;
  wire [10:0] trim_auto_in_ar_bits_user;
  wire  trim_auto_in_r_ready;
  wire  trim_auto_in_r_valid;
  wire [6:0] trim_auto_in_r_bits_id;
  wire [63:0] trim_auto_in_r_bits_data;
  wire [1:0] trim_auto_in_r_bits_resp;
  wire [10:0] trim_auto_in_r_bits_user;
  wire  trim_auto_in_r_bits_last;
  wire  trim_auto_out_aw_ready;
  wire  trim_auto_out_aw_valid;
  wire [3:0] trim_auto_out_aw_bits_id;
  wire [31:0] trim_auto_out_aw_bits_addr;
  wire [7:0] trim_auto_out_aw_bits_len;
  wire [2:0] trim_auto_out_aw_bits_size;
  wire [1:0] trim_auto_out_aw_bits_burst;
  wire  trim_auto_out_aw_bits_lock;
  wire [3:0] trim_auto_out_aw_bits_cache;
  wire [2:0] trim_auto_out_aw_bits_prot;
  wire [3:0] trim_auto_out_aw_bits_qos;
  wire [13:0] trim_auto_out_aw_bits_user;
  wire  trim_auto_out_w_ready;
  wire  trim_auto_out_w_valid;
  wire [63:0] trim_auto_out_w_bits_data;
  wire [7:0] trim_auto_out_w_bits_strb;
  wire  trim_auto_out_w_bits_last;
  wire  trim_auto_out_b_ready;
  wire  trim_auto_out_b_valid;
  wire [3:0] trim_auto_out_b_bits_id;
  wire [1:0] trim_auto_out_b_bits_resp;
  wire [13:0] trim_auto_out_b_bits_user;
  wire  trim_auto_out_ar_ready;
  wire  trim_auto_out_ar_valid;
  wire [3:0] trim_auto_out_ar_bits_id;
  wire [31:0] trim_auto_out_ar_bits_addr;
  wire [7:0] trim_auto_out_ar_bits_len;
  wire [2:0] trim_auto_out_ar_bits_size;
  wire [1:0] trim_auto_out_ar_bits_burst;
  wire  trim_auto_out_ar_bits_lock;
  wire [3:0] trim_auto_out_ar_bits_cache;
  wire [2:0] trim_auto_out_ar_bits_prot;
  wire [3:0] trim_auto_out_ar_bits_qos;
  wire [13:0] trim_auto_out_ar_bits_user;
  wire  trim_auto_out_r_ready;
  wire  trim_auto_out_r_valid;
  wire [3:0] trim_auto_out_r_bits_id;
  wire [63:0] trim_auto_out_r_bits_data;
  wire [1:0] trim_auto_out_r_bits_resp;
  wire [13:0] trim_auto_out_r_bits_user;
  wire  trim_auto_out_r_bits_last;
  wire  yank_clock;
  wire  yank_reset;
  wire  yank_auto_in_aw_ready;
  wire  yank_auto_in_aw_valid;
  wire [3:0] yank_auto_in_aw_bits_id;
  wire [31:0] yank_auto_in_aw_bits_addr;
  wire [7:0] yank_auto_in_aw_bits_len;
  wire [2:0] yank_auto_in_aw_bits_size;
  wire [1:0] yank_auto_in_aw_bits_burst;
  wire  yank_auto_in_aw_bits_lock;
  wire [3:0] yank_auto_in_aw_bits_cache;
  wire [2:0] yank_auto_in_aw_bits_prot;
  wire [3:0] yank_auto_in_aw_bits_qos;
  wire [13:0] yank_auto_in_aw_bits_user;
  wire  yank_auto_in_w_ready;
  wire  yank_auto_in_w_valid;
  wire [63:0] yank_auto_in_w_bits_data;
  wire [7:0] yank_auto_in_w_bits_strb;
  wire  yank_auto_in_w_bits_last;
  wire  yank_auto_in_b_ready;
  wire  yank_auto_in_b_valid;
  wire [3:0] yank_auto_in_b_bits_id;
  wire [1:0] yank_auto_in_b_bits_resp;
  wire [13:0] yank_auto_in_b_bits_user;
  wire  yank_auto_in_ar_ready;
  wire  yank_auto_in_ar_valid;
  wire [3:0] yank_auto_in_ar_bits_id;
  wire [31:0] yank_auto_in_ar_bits_addr;
  wire [7:0] yank_auto_in_ar_bits_len;
  wire [2:0] yank_auto_in_ar_bits_size;
  wire [1:0] yank_auto_in_ar_bits_burst;
  wire  yank_auto_in_ar_bits_lock;
  wire [3:0] yank_auto_in_ar_bits_cache;
  wire [2:0] yank_auto_in_ar_bits_prot;
  wire [3:0] yank_auto_in_ar_bits_qos;
  wire [13:0] yank_auto_in_ar_bits_user;
  wire  yank_auto_in_r_ready;
  wire  yank_auto_in_r_valid;
  wire [3:0] yank_auto_in_r_bits_id;
  wire [63:0] yank_auto_in_r_bits_data;
  wire [1:0] yank_auto_in_r_bits_resp;
  wire [13:0] yank_auto_in_r_bits_user;
  wire  yank_auto_in_r_bits_last;
  wire  yank_auto_out_aw_ready;
  wire  yank_auto_out_aw_valid;
  wire [3:0] yank_auto_out_aw_bits_id;
  wire [31:0] yank_auto_out_aw_bits_addr;
  wire [7:0] yank_auto_out_aw_bits_len;
  wire [2:0] yank_auto_out_aw_bits_size;
  wire [1:0] yank_auto_out_aw_bits_burst;
  wire  yank_auto_out_aw_bits_lock;
  wire [3:0] yank_auto_out_aw_bits_cache;
  wire [2:0] yank_auto_out_aw_bits_prot;
  wire [3:0] yank_auto_out_aw_bits_qos;
  wire  yank_auto_out_w_ready;
  wire  yank_auto_out_w_valid;
  wire [63:0] yank_auto_out_w_bits_data;
  wire [7:0] yank_auto_out_w_bits_strb;
  wire  yank_auto_out_w_bits_last;
  wire  yank_auto_out_b_ready;
  wire  yank_auto_out_b_valid;
  wire [3:0] yank_auto_out_b_bits_id;
  wire [1:0] yank_auto_out_b_bits_resp;
  wire  yank_auto_out_ar_ready;
  wire  yank_auto_out_ar_valid;
  wire [3:0] yank_auto_out_ar_bits_id;
  wire [31:0] yank_auto_out_ar_bits_addr;
  wire [7:0] yank_auto_out_ar_bits_len;
  wire [2:0] yank_auto_out_ar_bits_size;
  wire [1:0] yank_auto_out_ar_bits_burst;
  wire  yank_auto_out_ar_bits_lock;
  wire [3:0] yank_auto_out_ar_bits_cache;
  wire [2:0] yank_auto_out_ar_bits_prot;
  wire [3:0] yank_auto_out_ar_bits_qos;
  wire  yank_auto_out_r_ready;
  wire  yank_auto_out_r_valid;
  wire [3:0] yank_auto_out_r_bits_id;
  wire [63:0] yank_auto_out_r_bits_data;
  wire [1:0] yank_auto_out_r_bits_resp;
  wire  yank_auto_out_r_bits_last;
  wire  buffer_clock;
  wire  buffer_reset;
  wire  buffer_auto_in_aw_ready;
  wire  buffer_auto_in_aw_valid;
  wire [3:0] buffer_auto_in_aw_bits_id;
  wire [31:0] buffer_auto_in_aw_bits_addr;
  wire [7:0] buffer_auto_in_aw_bits_len;
  wire [2:0] buffer_auto_in_aw_bits_size;
  wire [1:0] buffer_auto_in_aw_bits_burst;
  wire  buffer_auto_in_aw_bits_lock;
  wire [3:0] buffer_auto_in_aw_bits_cache;
  wire [2:0] buffer_auto_in_aw_bits_prot;
  wire [3:0] buffer_auto_in_aw_bits_qos;
  wire  buffer_auto_in_w_ready;
  wire  buffer_auto_in_w_valid;
  wire [63:0] buffer_auto_in_w_bits_data;
  wire [7:0] buffer_auto_in_w_bits_strb;
  wire  buffer_auto_in_w_bits_last;
  wire  buffer_auto_in_b_ready;
  wire  buffer_auto_in_b_valid;
  wire [3:0] buffer_auto_in_b_bits_id;
  wire [1:0] buffer_auto_in_b_bits_resp;
  wire  buffer_auto_in_ar_ready;
  wire  buffer_auto_in_ar_valid;
  wire [3:0] buffer_auto_in_ar_bits_id;
  wire [31:0] buffer_auto_in_ar_bits_addr;
  wire [7:0] buffer_auto_in_ar_bits_len;
  wire [2:0] buffer_auto_in_ar_bits_size;
  wire [1:0] buffer_auto_in_ar_bits_burst;
  wire  buffer_auto_in_ar_bits_lock;
  wire [3:0] buffer_auto_in_ar_bits_cache;
  wire [2:0] buffer_auto_in_ar_bits_prot;
  wire [3:0] buffer_auto_in_ar_bits_qos;
  wire  buffer_auto_in_r_ready;
  wire  buffer_auto_in_r_valid;
  wire [3:0] buffer_auto_in_r_bits_id;
  wire [63:0] buffer_auto_in_r_bits_data;
  wire [1:0] buffer_auto_in_r_bits_resp;
  wire  buffer_auto_in_r_bits_last;
  wire  buffer_auto_out_aw_ready;
  wire  buffer_auto_out_aw_valid;
  wire [3:0] buffer_auto_out_aw_bits_id;
  wire [31:0] buffer_auto_out_aw_bits_addr;
  wire [7:0] buffer_auto_out_aw_bits_len;
  wire [2:0] buffer_auto_out_aw_bits_size;
  wire [1:0] buffer_auto_out_aw_bits_burst;
  wire  buffer_auto_out_aw_bits_lock;
  wire [3:0] buffer_auto_out_aw_bits_cache;
  wire [2:0] buffer_auto_out_aw_bits_prot;
  wire [3:0] buffer_auto_out_aw_bits_qos;
  wire  buffer_auto_out_w_ready;
  wire  buffer_auto_out_w_valid;
  wire [63:0] buffer_auto_out_w_bits_data;
  wire [7:0] buffer_auto_out_w_bits_strb;
  wire  buffer_auto_out_w_bits_last;
  wire  buffer_auto_out_b_ready;
  wire  buffer_auto_out_b_valid;
  wire [3:0] buffer_auto_out_b_bits_id;
  wire [1:0] buffer_auto_out_b_bits_resp;
  wire  buffer_auto_out_ar_ready;
  wire  buffer_auto_out_ar_valid;
  wire [3:0] buffer_auto_out_ar_bits_id;
  wire [31:0] buffer_auto_out_ar_bits_addr;
  wire [7:0] buffer_auto_out_ar_bits_len;
  wire [2:0] buffer_auto_out_ar_bits_size;
  wire [1:0] buffer_auto_out_ar_bits_burst;
  wire  buffer_auto_out_ar_bits_lock;
  wire [3:0] buffer_auto_out_ar_bits_cache;
  wire [2:0] buffer_auto_out_ar_bits_prot;
  wire [3:0] buffer_auto_out_ar_bits_qos;
  wire  buffer_auto_out_r_ready;
  wire  buffer_auto_out_r_valid;
  wire [3:0] buffer_auto_out_r_bits_id;
  wire [63:0] buffer_auto_out_r_bits_data;
  wire [1:0] buffer_auto_out_r_bits_resp;
  wire  buffer_auto_out_r_bits_last;
  wire  AXI4Buffer_clock;
  wire  AXI4Buffer_reset;
  wire  AXI4Buffer_auto_in_aw_ready;
  wire  AXI4Buffer_auto_in_aw_valid;
  wire [3:0] AXI4Buffer_auto_in_aw_bits_id;
  wire [30:0] AXI4Buffer_auto_in_aw_bits_addr;
  wire [7:0] AXI4Buffer_auto_in_aw_bits_len;
  wire [2:0] AXI4Buffer_auto_in_aw_bits_size;
  wire [1:0] AXI4Buffer_auto_in_aw_bits_burst;
  wire  AXI4Buffer_auto_in_aw_bits_lock;
  wire [3:0] AXI4Buffer_auto_in_aw_bits_cache;
  wire [2:0] AXI4Buffer_auto_in_aw_bits_prot;
  wire [3:0] AXI4Buffer_auto_in_aw_bits_qos;
  wire  AXI4Buffer_auto_in_w_ready;
  wire  AXI4Buffer_auto_in_w_valid;
  wire [63:0] AXI4Buffer_auto_in_w_bits_data;
  wire [7:0] AXI4Buffer_auto_in_w_bits_strb;
  wire  AXI4Buffer_auto_in_w_bits_last;
  wire  AXI4Buffer_auto_in_b_ready;
  wire  AXI4Buffer_auto_in_b_valid;
  wire [3:0] AXI4Buffer_auto_in_b_bits_id;
  wire [1:0] AXI4Buffer_auto_in_b_bits_resp;
  wire  AXI4Buffer_auto_in_ar_ready;
  wire  AXI4Buffer_auto_in_ar_valid;
  wire [3:0] AXI4Buffer_auto_in_ar_bits_id;
  wire [30:0] AXI4Buffer_auto_in_ar_bits_addr;
  wire [7:0] AXI4Buffer_auto_in_ar_bits_len;
  wire [2:0] AXI4Buffer_auto_in_ar_bits_size;
  wire [1:0] AXI4Buffer_auto_in_ar_bits_burst;
  wire  AXI4Buffer_auto_in_ar_bits_lock;
  wire [3:0] AXI4Buffer_auto_in_ar_bits_cache;
  wire [2:0] AXI4Buffer_auto_in_ar_bits_prot;
  wire [3:0] AXI4Buffer_auto_in_ar_bits_qos;
  wire  AXI4Buffer_auto_in_r_ready;
  wire  AXI4Buffer_auto_in_r_valid;
  wire [3:0] AXI4Buffer_auto_in_r_bits_id;
  wire [63:0] AXI4Buffer_auto_in_r_bits_data;
  wire [1:0] AXI4Buffer_auto_in_r_bits_resp;
  wire  AXI4Buffer_auto_in_r_bits_last;
  wire  AXI4Buffer_auto_out_aw_ready;
  wire  AXI4Buffer_auto_out_aw_valid;
  wire [3:0] AXI4Buffer_auto_out_aw_bits_id;
  wire [30:0] AXI4Buffer_auto_out_aw_bits_addr;
  wire [7:0] AXI4Buffer_auto_out_aw_bits_len;
  wire [2:0] AXI4Buffer_auto_out_aw_bits_size;
  wire [1:0] AXI4Buffer_auto_out_aw_bits_burst;
  wire  AXI4Buffer_auto_out_aw_bits_lock;
  wire [3:0] AXI4Buffer_auto_out_aw_bits_cache;
  wire [2:0] AXI4Buffer_auto_out_aw_bits_prot;
  wire [3:0] AXI4Buffer_auto_out_aw_bits_qos;
  wire  AXI4Buffer_auto_out_w_ready;
  wire  AXI4Buffer_auto_out_w_valid;
  wire [63:0] AXI4Buffer_auto_out_w_bits_data;
  wire [7:0] AXI4Buffer_auto_out_w_bits_strb;
  wire  AXI4Buffer_auto_out_w_bits_last;
  wire  AXI4Buffer_auto_out_b_ready;
  wire  AXI4Buffer_auto_out_b_valid;
  wire [3:0] AXI4Buffer_auto_out_b_bits_id;
  wire [1:0] AXI4Buffer_auto_out_b_bits_resp;
  wire  AXI4Buffer_auto_out_ar_ready;
  wire  AXI4Buffer_auto_out_ar_valid;
  wire [3:0] AXI4Buffer_auto_out_ar_bits_id;
  wire [30:0] AXI4Buffer_auto_out_ar_bits_addr;
  wire [7:0] AXI4Buffer_auto_out_ar_bits_len;
  wire [2:0] AXI4Buffer_auto_out_ar_bits_size;
  wire [1:0] AXI4Buffer_auto_out_ar_bits_burst;
  wire  AXI4Buffer_auto_out_ar_bits_lock;
  wire [3:0] AXI4Buffer_auto_out_ar_bits_cache;
  wire [2:0] AXI4Buffer_auto_out_ar_bits_prot;
  wire [3:0] AXI4Buffer_auto_out_ar_bits_qos;
  wire  AXI4Buffer_auto_out_r_ready;
  wire  AXI4Buffer_auto_out_r_valid;
  wire [3:0] AXI4Buffer_auto_out_r_bits_id;
  wire [63:0] AXI4Buffer_auto_out_r_bits_data;
  wire [1:0] AXI4Buffer_auto_out_r_bits_resp;
  wire  AXI4Buffer_auto_out_r_bits_last;
  wire  AXI4UserYanker_clock;
  wire  AXI4UserYanker_reset;
  wire  AXI4UserYanker_auto_in_aw_ready;
  wire  AXI4UserYanker_auto_in_aw_valid;
  wire [3:0] AXI4UserYanker_auto_in_aw_bits_id;
  wire [30:0] AXI4UserYanker_auto_in_aw_bits_addr;
  wire [7:0] AXI4UserYanker_auto_in_aw_bits_len;
  wire [2:0] AXI4UserYanker_auto_in_aw_bits_size;
  wire [1:0] AXI4UserYanker_auto_in_aw_bits_burst;
  wire  AXI4UserYanker_auto_in_aw_bits_lock;
  wire [3:0] AXI4UserYanker_auto_in_aw_bits_cache;
  wire [2:0] AXI4UserYanker_auto_in_aw_bits_prot;
  wire [3:0] AXI4UserYanker_auto_in_aw_bits_qos;
  wire [8:0] AXI4UserYanker_auto_in_aw_bits_user;
  wire  AXI4UserYanker_auto_in_w_ready;
  wire  AXI4UserYanker_auto_in_w_valid;
  wire [63:0] AXI4UserYanker_auto_in_w_bits_data;
  wire [7:0] AXI4UserYanker_auto_in_w_bits_strb;
  wire  AXI4UserYanker_auto_in_w_bits_last;
  wire  AXI4UserYanker_auto_in_b_ready;
  wire  AXI4UserYanker_auto_in_b_valid;
  wire [3:0] AXI4UserYanker_auto_in_b_bits_id;
  wire [1:0] AXI4UserYanker_auto_in_b_bits_resp;
  wire [8:0] AXI4UserYanker_auto_in_b_bits_user;
  wire  AXI4UserYanker_auto_in_ar_ready;
  wire  AXI4UserYanker_auto_in_ar_valid;
  wire [3:0] AXI4UserYanker_auto_in_ar_bits_id;
  wire [30:0] AXI4UserYanker_auto_in_ar_bits_addr;
  wire [7:0] AXI4UserYanker_auto_in_ar_bits_len;
  wire [2:0] AXI4UserYanker_auto_in_ar_bits_size;
  wire [1:0] AXI4UserYanker_auto_in_ar_bits_burst;
  wire  AXI4UserYanker_auto_in_ar_bits_lock;
  wire [3:0] AXI4UserYanker_auto_in_ar_bits_cache;
  wire [2:0] AXI4UserYanker_auto_in_ar_bits_prot;
  wire [3:0] AXI4UserYanker_auto_in_ar_bits_qos;
  wire [8:0] AXI4UserYanker_auto_in_ar_bits_user;
  wire  AXI4UserYanker_auto_in_r_ready;
  wire  AXI4UserYanker_auto_in_r_valid;
  wire [3:0] AXI4UserYanker_auto_in_r_bits_id;
  wire [63:0] AXI4UserYanker_auto_in_r_bits_data;
  wire [1:0] AXI4UserYanker_auto_in_r_bits_resp;
  wire [8:0] AXI4UserYanker_auto_in_r_bits_user;
  wire  AXI4UserYanker_auto_in_r_bits_last;
  wire  AXI4UserYanker_auto_out_aw_ready;
  wire  AXI4UserYanker_auto_out_aw_valid;
  wire [3:0] AXI4UserYanker_auto_out_aw_bits_id;
  wire [30:0] AXI4UserYanker_auto_out_aw_bits_addr;
  wire [7:0] AXI4UserYanker_auto_out_aw_bits_len;
  wire [2:0] AXI4UserYanker_auto_out_aw_bits_size;
  wire [1:0] AXI4UserYanker_auto_out_aw_bits_burst;
  wire  AXI4UserYanker_auto_out_aw_bits_lock;
  wire [3:0] AXI4UserYanker_auto_out_aw_bits_cache;
  wire [2:0] AXI4UserYanker_auto_out_aw_bits_prot;
  wire [3:0] AXI4UserYanker_auto_out_aw_bits_qos;
  wire  AXI4UserYanker_auto_out_w_ready;
  wire  AXI4UserYanker_auto_out_w_valid;
  wire [63:0] AXI4UserYanker_auto_out_w_bits_data;
  wire [7:0] AXI4UserYanker_auto_out_w_bits_strb;
  wire  AXI4UserYanker_auto_out_w_bits_last;
  wire  AXI4UserYanker_auto_out_b_ready;
  wire  AXI4UserYanker_auto_out_b_valid;
  wire [3:0] AXI4UserYanker_auto_out_b_bits_id;
  wire [1:0] AXI4UserYanker_auto_out_b_bits_resp;
  wire  AXI4UserYanker_auto_out_ar_ready;
  wire  AXI4UserYanker_auto_out_ar_valid;
  wire [3:0] AXI4UserYanker_auto_out_ar_bits_id;
  wire [30:0] AXI4UserYanker_auto_out_ar_bits_addr;
  wire [7:0] AXI4UserYanker_auto_out_ar_bits_len;
  wire [2:0] AXI4UserYanker_auto_out_ar_bits_size;
  wire [1:0] AXI4UserYanker_auto_out_ar_bits_burst;
  wire  AXI4UserYanker_auto_out_ar_bits_lock;
  wire [3:0] AXI4UserYanker_auto_out_ar_bits_cache;
  wire [2:0] AXI4UserYanker_auto_out_ar_bits_prot;
  wire [3:0] AXI4UserYanker_auto_out_ar_bits_qos;
  wire  AXI4UserYanker_auto_out_r_ready;
  wire  AXI4UserYanker_auto_out_r_valid;
  wire [3:0] AXI4UserYanker_auto_out_r_bits_id;
  wire [63:0] AXI4UserYanker_auto_out_r_bits_data;
  wire [1:0] AXI4UserYanker_auto_out_r_bits_resp;
  wire  AXI4UserYanker_auto_out_r_bits_last;
  wire  AXI4Deinterleaver_clock;
  wire  AXI4Deinterleaver_reset;
  wire  AXI4Deinterleaver_auto_in_aw_ready;
  wire  AXI4Deinterleaver_auto_in_aw_valid;
  wire [3:0] AXI4Deinterleaver_auto_in_aw_bits_id;
  wire [30:0] AXI4Deinterleaver_auto_in_aw_bits_addr;
  wire [7:0] AXI4Deinterleaver_auto_in_aw_bits_len;
  wire [2:0] AXI4Deinterleaver_auto_in_aw_bits_size;
  wire [1:0] AXI4Deinterleaver_auto_in_aw_bits_burst;
  wire  AXI4Deinterleaver_auto_in_aw_bits_lock;
  wire [3:0] AXI4Deinterleaver_auto_in_aw_bits_cache;
  wire [2:0] AXI4Deinterleaver_auto_in_aw_bits_prot;
  wire [3:0] AXI4Deinterleaver_auto_in_aw_bits_qos;
  wire [8:0] AXI4Deinterleaver_auto_in_aw_bits_user;
  wire  AXI4Deinterleaver_auto_in_w_ready;
  wire  AXI4Deinterleaver_auto_in_w_valid;
  wire [63:0] AXI4Deinterleaver_auto_in_w_bits_data;
  wire [7:0] AXI4Deinterleaver_auto_in_w_bits_strb;
  wire  AXI4Deinterleaver_auto_in_w_bits_last;
  wire  AXI4Deinterleaver_auto_in_b_ready;
  wire  AXI4Deinterleaver_auto_in_b_valid;
  wire [3:0] AXI4Deinterleaver_auto_in_b_bits_id;
  wire [1:0] AXI4Deinterleaver_auto_in_b_bits_resp;
  wire [8:0] AXI4Deinterleaver_auto_in_b_bits_user;
  wire  AXI4Deinterleaver_auto_in_ar_ready;
  wire  AXI4Deinterleaver_auto_in_ar_valid;
  wire [3:0] AXI4Deinterleaver_auto_in_ar_bits_id;
  wire [30:0] AXI4Deinterleaver_auto_in_ar_bits_addr;
  wire [7:0] AXI4Deinterleaver_auto_in_ar_bits_len;
  wire [2:0] AXI4Deinterleaver_auto_in_ar_bits_size;
  wire [1:0] AXI4Deinterleaver_auto_in_ar_bits_burst;
  wire  AXI4Deinterleaver_auto_in_ar_bits_lock;
  wire [3:0] AXI4Deinterleaver_auto_in_ar_bits_cache;
  wire [2:0] AXI4Deinterleaver_auto_in_ar_bits_prot;
  wire [3:0] AXI4Deinterleaver_auto_in_ar_bits_qos;
  wire [8:0] AXI4Deinterleaver_auto_in_ar_bits_user;
  wire  AXI4Deinterleaver_auto_in_r_ready;
  wire  AXI4Deinterleaver_auto_in_r_valid;
  wire [3:0] AXI4Deinterleaver_auto_in_r_bits_id;
  wire [63:0] AXI4Deinterleaver_auto_in_r_bits_data;
  wire [1:0] AXI4Deinterleaver_auto_in_r_bits_resp;
  wire [8:0] AXI4Deinterleaver_auto_in_r_bits_user;
  wire  AXI4Deinterleaver_auto_in_r_bits_last;
  wire  AXI4Deinterleaver_auto_out_aw_ready;
  wire  AXI4Deinterleaver_auto_out_aw_valid;
  wire [3:0] AXI4Deinterleaver_auto_out_aw_bits_id;
  wire [30:0] AXI4Deinterleaver_auto_out_aw_bits_addr;
  wire [7:0] AXI4Deinterleaver_auto_out_aw_bits_len;
  wire [2:0] AXI4Deinterleaver_auto_out_aw_bits_size;
  wire [1:0] AXI4Deinterleaver_auto_out_aw_bits_burst;
  wire  AXI4Deinterleaver_auto_out_aw_bits_lock;
  wire [3:0] AXI4Deinterleaver_auto_out_aw_bits_cache;
  wire [2:0] AXI4Deinterleaver_auto_out_aw_bits_prot;
  wire [3:0] AXI4Deinterleaver_auto_out_aw_bits_qos;
  wire [8:0] AXI4Deinterleaver_auto_out_aw_bits_user;
  wire  AXI4Deinterleaver_auto_out_w_ready;
  wire  AXI4Deinterleaver_auto_out_w_valid;
  wire [63:0] AXI4Deinterleaver_auto_out_w_bits_data;
  wire [7:0] AXI4Deinterleaver_auto_out_w_bits_strb;
  wire  AXI4Deinterleaver_auto_out_w_bits_last;
  wire  AXI4Deinterleaver_auto_out_b_ready;
  wire  AXI4Deinterleaver_auto_out_b_valid;
  wire [3:0] AXI4Deinterleaver_auto_out_b_bits_id;
  wire [1:0] AXI4Deinterleaver_auto_out_b_bits_resp;
  wire [8:0] AXI4Deinterleaver_auto_out_b_bits_user;
  wire  AXI4Deinterleaver_auto_out_ar_ready;
  wire  AXI4Deinterleaver_auto_out_ar_valid;
  wire [3:0] AXI4Deinterleaver_auto_out_ar_bits_id;
  wire [30:0] AXI4Deinterleaver_auto_out_ar_bits_addr;
  wire [7:0] AXI4Deinterleaver_auto_out_ar_bits_len;
  wire [2:0] AXI4Deinterleaver_auto_out_ar_bits_size;
  wire [1:0] AXI4Deinterleaver_auto_out_ar_bits_burst;
  wire  AXI4Deinterleaver_auto_out_ar_bits_lock;
  wire [3:0] AXI4Deinterleaver_auto_out_ar_bits_cache;
  wire [2:0] AXI4Deinterleaver_auto_out_ar_bits_prot;
  wire [3:0] AXI4Deinterleaver_auto_out_ar_bits_qos;
  wire [8:0] AXI4Deinterleaver_auto_out_ar_bits_user;
  wire  AXI4Deinterleaver_auto_out_r_ready;
  wire  AXI4Deinterleaver_auto_out_r_valid;
  wire [3:0] AXI4Deinterleaver_auto_out_r_bits_id;
  wire [63:0] AXI4Deinterleaver_auto_out_r_bits_data;
  wire [1:0] AXI4Deinterleaver_auto_out_r_bits_resp;
  wire [8:0] AXI4Deinterleaver_auto_out_r_bits_user;
  wire  AXI4Deinterleaver_auto_out_r_bits_last;
  wire  AXI4IdIndexer_auto_in_aw_ready;
  wire  AXI4IdIndexer_auto_in_aw_valid;
  wire [2:0] AXI4IdIndexer_auto_in_aw_bits_id;
  wire [30:0] AXI4IdIndexer_auto_in_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_auto_in_aw_bits_len;
  wire [2:0] AXI4IdIndexer_auto_in_aw_bits_size;
  wire [1:0] AXI4IdIndexer_auto_in_aw_bits_burst;
  wire  AXI4IdIndexer_auto_in_aw_bits_lock;
  wire [3:0] AXI4IdIndexer_auto_in_aw_bits_cache;
  wire [2:0] AXI4IdIndexer_auto_in_aw_bits_prot;
  wire [3:0] AXI4IdIndexer_auto_in_aw_bits_qos;
  wire [8:0] AXI4IdIndexer_auto_in_aw_bits_user;
  wire  AXI4IdIndexer_auto_in_w_ready;
  wire  AXI4IdIndexer_auto_in_w_valid;
  wire [63:0] AXI4IdIndexer_auto_in_w_bits_data;
  wire [7:0] AXI4IdIndexer_auto_in_w_bits_strb;
  wire  AXI4IdIndexer_auto_in_w_bits_last;
  wire  AXI4IdIndexer_auto_in_b_ready;
  wire  AXI4IdIndexer_auto_in_b_valid;
  wire [2:0] AXI4IdIndexer_auto_in_b_bits_id;
  wire [1:0] AXI4IdIndexer_auto_in_b_bits_resp;
  wire [8:0] AXI4IdIndexer_auto_in_b_bits_user;
  wire  AXI4IdIndexer_auto_in_ar_ready;
  wire  AXI4IdIndexer_auto_in_ar_valid;
  wire [2:0] AXI4IdIndexer_auto_in_ar_bits_id;
  wire [30:0] AXI4IdIndexer_auto_in_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_auto_in_ar_bits_len;
  wire [2:0] AXI4IdIndexer_auto_in_ar_bits_size;
  wire [1:0] AXI4IdIndexer_auto_in_ar_bits_burst;
  wire  AXI4IdIndexer_auto_in_ar_bits_lock;
  wire [3:0] AXI4IdIndexer_auto_in_ar_bits_cache;
  wire [2:0] AXI4IdIndexer_auto_in_ar_bits_prot;
  wire [3:0] AXI4IdIndexer_auto_in_ar_bits_qos;
  wire [8:0] AXI4IdIndexer_auto_in_ar_bits_user;
  wire  AXI4IdIndexer_auto_in_r_ready;
  wire  AXI4IdIndexer_auto_in_r_valid;
  wire [2:0] AXI4IdIndexer_auto_in_r_bits_id;
  wire [63:0] AXI4IdIndexer_auto_in_r_bits_data;
  wire [1:0] AXI4IdIndexer_auto_in_r_bits_resp;
  wire [8:0] AXI4IdIndexer_auto_in_r_bits_user;
  wire  AXI4IdIndexer_auto_in_r_bits_last;
  wire  AXI4IdIndexer_auto_out_aw_ready;
  wire  AXI4IdIndexer_auto_out_aw_valid;
  wire [3:0] AXI4IdIndexer_auto_out_aw_bits_id;
  wire [30:0] AXI4IdIndexer_auto_out_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_auto_out_aw_bits_len;
  wire [2:0] AXI4IdIndexer_auto_out_aw_bits_size;
  wire [1:0] AXI4IdIndexer_auto_out_aw_bits_burst;
  wire  AXI4IdIndexer_auto_out_aw_bits_lock;
  wire [3:0] AXI4IdIndexer_auto_out_aw_bits_cache;
  wire [2:0] AXI4IdIndexer_auto_out_aw_bits_prot;
  wire [3:0] AXI4IdIndexer_auto_out_aw_bits_qos;
  wire [8:0] AXI4IdIndexer_auto_out_aw_bits_user;
  wire  AXI4IdIndexer_auto_out_w_ready;
  wire  AXI4IdIndexer_auto_out_w_valid;
  wire [63:0] AXI4IdIndexer_auto_out_w_bits_data;
  wire [7:0] AXI4IdIndexer_auto_out_w_bits_strb;
  wire  AXI4IdIndexer_auto_out_w_bits_last;
  wire  AXI4IdIndexer_auto_out_b_ready;
  wire  AXI4IdIndexer_auto_out_b_valid;
  wire [3:0] AXI4IdIndexer_auto_out_b_bits_id;
  wire [1:0] AXI4IdIndexer_auto_out_b_bits_resp;
  wire [8:0] AXI4IdIndexer_auto_out_b_bits_user;
  wire  AXI4IdIndexer_auto_out_ar_ready;
  wire  AXI4IdIndexer_auto_out_ar_valid;
  wire [3:0] AXI4IdIndexer_auto_out_ar_bits_id;
  wire [30:0] AXI4IdIndexer_auto_out_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_auto_out_ar_bits_len;
  wire [2:0] AXI4IdIndexer_auto_out_ar_bits_size;
  wire [1:0] AXI4IdIndexer_auto_out_ar_bits_burst;
  wire  AXI4IdIndexer_auto_out_ar_bits_lock;
  wire [3:0] AXI4IdIndexer_auto_out_ar_bits_cache;
  wire [2:0] AXI4IdIndexer_auto_out_ar_bits_prot;
  wire [3:0] AXI4IdIndexer_auto_out_ar_bits_qos;
  wire [8:0] AXI4IdIndexer_auto_out_ar_bits_user;
  wire  AXI4IdIndexer_auto_out_r_ready;
  wire  AXI4IdIndexer_auto_out_r_valid;
  wire [3:0] AXI4IdIndexer_auto_out_r_bits_id;
  wire [63:0] AXI4IdIndexer_auto_out_r_bits_data;
  wire [1:0] AXI4IdIndexer_auto_out_r_bits_resp;
  wire [8:0] AXI4IdIndexer_auto_out_r_bits_user;
  wire  AXI4IdIndexer_auto_out_r_bits_last;
  wire  TLToAXI4_clock;
  wire  TLToAXI4_reset;
  wire  TLToAXI4_auto_in_a_ready;
  wire  TLToAXI4_auto_in_a_valid;
  wire [2:0] TLToAXI4_auto_in_a_bits_opcode;
  wire [3:0] TLToAXI4_auto_in_a_bits_size;
  wire [4:0] TLToAXI4_auto_in_a_bits_source;
  wire [30:0] TLToAXI4_auto_in_a_bits_address;
  wire [7:0] TLToAXI4_auto_in_a_bits_mask;
  wire [63:0] TLToAXI4_auto_in_a_bits_data;
  wire  TLToAXI4_auto_in_d_ready;
  wire  TLToAXI4_auto_in_d_valid;
  wire [2:0] TLToAXI4_auto_in_d_bits_opcode;
  wire [3:0] TLToAXI4_auto_in_d_bits_size;
  wire [4:0] TLToAXI4_auto_in_d_bits_source;
  wire [63:0] TLToAXI4_auto_in_d_bits_data;
  wire  TLToAXI4_auto_in_d_bits_error;
  wire  TLToAXI4_auto_out_aw_ready;
  wire  TLToAXI4_auto_out_aw_valid;
  wire [2:0] TLToAXI4_auto_out_aw_bits_id;
  wire [30:0] TLToAXI4_auto_out_aw_bits_addr;
  wire [7:0] TLToAXI4_auto_out_aw_bits_len;
  wire [2:0] TLToAXI4_auto_out_aw_bits_size;
  wire [1:0] TLToAXI4_auto_out_aw_bits_burst;
  wire  TLToAXI4_auto_out_aw_bits_lock;
  wire [3:0] TLToAXI4_auto_out_aw_bits_cache;
  wire [2:0] TLToAXI4_auto_out_aw_bits_prot;
  wire [3:0] TLToAXI4_auto_out_aw_bits_qos;
  wire [8:0] TLToAXI4_auto_out_aw_bits_user;
  wire  TLToAXI4_auto_out_w_ready;
  wire  TLToAXI4_auto_out_w_valid;
  wire [63:0] TLToAXI4_auto_out_w_bits_data;
  wire [7:0] TLToAXI4_auto_out_w_bits_strb;
  wire  TLToAXI4_auto_out_w_bits_last;
  wire  TLToAXI4_auto_out_b_ready;
  wire  TLToAXI4_auto_out_b_valid;
  wire [2:0] TLToAXI4_auto_out_b_bits_id;
  wire [1:0] TLToAXI4_auto_out_b_bits_resp;
  wire [8:0] TLToAXI4_auto_out_b_bits_user;
  wire  TLToAXI4_auto_out_ar_ready;
  wire  TLToAXI4_auto_out_ar_valid;
  wire [2:0] TLToAXI4_auto_out_ar_bits_id;
  wire [30:0] TLToAXI4_auto_out_ar_bits_addr;
  wire [7:0] TLToAXI4_auto_out_ar_bits_len;
  wire [2:0] TLToAXI4_auto_out_ar_bits_size;
  wire [1:0] TLToAXI4_auto_out_ar_bits_burst;
  wire  TLToAXI4_auto_out_ar_bits_lock;
  wire [3:0] TLToAXI4_auto_out_ar_bits_cache;
  wire [2:0] TLToAXI4_auto_out_ar_bits_prot;
  wire [3:0] TLToAXI4_auto_out_ar_bits_qos;
  wire [8:0] TLToAXI4_auto_out_ar_bits_user;
  wire  TLToAXI4_auto_out_r_ready;
  wire  TLToAXI4_auto_out_r_valid;
  wire [2:0] TLToAXI4_auto_out_r_bits_id;
  wire [63:0] TLToAXI4_auto_out_r_bits_data;
  wire [1:0] TLToAXI4_auto_out_r_bits_resp;
  wire [8:0] TLToAXI4_auto_out_r_bits_user;
  wire  TLToAXI4_auto_out_r_bits_last;
  wire  SystemBus_TLBuffer_clock;
  wire  SystemBus_TLBuffer_reset;
  wire  SystemBus_TLBuffer_auto_in_a_ready;
  wire  SystemBus_TLBuffer_auto_in_a_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_a_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_in_a_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_in_a_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_a_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_in_a_bits_address;
  wire [7:0] SystemBus_TLBuffer_auto_in_a_bits_mask;
  wire [63:0] SystemBus_TLBuffer_auto_in_a_bits_data;
  wire  SystemBus_TLBuffer_auto_in_d_ready;
  wire  SystemBus_TLBuffer_auto_in_d_valid;
  wire [2:0] SystemBus_TLBuffer_auto_in_d_bits_opcode;
  wire [3:0] SystemBus_TLBuffer_auto_in_d_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_in_d_bits_source;
  wire [63:0] SystemBus_TLBuffer_auto_in_d_bits_data;
  wire  SystemBus_TLBuffer_auto_in_d_bits_error;
  wire  SystemBus_TLBuffer_auto_out_a_ready;
  wire  SystemBus_TLBuffer_auto_out_a_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_a_bits_opcode;
  wire [2:0] SystemBus_TLBuffer_auto_out_a_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_a_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_a_bits_source;
  wire [31:0] SystemBus_TLBuffer_auto_out_a_bits_address;
  wire [7:0] SystemBus_TLBuffer_auto_out_a_bits_mask;
  wire [63:0] SystemBus_TLBuffer_auto_out_a_bits_data;
  wire  SystemBus_TLBuffer_auto_out_d_ready;
  wire  SystemBus_TLBuffer_auto_out_d_valid;
  wire [2:0] SystemBus_TLBuffer_auto_out_d_bits_opcode;
  wire [1:0] SystemBus_TLBuffer_auto_out_d_bits_param;
  wire [3:0] SystemBus_TLBuffer_auto_out_d_bits_size;
  wire [3:0] SystemBus_TLBuffer_auto_out_d_bits_source;
  wire [2:0] SystemBus_TLBuffer_auto_out_d_bits_sink;
  wire [63:0] SystemBus_TLBuffer_auto_out_d_bits_data;
  wire  SystemBus_TLBuffer_auto_out_d_bits_error;
  wire  SystemBus_TLWidthWidget_auto_in_a_ready;
  wire  SystemBus_TLWidthWidget_auto_in_a_valid;
  wire [2:0] SystemBus_TLWidthWidget_auto_in_a_bits_opcode;
  wire [2:0] SystemBus_TLWidthWidget_auto_in_a_bits_param;
  wire [3:0] SystemBus_TLWidthWidget_auto_in_a_bits_size;
  wire [3:0] SystemBus_TLWidthWidget_auto_in_a_bits_source;
  wire [31:0] SystemBus_TLWidthWidget_auto_in_a_bits_address;
  wire [7:0] SystemBus_TLWidthWidget_auto_in_a_bits_mask;
  wire [63:0] SystemBus_TLWidthWidget_auto_in_a_bits_data;
  wire  SystemBus_TLWidthWidget_auto_in_d_ready;
  wire  SystemBus_TLWidthWidget_auto_in_d_valid;
  wire [2:0] SystemBus_TLWidthWidget_auto_in_d_bits_opcode;
  wire [3:0] SystemBus_TLWidthWidget_auto_in_d_bits_size;
  wire [3:0] SystemBus_TLWidthWidget_auto_in_d_bits_source;
  wire [63:0] SystemBus_TLWidthWidget_auto_in_d_bits_data;
  wire  SystemBus_TLWidthWidget_auto_in_d_bits_error;
  wire  SystemBus_TLWidthWidget_auto_out_a_ready;
  wire  SystemBus_TLWidthWidget_auto_out_a_valid;
  wire [2:0] SystemBus_TLWidthWidget_auto_out_a_bits_opcode;
  wire [2:0] SystemBus_TLWidthWidget_auto_out_a_bits_param;
  wire [3:0] SystemBus_TLWidthWidget_auto_out_a_bits_size;
  wire [3:0] SystemBus_TLWidthWidget_auto_out_a_bits_source;
  wire [31:0] SystemBus_TLWidthWidget_auto_out_a_bits_address;
  wire [7:0] SystemBus_TLWidthWidget_auto_out_a_bits_mask;
  wire [63:0] SystemBus_TLWidthWidget_auto_out_a_bits_data;
  wire  SystemBus_TLWidthWidget_auto_out_d_ready;
  wire  SystemBus_TLWidthWidget_auto_out_d_valid;
  wire [2:0] SystemBus_TLWidthWidget_auto_out_d_bits_opcode;
  wire [3:0] SystemBus_TLWidthWidget_auto_out_d_bits_size;
  wire [3:0] SystemBus_TLWidthWidget_auto_out_d_bits_source;
  wire [63:0] SystemBus_TLWidthWidget_auto_out_d_bits_data;
  wire  SystemBus_TLWidthWidget_auto_out_d_bits_error;
  wire  AXI4ToTL_clock;
  wire  AXI4ToTL_reset;
  wire  AXI4ToTL_auto_in_aw_ready;
  wire  AXI4ToTL_auto_in_aw_valid;
  wire  AXI4ToTL_auto_in_aw_bits_id;
  wire [31:0] AXI4ToTL_auto_in_aw_bits_addr;
  wire [7:0] AXI4ToTL_auto_in_aw_bits_len;
  wire [2:0] AXI4ToTL_auto_in_aw_bits_size;
  wire  AXI4ToTL_auto_in_w_ready;
  wire  AXI4ToTL_auto_in_w_valid;
  wire [63:0] AXI4ToTL_auto_in_w_bits_data;
  wire [7:0] AXI4ToTL_auto_in_w_bits_strb;
  wire  AXI4ToTL_auto_in_w_bits_last;
  wire  AXI4ToTL_auto_in_b_ready;
  wire  AXI4ToTL_auto_in_b_valid;
  wire  AXI4ToTL_auto_in_b_bits_id;
  wire [1:0] AXI4ToTL_auto_in_b_bits_resp;
  wire  AXI4ToTL_auto_in_ar_ready;
  wire  AXI4ToTL_auto_in_ar_valid;
  wire  AXI4ToTL_auto_in_ar_bits_id;
  wire [31:0] AXI4ToTL_auto_in_ar_bits_addr;
  wire [7:0] AXI4ToTL_auto_in_ar_bits_len;
  wire [2:0] AXI4ToTL_auto_in_ar_bits_size;
  wire  AXI4ToTL_auto_in_r_ready;
  wire  AXI4ToTL_auto_in_r_valid;
  wire  AXI4ToTL_auto_in_r_bits_id;
  wire [63:0] AXI4ToTL_auto_in_r_bits_data;
  wire [1:0] AXI4ToTL_auto_in_r_bits_resp;
  wire  AXI4ToTL_auto_in_r_bits_last;
  wire  AXI4ToTL_auto_out_a_ready;
  wire  AXI4ToTL_auto_out_a_valid;
  wire [2:0] AXI4ToTL_auto_out_a_bits_opcode;
  wire [2:0] AXI4ToTL_auto_out_a_bits_param;
  wire [3:0] AXI4ToTL_auto_out_a_bits_size;
  wire [3:0] AXI4ToTL_auto_out_a_bits_source;
  wire [31:0] AXI4ToTL_auto_out_a_bits_address;
  wire [7:0] AXI4ToTL_auto_out_a_bits_mask;
  wire [63:0] AXI4ToTL_auto_out_a_bits_data;
  wire  AXI4ToTL_auto_out_d_ready;
  wire  AXI4ToTL_auto_out_d_valid;
  wire [2:0] AXI4ToTL_auto_out_d_bits_opcode;
  wire [3:0] AXI4ToTL_auto_out_d_bits_size;
  wire [3:0] AXI4ToTL_auto_out_d_bits_source;
  wire [63:0] AXI4ToTL_auto_out_d_bits_data;
  wire  AXI4ToTL_auto_out_d_bits_error;
  wire  AXI4UserYanker_1_clock;
  wire  AXI4UserYanker_1_reset;
  wire  AXI4UserYanker_1_auto_in_aw_ready;
  wire  AXI4UserYanker_1_auto_in_aw_valid;
  wire  AXI4UserYanker_1_auto_in_aw_bits_id;
  wire [31:0] AXI4UserYanker_1_auto_in_aw_bits_addr;
  wire [7:0] AXI4UserYanker_1_auto_in_aw_bits_len;
  wire [2:0] AXI4UserYanker_1_auto_in_aw_bits_size;
  wire [7:0] AXI4UserYanker_1_auto_in_aw_bits_user;
  wire  AXI4UserYanker_1_auto_in_w_ready;
  wire  AXI4UserYanker_1_auto_in_w_valid;
  wire [63:0] AXI4UserYanker_1_auto_in_w_bits_data;
  wire [7:0] AXI4UserYanker_1_auto_in_w_bits_strb;
  wire  AXI4UserYanker_1_auto_in_w_bits_last;
  wire  AXI4UserYanker_1_auto_in_b_ready;
  wire  AXI4UserYanker_1_auto_in_b_valid;
  wire  AXI4UserYanker_1_auto_in_b_bits_id;
  wire [1:0] AXI4UserYanker_1_auto_in_b_bits_resp;
  wire [7:0] AXI4UserYanker_1_auto_in_b_bits_user;
  wire  AXI4UserYanker_1_auto_in_ar_ready;
  wire  AXI4UserYanker_1_auto_in_ar_valid;
  wire  AXI4UserYanker_1_auto_in_ar_bits_id;
  wire [31:0] AXI4UserYanker_1_auto_in_ar_bits_addr;
  wire [7:0] AXI4UserYanker_1_auto_in_ar_bits_len;
  wire [2:0] AXI4UserYanker_1_auto_in_ar_bits_size;
  wire [7:0] AXI4UserYanker_1_auto_in_ar_bits_user;
  wire  AXI4UserYanker_1_auto_in_r_ready;
  wire  AXI4UserYanker_1_auto_in_r_valid;
  wire  AXI4UserYanker_1_auto_in_r_bits_id;
  wire [63:0] AXI4UserYanker_1_auto_in_r_bits_data;
  wire [1:0] AXI4UserYanker_1_auto_in_r_bits_resp;
  wire [7:0] AXI4UserYanker_1_auto_in_r_bits_user;
  wire  AXI4UserYanker_1_auto_in_r_bits_last;
  wire  AXI4UserYanker_1_auto_out_aw_ready;
  wire  AXI4UserYanker_1_auto_out_aw_valid;
  wire  AXI4UserYanker_1_auto_out_aw_bits_id;
  wire [31:0] AXI4UserYanker_1_auto_out_aw_bits_addr;
  wire [7:0] AXI4UserYanker_1_auto_out_aw_bits_len;
  wire [2:0] AXI4UserYanker_1_auto_out_aw_bits_size;
  wire  AXI4UserYanker_1_auto_out_w_ready;
  wire  AXI4UserYanker_1_auto_out_w_valid;
  wire [63:0] AXI4UserYanker_1_auto_out_w_bits_data;
  wire [7:0] AXI4UserYanker_1_auto_out_w_bits_strb;
  wire  AXI4UserYanker_1_auto_out_w_bits_last;
  wire  AXI4UserYanker_1_auto_out_b_ready;
  wire  AXI4UserYanker_1_auto_out_b_valid;
  wire  AXI4UserYanker_1_auto_out_b_bits_id;
  wire [1:0] AXI4UserYanker_1_auto_out_b_bits_resp;
  wire  AXI4UserYanker_1_auto_out_ar_ready;
  wire  AXI4UserYanker_1_auto_out_ar_valid;
  wire  AXI4UserYanker_1_auto_out_ar_bits_id;
  wire [31:0] AXI4UserYanker_1_auto_out_ar_bits_addr;
  wire [7:0] AXI4UserYanker_1_auto_out_ar_bits_len;
  wire [2:0] AXI4UserYanker_1_auto_out_ar_bits_size;
  wire  AXI4UserYanker_1_auto_out_r_ready;
  wire  AXI4UserYanker_1_auto_out_r_valid;
  wire  AXI4UserYanker_1_auto_out_r_bits_id;
  wire [63:0] AXI4UserYanker_1_auto_out_r_bits_data;
  wire [1:0] AXI4UserYanker_1_auto_out_r_bits_resp;
  wire  AXI4UserYanker_1_auto_out_r_bits_last;
  wire  AXI4Fragmenter_clock;
  wire  AXI4Fragmenter_reset;
  wire  AXI4Fragmenter_auto_in_aw_ready;
  wire  AXI4Fragmenter_auto_in_aw_valid;
  wire  AXI4Fragmenter_auto_in_aw_bits_id;
  wire [31:0] AXI4Fragmenter_auto_in_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_aw_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_aw_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_aw_bits_burst;
  wire [6:0] AXI4Fragmenter_auto_in_aw_bits_user;
  wire  AXI4Fragmenter_auto_in_w_ready;
  wire  AXI4Fragmenter_auto_in_w_valid;
  wire [63:0] AXI4Fragmenter_auto_in_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_in_w_bits_strb;
  wire  AXI4Fragmenter_auto_in_w_bits_last;
  wire  AXI4Fragmenter_auto_in_b_ready;
  wire  AXI4Fragmenter_auto_in_b_valid;
  wire  AXI4Fragmenter_auto_in_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_in_b_bits_resp;
  wire [6:0] AXI4Fragmenter_auto_in_b_bits_user;
  wire  AXI4Fragmenter_auto_in_ar_ready;
  wire  AXI4Fragmenter_auto_in_ar_valid;
  wire  AXI4Fragmenter_auto_in_ar_bits_id;
  wire [31:0] AXI4Fragmenter_auto_in_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_ar_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_ar_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_ar_bits_burst;
  wire [6:0] AXI4Fragmenter_auto_in_ar_bits_user;
  wire  AXI4Fragmenter_auto_in_r_ready;
  wire  AXI4Fragmenter_auto_in_r_valid;
  wire  AXI4Fragmenter_auto_in_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_in_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_in_r_bits_resp;
  wire [6:0] AXI4Fragmenter_auto_in_r_bits_user;
  wire  AXI4Fragmenter_auto_in_r_bits_last;
  wire  AXI4Fragmenter_auto_out_aw_ready;
  wire  AXI4Fragmenter_auto_out_aw_valid;
  wire  AXI4Fragmenter_auto_out_aw_bits_id;
  wire [31:0] AXI4Fragmenter_auto_out_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_out_aw_bits_len;
  wire [2:0] AXI4Fragmenter_auto_out_aw_bits_size;
  wire [7:0] AXI4Fragmenter_auto_out_aw_bits_user;
  wire  AXI4Fragmenter_auto_out_w_ready;
  wire  AXI4Fragmenter_auto_out_w_valid;
  wire [63:0] AXI4Fragmenter_auto_out_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_out_w_bits_strb;
  wire  AXI4Fragmenter_auto_out_w_bits_last;
  wire  AXI4Fragmenter_auto_out_b_ready;
  wire  AXI4Fragmenter_auto_out_b_valid;
  wire  AXI4Fragmenter_auto_out_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_out_b_bits_resp;
  wire [7:0] AXI4Fragmenter_auto_out_b_bits_user;
  wire  AXI4Fragmenter_auto_out_ar_ready;
  wire  AXI4Fragmenter_auto_out_ar_valid;
  wire  AXI4Fragmenter_auto_out_ar_bits_id;
  wire [31:0] AXI4Fragmenter_auto_out_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_out_ar_bits_len;
  wire [2:0] AXI4Fragmenter_auto_out_ar_bits_size;
  wire [7:0] AXI4Fragmenter_auto_out_ar_bits_user;
  wire  AXI4Fragmenter_auto_out_r_ready;
  wire  AXI4Fragmenter_auto_out_r_valid;
  wire  AXI4Fragmenter_auto_out_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_out_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_out_r_bits_resp;
  wire [7:0] AXI4Fragmenter_auto_out_r_bits_user;
  wire  AXI4Fragmenter_auto_out_r_bits_last;
  wire  AXI4IdIndexer_1_auto_in_aw_ready;
  wire  AXI4IdIndexer_1_auto_in_aw_valid;
  wire [7:0] AXI4IdIndexer_1_auto_in_aw_bits_id;
  wire [31:0] AXI4IdIndexer_1_auto_in_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_1_auto_in_aw_bits_len;
  wire [2:0] AXI4IdIndexer_1_auto_in_aw_bits_size;
  wire [1:0] AXI4IdIndexer_1_auto_in_aw_bits_burst;
  wire  AXI4IdIndexer_1_auto_in_w_ready;
  wire  AXI4IdIndexer_1_auto_in_w_valid;
  wire [63:0] AXI4IdIndexer_1_auto_in_w_bits_data;
  wire [7:0] AXI4IdIndexer_1_auto_in_w_bits_strb;
  wire  AXI4IdIndexer_1_auto_in_w_bits_last;
  wire  AXI4IdIndexer_1_auto_in_b_ready;
  wire  AXI4IdIndexer_1_auto_in_b_valid;
  wire [7:0] AXI4IdIndexer_1_auto_in_b_bits_id;
  wire [1:0] AXI4IdIndexer_1_auto_in_b_bits_resp;
  wire  AXI4IdIndexer_1_auto_in_ar_ready;
  wire  AXI4IdIndexer_1_auto_in_ar_valid;
  wire [7:0] AXI4IdIndexer_1_auto_in_ar_bits_id;
  wire [31:0] AXI4IdIndexer_1_auto_in_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_1_auto_in_ar_bits_len;
  wire [2:0] AXI4IdIndexer_1_auto_in_ar_bits_size;
  wire [1:0] AXI4IdIndexer_1_auto_in_ar_bits_burst;
  wire  AXI4IdIndexer_1_auto_in_r_ready;
  wire  AXI4IdIndexer_1_auto_in_r_valid;
  wire [7:0] AXI4IdIndexer_1_auto_in_r_bits_id;
  wire [63:0] AXI4IdIndexer_1_auto_in_r_bits_data;
  wire [1:0] AXI4IdIndexer_1_auto_in_r_bits_resp;
  wire  AXI4IdIndexer_1_auto_in_r_bits_last;
  wire  AXI4IdIndexer_1_auto_out_aw_ready;
  wire  AXI4IdIndexer_1_auto_out_aw_valid;
  wire  AXI4IdIndexer_1_auto_out_aw_bits_id;
  wire [31:0] AXI4IdIndexer_1_auto_out_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_1_auto_out_aw_bits_len;
  wire [2:0] AXI4IdIndexer_1_auto_out_aw_bits_size;
  wire [1:0] AXI4IdIndexer_1_auto_out_aw_bits_burst;
  wire [6:0] AXI4IdIndexer_1_auto_out_aw_bits_user;
  wire  AXI4IdIndexer_1_auto_out_w_ready;
  wire  AXI4IdIndexer_1_auto_out_w_valid;
  wire [63:0] AXI4IdIndexer_1_auto_out_w_bits_data;
  wire [7:0] AXI4IdIndexer_1_auto_out_w_bits_strb;
  wire  AXI4IdIndexer_1_auto_out_w_bits_last;
  wire  AXI4IdIndexer_1_auto_out_b_ready;
  wire  AXI4IdIndexer_1_auto_out_b_valid;
  wire  AXI4IdIndexer_1_auto_out_b_bits_id;
  wire [1:0] AXI4IdIndexer_1_auto_out_b_bits_resp;
  wire [6:0] AXI4IdIndexer_1_auto_out_b_bits_user;
  wire  AXI4IdIndexer_1_auto_out_ar_ready;
  wire  AXI4IdIndexer_1_auto_out_ar_valid;
  wire  AXI4IdIndexer_1_auto_out_ar_bits_id;
  wire [31:0] AXI4IdIndexer_1_auto_out_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_1_auto_out_ar_bits_len;
  wire [2:0] AXI4IdIndexer_1_auto_out_ar_bits_size;
  wire [1:0] AXI4IdIndexer_1_auto_out_ar_bits_burst;
  wire [6:0] AXI4IdIndexer_1_auto_out_ar_bits_user;
  wire  AXI4IdIndexer_1_auto_out_r_ready;
  wire  AXI4IdIndexer_1_auto_out_r_valid;
  wire  AXI4IdIndexer_1_auto_out_r_bits_id;
  wire [63:0] AXI4IdIndexer_1_auto_out_r_bits_data;
  wire [1:0] AXI4IdIndexer_1_auto_out_r_bits_resp;
  wire [6:0] AXI4IdIndexer_1_auto_out_r_bits_user;
  wire  AXI4IdIndexer_1_auto_out_r_bits_last;
  wire  bootrom_auto_in_a_ready;
  wire  bootrom_auto_in_a_valid;
  wire [1:0] bootrom_auto_in_a_bits_size;
  wire [8:0] bootrom_auto_in_a_bits_source;
  wire [16:0] bootrom_auto_in_a_bits_address;
  wire  bootrom_auto_in_d_ready;
  wire  bootrom_auto_in_d_valid;
  wire [1:0] bootrom_auto_in_d_bits_size;
  wire [8:0] bootrom_auto_in_d_bits_source;
  wire [63:0] bootrom_auto_in_d_bits_data;
  wire  error_clock;
  wire  error_reset;
  wire  error_auto_in_a_ready;
  wire  error_auto_in_a_valid;
  wire [2:0] error_auto_in_a_bits_opcode;
  wire [3:0] error_auto_in_a_bits_size;
  wire [4:0] error_auto_in_a_bits_source;
  wire  error_auto_in_c_ready;
  wire  error_auto_in_c_valid;
  wire [2:0] error_auto_in_c_bits_opcode;
  wire [2:0] error_auto_in_c_bits_param;
  wire [3:0] error_auto_in_c_bits_size;
  wire [4:0] error_auto_in_c_bits_source;
  wire  error_auto_in_d_ready;
  wire  error_auto_in_d_valid;
  wire [2:0] error_auto_in_d_bits_opcode;
  wire [1:0] error_auto_in_d_bits_param;
  wire [3:0] error_auto_in_d_bits_size;
  wire [4:0] error_auto_in_d_bits_source;
  wire  error_auto_in_d_bits_sink;
  wire [63:0] error_auto_in_d_bits_data;
  wire  error_auto_in_d_bits_error;
  wire  _T_5_0;
  wire  _T_5_1;
  wire  _T_39_aw_ready;
  wire  _T_39_aw_valid;
  wire [3:0] _T_39_aw_bits_id;
  wire [31:0] _T_39_aw_bits_addr;
  wire [7:0] _T_39_aw_bits_len;
  wire [2:0] _T_39_aw_bits_size;
  wire [1:0] _T_39_aw_bits_burst;
  wire  _T_39_aw_bits_lock;
  wire [3:0] _T_39_aw_bits_cache;
  wire [2:0] _T_39_aw_bits_prot;
  wire [3:0] _T_39_aw_bits_qos;
  wire  _T_39_w_ready;
  wire  _T_39_w_valid;
  wire [63:0] _T_39_w_bits_data;
  wire [7:0] _T_39_w_bits_strb;
  wire  _T_39_w_bits_last;
  wire  _T_39_b_ready;
  wire  _T_39_b_valid;
  wire [3:0] _T_39_b_bits_id;
  wire [1:0] _T_39_b_bits_resp;
  wire  _T_39_ar_ready;
  wire  _T_39_ar_valid;
  wire [3:0] _T_39_ar_bits_id;
  wire [31:0] _T_39_ar_bits_addr;
  wire [7:0] _T_39_ar_bits_len;
  wire [2:0] _T_39_ar_bits_size;
  wire [1:0] _T_39_ar_bits_burst;
  wire  _T_39_ar_bits_lock;
  wire [3:0] _T_39_ar_bits_cache;
  wire [2:0] _T_39_ar_bits_prot;
  wire [3:0] _T_39_ar_bits_qos;
  wire  _T_39_r_ready;
  wire  _T_39_r_valid;
  wire [3:0] _T_39_r_bits_id;
  wire [63:0] _T_39_r_bits_data;
  wire [1:0] _T_39_r_bits_resp;
  wire  _T_39_r_bits_last;
  wire  _T_97_aw_ready;
  wire  _T_97_aw_valid;
  wire [3:0] _T_97_aw_bits_id;
  wire [30:0] _T_97_aw_bits_addr;
  wire [7:0] _T_97_aw_bits_len;
  wire [2:0] _T_97_aw_bits_size;
  wire [1:0] _T_97_aw_bits_burst;
  wire  _T_97_aw_bits_lock;
  wire [3:0] _T_97_aw_bits_cache;
  wire [2:0] _T_97_aw_bits_prot;
  wire [3:0] _T_97_aw_bits_qos;
  wire  _T_97_w_ready;
  wire  _T_97_w_valid;
  wire [63:0] _T_97_w_bits_data;
  wire [7:0] _T_97_w_bits_strb;
  wire  _T_97_w_bits_last;
  wire  _T_97_b_ready;
  wire  _T_97_b_valid;
  wire [3:0] _T_97_b_bits_id;
  wire [1:0] _T_97_b_bits_resp;
  wire  _T_97_ar_ready;
  wire  _T_97_ar_valid;
  wire [3:0] _T_97_ar_bits_id;
  wire [30:0] _T_97_ar_bits_addr;
  wire [7:0] _T_97_ar_bits_len;
  wire [2:0] _T_97_ar_bits_size;
  wire [1:0] _T_97_ar_bits_burst;
  wire  _T_97_ar_bits_lock;
  wire [3:0] _T_97_ar_bits_cache;
  wire [2:0] _T_97_ar_bits_prot;
  wire [3:0] _T_97_ar_bits_qos;
  wire  _T_97_r_ready;
  wire  _T_97_r_valid;
  wire [3:0] _T_97_r_bits_id;
  wire [63:0] _T_97_r_bits_data;
  wire [1:0] _T_97_r_bits_resp;
  wire  _T_97_r_bits_last;
  wire  _T_155_aw_ready;
  wire  _T_155_aw_valid;
  wire [7:0] _T_155_aw_bits_id;
  wire [31:0] _T_155_aw_bits_addr;
  wire [7:0] _T_155_aw_bits_len;
  wire [2:0] _T_155_aw_bits_size;
  wire [1:0] _T_155_aw_bits_burst;
  wire  _T_155_w_ready;
  wire  _T_155_w_valid;
  wire [63:0] _T_155_w_bits_data;
  wire [7:0] _T_155_w_bits_strb;
  wire  _T_155_w_bits_last;
  wire  _T_155_b_ready;
  wire  _T_155_b_valid;
  wire [7:0] _T_155_b_bits_id;
  wire [1:0] _T_155_b_bits_resp;
  wire  _T_155_ar_ready;
  wire  _T_155_ar_valid;
  wire [7:0] _T_155_ar_bits_id;
  wire [31:0] _T_155_ar_bits_addr;
  wire [7:0] _T_155_ar_bits_len;
  wire [2:0] _T_155_ar_bits_size;
  wire [1:0] _T_155_ar_bits_burst;
  wire  _T_155_r_ready;
  wire  _T_155_r_valid;
  wire [7:0] _T_155_r_bits_id;
  wire [63:0] _T_155_r_bits_data;
  wire [1:0] _T_155_r_bits_resp;
  wire  _T_155_r_bits_last;
  wire  tile_inputs_0_clock;
  wire  tile_inputs_0_reset;
  reg [6:0] value;
  reg [31:0] _RAND_0;
  wire  int_rtc_tick;
  wire [7:0] _T_244;
  wire [6:0] _T_245;
  wire [6:0] _GEN_0;
  wire  _T_248;
  wire  _T_249;
  IntXbar IntXbar (
    .auto_int_in_0(IntXbar_auto_int_in_0),
    .auto_int_in_1(IntXbar_auto_int_in_1),
    .auto_int_out_0(IntXbar_auto_int_out_0),
    .auto_int_out_1(IntXbar_auto_int_out_1)
  );
  SystemBus_sbus sbus (
    .clock(sbus_clock),
    .reset(sbus_reset),
    .auto_SystemBusFromTiletile_anon_in_a_ready(sbus_auto_SystemBusFromTiletile_anon_in_a_ready),
    .auto_SystemBusFromTiletile_anon_in_a_valid(sbus_auto_SystemBusFromTiletile_anon_in_a_valid),
    .auto_SystemBusFromTiletile_anon_in_a_bits_opcode(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_opcode),
    .auto_SystemBusFromTiletile_anon_in_a_bits_param(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_param),
    .auto_SystemBusFromTiletile_anon_in_a_bits_size(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_size),
    .auto_SystemBusFromTiletile_anon_in_a_bits_source(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_source),
    .auto_SystemBusFromTiletile_anon_in_a_bits_address(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_address),
    .auto_SystemBusFromTiletile_anon_in_a_bits_mask(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_mask),
    .auto_SystemBusFromTiletile_anon_in_a_bits_data(sbus_auto_SystemBusFromTiletile_anon_in_a_bits_data),
    .auto_SystemBusFromTiletile_anon_in_b_ready(sbus_auto_SystemBusFromTiletile_anon_in_b_ready),
    .auto_SystemBusFromTiletile_anon_in_b_valid(sbus_auto_SystemBusFromTiletile_anon_in_b_valid),
    .auto_SystemBusFromTiletile_anon_in_b_bits_param(sbus_auto_SystemBusFromTiletile_anon_in_b_bits_param),
    .auto_SystemBusFromTiletile_anon_in_b_bits_size(sbus_auto_SystemBusFromTiletile_anon_in_b_bits_size),
    .auto_SystemBusFromTiletile_anon_in_b_bits_source(sbus_auto_SystemBusFromTiletile_anon_in_b_bits_source),
    .auto_SystemBusFromTiletile_anon_in_b_bits_address(sbus_auto_SystemBusFromTiletile_anon_in_b_bits_address),
    .auto_SystemBusFromTiletile_anon_in_c_ready(sbus_auto_SystemBusFromTiletile_anon_in_c_ready),
    .auto_SystemBusFromTiletile_anon_in_c_valid(sbus_auto_SystemBusFromTiletile_anon_in_c_valid),
    .auto_SystemBusFromTiletile_anon_in_c_bits_opcode(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_opcode),
    .auto_SystemBusFromTiletile_anon_in_c_bits_param(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_param),
    .auto_SystemBusFromTiletile_anon_in_c_bits_size(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_size),
    .auto_SystemBusFromTiletile_anon_in_c_bits_source(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_source),
    .auto_SystemBusFromTiletile_anon_in_c_bits_address(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_address),
    .auto_SystemBusFromTiletile_anon_in_c_bits_data(sbus_auto_SystemBusFromTiletile_anon_in_c_bits_data),
    .auto_SystemBusFromTiletile_anon_in_d_ready(sbus_auto_SystemBusFromTiletile_anon_in_d_ready),
    .auto_SystemBusFromTiletile_anon_in_d_valid(sbus_auto_SystemBusFromTiletile_anon_in_d_valid),
    .auto_SystemBusFromTiletile_anon_in_d_bits_opcode(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_opcode),
    .auto_SystemBusFromTiletile_anon_in_d_bits_param(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_param),
    .auto_SystemBusFromTiletile_anon_in_d_bits_size(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_size),
    .auto_SystemBusFromTiletile_anon_in_d_bits_source(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_source),
    .auto_SystemBusFromTiletile_anon_in_d_bits_sink(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_sink),
    .auto_SystemBusFromTiletile_anon_in_d_bits_data(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_data),
    .auto_SystemBusFromTiletile_anon_in_d_bits_error(sbus_auto_SystemBusFromTiletile_anon_in_d_bits_error),
    .auto_SystemBusFromTiletile_anon_in_e_ready(sbus_auto_SystemBusFromTiletile_anon_in_e_ready),
    .auto_SystemBusFromTiletile_anon_in_e_valid(sbus_auto_SystemBusFromTiletile_anon_in_e_valid),
    .auto_SystemBusFromTiletile_anon_in_e_bits_sink(sbus_auto_SystemBusFromTiletile_anon_in_e_bits_sink),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_ready(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_ready),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_valid(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_valid),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_opcode(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_opcode),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_param(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_param),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_size(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_size),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_source(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_source),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_address(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_address),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_mask(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_mask),
    .auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_data(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_data),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_ready(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_ready),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_valid(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_valid),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_opcode(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_opcode),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_param(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_param),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_size(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_size),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_source(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_source),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_sink(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_sink),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_data(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_data),
    .auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_error(sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_error),
    .auto_SystemBus_port_TLFIFOFixer_in_a_ready(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_ready),
    .auto_SystemBus_port_TLFIFOFixer_in_a_valid(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_valid),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_opcode(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_opcode),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_param(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_param),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_size(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_size),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_source(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_source),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_address(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_address),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_mask(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_mask),
    .auto_SystemBus_port_TLFIFOFixer_in_a_bits_data(sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_data),
    .auto_SystemBus_port_TLFIFOFixer_in_d_ready(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_ready),
    .auto_SystemBus_port_TLFIFOFixer_in_d_valid(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_valid),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_opcode(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_opcode),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_param(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_param),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_size(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_size),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_source(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_source),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_sink(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_sink),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_data(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_data),
    .auto_SystemBus_port_TLFIFOFixer_in_d_bits_error(sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_error),
    .auto_SystemBus_slave_TLWidthWidget_out_a_ready(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_ready),
    .auto_SystemBus_slave_TLWidthWidget_out_a_valid(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_valid),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_opcode(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_opcode),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_size(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_size),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_source(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_source),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_address(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_address),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_mask(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_mask),
    .auto_SystemBus_slave_TLWidthWidget_out_a_bits_data(sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_data),
    .auto_SystemBus_slave_TLWidthWidget_out_d_ready(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_ready),
    .auto_SystemBus_slave_TLWidthWidget_out_d_valid(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_valid),
    .auto_SystemBus_slave_TLWidthWidget_out_d_bits_opcode(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_opcode),
    .auto_SystemBus_slave_TLWidthWidget_out_d_bits_size(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_size),
    .auto_SystemBus_slave_TLWidthWidget_out_d_bits_source(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_source),
    .auto_SystemBus_slave_TLWidthWidget_out_d_bits_data(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_data),
    .auto_SystemBus_slave_TLWidthWidget_out_d_bits_error(sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_error),
    .auto_SystemBus_slave_TLBuffer_out_a_ready(sbus_auto_SystemBus_slave_TLBuffer_out_a_ready),
    .auto_SystemBus_slave_TLBuffer_out_a_valid(sbus_auto_SystemBus_slave_TLBuffer_out_a_valid),
    .auto_SystemBus_slave_TLBuffer_out_a_bits_opcode(sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_opcode),
    .auto_SystemBus_slave_TLBuffer_out_a_bits_size(sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_size),
    .auto_SystemBus_slave_TLBuffer_out_a_bits_source(sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_source),
    .auto_SystemBus_slave_TLBuffer_out_c_ready(sbus_auto_SystemBus_slave_TLBuffer_out_c_ready),
    .auto_SystemBus_slave_TLBuffer_out_c_valid(sbus_auto_SystemBus_slave_TLBuffer_out_c_valid),
    .auto_SystemBus_slave_TLBuffer_out_c_bits_opcode(sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_opcode),
    .auto_SystemBus_slave_TLBuffer_out_c_bits_param(sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_param),
    .auto_SystemBus_slave_TLBuffer_out_c_bits_size(sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_size),
    .auto_SystemBus_slave_TLBuffer_out_c_bits_source(sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_source),
    .auto_SystemBus_slave_TLBuffer_out_d_ready(sbus_auto_SystemBus_slave_TLBuffer_out_d_ready),
    .auto_SystemBus_slave_TLBuffer_out_d_valid(sbus_auto_SystemBus_slave_TLBuffer_out_d_valid),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_opcode(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_opcode),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_param(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_param),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_size(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_size),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_source(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_source),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_sink(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_sink),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_data(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_data),
    .auto_SystemBus_slave_TLBuffer_out_d_bits_error(sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_error),
    .auto_SystemBus_out_a_ready(sbus_auto_SystemBus_out_a_ready),
    .auto_SystemBus_out_a_valid(sbus_auto_SystemBus_out_a_valid),
    .auto_SystemBus_out_a_bits_opcode(sbus_auto_SystemBus_out_a_bits_opcode),
    .auto_SystemBus_out_a_bits_param(sbus_auto_SystemBus_out_a_bits_param),
    .auto_SystemBus_out_a_bits_size(sbus_auto_SystemBus_out_a_bits_size),
    .auto_SystemBus_out_a_bits_source(sbus_auto_SystemBus_out_a_bits_source),
    .auto_SystemBus_out_a_bits_address(sbus_auto_SystemBus_out_a_bits_address),
    .auto_SystemBus_out_a_bits_mask(sbus_auto_SystemBus_out_a_bits_mask),
    .auto_SystemBus_out_a_bits_data(sbus_auto_SystemBus_out_a_bits_data),
    .auto_SystemBus_out_b_ready(sbus_auto_SystemBus_out_b_ready),
    .auto_SystemBus_out_b_valid(sbus_auto_SystemBus_out_b_valid),
    .auto_SystemBus_out_b_bits_param(sbus_auto_SystemBus_out_b_bits_param),
    .auto_SystemBus_out_b_bits_address(sbus_auto_SystemBus_out_b_bits_address),
    .auto_SystemBus_out_c_ready(sbus_auto_SystemBus_out_c_ready),
    .auto_SystemBus_out_c_valid(sbus_auto_SystemBus_out_c_valid),
    .auto_SystemBus_out_c_bits_opcode(sbus_auto_SystemBus_out_c_bits_opcode),
    .auto_SystemBus_out_c_bits_size(sbus_auto_SystemBus_out_c_bits_size),
    .auto_SystemBus_out_c_bits_source(sbus_auto_SystemBus_out_c_bits_source),
    .auto_SystemBus_out_c_bits_address(sbus_auto_SystemBus_out_c_bits_address),
    .auto_SystemBus_out_c_bits_data(sbus_auto_SystemBus_out_c_bits_data),
    .auto_SystemBus_out_d_ready(sbus_auto_SystemBus_out_d_ready),
    .auto_SystemBus_out_d_valid(sbus_auto_SystemBus_out_d_valid),
    .auto_SystemBus_out_d_bits_opcode(sbus_auto_SystemBus_out_d_bits_opcode),
    .auto_SystemBus_out_d_bits_param(sbus_auto_SystemBus_out_d_bits_param),
    .auto_SystemBus_out_d_bits_size(sbus_auto_SystemBus_out_d_bits_size),
    .auto_SystemBus_out_d_bits_source(sbus_auto_SystemBus_out_d_bits_source),
    .auto_SystemBus_out_d_bits_sink(sbus_auto_SystemBus_out_d_bits_sink),
    .auto_SystemBus_out_d_bits_data(sbus_auto_SystemBus_out_d_bits_data),
    .auto_SystemBus_out_d_bits_error(sbus_auto_SystemBus_out_d_bits_error),
    .auto_SystemBus_out_e_valid(sbus_auto_SystemBus_out_e_valid),
    .auto_SystemBus_out_e_bits_sink(sbus_auto_SystemBus_out_e_bits_sink)
  );
  PeripheryBus_pbus pbus (
    .clock(pbus_clock),
    .reset(pbus_reset),
    .auto_anon_in_a_ready(pbus_auto_anon_in_a_ready),
    .auto_anon_in_a_valid(pbus_auto_anon_in_a_valid),
    .auto_anon_in_a_bits_opcode(pbus_auto_anon_in_a_bits_opcode),
    .auto_anon_in_a_bits_param(pbus_auto_anon_in_a_bits_param),
    .auto_anon_in_a_bits_size(pbus_auto_anon_in_a_bits_size),
    .auto_anon_in_a_bits_source(pbus_auto_anon_in_a_bits_source),
    .auto_anon_in_a_bits_address(pbus_auto_anon_in_a_bits_address),
    .auto_anon_in_a_bits_mask(pbus_auto_anon_in_a_bits_mask),
    .auto_anon_in_a_bits_data(pbus_auto_anon_in_a_bits_data),
    .auto_anon_in_d_ready(pbus_auto_anon_in_d_ready),
    .auto_anon_in_d_valid(pbus_auto_anon_in_d_valid),
    .auto_anon_in_d_bits_opcode(pbus_auto_anon_in_d_bits_opcode),
    .auto_anon_in_d_bits_param(pbus_auto_anon_in_d_bits_param),
    .auto_anon_in_d_bits_size(pbus_auto_anon_in_d_bits_size),
    .auto_anon_in_d_bits_source(pbus_auto_anon_in_d_bits_source),
    .auto_anon_in_d_bits_sink(pbus_auto_anon_in_d_bits_sink),
    .auto_anon_in_d_bits_data(pbus_auto_anon_in_d_bits_data),
    .auto_anon_in_d_bits_error(pbus_auto_anon_in_d_bits_error),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_a_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_a_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_address(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_address),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_d_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_d_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_address(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_address),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_mask(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_mask),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_address(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_address),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_mask(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_mask),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_address(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_address),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_mask(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_mask),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_data),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_ready(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_ready),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_valid(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_valid),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_opcode(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_opcode),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_size(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_size),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_source(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_source),
    .auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_data(pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_data)
  );
  TLBroadcast TLBroadcast (
    .clock(TLBroadcast_clock),
    .reset(TLBroadcast_reset),
    .auto_in_a_ready(TLBroadcast_auto_in_a_ready),
    .auto_in_a_valid(TLBroadcast_auto_in_a_valid),
    .auto_in_a_bits_opcode(TLBroadcast_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(TLBroadcast_auto_in_a_bits_param),
    .auto_in_a_bits_size(TLBroadcast_auto_in_a_bits_size),
    .auto_in_a_bits_source(TLBroadcast_auto_in_a_bits_source),
    .auto_in_a_bits_address(TLBroadcast_auto_in_a_bits_address),
    .auto_in_a_bits_mask(TLBroadcast_auto_in_a_bits_mask),
    .auto_in_a_bits_data(TLBroadcast_auto_in_a_bits_data),
    .auto_in_b_ready(TLBroadcast_auto_in_b_ready),
    .auto_in_b_valid(TLBroadcast_auto_in_b_valid),
    .auto_in_b_bits_param(TLBroadcast_auto_in_b_bits_param),
    .auto_in_b_bits_address(TLBroadcast_auto_in_b_bits_address),
    .auto_in_c_ready(TLBroadcast_auto_in_c_ready),
    .auto_in_c_valid(TLBroadcast_auto_in_c_valid),
    .auto_in_c_bits_opcode(TLBroadcast_auto_in_c_bits_opcode),
    .auto_in_c_bits_size(TLBroadcast_auto_in_c_bits_size),
    .auto_in_c_bits_source(TLBroadcast_auto_in_c_bits_source),
    .auto_in_c_bits_address(TLBroadcast_auto_in_c_bits_address),
    .auto_in_c_bits_data(TLBroadcast_auto_in_c_bits_data),
    .auto_in_d_ready(TLBroadcast_auto_in_d_ready),
    .auto_in_d_valid(TLBroadcast_auto_in_d_valid),
    .auto_in_d_bits_opcode(TLBroadcast_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(TLBroadcast_auto_in_d_bits_param),
    .auto_in_d_bits_size(TLBroadcast_auto_in_d_bits_size),
    .auto_in_d_bits_source(TLBroadcast_auto_in_d_bits_source),
    .auto_in_d_bits_sink(TLBroadcast_auto_in_d_bits_sink),
    .auto_in_d_bits_data(TLBroadcast_auto_in_d_bits_data),
    .auto_in_d_bits_error(TLBroadcast_auto_in_d_bits_error),
    .auto_in_e_valid(TLBroadcast_auto_in_e_valid),
    .auto_in_e_bits_sink(TLBroadcast_auto_in_e_bits_sink),
    .auto_out_a_ready(TLBroadcast_auto_out_a_ready),
    .auto_out_a_valid(TLBroadcast_auto_out_a_valid),
    .auto_out_a_bits_opcode(TLBroadcast_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(TLBroadcast_auto_out_a_bits_size),
    .auto_out_a_bits_source(TLBroadcast_auto_out_a_bits_source),
    .auto_out_a_bits_address(TLBroadcast_auto_out_a_bits_address),
    .auto_out_a_bits_mask(TLBroadcast_auto_out_a_bits_mask),
    .auto_out_a_bits_data(TLBroadcast_auto_out_a_bits_data),
    .auto_out_d_ready(TLBroadcast_auto_out_d_ready),
    .auto_out_d_valid(TLBroadcast_auto_out_d_valid),
    .auto_out_d_bits_opcode(TLBroadcast_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(TLBroadcast_auto_out_d_bits_param),
    .auto_out_d_bits_size(TLBroadcast_auto_out_d_bits_size),
    .auto_out_d_bits_source(TLBroadcast_auto_out_d_bits_source),
    .auto_out_d_bits_data(TLBroadcast_auto_out_d_bits_data),
    .auto_out_d_bits_error(TLBroadcast_auto_out_d_bits_error)
  );
  TLWidthWidget TLWidthWidget (
    .auto_in_a_ready(TLWidthWidget_auto_in_a_ready),
    .auto_in_a_valid(TLWidthWidget_auto_in_a_valid),
    .auto_in_a_bits_opcode(TLWidthWidget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(TLWidthWidget_auto_in_a_bits_size),
    .auto_in_a_bits_source(TLWidthWidget_auto_in_a_bits_source),
    .auto_in_a_bits_address(TLWidthWidget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(TLWidthWidget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(TLWidthWidget_auto_in_a_bits_data),
    .auto_in_d_ready(TLWidthWidget_auto_in_d_ready),
    .auto_in_d_valid(TLWidthWidget_auto_in_d_valid),
    .auto_in_d_bits_opcode(TLWidthWidget_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(TLWidthWidget_auto_in_d_bits_param),
    .auto_in_d_bits_size(TLWidthWidget_auto_in_d_bits_size),
    .auto_in_d_bits_source(TLWidthWidget_auto_in_d_bits_source),
    .auto_in_d_bits_data(TLWidthWidget_auto_in_d_bits_data),
    .auto_in_d_bits_error(TLWidthWidget_auto_in_d_bits_error),
    .auto_out_a_ready(TLWidthWidget_auto_out_a_ready),
    .auto_out_a_valid(TLWidthWidget_auto_out_a_valid),
    .auto_out_a_bits_opcode(TLWidthWidget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(TLWidthWidget_auto_out_a_bits_size),
    .auto_out_a_bits_source(TLWidthWidget_auto_out_a_bits_source),
    .auto_out_a_bits_address(TLWidthWidget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(TLWidthWidget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(TLWidthWidget_auto_out_a_bits_data),
    .auto_out_d_ready(TLWidthWidget_auto_out_d_ready),
    .auto_out_d_valid(TLWidthWidget_auto_out_d_valid),
    .auto_out_d_bits_opcode(TLWidthWidget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(TLWidthWidget_auto_out_d_bits_param),
    .auto_out_d_bits_size(TLWidthWidget_auto_out_d_bits_size),
    .auto_out_d_bits_source(TLWidthWidget_auto_out_d_bits_source),
    .auto_out_d_bits_data(TLWidthWidget_auto_out_d_bits_data),
    .auto_out_d_bits_error(TLWidthWidget_auto_out_d_bits_error)
  );
  MemoryBus_memBuses_0 memBuses_0 (
    .clock(memBuses_0_clock),
    .reset(memBuses_0_reset),
    .auto_MemoryBus_slave_TLBuffer_out_a_ready(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_ready),
    .auto_MemoryBus_slave_TLBuffer_out_a_valid(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_valid),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_opcode(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_opcode),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_size(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_size),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_source(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_source),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_address(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_address),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_mask(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_mask),
    .auto_MemoryBus_slave_TLBuffer_out_a_bits_data(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_data),
    .auto_MemoryBus_slave_TLBuffer_out_d_ready(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_ready),
    .auto_MemoryBus_slave_TLBuffer_out_d_valid(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_valid),
    .auto_MemoryBus_slave_TLBuffer_out_d_bits_opcode(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_opcode),
    .auto_MemoryBus_slave_TLBuffer_out_d_bits_size(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_size),
    .auto_MemoryBus_slave_TLBuffer_out_d_bits_source(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_source),
    .auto_MemoryBus_slave_TLBuffer_out_d_bits_data(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_data),
    .auto_MemoryBus_slave_TLBuffer_out_d_bits_error(memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_error),
    .auto_MemoryBus_master_TLBuffer_in_a_ready(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_ready),
    .auto_MemoryBus_master_TLBuffer_in_a_valid(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_valid),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_opcode(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_opcode),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_size(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_size),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_source(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_source),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_address(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_address),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_mask(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_mask),
    .auto_MemoryBus_master_TLBuffer_in_a_bits_data(memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_data),
    .auto_MemoryBus_master_TLBuffer_in_d_ready(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_ready),
    .auto_MemoryBus_master_TLBuffer_in_d_valid(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_valid),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_opcode(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_opcode),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_param(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_param),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_size(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_size),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_source(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_source),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_data(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_data),
    .auto_MemoryBus_master_TLBuffer_in_d_bits_error(memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_error)
  );
  TLFilter TLFilter (
    .auto_in_a_ready(TLFilter_auto_in_a_ready),
    .auto_in_a_valid(TLFilter_auto_in_a_valid),
    .auto_in_a_bits_opcode(TLFilter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(TLFilter_auto_in_a_bits_size),
    .auto_in_a_bits_source(TLFilter_auto_in_a_bits_source),
    .auto_in_a_bits_address(TLFilter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(TLFilter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(TLFilter_auto_in_a_bits_data),
    .auto_in_d_ready(TLFilter_auto_in_d_ready),
    .auto_in_d_valid(TLFilter_auto_in_d_valid),
    .auto_in_d_bits_opcode(TLFilter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(TLFilter_auto_in_d_bits_param),
    .auto_in_d_bits_size(TLFilter_auto_in_d_bits_size),
    .auto_in_d_bits_source(TLFilter_auto_in_d_bits_source),
    .auto_in_d_bits_data(TLFilter_auto_in_d_bits_data),
    .auto_in_d_bits_error(TLFilter_auto_in_d_bits_error),
    .auto_out_a_ready(TLFilter_auto_out_a_ready),
    .auto_out_a_valid(TLFilter_auto_out_a_valid),
    .auto_out_a_bits_opcode(TLFilter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(TLFilter_auto_out_a_bits_size),
    .auto_out_a_bits_source(TLFilter_auto_out_a_bits_source),
    .auto_out_a_bits_address(TLFilter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(TLFilter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(TLFilter_auto_out_a_bits_data),
    .auto_out_d_ready(TLFilter_auto_out_d_ready),
    .auto_out_d_valid(TLFilter_auto_out_d_valid),
    .auto_out_d_bits_opcode(TLFilter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(TLFilter_auto_out_d_bits_param),
    .auto_out_d_bits_size(TLFilter_auto_out_d_bits_size),
    .auto_out_d_bits_source(TLFilter_auto_out_d_bits_source),
    .auto_out_d_bits_data(TLFilter_auto_out_d_bits_data),
    .auto_out_d_bits_error(TLFilter_auto_out_d_bits_error)
  );
  TLPLIC_plic plic (
    .clock(plic_clock),
    .reset(plic_reset),
    .auto_int_in_0(plic_auto_int_in_0),
    .auto_int_in_1(plic_auto_int_in_1),
    .auto_int_out_1_0(plic_auto_int_out_1_0),
    .auto_int_out_0_0(plic_auto_int_out_0_0),
    .auto_in_a_ready(plic_auto_in_a_ready),
    .auto_in_a_valid(plic_auto_in_a_valid),
    .auto_in_a_bits_opcode(plic_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(plic_auto_in_a_bits_size),
    .auto_in_a_bits_source(plic_auto_in_a_bits_source),
    .auto_in_a_bits_address(plic_auto_in_a_bits_address),
    .auto_in_a_bits_mask(plic_auto_in_a_bits_mask),
    .auto_in_a_bits_data(plic_auto_in_a_bits_data),
    .auto_in_d_ready(plic_auto_in_d_ready),
    .auto_in_d_valid(plic_auto_in_d_valid),
    .auto_in_d_bits_opcode(plic_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(plic_auto_in_d_bits_size),
    .auto_in_d_bits_source(plic_auto_in_d_bits_source),
    .auto_in_d_bits_data(plic_auto_in_d_bits_data)
  );
  CoreplexLocalInterrupter_clint clint (
    .clock(clint_clock),
    .reset(clint_reset),
    .auto_int_out_0(clint_auto_int_out_0),
    .auto_int_out_1(clint_auto_int_out_1),
    .auto_in_a_ready(clint_auto_in_a_ready),
    .auto_in_a_valid(clint_auto_in_a_valid),
    .auto_in_a_bits_opcode(clint_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(clint_auto_in_a_bits_size),
    .auto_in_a_bits_source(clint_auto_in_a_bits_source),
    .auto_in_a_bits_address(clint_auto_in_a_bits_address),
    .auto_in_a_bits_mask(clint_auto_in_a_bits_mask),
    .auto_in_a_bits_data(clint_auto_in_a_bits_data),
    .auto_in_d_ready(clint_auto_in_d_ready),
    .auto_in_d_valid(clint_auto_in_d_valid),
    .auto_in_d_bits_opcode(clint_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(clint_auto_in_d_bits_size),
    .auto_in_d_bits_source(clint_auto_in_d_bits_source),
    .auto_in_d_bits_data(clint_auto_in_d_bits_data),
    .io_rtcTick(clint_io_rtcTick)
  );
  TLDebugModule_debug debug_1 (
    .clock(debug_1_clock),
    .reset(debug_1_reset),
    .auto_dmInner_dmInner_tl_in_a_ready(debug_1_auto_dmInner_dmInner_tl_in_a_ready),
    .auto_dmInner_dmInner_tl_in_a_valid(debug_1_auto_dmInner_dmInner_tl_in_a_valid),
    .auto_dmInner_dmInner_tl_in_a_bits_opcode(debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode),
    .auto_dmInner_dmInner_tl_in_a_bits_size(debug_1_auto_dmInner_dmInner_tl_in_a_bits_size),
    .auto_dmInner_dmInner_tl_in_a_bits_source(debug_1_auto_dmInner_dmInner_tl_in_a_bits_source),
    .auto_dmInner_dmInner_tl_in_a_bits_address(debug_1_auto_dmInner_dmInner_tl_in_a_bits_address),
    .auto_dmInner_dmInner_tl_in_a_bits_mask(debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask),
    .auto_dmInner_dmInner_tl_in_a_bits_data(debug_1_auto_dmInner_dmInner_tl_in_a_bits_data),
    .auto_dmInner_dmInner_tl_in_d_ready(debug_1_auto_dmInner_dmInner_tl_in_d_ready),
    .auto_dmInner_dmInner_tl_in_d_valid(debug_1_auto_dmInner_dmInner_tl_in_d_valid),
    .auto_dmInner_dmInner_tl_in_d_bits_opcode(debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode),
    .auto_dmInner_dmInner_tl_in_d_bits_size(debug_1_auto_dmInner_dmInner_tl_in_d_bits_size),
    .auto_dmInner_dmInner_tl_in_d_bits_source(debug_1_auto_dmInner_dmInner_tl_in_d_bits_source),
    .auto_dmInner_dmInner_tl_in_d_bits_data(debug_1_auto_dmInner_dmInner_tl_in_d_bits_data),
    .auto_dmOuter_anon_out_sync_0(debug_1_auto_dmOuter_anon_out_sync_0),
    .io_ctrl_ndreset(debug_1_io_ctrl_ndreset),
    .io_ctrl_dmactive(debug_1_io_ctrl_dmactive),
    .io_dmi_dmi_req_ready(debug_1_io_dmi_dmi_req_ready),
    .io_dmi_dmi_req_valid(debug_1_io_dmi_dmi_req_valid),
    .io_dmi_dmi_req_bits_addr(debug_1_io_dmi_dmi_req_bits_addr),
    .io_dmi_dmi_req_bits_data(debug_1_io_dmi_dmi_req_bits_data),
    .io_dmi_dmi_req_bits_op(debug_1_io_dmi_dmi_req_bits_op),
    .io_dmi_dmi_resp_ready(debug_1_io_dmi_dmi_resp_ready),
    .io_dmi_dmi_resp_valid(debug_1_io_dmi_dmi_resp_valid),
    .io_dmi_dmi_resp_bits_data(debug_1_io_dmi_dmi_resp_bits_data),
    .io_dmi_dmi_resp_bits_resp(debug_1_io_dmi_dmi_resp_bits_resp),
    .io_dmi_dmiClock(debug_1_io_dmi_dmiClock),
    .io_dmi_dmiReset(debug_1_io_dmi_dmiReset)
  );
  BoomTileWrapper_tile tile (
    .clock(tile_clock),
    .reset(tile_reset),
    .auto_anon_in_3_sync_0(tile_auto_anon_in_3_sync_0),
    .auto_anon_in_2_sync_0(tile_auto_anon_in_2_sync_0),
    .auto_anon_in_1_sync_0(tile_auto_anon_in_1_sync_0),
    .auto_anon_in_1_sync_1(tile_auto_anon_in_1_sync_1),
    .auto_anon_in_0_sync_0(tile_auto_anon_in_0_sync_0),
    .auto_anon_out_a_ready(tile_auto_anon_out_a_ready),
    .auto_anon_out_a_valid(tile_auto_anon_out_a_valid),
    .auto_anon_out_a_bits_opcode(tile_auto_anon_out_a_bits_opcode),
    .auto_anon_out_a_bits_param(tile_auto_anon_out_a_bits_param),
    .auto_anon_out_a_bits_size(tile_auto_anon_out_a_bits_size),
    .auto_anon_out_a_bits_source(tile_auto_anon_out_a_bits_source),
    .auto_anon_out_a_bits_address(tile_auto_anon_out_a_bits_address),
    .auto_anon_out_a_bits_mask(tile_auto_anon_out_a_bits_mask),
    .auto_anon_out_a_bits_data(tile_auto_anon_out_a_bits_data),
    .auto_anon_out_b_ready(tile_auto_anon_out_b_ready),
    .auto_anon_out_b_valid(tile_auto_anon_out_b_valid),
    .auto_anon_out_b_bits_param(tile_auto_anon_out_b_bits_param),
    .auto_anon_out_b_bits_size(tile_auto_anon_out_b_bits_size),
    .auto_anon_out_b_bits_source(tile_auto_anon_out_b_bits_source),
    .auto_anon_out_b_bits_address(tile_auto_anon_out_b_bits_address),
    .auto_anon_out_c_ready(tile_auto_anon_out_c_ready),
    .auto_anon_out_c_valid(tile_auto_anon_out_c_valid),
    .auto_anon_out_c_bits_opcode(tile_auto_anon_out_c_bits_opcode),
    .auto_anon_out_c_bits_param(tile_auto_anon_out_c_bits_param),
    .auto_anon_out_c_bits_size(tile_auto_anon_out_c_bits_size),
    .auto_anon_out_c_bits_source(tile_auto_anon_out_c_bits_source),
    .auto_anon_out_c_bits_address(tile_auto_anon_out_c_bits_address),
    .auto_anon_out_c_bits_data(tile_auto_anon_out_c_bits_data),
    .auto_anon_out_d_ready(tile_auto_anon_out_d_ready),
    .auto_anon_out_d_valid(tile_auto_anon_out_d_valid),
    .auto_anon_out_d_bits_opcode(tile_auto_anon_out_d_bits_opcode),
    .auto_anon_out_d_bits_param(tile_auto_anon_out_d_bits_param),
    .auto_anon_out_d_bits_size(tile_auto_anon_out_d_bits_size),
    .auto_anon_out_d_bits_source(tile_auto_anon_out_d_bits_source),
    .auto_anon_out_d_bits_sink(tile_auto_anon_out_d_bits_sink),
    .auto_anon_out_d_bits_data(tile_auto_anon_out_d_bits_data),
    .auto_anon_out_d_bits_error(tile_auto_anon_out_d_bits_error),
    .auto_anon_out_e_ready(tile_auto_anon_out_e_ready),
    .auto_anon_out_e_valid(tile_auto_anon_out_e_valid),
    .auto_anon_out_e_bits_sink(tile_auto_anon_out_e_bits_sink)
  );
  IntSyncCrossingSource_1 IntSyncCrossingSource (
    .clock(IntSyncCrossingSource_clock),
    .reset(IntSyncCrossingSource_reset),
    .auto_in_2_0(IntSyncCrossingSource_auto_in_2_0),
    .auto_in_1_0(IntSyncCrossingSource_auto_in_1_0),
    .auto_in_0_0(IntSyncCrossingSource_auto_in_0_0),
    .auto_in_0_1(IntSyncCrossingSource_auto_in_0_1),
    .auto_out_2_sync_0(IntSyncCrossingSource_auto_out_2_sync_0),
    .auto_out_1_sync_0(IntSyncCrossingSource_auto_out_1_sync_0),
    .auto_out_0_sync_0(IntSyncCrossingSource_auto_out_0_sync_0),
    .auto_out_0_sync_1(IntSyncCrossingSource_auto_out_0_sync_1)
  );
  IntXing IntXing (
    .clock(IntXing_clock),
    .auto_int_in_0(IntXing_auto_int_in_0),
    .auto_int_in_1(IntXing_auto_int_in_1),
    .auto_int_out_0(IntXing_auto_int_out_0),
    .auto_int_out_1(IntXing_auto_int_out_1)
  );
  TLToAXI4_converter converter (
    .clock(converter_clock),
    .reset(converter_reset),
    .auto_in_a_ready(converter_auto_in_a_ready),
    .auto_in_a_valid(converter_auto_in_a_valid),
    .auto_in_a_bits_opcode(converter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(converter_auto_in_a_bits_size),
    .auto_in_a_bits_source(converter_auto_in_a_bits_source),
    .auto_in_a_bits_address(converter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(converter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(converter_auto_in_a_bits_data),
    .auto_in_d_ready(converter_auto_in_d_ready),
    .auto_in_d_valid(converter_auto_in_d_valid),
    .auto_in_d_bits_opcode(converter_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(converter_auto_in_d_bits_size),
    .auto_in_d_bits_source(converter_auto_in_d_bits_source),
    .auto_in_d_bits_data(converter_auto_in_d_bits_data),
    .auto_in_d_bits_error(converter_auto_in_d_bits_error),
    .auto_out_aw_ready(converter_auto_out_aw_ready),
    .auto_out_aw_valid(converter_auto_out_aw_valid),
    .auto_out_aw_bits_id(converter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(converter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(converter_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(converter_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(converter_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(converter_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(converter_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(converter_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(converter_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(converter_auto_out_aw_bits_user),
    .auto_out_w_ready(converter_auto_out_w_ready),
    .auto_out_w_valid(converter_auto_out_w_valid),
    .auto_out_w_bits_data(converter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(converter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(converter_auto_out_w_bits_last),
    .auto_out_b_ready(converter_auto_out_b_ready),
    .auto_out_b_valid(converter_auto_out_b_valid),
    .auto_out_b_bits_id(converter_auto_out_b_bits_id),
    .auto_out_b_bits_resp(converter_auto_out_b_bits_resp),
    .auto_out_b_bits_user(converter_auto_out_b_bits_user),
    .auto_out_ar_ready(converter_auto_out_ar_ready),
    .auto_out_ar_valid(converter_auto_out_ar_valid),
    .auto_out_ar_bits_id(converter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(converter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(converter_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(converter_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(converter_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(converter_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(converter_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(converter_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(converter_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(converter_auto_out_ar_bits_user),
    .auto_out_r_ready(converter_auto_out_r_ready),
    .auto_out_r_valid(converter_auto_out_r_valid),
    .auto_out_r_bits_id(converter_auto_out_r_bits_id),
    .auto_out_r_bits_data(converter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(converter_auto_out_r_bits_resp),
    .auto_out_r_bits_user(converter_auto_out_r_bits_user),
    .auto_out_r_bits_last(converter_auto_out_r_bits_last)
  );
  AXI4IdIndexer_trim trim (
    .auto_in_aw_ready(trim_auto_in_aw_ready),
    .auto_in_aw_valid(trim_auto_in_aw_valid),
    .auto_in_aw_bits_id(trim_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(trim_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(trim_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(trim_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(trim_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(trim_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(trim_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(trim_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(trim_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(trim_auto_in_aw_bits_user),
    .auto_in_w_ready(trim_auto_in_w_ready),
    .auto_in_w_valid(trim_auto_in_w_valid),
    .auto_in_w_bits_data(trim_auto_in_w_bits_data),
    .auto_in_w_bits_strb(trim_auto_in_w_bits_strb),
    .auto_in_w_bits_last(trim_auto_in_w_bits_last),
    .auto_in_b_ready(trim_auto_in_b_ready),
    .auto_in_b_valid(trim_auto_in_b_valid),
    .auto_in_b_bits_id(trim_auto_in_b_bits_id),
    .auto_in_b_bits_resp(trim_auto_in_b_bits_resp),
    .auto_in_b_bits_user(trim_auto_in_b_bits_user),
    .auto_in_ar_ready(trim_auto_in_ar_ready),
    .auto_in_ar_valid(trim_auto_in_ar_valid),
    .auto_in_ar_bits_id(trim_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(trim_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(trim_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(trim_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(trim_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(trim_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(trim_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(trim_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(trim_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(trim_auto_in_ar_bits_user),
    .auto_in_r_ready(trim_auto_in_r_ready),
    .auto_in_r_valid(trim_auto_in_r_valid),
    .auto_in_r_bits_id(trim_auto_in_r_bits_id),
    .auto_in_r_bits_data(trim_auto_in_r_bits_data),
    .auto_in_r_bits_resp(trim_auto_in_r_bits_resp),
    .auto_in_r_bits_user(trim_auto_in_r_bits_user),
    .auto_in_r_bits_last(trim_auto_in_r_bits_last),
    .auto_out_aw_ready(trim_auto_out_aw_ready),
    .auto_out_aw_valid(trim_auto_out_aw_valid),
    .auto_out_aw_bits_id(trim_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(trim_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(trim_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(trim_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(trim_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(trim_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(trim_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(trim_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(trim_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(trim_auto_out_aw_bits_user),
    .auto_out_w_ready(trim_auto_out_w_ready),
    .auto_out_w_valid(trim_auto_out_w_valid),
    .auto_out_w_bits_data(trim_auto_out_w_bits_data),
    .auto_out_w_bits_strb(trim_auto_out_w_bits_strb),
    .auto_out_w_bits_last(trim_auto_out_w_bits_last),
    .auto_out_b_ready(trim_auto_out_b_ready),
    .auto_out_b_valid(trim_auto_out_b_valid),
    .auto_out_b_bits_id(trim_auto_out_b_bits_id),
    .auto_out_b_bits_resp(trim_auto_out_b_bits_resp),
    .auto_out_b_bits_user(trim_auto_out_b_bits_user),
    .auto_out_ar_ready(trim_auto_out_ar_ready),
    .auto_out_ar_valid(trim_auto_out_ar_valid),
    .auto_out_ar_bits_id(trim_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(trim_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(trim_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(trim_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(trim_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(trim_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(trim_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(trim_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(trim_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(trim_auto_out_ar_bits_user),
    .auto_out_r_ready(trim_auto_out_r_ready),
    .auto_out_r_valid(trim_auto_out_r_valid),
    .auto_out_r_bits_id(trim_auto_out_r_bits_id),
    .auto_out_r_bits_data(trim_auto_out_r_bits_data),
    .auto_out_r_bits_resp(trim_auto_out_r_bits_resp),
    .auto_out_r_bits_user(trim_auto_out_r_bits_user),
    .auto_out_r_bits_last(trim_auto_out_r_bits_last)
  );
  AXI4UserYanker_yank yank (
    .clock(yank_clock),
    .reset(yank_reset),
    .auto_in_aw_ready(yank_auto_in_aw_ready),
    .auto_in_aw_valid(yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(yank_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(yank_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(yank_auto_in_aw_bits_user),
    .auto_in_w_ready(yank_auto_in_w_ready),
    .auto_in_w_valid(yank_auto_in_w_valid),
    .auto_in_w_bits_data(yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(yank_auto_in_w_bits_last),
    .auto_in_b_ready(yank_auto_in_b_ready),
    .auto_in_b_valid(yank_auto_in_b_valid),
    .auto_in_b_bits_id(yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(yank_auto_in_b_bits_resp),
    .auto_in_b_bits_user(yank_auto_in_b_bits_user),
    .auto_in_ar_ready(yank_auto_in_ar_ready),
    .auto_in_ar_valid(yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(yank_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(yank_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(yank_auto_in_ar_bits_user),
    .auto_in_r_ready(yank_auto_in_r_ready),
    .auto_in_r_valid(yank_auto_in_r_valid),
    .auto_in_r_bits_id(yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(yank_auto_in_r_bits_resp),
    .auto_in_r_bits_user(yank_auto_in_r_bits_user),
    .auto_in_r_bits_last(yank_auto_in_r_bits_last),
    .auto_out_aw_ready(yank_auto_out_aw_ready),
    .auto_out_aw_valid(yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(yank_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(yank_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(yank_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(yank_auto_out_aw_bits_qos),
    .auto_out_w_ready(yank_auto_out_w_ready),
    .auto_out_w_valid(yank_auto_out_w_valid),
    .auto_out_w_bits_data(yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(yank_auto_out_w_bits_last),
    .auto_out_b_ready(yank_auto_out_b_ready),
    .auto_out_b_valid(yank_auto_out_b_valid),
    .auto_out_b_bits_id(yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(yank_auto_out_ar_ready),
    .auto_out_ar_valid(yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(yank_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(yank_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(yank_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(yank_auto_out_ar_bits_qos),
    .auto_out_r_ready(yank_auto_out_r_ready),
    .auto_out_r_valid(yank_auto_out_r_valid),
    .auto_out_r_bits_id(yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(yank_auto_out_r_bits_last)
  );
  AXI4Buffer_buffer buffer (
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_aw_ready(buffer_auto_in_aw_ready),
    .auto_in_aw_valid(buffer_auto_in_aw_valid),
    .auto_in_aw_bits_id(buffer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(buffer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(buffer_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(buffer_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(buffer_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(buffer_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(buffer_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(buffer_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(buffer_auto_in_aw_bits_qos),
    .auto_in_w_ready(buffer_auto_in_w_ready),
    .auto_in_w_valid(buffer_auto_in_w_valid),
    .auto_in_w_bits_data(buffer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(buffer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(buffer_auto_in_w_bits_last),
    .auto_in_b_ready(buffer_auto_in_b_ready),
    .auto_in_b_valid(buffer_auto_in_b_valid),
    .auto_in_b_bits_id(buffer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(buffer_auto_in_b_bits_resp),
    .auto_in_ar_ready(buffer_auto_in_ar_ready),
    .auto_in_ar_valid(buffer_auto_in_ar_valid),
    .auto_in_ar_bits_id(buffer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(buffer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(buffer_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(buffer_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(buffer_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(buffer_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(buffer_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(buffer_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(buffer_auto_in_ar_bits_qos),
    .auto_in_r_ready(buffer_auto_in_r_ready),
    .auto_in_r_valid(buffer_auto_in_r_valid),
    .auto_in_r_bits_id(buffer_auto_in_r_bits_id),
    .auto_in_r_bits_data(buffer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(buffer_auto_in_r_bits_resp),
    .auto_in_r_bits_last(buffer_auto_in_r_bits_last),
    .auto_out_aw_ready(buffer_auto_out_aw_ready),
    .auto_out_aw_valid(buffer_auto_out_aw_valid),
    .auto_out_aw_bits_id(buffer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(buffer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(buffer_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(buffer_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(buffer_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(buffer_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(buffer_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(buffer_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(buffer_auto_out_aw_bits_qos),
    .auto_out_w_ready(buffer_auto_out_w_ready),
    .auto_out_w_valid(buffer_auto_out_w_valid),
    .auto_out_w_bits_data(buffer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(buffer_auto_out_w_bits_strb),
    .auto_out_w_bits_last(buffer_auto_out_w_bits_last),
    .auto_out_b_ready(buffer_auto_out_b_ready),
    .auto_out_b_valid(buffer_auto_out_b_valid),
    .auto_out_b_bits_id(buffer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(buffer_auto_out_b_bits_resp),
    .auto_out_ar_ready(buffer_auto_out_ar_ready),
    .auto_out_ar_valid(buffer_auto_out_ar_valid),
    .auto_out_ar_bits_id(buffer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(buffer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(buffer_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(buffer_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(buffer_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(buffer_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(buffer_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(buffer_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(buffer_auto_out_ar_bits_qos),
    .auto_out_r_ready(buffer_auto_out_r_ready),
    .auto_out_r_valid(buffer_auto_out_r_valid),
    .auto_out_r_bits_id(buffer_auto_out_r_bits_id),
    .auto_out_r_bits_data(buffer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(buffer_auto_out_r_bits_resp),
    .auto_out_r_bits_last(buffer_auto_out_r_bits_last)
  );
  AXI4Buffer AXI4Buffer (
    .clock(AXI4Buffer_clock),
    .reset(AXI4Buffer_reset),
    .auto_in_aw_ready(AXI4Buffer_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Buffer_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Buffer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Buffer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4Buffer_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4Buffer_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4Buffer_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(AXI4Buffer_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(AXI4Buffer_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(AXI4Buffer_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(AXI4Buffer_auto_in_aw_bits_qos),
    .auto_in_w_ready(AXI4Buffer_auto_in_w_ready),
    .auto_in_w_valid(AXI4Buffer_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Buffer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Buffer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Buffer_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Buffer_auto_in_b_ready),
    .auto_in_b_valid(AXI4Buffer_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Buffer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Buffer_auto_in_b_bits_resp),
    .auto_in_ar_ready(AXI4Buffer_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Buffer_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Buffer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Buffer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4Buffer_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4Buffer_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4Buffer_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(AXI4Buffer_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(AXI4Buffer_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(AXI4Buffer_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(AXI4Buffer_auto_in_ar_bits_qos),
    .auto_in_r_ready(AXI4Buffer_auto_in_r_ready),
    .auto_in_r_valid(AXI4Buffer_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Buffer_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Buffer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Buffer_auto_in_r_bits_resp),
    .auto_in_r_bits_last(AXI4Buffer_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Buffer_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Buffer_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Buffer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Buffer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4Buffer_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4Buffer_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(AXI4Buffer_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(AXI4Buffer_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(AXI4Buffer_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(AXI4Buffer_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(AXI4Buffer_auto_out_aw_bits_qos),
    .auto_out_w_ready(AXI4Buffer_auto_out_w_ready),
    .auto_out_w_valid(AXI4Buffer_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Buffer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Buffer_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4Buffer_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4Buffer_auto_out_b_ready),
    .auto_out_b_valid(AXI4Buffer_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Buffer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Buffer_auto_out_b_bits_resp),
    .auto_out_ar_ready(AXI4Buffer_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Buffer_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Buffer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Buffer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4Buffer_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4Buffer_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(AXI4Buffer_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(AXI4Buffer_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(AXI4Buffer_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(AXI4Buffer_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(AXI4Buffer_auto_out_ar_bits_qos),
    .auto_out_r_ready(AXI4Buffer_auto_out_r_ready),
    .auto_out_r_valid(AXI4Buffer_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Buffer_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Buffer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Buffer_auto_out_r_bits_resp),
    .auto_out_r_bits_last(AXI4Buffer_auto_out_r_bits_last)
  );
  AXI4UserYanker AXI4UserYanker (
    .clock(AXI4UserYanker_clock),
    .reset(AXI4UserYanker_reset),
    .auto_in_aw_ready(AXI4UserYanker_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4UserYanker_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4UserYanker_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4UserYanker_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4UserYanker_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4UserYanker_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4UserYanker_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(AXI4UserYanker_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(AXI4UserYanker_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(AXI4UserYanker_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(AXI4UserYanker_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(AXI4UserYanker_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4UserYanker_auto_in_w_ready),
    .auto_in_w_valid(AXI4UserYanker_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4UserYanker_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4UserYanker_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4UserYanker_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4UserYanker_auto_in_b_ready),
    .auto_in_b_valid(AXI4UserYanker_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4UserYanker_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4UserYanker_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4UserYanker_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4UserYanker_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4UserYanker_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4UserYanker_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4UserYanker_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4UserYanker_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4UserYanker_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4UserYanker_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(AXI4UserYanker_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(AXI4UserYanker_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(AXI4UserYanker_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(AXI4UserYanker_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(AXI4UserYanker_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4UserYanker_auto_in_r_ready),
    .auto_in_r_valid(AXI4UserYanker_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4UserYanker_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4UserYanker_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4UserYanker_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4UserYanker_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4UserYanker_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4UserYanker_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4UserYanker_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4UserYanker_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4UserYanker_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4UserYanker_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4UserYanker_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(AXI4UserYanker_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(AXI4UserYanker_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(AXI4UserYanker_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(AXI4UserYanker_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(AXI4UserYanker_auto_out_aw_bits_qos),
    .auto_out_w_ready(AXI4UserYanker_auto_out_w_ready),
    .auto_out_w_valid(AXI4UserYanker_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4UserYanker_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4UserYanker_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4UserYanker_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4UserYanker_auto_out_b_ready),
    .auto_out_b_valid(AXI4UserYanker_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4UserYanker_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4UserYanker_auto_out_b_bits_resp),
    .auto_out_ar_ready(AXI4UserYanker_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4UserYanker_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4UserYanker_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4UserYanker_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4UserYanker_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4UserYanker_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(AXI4UserYanker_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(AXI4UserYanker_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(AXI4UserYanker_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(AXI4UserYanker_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(AXI4UserYanker_auto_out_ar_bits_qos),
    .auto_out_r_ready(AXI4UserYanker_auto_out_r_ready),
    .auto_out_r_valid(AXI4UserYanker_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4UserYanker_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4UserYanker_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4UserYanker_auto_out_r_bits_resp),
    .auto_out_r_bits_last(AXI4UserYanker_auto_out_r_bits_last)
  );
  AXI4Deinterleaver AXI4Deinterleaver (
    .clock(AXI4Deinterleaver_clock),
    .reset(AXI4Deinterleaver_reset),
    .auto_in_aw_ready(AXI4Deinterleaver_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Deinterleaver_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Deinterleaver_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Deinterleaver_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4Deinterleaver_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4Deinterleaver_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4Deinterleaver_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(AXI4Deinterleaver_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(AXI4Deinterleaver_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(AXI4Deinterleaver_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(AXI4Deinterleaver_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(AXI4Deinterleaver_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4Deinterleaver_auto_in_w_ready),
    .auto_in_w_valid(AXI4Deinterleaver_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Deinterleaver_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Deinterleaver_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Deinterleaver_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Deinterleaver_auto_in_b_ready),
    .auto_in_b_valid(AXI4Deinterleaver_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Deinterleaver_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Deinterleaver_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4Deinterleaver_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4Deinterleaver_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Deinterleaver_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Deinterleaver_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Deinterleaver_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4Deinterleaver_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4Deinterleaver_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4Deinterleaver_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(AXI4Deinterleaver_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(AXI4Deinterleaver_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(AXI4Deinterleaver_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(AXI4Deinterleaver_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(AXI4Deinterleaver_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4Deinterleaver_auto_in_r_ready),
    .auto_in_r_valid(AXI4Deinterleaver_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Deinterleaver_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Deinterleaver_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Deinterleaver_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4Deinterleaver_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4Deinterleaver_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Deinterleaver_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Deinterleaver_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Deinterleaver_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Deinterleaver_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4Deinterleaver_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4Deinterleaver_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(AXI4Deinterleaver_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(AXI4Deinterleaver_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(AXI4Deinterleaver_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(AXI4Deinterleaver_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(AXI4Deinterleaver_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(AXI4Deinterleaver_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Deinterleaver_auto_out_w_ready),
    .auto_out_w_valid(AXI4Deinterleaver_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Deinterleaver_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Deinterleaver_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4Deinterleaver_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4Deinterleaver_auto_out_b_ready),
    .auto_out_b_valid(AXI4Deinterleaver_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Deinterleaver_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Deinterleaver_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Deinterleaver_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Deinterleaver_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Deinterleaver_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Deinterleaver_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Deinterleaver_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4Deinterleaver_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4Deinterleaver_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(AXI4Deinterleaver_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(AXI4Deinterleaver_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(AXI4Deinterleaver_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(AXI4Deinterleaver_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(AXI4Deinterleaver_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(AXI4Deinterleaver_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Deinterleaver_auto_out_r_ready),
    .auto_out_r_valid(AXI4Deinterleaver_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Deinterleaver_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Deinterleaver_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Deinterleaver_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Deinterleaver_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4Deinterleaver_auto_out_r_bits_last)
  );
  AXI4IdIndexer AXI4IdIndexer (
    .auto_in_aw_ready(AXI4IdIndexer_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4IdIndexer_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4IdIndexer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4IdIndexer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4IdIndexer_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4IdIndexer_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4IdIndexer_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(AXI4IdIndexer_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(AXI4IdIndexer_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(AXI4IdIndexer_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(AXI4IdIndexer_auto_in_aw_bits_qos),
    .auto_in_aw_bits_user(AXI4IdIndexer_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4IdIndexer_auto_in_w_ready),
    .auto_in_w_valid(AXI4IdIndexer_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4IdIndexer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4IdIndexer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4IdIndexer_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4IdIndexer_auto_in_b_ready),
    .auto_in_b_valid(AXI4IdIndexer_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4IdIndexer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4IdIndexer_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4IdIndexer_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4IdIndexer_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4IdIndexer_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4IdIndexer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4IdIndexer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4IdIndexer_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4IdIndexer_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4IdIndexer_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(AXI4IdIndexer_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(AXI4IdIndexer_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(AXI4IdIndexer_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(AXI4IdIndexer_auto_in_ar_bits_qos),
    .auto_in_ar_bits_user(AXI4IdIndexer_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4IdIndexer_auto_in_r_ready),
    .auto_in_r_valid(AXI4IdIndexer_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4IdIndexer_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4IdIndexer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4IdIndexer_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4IdIndexer_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4IdIndexer_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4IdIndexer_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4IdIndexer_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4IdIndexer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4IdIndexer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4IdIndexer_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4IdIndexer_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(AXI4IdIndexer_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(AXI4IdIndexer_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(AXI4IdIndexer_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(AXI4IdIndexer_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(AXI4IdIndexer_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(AXI4IdIndexer_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4IdIndexer_auto_out_w_ready),
    .auto_out_w_valid(AXI4IdIndexer_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4IdIndexer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4IdIndexer_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4IdIndexer_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4IdIndexer_auto_out_b_ready),
    .auto_out_b_valid(AXI4IdIndexer_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4IdIndexer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4IdIndexer_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4IdIndexer_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4IdIndexer_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4IdIndexer_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4IdIndexer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4IdIndexer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4IdIndexer_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4IdIndexer_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(AXI4IdIndexer_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(AXI4IdIndexer_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(AXI4IdIndexer_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(AXI4IdIndexer_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(AXI4IdIndexer_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(AXI4IdIndexer_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4IdIndexer_auto_out_r_ready),
    .auto_out_r_valid(AXI4IdIndexer_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4IdIndexer_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4IdIndexer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4IdIndexer_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4IdIndexer_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4IdIndexer_auto_out_r_bits_last)
  );
  TLToAXI4 TLToAXI4 (
    .clock(TLToAXI4_clock),
    .reset(TLToAXI4_reset),
    .auto_in_a_ready(TLToAXI4_auto_in_a_ready),
    .auto_in_a_valid(TLToAXI4_auto_in_a_valid),
    .auto_in_a_bits_opcode(TLToAXI4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(TLToAXI4_auto_in_a_bits_size),
    .auto_in_a_bits_source(TLToAXI4_auto_in_a_bits_source),
    .auto_in_a_bits_address(TLToAXI4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(TLToAXI4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(TLToAXI4_auto_in_a_bits_data),
    .auto_in_d_ready(TLToAXI4_auto_in_d_ready),
    .auto_in_d_valid(TLToAXI4_auto_in_d_valid),
    .auto_in_d_bits_opcode(TLToAXI4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(TLToAXI4_auto_in_d_bits_size),
    .auto_in_d_bits_source(TLToAXI4_auto_in_d_bits_source),
    .auto_in_d_bits_data(TLToAXI4_auto_in_d_bits_data),
    .auto_in_d_bits_error(TLToAXI4_auto_in_d_bits_error),
    .auto_out_aw_ready(TLToAXI4_auto_out_aw_ready),
    .auto_out_aw_valid(TLToAXI4_auto_out_aw_valid),
    .auto_out_aw_bits_id(TLToAXI4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(TLToAXI4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(TLToAXI4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(TLToAXI4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(TLToAXI4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(TLToAXI4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(TLToAXI4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(TLToAXI4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(TLToAXI4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_user(TLToAXI4_auto_out_aw_bits_user),
    .auto_out_w_ready(TLToAXI4_auto_out_w_ready),
    .auto_out_w_valid(TLToAXI4_auto_out_w_valid),
    .auto_out_w_bits_data(TLToAXI4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(TLToAXI4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(TLToAXI4_auto_out_w_bits_last),
    .auto_out_b_ready(TLToAXI4_auto_out_b_ready),
    .auto_out_b_valid(TLToAXI4_auto_out_b_valid),
    .auto_out_b_bits_id(TLToAXI4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(TLToAXI4_auto_out_b_bits_resp),
    .auto_out_b_bits_user(TLToAXI4_auto_out_b_bits_user),
    .auto_out_ar_ready(TLToAXI4_auto_out_ar_ready),
    .auto_out_ar_valid(TLToAXI4_auto_out_ar_valid),
    .auto_out_ar_bits_id(TLToAXI4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(TLToAXI4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(TLToAXI4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(TLToAXI4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(TLToAXI4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(TLToAXI4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(TLToAXI4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(TLToAXI4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(TLToAXI4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_user(TLToAXI4_auto_out_ar_bits_user),
    .auto_out_r_ready(TLToAXI4_auto_out_r_ready),
    .auto_out_r_valid(TLToAXI4_auto_out_r_valid),
    .auto_out_r_bits_id(TLToAXI4_auto_out_r_bits_id),
    .auto_out_r_bits_data(TLToAXI4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(TLToAXI4_auto_out_r_bits_resp),
    .auto_out_r_bits_user(TLToAXI4_auto_out_r_bits_user),
    .auto_out_r_bits_last(TLToAXI4_auto_out_r_bits_last)
  );
  TLBuffer_SystemBus_1 SystemBus_TLBuffer (
    .clock(SystemBus_TLBuffer_clock),
    .reset(SystemBus_TLBuffer_reset),
    .auto_in_a_ready(SystemBus_TLBuffer_auto_in_a_ready),
    .auto_in_a_valid(SystemBus_TLBuffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(SystemBus_TLBuffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(SystemBus_TLBuffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(SystemBus_TLBuffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(SystemBus_TLBuffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(SystemBus_TLBuffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(SystemBus_TLBuffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(SystemBus_TLBuffer_auto_in_a_bits_data),
    .auto_in_d_ready(SystemBus_TLBuffer_auto_in_d_ready),
    .auto_in_d_valid(SystemBus_TLBuffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(SystemBus_TLBuffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(SystemBus_TLBuffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(SystemBus_TLBuffer_auto_in_d_bits_source),
    .auto_in_d_bits_data(SystemBus_TLBuffer_auto_in_d_bits_data),
    .auto_in_d_bits_error(SystemBus_TLBuffer_auto_in_d_bits_error),
    .auto_out_a_ready(SystemBus_TLBuffer_auto_out_a_ready),
    .auto_out_a_valid(SystemBus_TLBuffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(SystemBus_TLBuffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(SystemBus_TLBuffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(SystemBus_TLBuffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(SystemBus_TLBuffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(SystemBus_TLBuffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(SystemBus_TLBuffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(SystemBus_TLBuffer_auto_out_a_bits_data),
    .auto_out_d_ready(SystemBus_TLBuffer_auto_out_d_ready),
    .auto_out_d_valid(SystemBus_TLBuffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(SystemBus_TLBuffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(SystemBus_TLBuffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(SystemBus_TLBuffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(SystemBus_TLBuffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(SystemBus_TLBuffer_auto_out_d_bits_sink),
    .auto_out_d_bits_data(SystemBus_TLBuffer_auto_out_d_bits_data),
    .auto_out_d_bits_error(SystemBus_TLBuffer_auto_out_d_bits_error)
  );
  TLWidthWidget_SystemBus SystemBus_TLWidthWidget (
    .auto_in_a_ready(SystemBus_TLWidthWidget_auto_in_a_ready),
    .auto_in_a_valid(SystemBus_TLWidthWidget_auto_in_a_valid),
    .auto_in_a_bits_opcode(SystemBus_TLWidthWidget_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(SystemBus_TLWidthWidget_auto_in_a_bits_param),
    .auto_in_a_bits_size(SystemBus_TLWidthWidget_auto_in_a_bits_size),
    .auto_in_a_bits_source(SystemBus_TLWidthWidget_auto_in_a_bits_source),
    .auto_in_a_bits_address(SystemBus_TLWidthWidget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(SystemBus_TLWidthWidget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(SystemBus_TLWidthWidget_auto_in_a_bits_data),
    .auto_in_d_ready(SystemBus_TLWidthWidget_auto_in_d_ready),
    .auto_in_d_valid(SystemBus_TLWidthWidget_auto_in_d_valid),
    .auto_in_d_bits_opcode(SystemBus_TLWidthWidget_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(SystemBus_TLWidthWidget_auto_in_d_bits_size),
    .auto_in_d_bits_source(SystemBus_TLWidthWidget_auto_in_d_bits_source),
    .auto_in_d_bits_data(SystemBus_TLWidthWidget_auto_in_d_bits_data),
    .auto_in_d_bits_error(SystemBus_TLWidthWidget_auto_in_d_bits_error),
    .auto_out_a_ready(SystemBus_TLWidthWidget_auto_out_a_ready),
    .auto_out_a_valid(SystemBus_TLWidthWidget_auto_out_a_valid),
    .auto_out_a_bits_opcode(SystemBus_TLWidthWidget_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(SystemBus_TLWidthWidget_auto_out_a_bits_param),
    .auto_out_a_bits_size(SystemBus_TLWidthWidget_auto_out_a_bits_size),
    .auto_out_a_bits_source(SystemBus_TLWidthWidget_auto_out_a_bits_source),
    .auto_out_a_bits_address(SystemBus_TLWidthWidget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(SystemBus_TLWidthWidget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(SystemBus_TLWidthWidget_auto_out_a_bits_data),
    .auto_out_d_ready(SystemBus_TLWidthWidget_auto_out_d_ready),
    .auto_out_d_valid(SystemBus_TLWidthWidget_auto_out_d_valid),
    .auto_out_d_bits_opcode(SystemBus_TLWidthWidget_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(SystemBus_TLWidthWidget_auto_out_d_bits_size),
    .auto_out_d_bits_source(SystemBus_TLWidthWidget_auto_out_d_bits_source),
    .auto_out_d_bits_data(SystemBus_TLWidthWidget_auto_out_d_bits_data),
    .auto_out_d_bits_error(SystemBus_TLWidthWidget_auto_out_d_bits_error)
  );
  AXI4ToTL AXI4ToTL (
    .clock(AXI4ToTL_clock),
    .reset(AXI4ToTL_reset),
    .auto_in_aw_ready(AXI4ToTL_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4ToTL_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4ToTL_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4ToTL_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4ToTL_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4ToTL_auto_in_aw_bits_size),
    .auto_in_w_ready(AXI4ToTL_auto_in_w_ready),
    .auto_in_w_valid(AXI4ToTL_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4ToTL_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4ToTL_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4ToTL_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4ToTL_auto_in_b_ready),
    .auto_in_b_valid(AXI4ToTL_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4ToTL_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4ToTL_auto_in_b_bits_resp),
    .auto_in_ar_ready(AXI4ToTL_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4ToTL_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4ToTL_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4ToTL_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4ToTL_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4ToTL_auto_in_ar_bits_size),
    .auto_in_r_ready(AXI4ToTL_auto_in_r_ready),
    .auto_in_r_valid(AXI4ToTL_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4ToTL_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4ToTL_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4ToTL_auto_in_r_bits_resp),
    .auto_in_r_bits_last(AXI4ToTL_auto_in_r_bits_last),
    .auto_out_a_ready(AXI4ToTL_auto_out_a_ready),
    .auto_out_a_valid(AXI4ToTL_auto_out_a_valid),
    .auto_out_a_bits_opcode(AXI4ToTL_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(AXI4ToTL_auto_out_a_bits_param),
    .auto_out_a_bits_size(AXI4ToTL_auto_out_a_bits_size),
    .auto_out_a_bits_source(AXI4ToTL_auto_out_a_bits_source),
    .auto_out_a_bits_address(AXI4ToTL_auto_out_a_bits_address),
    .auto_out_a_bits_mask(AXI4ToTL_auto_out_a_bits_mask),
    .auto_out_a_bits_data(AXI4ToTL_auto_out_a_bits_data),
    .auto_out_d_ready(AXI4ToTL_auto_out_d_ready),
    .auto_out_d_valid(AXI4ToTL_auto_out_d_valid),
    .auto_out_d_bits_opcode(AXI4ToTL_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(AXI4ToTL_auto_out_d_bits_size),
    .auto_out_d_bits_source(AXI4ToTL_auto_out_d_bits_source),
    .auto_out_d_bits_data(AXI4ToTL_auto_out_d_bits_data),
    .auto_out_d_bits_error(AXI4ToTL_auto_out_d_bits_error)
  );
  AXI4UserYanker_1 AXI4UserYanker_1 (
    .clock(AXI4UserYanker_1_clock),
    .reset(AXI4UserYanker_1_reset),
    .auto_in_aw_ready(AXI4UserYanker_1_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4UserYanker_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4UserYanker_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4UserYanker_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4UserYanker_1_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4UserYanker_1_auto_in_aw_bits_size),
    .auto_in_aw_bits_user(AXI4UserYanker_1_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4UserYanker_1_auto_in_w_ready),
    .auto_in_w_valid(AXI4UserYanker_1_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4UserYanker_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4UserYanker_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4UserYanker_1_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4UserYanker_1_auto_in_b_ready),
    .auto_in_b_valid(AXI4UserYanker_1_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4UserYanker_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4UserYanker_1_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4UserYanker_1_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4UserYanker_1_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4UserYanker_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4UserYanker_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4UserYanker_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4UserYanker_1_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4UserYanker_1_auto_in_ar_bits_size),
    .auto_in_ar_bits_user(AXI4UserYanker_1_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4UserYanker_1_auto_in_r_ready),
    .auto_in_r_valid(AXI4UserYanker_1_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4UserYanker_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4UserYanker_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4UserYanker_1_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4UserYanker_1_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4UserYanker_1_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4UserYanker_1_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4UserYanker_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4UserYanker_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4UserYanker_1_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4UserYanker_1_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4UserYanker_1_auto_out_aw_bits_size),
    .auto_out_w_ready(AXI4UserYanker_1_auto_out_w_ready),
    .auto_out_w_valid(AXI4UserYanker_1_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4UserYanker_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4UserYanker_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4UserYanker_1_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4UserYanker_1_auto_out_b_ready),
    .auto_out_b_valid(AXI4UserYanker_1_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4UserYanker_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4UserYanker_1_auto_out_b_bits_resp),
    .auto_out_ar_ready(AXI4UserYanker_1_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4UserYanker_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4UserYanker_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4UserYanker_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4UserYanker_1_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4UserYanker_1_auto_out_ar_bits_size),
    .auto_out_r_ready(AXI4UserYanker_1_auto_out_r_ready),
    .auto_out_r_valid(AXI4UserYanker_1_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4UserYanker_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4UserYanker_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4UserYanker_1_auto_out_r_bits_resp),
    .auto_out_r_bits_last(AXI4UserYanker_1_auto_out_r_bits_last)
  );
  AXI4Fragmenter AXI4Fragmenter (
    .clock(AXI4Fragmenter_clock),
    .reset(AXI4Fragmenter_reset),
    .auto_in_aw_ready(AXI4Fragmenter_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Fragmenter_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Fragmenter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Fragmenter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4Fragmenter_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4Fragmenter_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4Fragmenter_auto_in_aw_bits_burst),
    .auto_in_aw_bits_user(AXI4Fragmenter_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4Fragmenter_auto_in_w_ready),
    .auto_in_w_valid(AXI4Fragmenter_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Fragmenter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Fragmenter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Fragmenter_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Fragmenter_auto_in_b_ready),
    .auto_in_b_valid(AXI4Fragmenter_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Fragmenter_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Fragmenter_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4Fragmenter_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4Fragmenter_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Fragmenter_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Fragmenter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Fragmenter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4Fragmenter_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4Fragmenter_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4Fragmenter_auto_in_ar_bits_burst),
    .auto_in_ar_bits_user(AXI4Fragmenter_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4Fragmenter_auto_in_r_ready),
    .auto_in_r_valid(AXI4Fragmenter_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Fragmenter_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Fragmenter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Fragmenter_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4Fragmenter_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4Fragmenter_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Fragmenter_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Fragmenter_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Fragmenter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Fragmenter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4Fragmenter_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4Fragmenter_auto_out_aw_bits_size),
    .auto_out_aw_bits_user(AXI4Fragmenter_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Fragmenter_auto_out_w_ready),
    .auto_out_w_valid(AXI4Fragmenter_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Fragmenter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Fragmenter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4Fragmenter_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4Fragmenter_auto_out_b_ready),
    .auto_out_b_valid(AXI4Fragmenter_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Fragmenter_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Fragmenter_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Fragmenter_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Fragmenter_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Fragmenter_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Fragmenter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Fragmenter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4Fragmenter_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4Fragmenter_auto_out_ar_bits_size),
    .auto_out_ar_bits_user(AXI4Fragmenter_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Fragmenter_auto_out_r_ready),
    .auto_out_r_valid(AXI4Fragmenter_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Fragmenter_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Fragmenter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Fragmenter_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Fragmenter_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4Fragmenter_auto_out_r_bits_last)
  );
  AXI4IdIndexer_1 AXI4IdIndexer_1 (
    .auto_in_aw_ready(AXI4IdIndexer_1_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4IdIndexer_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4IdIndexer_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4IdIndexer_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4IdIndexer_1_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4IdIndexer_1_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4IdIndexer_1_auto_in_aw_bits_burst),
    .auto_in_w_ready(AXI4IdIndexer_1_auto_in_w_ready),
    .auto_in_w_valid(AXI4IdIndexer_1_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4IdIndexer_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4IdIndexer_1_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4IdIndexer_1_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4IdIndexer_1_auto_in_b_ready),
    .auto_in_b_valid(AXI4IdIndexer_1_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4IdIndexer_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4IdIndexer_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(AXI4IdIndexer_1_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4IdIndexer_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4IdIndexer_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4IdIndexer_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4IdIndexer_1_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4IdIndexer_1_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4IdIndexer_1_auto_in_ar_bits_burst),
    .auto_in_r_ready(AXI4IdIndexer_1_auto_in_r_ready),
    .auto_in_r_valid(AXI4IdIndexer_1_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4IdIndexer_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4IdIndexer_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4IdIndexer_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(AXI4IdIndexer_1_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4IdIndexer_1_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4IdIndexer_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4IdIndexer_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4IdIndexer_1_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(AXI4IdIndexer_1_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(AXI4IdIndexer_1_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(AXI4IdIndexer_1_auto_out_aw_bits_burst),
    .auto_out_aw_bits_user(AXI4IdIndexer_1_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4IdIndexer_1_auto_out_w_ready),
    .auto_out_w_valid(AXI4IdIndexer_1_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4IdIndexer_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4IdIndexer_1_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4IdIndexer_1_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4IdIndexer_1_auto_out_b_ready),
    .auto_out_b_valid(AXI4IdIndexer_1_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4IdIndexer_1_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4IdIndexer_1_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4IdIndexer_1_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4IdIndexer_1_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4IdIndexer_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4IdIndexer_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4IdIndexer_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(AXI4IdIndexer_1_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(AXI4IdIndexer_1_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(AXI4IdIndexer_1_auto_out_ar_bits_burst),
    .auto_out_ar_bits_user(AXI4IdIndexer_1_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4IdIndexer_1_auto_out_r_ready),
    .auto_out_r_valid(AXI4IdIndexer_1_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4IdIndexer_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4IdIndexer_1_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4IdIndexer_1_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4IdIndexer_1_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4IdIndexer_1_auto_out_r_bits_last)
  );
  TLROM_bootrom bootrom (
    .auto_in_a_ready(bootrom_auto_in_a_ready),
    .auto_in_a_valid(bootrom_auto_in_a_valid),
    .auto_in_a_bits_size(bootrom_auto_in_a_bits_size),
    .auto_in_a_bits_source(bootrom_auto_in_a_bits_source),
    .auto_in_a_bits_address(bootrom_auto_in_a_bits_address),
    .auto_in_d_ready(bootrom_auto_in_d_ready),
    .auto_in_d_valid(bootrom_auto_in_d_valid),
    .auto_in_d_bits_size(bootrom_auto_in_d_bits_size),
    .auto_in_d_bits_source(bootrom_auto_in_d_bits_source),
    .auto_in_d_bits_data(bootrom_auto_in_d_bits_data)
  );
  TLError_error error (
    .clock(error_clock),
    .reset(error_reset),
    .auto_in_a_ready(error_auto_in_a_ready),
    .auto_in_a_valid(error_auto_in_a_valid),
    .auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(error_auto_in_a_bits_size),
    .auto_in_a_bits_source(error_auto_in_a_bits_source),
    .auto_in_c_ready(error_auto_in_c_ready),
    .auto_in_c_valid(error_auto_in_c_valid),
    .auto_in_c_bits_opcode(error_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(error_auto_in_c_bits_param),
    .auto_in_c_bits_size(error_auto_in_c_bits_size),
    .auto_in_c_bits_source(error_auto_in_c_bits_source),
    .auto_in_d_ready(error_auto_in_d_ready),
    .auto_in_d_valid(error_auto_in_d_valid),
    .auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(error_auto_in_d_bits_param),
    .auto_in_d_bits_size(error_auto_in_d_bits_size),
    .auto_in_d_bits_source(error_auto_in_d_bits_source),
    .auto_in_d_bits_sink(error_auto_in_d_bits_sink),
    .auto_in_d_bits_data(error_auto_in_d_bits_data),
    .auto_in_d_bits_error(error_auto_in_d_bits_error)
  );
  assign int_rtc_tick = value == 7'h63;
  assign _T_244 = value + 7'h1;
  assign _T_245 = _T_244[6:0];
  assign _GEN_0 = int_rtc_tick ? 7'h0 : _T_245;
  assign _T_248 = interrupts[0];
  assign _T_249 = interrupts[1];
  assign debug_clockeddmi_dmi_req_ready = debug_1_io_dmi_dmi_req_ready;
  assign debug_clockeddmi_dmi_resp_valid = debug_1_io_dmi_dmi_resp_valid;
  assign debug_clockeddmi_dmi_resp_bits_data = debug_1_io_dmi_dmi_resp_bits_data;
  assign debug_clockeddmi_dmi_resp_bits_resp = debug_1_io_dmi_dmi_resp_bits_resp;
  assign debug_ndreset = debug_1_io_ctrl_ndreset;
  assign debug_dmactive = debug_1_io_ctrl_dmactive;
  assign mem_axi4_0_aw_valid = _T_39_aw_valid;
  assign mem_axi4_0_aw_bits_id = _T_39_aw_bits_id;
  assign mem_axi4_0_aw_bits_addr = _T_39_aw_bits_addr;
  assign mem_axi4_0_aw_bits_len = _T_39_aw_bits_len;
  assign mem_axi4_0_aw_bits_size = _T_39_aw_bits_size;
  assign mem_axi4_0_aw_bits_burst = _T_39_aw_bits_burst;
  assign mem_axi4_0_aw_bits_lock = _T_39_aw_bits_lock;
  assign mem_axi4_0_aw_bits_cache = _T_39_aw_bits_cache;
  assign mem_axi4_0_aw_bits_prot = _T_39_aw_bits_prot;
  assign mem_axi4_0_aw_bits_qos = _T_39_aw_bits_qos;
  assign mem_axi4_0_w_valid = _T_39_w_valid;
  assign mem_axi4_0_w_bits_data = _T_39_w_bits_data;
  assign mem_axi4_0_w_bits_strb = _T_39_w_bits_strb;
  assign mem_axi4_0_w_bits_last = _T_39_w_bits_last;
  assign mem_axi4_0_b_ready = _T_39_b_ready;
  assign mem_axi4_0_ar_valid = _T_39_ar_valid;
  assign mem_axi4_0_ar_bits_id = _T_39_ar_bits_id;
  assign mem_axi4_0_ar_bits_addr = _T_39_ar_bits_addr;
  assign mem_axi4_0_ar_bits_len = _T_39_ar_bits_len;
  assign mem_axi4_0_ar_bits_size = _T_39_ar_bits_size;
  assign mem_axi4_0_ar_bits_burst = _T_39_ar_bits_burst;
  assign mem_axi4_0_ar_bits_lock = _T_39_ar_bits_lock;
  assign mem_axi4_0_ar_bits_cache = _T_39_ar_bits_cache;
  assign mem_axi4_0_ar_bits_prot = _T_39_ar_bits_prot;
  assign mem_axi4_0_ar_bits_qos = _T_39_ar_bits_qos;
  assign mem_axi4_0_r_ready = _T_39_r_ready;
  assign mmio_axi4_0_aw_valid = _T_97_aw_valid;
  assign mmio_axi4_0_aw_bits_id = _T_97_aw_bits_id;
  assign mmio_axi4_0_aw_bits_addr = _T_97_aw_bits_addr;
  assign mmio_axi4_0_aw_bits_len = _T_97_aw_bits_len;
  assign mmio_axi4_0_aw_bits_size = _T_97_aw_bits_size;
  assign mmio_axi4_0_aw_bits_burst = _T_97_aw_bits_burst;
  assign mmio_axi4_0_aw_bits_lock = _T_97_aw_bits_lock;
  assign mmio_axi4_0_aw_bits_cache = _T_97_aw_bits_cache;
  assign mmio_axi4_0_aw_bits_prot = _T_97_aw_bits_prot;
  assign mmio_axi4_0_aw_bits_qos = _T_97_aw_bits_qos;
  assign mmio_axi4_0_w_valid = _T_97_w_valid;
  assign mmio_axi4_0_w_bits_data = _T_97_w_bits_data;
  assign mmio_axi4_0_w_bits_strb = _T_97_w_bits_strb;
  assign mmio_axi4_0_w_bits_last = _T_97_w_bits_last;
  assign mmio_axi4_0_b_ready = _T_97_b_ready;
  assign mmio_axi4_0_ar_valid = _T_97_ar_valid;
  assign mmio_axi4_0_ar_bits_id = _T_97_ar_bits_id;
  assign mmio_axi4_0_ar_bits_addr = _T_97_ar_bits_addr;
  assign mmio_axi4_0_ar_bits_len = _T_97_ar_bits_len;
  assign mmio_axi4_0_ar_bits_size = _T_97_ar_bits_size;
  assign mmio_axi4_0_ar_bits_burst = _T_97_ar_bits_burst;
  assign mmio_axi4_0_ar_bits_lock = _T_97_ar_bits_lock;
  assign mmio_axi4_0_ar_bits_cache = _T_97_ar_bits_cache;
  assign mmio_axi4_0_ar_bits_prot = _T_97_ar_bits_prot;
  assign mmio_axi4_0_ar_bits_qos = _T_97_ar_bits_qos;
  assign mmio_axi4_0_r_ready = _T_97_r_ready;
  assign l2_frontend_bus_axi4_0_aw_ready = _T_155_aw_ready;
  assign l2_frontend_bus_axi4_0_w_ready = _T_155_w_ready;
  assign l2_frontend_bus_axi4_0_b_valid = _T_155_b_valid;
  assign l2_frontend_bus_axi4_0_b_bits_id = _T_155_b_bits_id;
  assign l2_frontend_bus_axi4_0_b_bits_resp = _T_155_b_bits_resp;
  assign l2_frontend_bus_axi4_0_ar_ready = _T_155_ar_ready;
  assign l2_frontend_bus_axi4_0_r_valid = _T_155_r_valid;
  assign l2_frontend_bus_axi4_0_r_bits_id = _T_155_r_bits_id;
  assign l2_frontend_bus_axi4_0_r_bits_data = _T_155_r_bits_data;
  assign l2_frontend_bus_axi4_0_r_bits_resp = _T_155_r_bits_resp;
  assign l2_frontend_bus_axi4_0_r_bits_last = _T_155_r_bits_last;
  assign IntXbar_auto_int_in_0 = IntXing_auto_int_out_0;
  assign IntXbar_auto_int_in_1 = IntXing_auto_int_out_1;
  assign sbus_clock = clock;
  assign sbus_reset = reset;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_valid = tile_auto_anon_out_a_valid;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_opcode = tile_auto_anon_out_a_bits_opcode;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_param = tile_auto_anon_out_a_bits_param;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_size = tile_auto_anon_out_a_bits_size;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_source = tile_auto_anon_out_a_bits_source;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_address = tile_auto_anon_out_a_bits_address;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_mask = tile_auto_anon_out_a_bits_mask;
  assign sbus_auto_SystemBusFromTiletile_anon_in_a_bits_data = tile_auto_anon_out_a_bits_data;
  assign sbus_auto_SystemBusFromTiletile_anon_in_b_ready = tile_auto_anon_out_b_ready;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_valid = tile_auto_anon_out_c_valid;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_opcode = tile_auto_anon_out_c_bits_opcode;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_param = tile_auto_anon_out_c_bits_param;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_size = tile_auto_anon_out_c_bits_size;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_source = tile_auto_anon_out_c_bits_source;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_address = tile_auto_anon_out_c_bits_address;
  assign sbus_auto_SystemBusFromTiletile_anon_in_c_bits_data = tile_auto_anon_out_c_bits_data;
  assign sbus_auto_SystemBusFromTiletile_anon_in_d_ready = tile_auto_anon_out_d_ready;
  assign sbus_auto_SystemBusFromTiletile_anon_in_e_valid = tile_auto_anon_out_e_valid;
  assign sbus_auto_SystemBusFromTiletile_anon_in_e_bits_sink = tile_auto_anon_out_e_bits_sink;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_ready = pbus_auto_anon_in_a_ready;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_valid = pbus_auto_anon_in_d_valid;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_opcode = pbus_auto_anon_in_d_bits_opcode;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_param = pbus_auto_anon_in_d_bits_param;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_size = pbus_auto_anon_in_d_bits_size;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_source = pbus_auto_anon_in_d_bits_source;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_sink = pbus_auto_anon_in_d_bits_sink;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_data = pbus_auto_anon_in_d_bits_data;
  assign sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_bits_error = pbus_auto_anon_in_d_bits_error;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_valid = SystemBus_TLBuffer_auto_out_a_valid;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_opcode = SystemBus_TLBuffer_auto_out_a_bits_opcode;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_param = SystemBus_TLBuffer_auto_out_a_bits_param;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_size = SystemBus_TLBuffer_auto_out_a_bits_size;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_source = SystemBus_TLBuffer_auto_out_a_bits_source;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_address = SystemBus_TLBuffer_auto_out_a_bits_address;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_mask = SystemBus_TLBuffer_auto_out_a_bits_mask;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_a_bits_data = SystemBus_TLBuffer_auto_out_a_bits_data;
  assign sbus_auto_SystemBus_port_TLFIFOFixer_in_d_ready = SystemBus_TLBuffer_auto_out_d_ready;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_a_ready = TLToAXI4_auto_in_a_ready;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_valid = TLToAXI4_auto_in_d_valid;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_opcode = TLToAXI4_auto_in_d_bits_opcode;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_size = TLToAXI4_auto_in_d_bits_size;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_source = TLToAXI4_auto_in_d_bits_source;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_data = TLToAXI4_auto_in_d_bits_data;
  assign sbus_auto_SystemBus_slave_TLWidthWidget_out_d_bits_error = TLToAXI4_auto_in_d_bits_error;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_a_ready = error_auto_in_a_ready;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_c_ready = error_auto_in_c_ready;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_valid = error_auto_in_d_valid;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_opcode = error_auto_in_d_bits_opcode;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_param = error_auto_in_d_bits_param;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_size = error_auto_in_d_bits_size;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_source = error_auto_in_d_bits_source;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_sink = error_auto_in_d_bits_sink;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_data = error_auto_in_d_bits_data;
  assign sbus_auto_SystemBus_slave_TLBuffer_out_d_bits_error = error_auto_in_d_bits_error;
  assign sbus_auto_SystemBus_out_a_ready = TLBroadcast_auto_in_a_ready;
  assign sbus_auto_SystemBus_out_b_valid = TLBroadcast_auto_in_b_valid;
  assign sbus_auto_SystemBus_out_b_bits_param = TLBroadcast_auto_in_b_bits_param;
  assign sbus_auto_SystemBus_out_b_bits_address = TLBroadcast_auto_in_b_bits_address;
  assign sbus_auto_SystemBus_out_c_ready = TLBroadcast_auto_in_c_ready;
  assign sbus_auto_SystemBus_out_d_valid = TLBroadcast_auto_in_d_valid;
  assign sbus_auto_SystemBus_out_d_bits_opcode = TLBroadcast_auto_in_d_bits_opcode;
  assign sbus_auto_SystemBus_out_d_bits_param = TLBroadcast_auto_in_d_bits_param;
  assign sbus_auto_SystemBus_out_d_bits_size = TLBroadcast_auto_in_d_bits_size;
  assign sbus_auto_SystemBus_out_d_bits_source = TLBroadcast_auto_in_d_bits_source;
  assign sbus_auto_SystemBus_out_d_bits_sink = TLBroadcast_auto_in_d_bits_sink;
  assign sbus_auto_SystemBus_out_d_bits_data = TLBroadcast_auto_in_d_bits_data;
  assign sbus_auto_SystemBus_out_d_bits_error = TLBroadcast_auto_in_d_bits_error;
  assign pbus_clock = clock;
  assign pbus_reset = reset;
  assign pbus_auto_anon_in_a_valid = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_valid;
  assign pbus_auto_anon_in_a_bits_opcode = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_opcode;
  assign pbus_auto_anon_in_a_bits_param = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_param;
  assign pbus_auto_anon_in_a_bits_size = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_size;
  assign pbus_auto_anon_in_a_bits_source = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_source;
  assign pbus_auto_anon_in_a_bits_address = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_address;
  assign pbus_auto_anon_in_a_bits_mask = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_mask;
  assign pbus_auto_anon_in_a_bits_data = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_a_bits_data;
  assign pbus_auto_anon_in_d_ready = sbus_auto_SystemBus_pbus_TLFIFOFixer_out_d_ready;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_ready = bootrom_auto_in_a_ready;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_valid = bootrom_auto_in_d_valid;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_size = bootrom_auto_in_d_bits_size;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_source = bootrom_auto_in_d_bits_source;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_bits_data = bootrom_auto_in_d_bits_data;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_ready = debug_1_auto_dmInner_dmInner_tl_in_a_ready;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_valid = debug_1_auto_dmInner_dmInner_tl_in_d_valid;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_opcode = debug_1_auto_dmInner_dmInner_tl_in_d_bits_opcode;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_size = debug_1_auto_dmInner_dmInner_tl_in_d_bits_size;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_source = debug_1_auto_dmInner_dmInner_tl_in_d_bits_source;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_bits_data = debug_1_auto_dmInner_dmInner_tl_in_d_bits_data;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_ready = clint_auto_in_a_ready;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_valid = clint_auto_in_d_valid;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_opcode = clint_auto_in_d_bits_opcode;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_size = clint_auto_in_d_bits_size;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_source = clint_auto_in_d_bits_source;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_bits_data = clint_auto_in_d_bits_data;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_ready = plic_auto_in_a_ready;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_valid = plic_auto_in_d_valid;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_opcode = plic_auto_in_d_bits_opcode;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_size = plic_auto_in_d_bits_size;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_source = plic_auto_in_d_bits_source;
  assign pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_bits_data = plic_auto_in_d_bits_data;
  assign TLBroadcast_clock = clock;
  assign TLBroadcast_reset = reset;
  assign TLBroadcast_auto_in_a_valid = sbus_auto_SystemBus_out_a_valid;
  assign TLBroadcast_auto_in_a_bits_opcode = sbus_auto_SystemBus_out_a_bits_opcode;
  assign TLBroadcast_auto_in_a_bits_param = sbus_auto_SystemBus_out_a_bits_param;
  assign TLBroadcast_auto_in_a_bits_size = sbus_auto_SystemBus_out_a_bits_size;
  assign TLBroadcast_auto_in_a_bits_source = sbus_auto_SystemBus_out_a_bits_source;
  assign TLBroadcast_auto_in_a_bits_address = sbus_auto_SystemBus_out_a_bits_address;
  assign TLBroadcast_auto_in_a_bits_mask = sbus_auto_SystemBus_out_a_bits_mask;
  assign TLBroadcast_auto_in_a_bits_data = sbus_auto_SystemBus_out_a_bits_data;
  assign TLBroadcast_auto_in_b_ready = sbus_auto_SystemBus_out_b_ready;
  assign TLBroadcast_auto_in_c_valid = sbus_auto_SystemBus_out_c_valid;
  assign TLBroadcast_auto_in_c_bits_opcode = sbus_auto_SystemBus_out_c_bits_opcode;
  assign TLBroadcast_auto_in_c_bits_size = sbus_auto_SystemBus_out_c_bits_size;
  assign TLBroadcast_auto_in_c_bits_source = sbus_auto_SystemBus_out_c_bits_source;
  assign TLBroadcast_auto_in_c_bits_address = sbus_auto_SystemBus_out_c_bits_address;
  assign TLBroadcast_auto_in_c_bits_data = sbus_auto_SystemBus_out_c_bits_data;
  assign TLBroadcast_auto_in_d_ready = sbus_auto_SystemBus_out_d_ready;
  assign TLBroadcast_auto_in_e_valid = sbus_auto_SystemBus_out_e_valid;
  assign TLBroadcast_auto_in_e_bits_sink = sbus_auto_SystemBus_out_e_bits_sink;
  assign TLBroadcast_auto_out_a_ready = TLWidthWidget_auto_in_a_ready;
  assign TLBroadcast_auto_out_d_valid = TLWidthWidget_auto_in_d_valid;
  assign TLBroadcast_auto_out_d_bits_opcode = TLWidthWidget_auto_in_d_bits_opcode;
  assign TLBroadcast_auto_out_d_bits_param = TLWidthWidget_auto_in_d_bits_param;
  assign TLBroadcast_auto_out_d_bits_size = TLWidthWidget_auto_in_d_bits_size;
  assign TLBroadcast_auto_out_d_bits_source = TLWidthWidget_auto_in_d_bits_source;
  assign TLBroadcast_auto_out_d_bits_data = TLWidthWidget_auto_in_d_bits_data;
  assign TLBroadcast_auto_out_d_bits_error = TLWidthWidget_auto_in_d_bits_error;
  assign TLWidthWidget_auto_in_a_valid = TLBroadcast_auto_out_a_valid;
  assign TLWidthWidget_auto_in_a_bits_opcode = TLBroadcast_auto_out_a_bits_opcode;
  assign TLWidthWidget_auto_in_a_bits_size = TLBroadcast_auto_out_a_bits_size;
  assign TLWidthWidget_auto_in_a_bits_source = TLBroadcast_auto_out_a_bits_source;
  assign TLWidthWidget_auto_in_a_bits_address = TLBroadcast_auto_out_a_bits_address;
  assign TLWidthWidget_auto_in_a_bits_mask = TLBroadcast_auto_out_a_bits_mask;
  assign TLWidthWidget_auto_in_a_bits_data = TLBroadcast_auto_out_a_bits_data;
  assign TLWidthWidget_auto_in_d_ready = TLBroadcast_auto_out_d_ready;
  assign TLWidthWidget_auto_out_a_ready = TLFilter_auto_in_a_ready;
  assign TLWidthWidget_auto_out_d_valid = TLFilter_auto_in_d_valid;
  assign TLWidthWidget_auto_out_d_bits_opcode = TLFilter_auto_in_d_bits_opcode;
  assign TLWidthWidget_auto_out_d_bits_param = TLFilter_auto_in_d_bits_param;
  assign TLWidthWidget_auto_out_d_bits_size = TLFilter_auto_in_d_bits_size;
  assign TLWidthWidget_auto_out_d_bits_source = TLFilter_auto_in_d_bits_source;
  assign TLWidthWidget_auto_out_d_bits_data = TLFilter_auto_in_d_bits_data;
  assign TLWidthWidget_auto_out_d_bits_error = TLFilter_auto_in_d_bits_error;
  assign memBuses_0_clock = clock;
  assign memBuses_0_reset = reset;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_ready = converter_auto_in_a_ready;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_valid = converter_auto_in_d_valid;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_opcode = converter_auto_in_d_bits_opcode;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_size = converter_auto_in_d_bits_size;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_source = converter_auto_in_d_bits_source;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_data = converter_auto_in_d_bits_data;
  assign memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_bits_error = converter_auto_in_d_bits_error;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_valid = TLFilter_auto_out_a_valid;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_opcode = TLFilter_auto_out_a_bits_opcode;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_size = TLFilter_auto_out_a_bits_size;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_source = TLFilter_auto_out_a_bits_source;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_address = TLFilter_auto_out_a_bits_address;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_mask = TLFilter_auto_out_a_bits_mask;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_bits_data = TLFilter_auto_out_a_bits_data;
  assign memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_ready = TLFilter_auto_out_d_ready;
  assign TLFilter_auto_in_a_valid = TLWidthWidget_auto_out_a_valid;
  assign TLFilter_auto_in_a_bits_opcode = TLWidthWidget_auto_out_a_bits_opcode;
  assign TLFilter_auto_in_a_bits_size = TLWidthWidget_auto_out_a_bits_size;
  assign TLFilter_auto_in_a_bits_source = TLWidthWidget_auto_out_a_bits_source;
  assign TLFilter_auto_in_a_bits_address = TLWidthWidget_auto_out_a_bits_address;
  assign TLFilter_auto_in_a_bits_mask = TLWidthWidget_auto_out_a_bits_mask;
  assign TLFilter_auto_in_a_bits_data = TLWidthWidget_auto_out_a_bits_data;
  assign TLFilter_auto_in_d_ready = TLWidthWidget_auto_out_d_ready;
  assign TLFilter_auto_out_a_ready = memBuses_0_auto_MemoryBus_master_TLBuffer_in_a_ready;
  assign TLFilter_auto_out_d_valid = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_valid;
  assign TLFilter_auto_out_d_bits_opcode = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_opcode;
  assign TLFilter_auto_out_d_bits_param = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_param;
  assign TLFilter_auto_out_d_bits_size = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_size;
  assign TLFilter_auto_out_d_bits_source = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_source;
  assign TLFilter_auto_out_d_bits_data = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_data;
  assign TLFilter_auto_out_d_bits_error = memBuses_0_auto_MemoryBus_master_TLBuffer_in_d_bits_error;
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_auto_int_in_0 = IntXbar_auto_int_out_0;
  assign plic_auto_int_in_1 = IntXbar_auto_int_out_1;
  assign plic_auto_in_a_valid = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_valid;
  assign plic_auto_in_a_bits_opcode = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_opcode;
  assign plic_auto_in_a_bits_size = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_size;
  assign plic_auto_in_a_bits_source = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_source;
  assign plic_auto_in_a_bits_address = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_address;
  assign plic_auto_in_a_bits_mask = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_mask;
  assign plic_auto_in_a_bits_data = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_a_bits_data;
  assign plic_auto_in_d_ready = pbus_auto_PeripheryBus_slave_TLFragmenter_out_0_d_ready;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_auto_in_a_valid = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_valid;
  assign clint_auto_in_a_bits_opcode = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_opcode;
  assign clint_auto_in_a_bits_size = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_size;
  assign clint_auto_in_a_bits_source = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_source;
  assign clint_auto_in_a_bits_address = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_address;
  assign clint_auto_in_a_bits_mask = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_mask;
  assign clint_auto_in_a_bits_data = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_a_bits_data;
  assign clint_auto_in_d_ready = pbus_auto_PeripheryBus_slave_TLFragmenter_out_1_d_ready;
  assign clint_io_rtcTick = int_rtc_tick;
  assign debug_1_clock = clock;
  assign debug_1_reset = reset;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_valid = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_valid;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_opcode = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_opcode;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_size = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_size;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_source = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_source;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_address = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_address;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_mask = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_mask;
  assign debug_1_auto_dmInner_dmInner_tl_in_a_bits_data = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_a_bits_data;
  assign debug_1_auto_dmInner_dmInner_tl_in_d_ready = pbus_auto_PeripheryBus_slave_TLFragmenter_out_2_d_ready;
  assign debug_1_io_dmi_dmi_req_valid = debug_clockeddmi_dmi_req_valid;
  assign debug_1_io_dmi_dmi_req_bits_addr = debug_clockeddmi_dmi_req_bits_addr;
  assign debug_1_io_dmi_dmi_req_bits_data = debug_clockeddmi_dmi_req_bits_data;
  assign debug_1_io_dmi_dmi_req_bits_op = debug_clockeddmi_dmi_req_bits_op;
  assign debug_1_io_dmi_dmi_resp_ready = debug_clockeddmi_dmi_resp_ready;
  assign debug_1_io_dmi_dmiClock = debug_clockeddmi_dmiClock;
  assign debug_1_io_dmi_dmiReset = debug_clockeddmi_dmiReset;
  assign tile_clock = tile_inputs_0_clock;
  assign tile_reset = tile_inputs_0_reset;
  assign tile_auto_anon_in_3_sync_0 = IntSyncCrossingSource_auto_out_2_sync_0;
  assign tile_auto_anon_in_2_sync_0 = IntSyncCrossingSource_auto_out_1_sync_0;
  assign tile_auto_anon_in_1_sync_0 = IntSyncCrossingSource_auto_out_0_sync_0;
  assign tile_auto_anon_in_1_sync_1 = IntSyncCrossingSource_auto_out_0_sync_1;
  assign tile_auto_anon_in_0_sync_0 = debug_1_auto_dmOuter_anon_out_sync_0;
  assign tile_auto_anon_out_a_ready = sbus_auto_SystemBusFromTiletile_anon_in_a_ready;
  assign tile_auto_anon_out_b_valid = sbus_auto_SystemBusFromTiletile_anon_in_b_valid;
  assign tile_auto_anon_out_b_bits_param = sbus_auto_SystemBusFromTiletile_anon_in_b_bits_param;
  assign tile_auto_anon_out_b_bits_size = sbus_auto_SystemBusFromTiletile_anon_in_b_bits_size;
  assign tile_auto_anon_out_b_bits_source = sbus_auto_SystemBusFromTiletile_anon_in_b_bits_source;
  assign tile_auto_anon_out_b_bits_address = sbus_auto_SystemBusFromTiletile_anon_in_b_bits_address;
  assign tile_auto_anon_out_c_ready = sbus_auto_SystemBusFromTiletile_anon_in_c_ready;
  assign tile_auto_anon_out_d_valid = sbus_auto_SystemBusFromTiletile_anon_in_d_valid;
  assign tile_auto_anon_out_d_bits_opcode = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_opcode;
  assign tile_auto_anon_out_d_bits_param = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_param;
  assign tile_auto_anon_out_d_bits_size = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_size;
  assign tile_auto_anon_out_d_bits_source = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_source;
  assign tile_auto_anon_out_d_bits_sink = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_sink;
  assign tile_auto_anon_out_d_bits_data = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_data;
  assign tile_auto_anon_out_d_bits_error = sbus_auto_SystemBusFromTiletile_anon_in_d_bits_error;
  assign tile_auto_anon_out_e_ready = sbus_auto_SystemBusFromTiletile_anon_in_e_ready;
  assign IntSyncCrossingSource_clock = clock;
  assign IntSyncCrossingSource_reset = reset;
  assign IntSyncCrossingSource_auto_in_2_0 = plic_auto_int_out_1_0;
  assign IntSyncCrossingSource_auto_in_1_0 = plic_auto_int_out_0_0;
  assign IntSyncCrossingSource_auto_in_0_0 = clint_auto_int_out_0;
  assign IntSyncCrossingSource_auto_in_0_1 = clint_auto_int_out_1;
  assign IntXing_clock = clock;
  assign IntXing_auto_int_in_0 = _T_5_0;
  assign IntXing_auto_int_in_1 = _T_5_1;
  assign converter_clock = clock;
  assign converter_reset = reset;
  assign converter_auto_in_a_valid = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_valid;
  assign converter_auto_in_a_bits_opcode = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_opcode;
  assign converter_auto_in_a_bits_size = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_size;
  assign converter_auto_in_a_bits_source = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_source;
  assign converter_auto_in_a_bits_address = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_address;
  assign converter_auto_in_a_bits_mask = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_mask;
  assign converter_auto_in_a_bits_data = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_a_bits_data;
  assign converter_auto_in_d_ready = memBuses_0_auto_MemoryBus_slave_TLBuffer_out_d_ready;
  assign converter_auto_out_aw_ready = trim_auto_in_aw_ready;
  assign converter_auto_out_w_ready = trim_auto_in_w_ready;
  assign converter_auto_out_b_valid = trim_auto_in_b_valid;
  assign converter_auto_out_b_bits_id = trim_auto_in_b_bits_id;
  assign converter_auto_out_b_bits_resp = trim_auto_in_b_bits_resp;
  assign converter_auto_out_b_bits_user = trim_auto_in_b_bits_user;
  assign converter_auto_out_ar_ready = trim_auto_in_ar_ready;
  assign converter_auto_out_r_valid = trim_auto_in_r_valid;
  assign converter_auto_out_r_bits_id = trim_auto_in_r_bits_id;
  assign converter_auto_out_r_bits_data = trim_auto_in_r_bits_data;
  assign converter_auto_out_r_bits_resp = trim_auto_in_r_bits_resp;
  assign converter_auto_out_r_bits_user = trim_auto_in_r_bits_user;
  assign converter_auto_out_r_bits_last = trim_auto_in_r_bits_last;
  assign trim_auto_in_aw_valid = converter_auto_out_aw_valid;
  assign trim_auto_in_aw_bits_id = converter_auto_out_aw_bits_id;
  assign trim_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr;
  assign trim_auto_in_aw_bits_len = converter_auto_out_aw_bits_len;
  assign trim_auto_in_aw_bits_size = converter_auto_out_aw_bits_size;
  assign trim_auto_in_aw_bits_burst = converter_auto_out_aw_bits_burst;
  assign trim_auto_in_aw_bits_lock = converter_auto_out_aw_bits_lock;
  assign trim_auto_in_aw_bits_cache = converter_auto_out_aw_bits_cache;
  assign trim_auto_in_aw_bits_prot = converter_auto_out_aw_bits_prot;
  assign trim_auto_in_aw_bits_qos = converter_auto_out_aw_bits_qos;
  assign trim_auto_in_aw_bits_user = converter_auto_out_aw_bits_user;
  assign trim_auto_in_w_valid = converter_auto_out_w_valid;
  assign trim_auto_in_w_bits_data = converter_auto_out_w_bits_data;
  assign trim_auto_in_w_bits_strb = converter_auto_out_w_bits_strb;
  assign trim_auto_in_w_bits_last = converter_auto_out_w_bits_last;
  assign trim_auto_in_b_ready = converter_auto_out_b_ready;
  assign trim_auto_in_ar_valid = converter_auto_out_ar_valid;
  assign trim_auto_in_ar_bits_id = converter_auto_out_ar_bits_id;
  assign trim_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr;
  assign trim_auto_in_ar_bits_len = converter_auto_out_ar_bits_len;
  assign trim_auto_in_ar_bits_size = converter_auto_out_ar_bits_size;
  assign trim_auto_in_ar_bits_burst = converter_auto_out_ar_bits_burst;
  assign trim_auto_in_ar_bits_lock = converter_auto_out_ar_bits_lock;
  assign trim_auto_in_ar_bits_cache = converter_auto_out_ar_bits_cache;
  assign trim_auto_in_ar_bits_prot = converter_auto_out_ar_bits_prot;
  assign trim_auto_in_ar_bits_qos = converter_auto_out_ar_bits_qos;
  assign trim_auto_in_ar_bits_user = converter_auto_out_ar_bits_user;
  assign trim_auto_in_r_ready = converter_auto_out_r_ready;
  assign trim_auto_out_aw_ready = yank_auto_in_aw_ready;
  assign trim_auto_out_w_ready = yank_auto_in_w_ready;
  assign trim_auto_out_b_valid = yank_auto_in_b_valid;
  assign trim_auto_out_b_bits_id = yank_auto_in_b_bits_id;
  assign trim_auto_out_b_bits_resp = yank_auto_in_b_bits_resp;
  assign trim_auto_out_b_bits_user = yank_auto_in_b_bits_user;
  assign trim_auto_out_ar_ready = yank_auto_in_ar_ready;
  assign trim_auto_out_r_valid = yank_auto_in_r_valid;
  assign trim_auto_out_r_bits_id = yank_auto_in_r_bits_id;
  assign trim_auto_out_r_bits_data = yank_auto_in_r_bits_data;
  assign trim_auto_out_r_bits_resp = yank_auto_in_r_bits_resp;
  assign trim_auto_out_r_bits_user = yank_auto_in_r_bits_user;
  assign trim_auto_out_r_bits_last = yank_auto_in_r_bits_last;
  assign yank_clock = clock;
  assign yank_reset = reset;
  assign yank_auto_in_aw_valid = trim_auto_out_aw_valid;
  assign yank_auto_in_aw_bits_id = trim_auto_out_aw_bits_id;
  assign yank_auto_in_aw_bits_addr = trim_auto_out_aw_bits_addr;
  assign yank_auto_in_aw_bits_len = trim_auto_out_aw_bits_len;
  assign yank_auto_in_aw_bits_size = trim_auto_out_aw_bits_size;
  assign yank_auto_in_aw_bits_burst = trim_auto_out_aw_bits_burst;
  assign yank_auto_in_aw_bits_lock = trim_auto_out_aw_bits_lock;
  assign yank_auto_in_aw_bits_cache = trim_auto_out_aw_bits_cache;
  assign yank_auto_in_aw_bits_prot = trim_auto_out_aw_bits_prot;
  assign yank_auto_in_aw_bits_qos = trim_auto_out_aw_bits_qos;
  assign yank_auto_in_aw_bits_user = trim_auto_out_aw_bits_user;
  assign yank_auto_in_w_valid = trim_auto_out_w_valid;
  assign yank_auto_in_w_bits_data = trim_auto_out_w_bits_data;
  assign yank_auto_in_w_bits_strb = trim_auto_out_w_bits_strb;
  assign yank_auto_in_w_bits_last = trim_auto_out_w_bits_last;
  assign yank_auto_in_b_ready = trim_auto_out_b_ready;
  assign yank_auto_in_ar_valid = trim_auto_out_ar_valid;
  assign yank_auto_in_ar_bits_id = trim_auto_out_ar_bits_id;
  assign yank_auto_in_ar_bits_addr = trim_auto_out_ar_bits_addr;
  assign yank_auto_in_ar_bits_len = trim_auto_out_ar_bits_len;
  assign yank_auto_in_ar_bits_size = trim_auto_out_ar_bits_size;
  assign yank_auto_in_ar_bits_burst = trim_auto_out_ar_bits_burst;
  assign yank_auto_in_ar_bits_lock = trim_auto_out_ar_bits_lock;
  assign yank_auto_in_ar_bits_cache = trim_auto_out_ar_bits_cache;
  assign yank_auto_in_ar_bits_prot = trim_auto_out_ar_bits_prot;
  assign yank_auto_in_ar_bits_qos = trim_auto_out_ar_bits_qos;
  assign yank_auto_in_ar_bits_user = trim_auto_out_ar_bits_user;
  assign yank_auto_in_r_ready = trim_auto_out_r_ready;
  assign yank_auto_out_aw_ready = buffer_auto_in_aw_ready;
  assign yank_auto_out_w_ready = buffer_auto_in_w_ready;
  assign yank_auto_out_b_valid = buffer_auto_in_b_valid;
  assign yank_auto_out_b_bits_id = buffer_auto_in_b_bits_id;
  assign yank_auto_out_b_bits_resp = buffer_auto_in_b_bits_resp;
  assign yank_auto_out_ar_ready = buffer_auto_in_ar_ready;
  assign yank_auto_out_r_valid = buffer_auto_in_r_valid;
  assign yank_auto_out_r_bits_id = buffer_auto_in_r_bits_id;
  assign yank_auto_out_r_bits_data = buffer_auto_in_r_bits_data;
  assign yank_auto_out_r_bits_resp = buffer_auto_in_r_bits_resp;
  assign yank_auto_out_r_bits_last = buffer_auto_in_r_bits_last;
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_aw_valid = yank_auto_out_aw_valid;
  assign buffer_auto_in_aw_bits_id = yank_auto_out_aw_bits_id;
  assign buffer_auto_in_aw_bits_addr = yank_auto_out_aw_bits_addr;
  assign buffer_auto_in_aw_bits_len = yank_auto_out_aw_bits_len;
  assign buffer_auto_in_aw_bits_size = yank_auto_out_aw_bits_size;
  assign buffer_auto_in_aw_bits_burst = yank_auto_out_aw_bits_burst;
  assign buffer_auto_in_aw_bits_lock = yank_auto_out_aw_bits_lock;
  assign buffer_auto_in_aw_bits_cache = yank_auto_out_aw_bits_cache;
  assign buffer_auto_in_aw_bits_prot = yank_auto_out_aw_bits_prot;
  assign buffer_auto_in_aw_bits_qos = yank_auto_out_aw_bits_qos;
  assign buffer_auto_in_w_valid = yank_auto_out_w_valid;
  assign buffer_auto_in_w_bits_data = yank_auto_out_w_bits_data;
  assign buffer_auto_in_w_bits_strb = yank_auto_out_w_bits_strb;
  assign buffer_auto_in_w_bits_last = yank_auto_out_w_bits_last;
  assign buffer_auto_in_b_ready = yank_auto_out_b_ready;
  assign buffer_auto_in_ar_valid = yank_auto_out_ar_valid;
  assign buffer_auto_in_ar_bits_id = yank_auto_out_ar_bits_id;
  assign buffer_auto_in_ar_bits_addr = yank_auto_out_ar_bits_addr;
  assign buffer_auto_in_ar_bits_len = yank_auto_out_ar_bits_len;
  assign buffer_auto_in_ar_bits_size = yank_auto_out_ar_bits_size;
  assign buffer_auto_in_ar_bits_burst = yank_auto_out_ar_bits_burst;
  assign buffer_auto_in_ar_bits_lock = yank_auto_out_ar_bits_lock;
  assign buffer_auto_in_ar_bits_cache = yank_auto_out_ar_bits_cache;
  assign buffer_auto_in_ar_bits_prot = yank_auto_out_ar_bits_prot;
  assign buffer_auto_in_ar_bits_qos = yank_auto_out_ar_bits_qos;
  assign buffer_auto_in_r_ready = yank_auto_out_r_ready;
  assign buffer_auto_out_aw_ready = _T_39_aw_ready;
  assign buffer_auto_out_w_ready = _T_39_w_ready;
  assign buffer_auto_out_b_valid = _T_39_b_valid;
  assign buffer_auto_out_b_bits_id = _T_39_b_bits_id;
  assign buffer_auto_out_b_bits_resp = _T_39_b_bits_resp;
  assign buffer_auto_out_ar_ready = _T_39_ar_ready;
  assign buffer_auto_out_r_valid = _T_39_r_valid;
  assign buffer_auto_out_r_bits_id = _T_39_r_bits_id;
  assign buffer_auto_out_r_bits_data = _T_39_r_bits_data;
  assign buffer_auto_out_r_bits_resp = _T_39_r_bits_resp;
  assign buffer_auto_out_r_bits_last = _T_39_r_bits_last;
  assign AXI4Buffer_clock = clock;
  assign AXI4Buffer_reset = reset;
  assign AXI4Buffer_auto_in_aw_valid = AXI4UserYanker_auto_out_aw_valid;
  assign AXI4Buffer_auto_in_aw_bits_id = AXI4UserYanker_auto_out_aw_bits_id;
  assign AXI4Buffer_auto_in_aw_bits_addr = AXI4UserYanker_auto_out_aw_bits_addr;
  assign AXI4Buffer_auto_in_aw_bits_len = AXI4UserYanker_auto_out_aw_bits_len;
  assign AXI4Buffer_auto_in_aw_bits_size = AXI4UserYanker_auto_out_aw_bits_size;
  assign AXI4Buffer_auto_in_aw_bits_burst = AXI4UserYanker_auto_out_aw_bits_burst;
  assign AXI4Buffer_auto_in_aw_bits_lock = AXI4UserYanker_auto_out_aw_bits_lock;
  assign AXI4Buffer_auto_in_aw_bits_cache = AXI4UserYanker_auto_out_aw_bits_cache;
  assign AXI4Buffer_auto_in_aw_bits_prot = AXI4UserYanker_auto_out_aw_bits_prot;
  assign AXI4Buffer_auto_in_aw_bits_qos = AXI4UserYanker_auto_out_aw_bits_qos;
  assign AXI4Buffer_auto_in_w_valid = AXI4UserYanker_auto_out_w_valid;
  assign AXI4Buffer_auto_in_w_bits_data = AXI4UserYanker_auto_out_w_bits_data;
  assign AXI4Buffer_auto_in_w_bits_strb = AXI4UserYanker_auto_out_w_bits_strb;
  assign AXI4Buffer_auto_in_w_bits_last = AXI4UserYanker_auto_out_w_bits_last;
  assign AXI4Buffer_auto_in_b_ready = AXI4UserYanker_auto_out_b_ready;
  assign AXI4Buffer_auto_in_ar_valid = AXI4UserYanker_auto_out_ar_valid;
  assign AXI4Buffer_auto_in_ar_bits_id = AXI4UserYanker_auto_out_ar_bits_id;
  assign AXI4Buffer_auto_in_ar_bits_addr = AXI4UserYanker_auto_out_ar_bits_addr;
  assign AXI4Buffer_auto_in_ar_bits_len = AXI4UserYanker_auto_out_ar_bits_len;
  assign AXI4Buffer_auto_in_ar_bits_size = AXI4UserYanker_auto_out_ar_bits_size;
  assign AXI4Buffer_auto_in_ar_bits_burst = AXI4UserYanker_auto_out_ar_bits_burst;
  assign AXI4Buffer_auto_in_ar_bits_lock = AXI4UserYanker_auto_out_ar_bits_lock;
  assign AXI4Buffer_auto_in_ar_bits_cache = AXI4UserYanker_auto_out_ar_bits_cache;
  assign AXI4Buffer_auto_in_ar_bits_prot = AXI4UserYanker_auto_out_ar_bits_prot;
  assign AXI4Buffer_auto_in_ar_bits_qos = AXI4UserYanker_auto_out_ar_bits_qos;
  assign AXI4Buffer_auto_in_r_ready = AXI4UserYanker_auto_out_r_ready;
  assign AXI4Buffer_auto_out_aw_ready = _T_97_aw_ready;
  assign AXI4Buffer_auto_out_w_ready = _T_97_w_ready;
  assign AXI4Buffer_auto_out_b_valid = _T_97_b_valid;
  assign AXI4Buffer_auto_out_b_bits_id = _T_97_b_bits_id;
  assign AXI4Buffer_auto_out_b_bits_resp = _T_97_b_bits_resp;
  assign AXI4Buffer_auto_out_ar_ready = _T_97_ar_ready;
  assign AXI4Buffer_auto_out_r_valid = _T_97_r_valid;
  assign AXI4Buffer_auto_out_r_bits_id = _T_97_r_bits_id;
  assign AXI4Buffer_auto_out_r_bits_data = _T_97_r_bits_data;
  assign AXI4Buffer_auto_out_r_bits_resp = _T_97_r_bits_resp;
  assign AXI4Buffer_auto_out_r_bits_last = _T_97_r_bits_last;
  assign AXI4UserYanker_clock = clock;
  assign AXI4UserYanker_reset = reset;
  assign AXI4UserYanker_auto_in_aw_valid = AXI4Deinterleaver_auto_out_aw_valid;
  assign AXI4UserYanker_auto_in_aw_bits_id = AXI4Deinterleaver_auto_out_aw_bits_id;
  assign AXI4UserYanker_auto_in_aw_bits_addr = AXI4Deinterleaver_auto_out_aw_bits_addr;
  assign AXI4UserYanker_auto_in_aw_bits_len = AXI4Deinterleaver_auto_out_aw_bits_len;
  assign AXI4UserYanker_auto_in_aw_bits_size = AXI4Deinterleaver_auto_out_aw_bits_size;
  assign AXI4UserYanker_auto_in_aw_bits_burst = AXI4Deinterleaver_auto_out_aw_bits_burst;
  assign AXI4UserYanker_auto_in_aw_bits_lock = AXI4Deinterleaver_auto_out_aw_bits_lock;
  assign AXI4UserYanker_auto_in_aw_bits_cache = AXI4Deinterleaver_auto_out_aw_bits_cache;
  assign AXI4UserYanker_auto_in_aw_bits_prot = AXI4Deinterleaver_auto_out_aw_bits_prot;
  assign AXI4UserYanker_auto_in_aw_bits_qos = AXI4Deinterleaver_auto_out_aw_bits_qos;
  assign AXI4UserYanker_auto_in_aw_bits_user = AXI4Deinterleaver_auto_out_aw_bits_user;
  assign AXI4UserYanker_auto_in_w_valid = AXI4Deinterleaver_auto_out_w_valid;
  assign AXI4UserYanker_auto_in_w_bits_data = AXI4Deinterleaver_auto_out_w_bits_data;
  assign AXI4UserYanker_auto_in_w_bits_strb = AXI4Deinterleaver_auto_out_w_bits_strb;
  assign AXI4UserYanker_auto_in_w_bits_last = AXI4Deinterleaver_auto_out_w_bits_last;
  assign AXI4UserYanker_auto_in_b_ready = AXI4Deinterleaver_auto_out_b_ready;
  assign AXI4UserYanker_auto_in_ar_valid = AXI4Deinterleaver_auto_out_ar_valid;
  assign AXI4UserYanker_auto_in_ar_bits_id = AXI4Deinterleaver_auto_out_ar_bits_id;
  assign AXI4UserYanker_auto_in_ar_bits_addr = AXI4Deinterleaver_auto_out_ar_bits_addr;
  assign AXI4UserYanker_auto_in_ar_bits_len = AXI4Deinterleaver_auto_out_ar_bits_len;
  assign AXI4UserYanker_auto_in_ar_bits_size = AXI4Deinterleaver_auto_out_ar_bits_size;
  assign AXI4UserYanker_auto_in_ar_bits_burst = AXI4Deinterleaver_auto_out_ar_bits_burst;
  assign AXI4UserYanker_auto_in_ar_bits_lock = AXI4Deinterleaver_auto_out_ar_bits_lock;
  assign AXI4UserYanker_auto_in_ar_bits_cache = AXI4Deinterleaver_auto_out_ar_bits_cache;
  assign AXI4UserYanker_auto_in_ar_bits_prot = AXI4Deinterleaver_auto_out_ar_bits_prot;
  assign AXI4UserYanker_auto_in_ar_bits_qos = AXI4Deinterleaver_auto_out_ar_bits_qos;
  assign AXI4UserYanker_auto_in_ar_bits_user = AXI4Deinterleaver_auto_out_ar_bits_user;
  assign AXI4UserYanker_auto_in_r_ready = AXI4Deinterleaver_auto_out_r_ready;
  assign AXI4UserYanker_auto_out_aw_ready = AXI4Buffer_auto_in_aw_ready;
  assign AXI4UserYanker_auto_out_w_ready = AXI4Buffer_auto_in_w_ready;
  assign AXI4UserYanker_auto_out_b_valid = AXI4Buffer_auto_in_b_valid;
  assign AXI4UserYanker_auto_out_b_bits_id = AXI4Buffer_auto_in_b_bits_id;
  assign AXI4UserYanker_auto_out_b_bits_resp = AXI4Buffer_auto_in_b_bits_resp;
  assign AXI4UserYanker_auto_out_ar_ready = AXI4Buffer_auto_in_ar_ready;
  assign AXI4UserYanker_auto_out_r_valid = AXI4Buffer_auto_in_r_valid;
  assign AXI4UserYanker_auto_out_r_bits_id = AXI4Buffer_auto_in_r_bits_id;
  assign AXI4UserYanker_auto_out_r_bits_data = AXI4Buffer_auto_in_r_bits_data;
  assign AXI4UserYanker_auto_out_r_bits_resp = AXI4Buffer_auto_in_r_bits_resp;
  assign AXI4UserYanker_auto_out_r_bits_last = AXI4Buffer_auto_in_r_bits_last;
  assign AXI4Deinterleaver_clock = clock;
  assign AXI4Deinterleaver_reset = reset;
  assign AXI4Deinterleaver_auto_in_aw_valid = AXI4IdIndexer_auto_out_aw_valid;
  assign AXI4Deinterleaver_auto_in_aw_bits_id = AXI4IdIndexer_auto_out_aw_bits_id;
  assign AXI4Deinterleaver_auto_in_aw_bits_addr = AXI4IdIndexer_auto_out_aw_bits_addr;
  assign AXI4Deinterleaver_auto_in_aw_bits_len = AXI4IdIndexer_auto_out_aw_bits_len;
  assign AXI4Deinterleaver_auto_in_aw_bits_size = AXI4IdIndexer_auto_out_aw_bits_size;
  assign AXI4Deinterleaver_auto_in_aw_bits_burst = AXI4IdIndexer_auto_out_aw_bits_burst;
  assign AXI4Deinterleaver_auto_in_aw_bits_lock = AXI4IdIndexer_auto_out_aw_bits_lock;
  assign AXI4Deinterleaver_auto_in_aw_bits_cache = AXI4IdIndexer_auto_out_aw_bits_cache;
  assign AXI4Deinterleaver_auto_in_aw_bits_prot = AXI4IdIndexer_auto_out_aw_bits_prot;
  assign AXI4Deinterleaver_auto_in_aw_bits_qos = AXI4IdIndexer_auto_out_aw_bits_qos;
  assign AXI4Deinterleaver_auto_in_aw_bits_user = AXI4IdIndexer_auto_out_aw_bits_user;
  assign AXI4Deinterleaver_auto_in_w_valid = AXI4IdIndexer_auto_out_w_valid;
  assign AXI4Deinterleaver_auto_in_w_bits_data = AXI4IdIndexer_auto_out_w_bits_data;
  assign AXI4Deinterleaver_auto_in_w_bits_strb = AXI4IdIndexer_auto_out_w_bits_strb;
  assign AXI4Deinterleaver_auto_in_w_bits_last = AXI4IdIndexer_auto_out_w_bits_last;
  assign AXI4Deinterleaver_auto_in_b_ready = AXI4IdIndexer_auto_out_b_ready;
  assign AXI4Deinterleaver_auto_in_ar_valid = AXI4IdIndexer_auto_out_ar_valid;
  assign AXI4Deinterleaver_auto_in_ar_bits_id = AXI4IdIndexer_auto_out_ar_bits_id;
  assign AXI4Deinterleaver_auto_in_ar_bits_addr = AXI4IdIndexer_auto_out_ar_bits_addr;
  assign AXI4Deinterleaver_auto_in_ar_bits_len = AXI4IdIndexer_auto_out_ar_bits_len;
  assign AXI4Deinterleaver_auto_in_ar_bits_size = AXI4IdIndexer_auto_out_ar_bits_size;
  assign AXI4Deinterleaver_auto_in_ar_bits_burst = AXI4IdIndexer_auto_out_ar_bits_burst;
  assign AXI4Deinterleaver_auto_in_ar_bits_lock = AXI4IdIndexer_auto_out_ar_bits_lock;
  assign AXI4Deinterleaver_auto_in_ar_bits_cache = AXI4IdIndexer_auto_out_ar_bits_cache;
  assign AXI4Deinterleaver_auto_in_ar_bits_prot = AXI4IdIndexer_auto_out_ar_bits_prot;
  assign AXI4Deinterleaver_auto_in_ar_bits_qos = AXI4IdIndexer_auto_out_ar_bits_qos;
  assign AXI4Deinterleaver_auto_in_ar_bits_user = AXI4IdIndexer_auto_out_ar_bits_user;
  assign AXI4Deinterleaver_auto_in_r_ready = AXI4IdIndexer_auto_out_r_ready;
  assign AXI4Deinterleaver_auto_out_aw_ready = AXI4UserYanker_auto_in_aw_ready;
  assign AXI4Deinterleaver_auto_out_w_ready = AXI4UserYanker_auto_in_w_ready;
  assign AXI4Deinterleaver_auto_out_b_valid = AXI4UserYanker_auto_in_b_valid;
  assign AXI4Deinterleaver_auto_out_b_bits_id = AXI4UserYanker_auto_in_b_bits_id;
  assign AXI4Deinterleaver_auto_out_b_bits_resp = AXI4UserYanker_auto_in_b_bits_resp;
  assign AXI4Deinterleaver_auto_out_b_bits_user = AXI4UserYanker_auto_in_b_bits_user;
  assign AXI4Deinterleaver_auto_out_ar_ready = AXI4UserYanker_auto_in_ar_ready;
  assign AXI4Deinterleaver_auto_out_r_valid = AXI4UserYanker_auto_in_r_valid;
  assign AXI4Deinterleaver_auto_out_r_bits_id = AXI4UserYanker_auto_in_r_bits_id;
  assign AXI4Deinterleaver_auto_out_r_bits_data = AXI4UserYanker_auto_in_r_bits_data;
  assign AXI4Deinterleaver_auto_out_r_bits_resp = AXI4UserYanker_auto_in_r_bits_resp;
  assign AXI4Deinterleaver_auto_out_r_bits_user = AXI4UserYanker_auto_in_r_bits_user;
  assign AXI4Deinterleaver_auto_out_r_bits_last = AXI4UserYanker_auto_in_r_bits_last;
  assign AXI4IdIndexer_auto_in_aw_valid = TLToAXI4_auto_out_aw_valid;
  assign AXI4IdIndexer_auto_in_aw_bits_id = TLToAXI4_auto_out_aw_bits_id;
  assign AXI4IdIndexer_auto_in_aw_bits_addr = TLToAXI4_auto_out_aw_bits_addr;
  assign AXI4IdIndexer_auto_in_aw_bits_len = TLToAXI4_auto_out_aw_bits_len;
  assign AXI4IdIndexer_auto_in_aw_bits_size = TLToAXI4_auto_out_aw_bits_size;
  assign AXI4IdIndexer_auto_in_aw_bits_burst = TLToAXI4_auto_out_aw_bits_burst;
  assign AXI4IdIndexer_auto_in_aw_bits_lock = TLToAXI4_auto_out_aw_bits_lock;
  assign AXI4IdIndexer_auto_in_aw_bits_cache = TLToAXI4_auto_out_aw_bits_cache;
  assign AXI4IdIndexer_auto_in_aw_bits_prot = TLToAXI4_auto_out_aw_bits_prot;
  assign AXI4IdIndexer_auto_in_aw_bits_qos = TLToAXI4_auto_out_aw_bits_qos;
  assign AXI4IdIndexer_auto_in_aw_bits_user = TLToAXI4_auto_out_aw_bits_user;
  assign AXI4IdIndexer_auto_in_w_valid = TLToAXI4_auto_out_w_valid;
  assign AXI4IdIndexer_auto_in_w_bits_data = TLToAXI4_auto_out_w_bits_data;
  assign AXI4IdIndexer_auto_in_w_bits_strb = TLToAXI4_auto_out_w_bits_strb;
  assign AXI4IdIndexer_auto_in_w_bits_last = TLToAXI4_auto_out_w_bits_last;
  assign AXI4IdIndexer_auto_in_b_ready = TLToAXI4_auto_out_b_ready;
  assign AXI4IdIndexer_auto_in_ar_valid = TLToAXI4_auto_out_ar_valid;
  assign AXI4IdIndexer_auto_in_ar_bits_id = TLToAXI4_auto_out_ar_bits_id;
  assign AXI4IdIndexer_auto_in_ar_bits_addr = TLToAXI4_auto_out_ar_bits_addr;
  assign AXI4IdIndexer_auto_in_ar_bits_len = TLToAXI4_auto_out_ar_bits_len;
  assign AXI4IdIndexer_auto_in_ar_bits_size = TLToAXI4_auto_out_ar_bits_size;
  assign AXI4IdIndexer_auto_in_ar_bits_burst = TLToAXI4_auto_out_ar_bits_burst;
  assign AXI4IdIndexer_auto_in_ar_bits_lock = TLToAXI4_auto_out_ar_bits_lock;
  assign AXI4IdIndexer_auto_in_ar_bits_cache = TLToAXI4_auto_out_ar_bits_cache;
  assign AXI4IdIndexer_auto_in_ar_bits_prot = TLToAXI4_auto_out_ar_bits_prot;
  assign AXI4IdIndexer_auto_in_ar_bits_qos = TLToAXI4_auto_out_ar_bits_qos;
  assign AXI4IdIndexer_auto_in_ar_bits_user = TLToAXI4_auto_out_ar_bits_user;
  assign AXI4IdIndexer_auto_in_r_ready = TLToAXI4_auto_out_r_ready;
  assign AXI4IdIndexer_auto_out_aw_ready = AXI4Deinterleaver_auto_in_aw_ready;
  assign AXI4IdIndexer_auto_out_w_ready = AXI4Deinterleaver_auto_in_w_ready;
  assign AXI4IdIndexer_auto_out_b_valid = AXI4Deinterleaver_auto_in_b_valid;
  assign AXI4IdIndexer_auto_out_b_bits_id = AXI4Deinterleaver_auto_in_b_bits_id;
  assign AXI4IdIndexer_auto_out_b_bits_resp = AXI4Deinterleaver_auto_in_b_bits_resp;
  assign AXI4IdIndexer_auto_out_b_bits_user = AXI4Deinterleaver_auto_in_b_bits_user;
  assign AXI4IdIndexer_auto_out_ar_ready = AXI4Deinterleaver_auto_in_ar_ready;
  assign AXI4IdIndexer_auto_out_r_valid = AXI4Deinterleaver_auto_in_r_valid;
  assign AXI4IdIndexer_auto_out_r_bits_id = AXI4Deinterleaver_auto_in_r_bits_id;
  assign AXI4IdIndexer_auto_out_r_bits_data = AXI4Deinterleaver_auto_in_r_bits_data;
  assign AXI4IdIndexer_auto_out_r_bits_resp = AXI4Deinterleaver_auto_in_r_bits_resp;
  assign AXI4IdIndexer_auto_out_r_bits_user = AXI4Deinterleaver_auto_in_r_bits_user;
  assign AXI4IdIndexer_auto_out_r_bits_last = AXI4Deinterleaver_auto_in_r_bits_last;
  assign TLToAXI4_clock = clock;
  assign TLToAXI4_reset = reset;
  assign TLToAXI4_auto_in_a_valid = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_valid;
  assign TLToAXI4_auto_in_a_bits_opcode = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_opcode;
  assign TLToAXI4_auto_in_a_bits_size = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_size;
  assign TLToAXI4_auto_in_a_bits_source = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_source;
  assign TLToAXI4_auto_in_a_bits_address = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_address;
  assign TLToAXI4_auto_in_a_bits_mask = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_mask;
  assign TLToAXI4_auto_in_a_bits_data = sbus_auto_SystemBus_slave_TLWidthWidget_out_a_bits_data;
  assign TLToAXI4_auto_in_d_ready = sbus_auto_SystemBus_slave_TLWidthWidget_out_d_ready;
  assign TLToAXI4_auto_out_aw_ready = AXI4IdIndexer_auto_in_aw_ready;
  assign TLToAXI4_auto_out_w_ready = AXI4IdIndexer_auto_in_w_ready;
  assign TLToAXI4_auto_out_b_valid = AXI4IdIndexer_auto_in_b_valid;
  assign TLToAXI4_auto_out_b_bits_id = AXI4IdIndexer_auto_in_b_bits_id;
  assign TLToAXI4_auto_out_b_bits_resp = AXI4IdIndexer_auto_in_b_bits_resp;
  assign TLToAXI4_auto_out_b_bits_user = AXI4IdIndexer_auto_in_b_bits_user;
  assign TLToAXI4_auto_out_ar_ready = AXI4IdIndexer_auto_in_ar_ready;
  assign TLToAXI4_auto_out_r_valid = AXI4IdIndexer_auto_in_r_valid;
  assign TLToAXI4_auto_out_r_bits_id = AXI4IdIndexer_auto_in_r_bits_id;
  assign TLToAXI4_auto_out_r_bits_data = AXI4IdIndexer_auto_in_r_bits_data;
  assign TLToAXI4_auto_out_r_bits_resp = AXI4IdIndexer_auto_in_r_bits_resp;
  assign TLToAXI4_auto_out_r_bits_user = AXI4IdIndexer_auto_in_r_bits_user;
  assign TLToAXI4_auto_out_r_bits_last = AXI4IdIndexer_auto_in_r_bits_last;
  assign SystemBus_TLBuffer_clock = clock;
  assign SystemBus_TLBuffer_reset = reset;
  assign SystemBus_TLBuffer_auto_in_a_valid = SystemBus_TLWidthWidget_auto_out_a_valid;
  assign SystemBus_TLBuffer_auto_in_a_bits_opcode = SystemBus_TLWidthWidget_auto_out_a_bits_opcode;
  assign SystemBus_TLBuffer_auto_in_a_bits_param = SystemBus_TLWidthWidget_auto_out_a_bits_param;
  assign SystemBus_TLBuffer_auto_in_a_bits_size = SystemBus_TLWidthWidget_auto_out_a_bits_size;
  assign SystemBus_TLBuffer_auto_in_a_bits_source = SystemBus_TLWidthWidget_auto_out_a_bits_source;
  assign SystemBus_TLBuffer_auto_in_a_bits_address = SystemBus_TLWidthWidget_auto_out_a_bits_address;
  assign SystemBus_TLBuffer_auto_in_a_bits_mask = SystemBus_TLWidthWidget_auto_out_a_bits_mask;
  assign SystemBus_TLBuffer_auto_in_a_bits_data = SystemBus_TLWidthWidget_auto_out_a_bits_data;
  assign SystemBus_TLBuffer_auto_in_d_ready = SystemBus_TLWidthWidget_auto_out_d_ready;
  assign SystemBus_TLBuffer_auto_out_a_ready = sbus_auto_SystemBus_port_TLFIFOFixer_in_a_ready;
  assign SystemBus_TLBuffer_auto_out_d_valid = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_valid;
  assign SystemBus_TLBuffer_auto_out_d_bits_opcode = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_opcode;
  assign SystemBus_TLBuffer_auto_out_d_bits_param = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_param;
  assign SystemBus_TLBuffer_auto_out_d_bits_size = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_size;
  assign SystemBus_TLBuffer_auto_out_d_bits_source = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_source;
  assign SystemBus_TLBuffer_auto_out_d_bits_sink = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_sink;
  assign SystemBus_TLBuffer_auto_out_d_bits_data = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_data;
  assign SystemBus_TLBuffer_auto_out_d_bits_error = sbus_auto_SystemBus_port_TLFIFOFixer_in_d_bits_error;
  assign SystemBus_TLWidthWidget_auto_in_a_valid = AXI4ToTL_auto_out_a_valid;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_opcode = AXI4ToTL_auto_out_a_bits_opcode;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_param = AXI4ToTL_auto_out_a_bits_param;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_size = AXI4ToTL_auto_out_a_bits_size;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_source = AXI4ToTL_auto_out_a_bits_source;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_address = AXI4ToTL_auto_out_a_bits_address;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_mask = AXI4ToTL_auto_out_a_bits_mask;
  assign SystemBus_TLWidthWidget_auto_in_a_bits_data = AXI4ToTL_auto_out_a_bits_data;
  assign SystemBus_TLWidthWidget_auto_in_d_ready = AXI4ToTL_auto_out_d_ready;
  assign SystemBus_TLWidthWidget_auto_out_a_ready = SystemBus_TLBuffer_auto_in_a_ready;
  assign SystemBus_TLWidthWidget_auto_out_d_valid = SystemBus_TLBuffer_auto_in_d_valid;
  assign SystemBus_TLWidthWidget_auto_out_d_bits_opcode = SystemBus_TLBuffer_auto_in_d_bits_opcode;
  assign SystemBus_TLWidthWidget_auto_out_d_bits_size = SystemBus_TLBuffer_auto_in_d_bits_size;
  assign SystemBus_TLWidthWidget_auto_out_d_bits_source = SystemBus_TLBuffer_auto_in_d_bits_source;
  assign SystemBus_TLWidthWidget_auto_out_d_bits_data = SystemBus_TLBuffer_auto_in_d_bits_data;
  assign SystemBus_TLWidthWidget_auto_out_d_bits_error = SystemBus_TLBuffer_auto_in_d_bits_error;
  assign AXI4ToTL_clock = clock;
  assign AXI4ToTL_reset = reset;
  assign AXI4ToTL_auto_in_aw_valid = AXI4UserYanker_1_auto_out_aw_valid;
  assign AXI4ToTL_auto_in_aw_bits_id = AXI4UserYanker_1_auto_out_aw_bits_id;
  assign AXI4ToTL_auto_in_aw_bits_addr = AXI4UserYanker_1_auto_out_aw_bits_addr;
  assign AXI4ToTL_auto_in_aw_bits_len = AXI4UserYanker_1_auto_out_aw_bits_len;
  assign AXI4ToTL_auto_in_aw_bits_size = AXI4UserYanker_1_auto_out_aw_bits_size;
  assign AXI4ToTL_auto_in_w_valid = AXI4UserYanker_1_auto_out_w_valid;
  assign AXI4ToTL_auto_in_w_bits_data = AXI4UserYanker_1_auto_out_w_bits_data;
  assign AXI4ToTL_auto_in_w_bits_strb = AXI4UserYanker_1_auto_out_w_bits_strb;
  assign AXI4ToTL_auto_in_w_bits_last = AXI4UserYanker_1_auto_out_w_bits_last;
  assign AXI4ToTL_auto_in_b_ready = AXI4UserYanker_1_auto_out_b_ready;
  assign AXI4ToTL_auto_in_ar_valid = AXI4UserYanker_1_auto_out_ar_valid;
  assign AXI4ToTL_auto_in_ar_bits_id = AXI4UserYanker_1_auto_out_ar_bits_id;
  assign AXI4ToTL_auto_in_ar_bits_addr = AXI4UserYanker_1_auto_out_ar_bits_addr;
  assign AXI4ToTL_auto_in_ar_bits_len = AXI4UserYanker_1_auto_out_ar_bits_len;
  assign AXI4ToTL_auto_in_ar_bits_size = AXI4UserYanker_1_auto_out_ar_bits_size;
  assign AXI4ToTL_auto_in_r_ready = AXI4UserYanker_1_auto_out_r_ready;
  assign AXI4ToTL_auto_out_a_ready = SystemBus_TLWidthWidget_auto_in_a_ready;
  assign AXI4ToTL_auto_out_d_valid = SystemBus_TLWidthWidget_auto_in_d_valid;
  assign AXI4ToTL_auto_out_d_bits_opcode = SystemBus_TLWidthWidget_auto_in_d_bits_opcode;
  assign AXI4ToTL_auto_out_d_bits_size = SystemBus_TLWidthWidget_auto_in_d_bits_size;
  assign AXI4ToTL_auto_out_d_bits_source = SystemBus_TLWidthWidget_auto_in_d_bits_source;
  assign AXI4ToTL_auto_out_d_bits_data = SystemBus_TLWidthWidget_auto_in_d_bits_data;
  assign AXI4ToTL_auto_out_d_bits_error = SystemBus_TLWidthWidget_auto_in_d_bits_error;
  assign AXI4UserYanker_1_clock = clock;
  assign AXI4UserYanker_1_reset = reset;
  assign AXI4UserYanker_1_auto_in_aw_valid = AXI4Fragmenter_auto_out_aw_valid;
  assign AXI4UserYanker_1_auto_in_aw_bits_id = AXI4Fragmenter_auto_out_aw_bits_id;
  assign AXI4UserYanker_1_auto_in_aw_bits_addr = AXI4Fragmenter_auto_out_aw_bits_addr;
  assign AXI4UserYanker_1_auto_in_aw_bits_len = AXI4Fragmenter_auto_out_aw_bits_len;
  assign AXI4UserYanker_1_auto_in_aw_bits_size = AXI4Fragmenter_auto_out_aw_bits_size;
  assign AXI4UserYanker_1_auto_in_aw_bits_user = AXI4Fragmenter_auto_out_aw_bits_user;
  assign AXI4UserYanker_1_auto_in_w_valid = AXI4Fragmenter_auto_out_w_valid;
  assign AXI4UserYanker_1_auto_in_w_bits_data = AXI4Fragmenter_auto_out_w_bits_data;
  assign AXI4UserYanker_1_auto_in_w_bits_strb = AXI4Fragmenter_auto_out_w_bits_strb;
  assign AXI4UserYanker_1_auto_in_w_bits_last = AXI4Fragmenter_auto_out_w_bits_last;
  assign AXI4UserYanker_1_auto_in_b_ready = AXI4Fragmenter_auto_out_b_ready;
  assign AXI4UserYanker_1_auto_in_ar_valid = AXI4Fragmenter_auto_out_ar_valid;
  assign AXI4UserYanker_1_auto_in_ar_bits_id = AXI4Fragmenter_auto_out_ar_bits_id;
  assign AXI4UserYanker_1_auto_in_ar_bits_addr = AXI4Fragmenter_auto_out_ar_bits_addr;
  assign AXI4UserYanker_1_auto_in_ar_bits_len = AXI4Fragmenter_auto_out_ar_bits_len;
  assign AXI4UserYanker_1_auto_in_ar_bits_size = AXI4Fragmenter_auto_out_ar_bits_size;
  assign AXI4UserYanker_1_auto_in_ar_bits_user = AXI4Fragmenter_auto_out_ar_bits_user;
  assign AXI4UserYanker_1_auto_in_r_ready = AXI4Fragmenter_auto_out_r_ready;
  assign AXI4UserYanker_1_auto_out_aw_ready = AXI4ToTL_auto_in_aw_ready;
  assign AXI4UserYanker_1_auto_out_w_ready = AXI4ToTL_auto_in_w_ready;
  assign AXI4UserYanker_1_auto_out_b_valid = AXI4ToTL_auto_in_b_valid;
  assign AXI4UserYanker_1_auto_out_b_bits_id = AXI4ToTL_auto_in_b_bits_id;
  assign AXI4UserYanker_1_auto_out_b_bits_resp = AXI4ToTL_auto_in_b_bits_resp;
  assign AXI4UserYanker_1_auto_out_ar_ready = AXI4ToTL_auto_in_ar_ready;
  assign AXI4UserYanker_1_auto_out_r_valid = AXI4ToTL_auto_in_r_valid;
  assign AXI4UserYanker_1_auto_out_r_bits_id = AXI4ToTL_auto_in_r_bits_id;
  assign AXI4UserYanker_1_auto_out_r_bits_data = AXI4ToTL_auto_in_r_bits_data;
  assign AXI4UserYanker_1_auto_out_r_bits_resp = AXI4ToTL_auto_in_r_bits_resp;
  assign AXI4UserYanker_1_auto_out_r_bits_last = AXI4ToTL_auto_in_r_bits_last;
  assign AXI4Fragmenter_clock = clock;
  assign AXI4Fragmenter_reset = reset;
  assign AXI4Fragmenter_auto_in_aw_valid = AXI4IdIndexer_1_auto_out_aw_valid;
  assign AXI4Fragmenter_auto_in_aw_bits_id = AXI4IdIndexer_1_auto_out_aw_bits_id;
  assign AXI4Fragmenter_auto_in_aw_bits_addr = AXI4IdIndexer_1_auto_out_aw_bits_addr;
  assign AXI4Fragmenter_auto_in_aw_bits_len = AXI4IdIndexer_1_auto_out_aw_bits_len;
  assign AXI4Fragmenter_auto_in_aw_bits_size = AXI4IdIndexer_1_auto_out_aw_bits_size;
  assign AXI4Fragmenter_auto_in_aw_bits_burst = AXI4IdIndexer_1_auto_out_aw_bits_burst;
  assign AXI4Fragmenter_auto_in_aw_bits_user = AXI4IdIndexer_1_auto_out_aw_bits_user;
  assign AXI4Fragmenter_auto_in_w_valid = AXI4IdIndexer_1_auto_out_w_valid;
  assign AXI4Fragmenter_auto_in_w_bits_data = AXI4IdIndexer_1_auto_out_w_bits_data;
  assign AXI4Fragmenter_auto_in_w_bits_strb = AXI4IdIndexer_1_auto_out_w_bits_strb;
  assign AXI4Fragmenter_auto_in_w_bits_last = AXI4IdIndexer_1_auto_out_w_bits_last;
  assign AXI4Fragmenter_auto_in_b_ready = AXI4IdIndexer_1_auto_out_b_ready;
  assign AXI4Fragmenter_auto_in_ar_valid = AXI4IdIndexer_1_auto_out_ar_valid;
  assign AXI4Fragmenter_auto_in_ar_bits_id = AXI4IdIndexer_1_auto_out_ar_bits_id;
  assign AXI4Fragmenter_auto_in_ar_bits_addr = AXI4IdIndexer_1_auto_out_ar_bits_addr;
  assign AXI4Fragmenter_auto_in_ar_bits_len = AXI4IdIndexer_1_auto_out_ar_bits_len;
  assign AXI4Fragmenter_auto_in_ar_bits_size = AXI4IdIndexer_1_auto_out_ar_bits_size;
  assign AXI4Fragmenter_auto_in_ar_bits_burst = AXI4IdIndexer_1_auto_out_ar_bits_burst;
  assign AXI4Fragmenter_auto_in_ar_bits_user = AXI4IdIndexer_1_auto_out_ar_bits_user;
  assign AXI4Fragmenter_auto_in_r_ready = AXI4IdIndexer_1_auto_out_r_ready;
  assign AXI4Fragmenter_auto_out_aw_ready = AXI4UserYanker_1_auto_in_aw_ready;
  assign AXI4Fragmenter_auto_out_w_ready = AXI4UserYanker_1_auto_in_w_ready;
  assign AXI4Fragmenter_auto_out_b_valid = AXI4UserYanker_1_auto_in_b_valid;
  assign AXI4Fragmenter_auto_out_b_bits_id = AXI4UserYanker_1_auto_in_b_bits_id;
  assign AXI4Fragmenter_auto_out_b_bits_resp = AXI4UserYanker_1_auto_in_b_bits_resp;
  assign AXI4Fragmenter_auto_out_b_bits_user = AXI4UserYanker_1_auto_in_b_bits_user;
  assign AXI4Fragmenter_auto_out_ar_ready = AXI4UserYanker_1_auto_in_ar_ready;
  assign AXI4Fragmenter_auto_out_r_valid = AXI4UserYanker_1_auto_in_r_valid;
  assign AXI4Fragmenter_auto_out_r_bits_id = AXI4UserYanker_1_auto_in_r_bits_id;
  assign AXI4Fragmenter_auto_out_r_bits_data = AXI4UserYanker_1_auto_in_r_bits_data;
  assign AXI4Fragmenter_auto_out_r_bits_resp = AXI4UserYanker_1_auto_in_r_bits_resp;
  assign AXI4Fragmenter_auto_out_r_bits_user = AXI4UserYanker_1_auto_in_r_bits_user;
  assign AXI4Fragmenter_auto_out_r_bits_last = AXI4UserYanker_1_auto_in_r_bits_last;
  assign AXI4IdIndexer_1_auto_in_aw_valid = _T_155_aw_valid;
  assign AXI4IdIndexer_1_auto_in_aw_bits_id = _T_155_aw_bits_id;
  assign AXI4IdIndexer_1_auto_in_aw_bits_addr = _T_155_aw_bits_addr;
  assign AXI4IdIndexer_1_auto_in_aw_bits_len = _T_155_aw_bits_len;
  assign AXI4IdIndexer_1_auto_in_aw_bits_size = _T_155_aw_bits_size;
  assign AXI4IdIndexer_1_auto_in_aw_bits_burst = _T_155_aw_bits_burst;
  assign AXI4IdIndexer_1_auto_in_w_valid = _T_155_w_valid;
  assign AXI4IdIndexer_1_auto_in_w_bits_data = _T_155_w_bits_data;
  assign AXI4IdIndexer_1_auto_in_w_bits_strb = _T_155_w_bits_strb;
  assign AXI4IdIndexer_1_auto_in_w_bits_last = _T_155_w_bits_last;
  assign AXI4IdIndexer_1_auto_in_b_ready = _T_155_b_ready;
  assign AXI4IdIndexer_1_auto_in_ar_valid = _T_155_ar_valid;
  assign AXI4IdIndexer_1_auto_in_ar_bits_id = _T_155_ar_bits_id;
  assign AXI4IdIndexer_1_auto_in_ar_bits_addr = _T_155_ar_bits_addr;
  assign AXI4IdIndexer_1_auto_in_ar_bits_len = _T_155_ar_bits_len;
  assign AXI4IdIndexer_1_auto_in_ar_bits_size = _T_155_ar_bits_size;
  assign AXI4IdIndexer_1_auto_in_ar_bits_burst = _T_155_ar_bits_burst;
  assign AXI4IdIndexer_1_auto_in_r_ready = _T_155_r_ready;
  assign AXI4IdIndexer_1_auto_out_aw_ready = AXI4Fragmenter_auto_in_aw_ready;
  assign AXI4IdIndexer_1_auto_out_w_ready = AXI4Fragmenter_auto_in_w_ready;
  assign AXI4IdIndexer_1_auto_out_b_valid = AXI4Fragmenter_auto_in_b_valid;
  assign AXI4IdIndexer_1_auto_out_b_bits_id = AXI4Fragmenter_auto_in_b_bits_id;
  assign AXI4IdIndexer_1_auto_out_b_bits_resp = AXI4Fragmenter_auto_in_b_bits_resp;
  assign AXI4IdIndexer_1_auto_out_b_bits_user = AXI4Fragmenter_auto_in_b_bits_user;
  assign AXI4IdIndexer_1_auto_out_ar_ready = AXI4Fragmenter_auto_in_ar_ready;
  assign AXI4IdIndexer_1_auto_out_r_valid = AXI4Fragmenter_auto_in_r_valid;
  assign AXI4IdIndexer_1_auto_out_r_bits_id = AXI4Fragmenter_auto_in_r_bits_id;
  assign AXI4IdIndexer_1_auto_out_r_bits_data = AXI4Fragmenter_auto_in_r_bits_data;
  assign AXI4IdIndexer_1_auto_out_r_bits_resp = AXI4Fragmenter_auto_in_r_bits_resp;
  assign AXI4IdIndexer_1_auto_out_r_bits_user = AXI4Fragmenter_auto_in_r_bits_user;
  assign AXI4IdIndexer_1_auto_out_r_bits_last = AXI4Fragmenter_auto_in_r_bits_last;
  assign bootrom_auto_in_a_valid = pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_valid;
  assign bootrom_auto_in_a_bits_size = pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_size;
  assign bootrom_auto_in_a_bits_source = pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_source;
  assign bootrom_auto_in_a_bits_address = pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_a_bits_address;
  assign bootrom_auto_in_d_ready = pbus_auto_PeripheryBus_slave_TLFragmenter_out_3_d_ready;
  assign error_clock = clock;
  assign error_reset = reset;
  assign error_auto_in_a_valid = sbus_auto_SystemBus_slave_TLBuffer_out_a_valid;
  assign error_auto_in_a_bits_opcode = sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_opcode;
  assign error_auto_in_a_bits_size = sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_size;
  assign error_auto_in_a_bits_source = sbus_auto_SystemBus_slave_TLBuffer_out_a_bits_source;
  assign error_auto_in_c_valid = sbus_auto_SystemBus_slave_TLBuffer_out_c_valid;
  assign error_auto_in_c_bits_opcode = sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_opcode;
  assign error_auto_in_c_bits_param = sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_param;
  assign error_auto_in_c_bits_size = sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_size;
  assign error_auto_in_c_bits_source = sbus_auto_SystemBus_slave_TLBuffer_out_c_bits_source;
  assign error_auto_in_d_ready = sbus_auto_SystemBus_slave_TLBuffer_out_d_ready;
  assign _T_5_0 = _T_248;
  assign _T_5_1 = _T_249;
  assign _T_39_aw_ready = mem_axi4_0_aw_ready;
  assign _T_39_aw_valid = buffer_auto_out_aw_valid;
  assign _T_39_aw_bits_id = buffer_auto_out_aw_bits_id;
  assign _T_39_aw_bits_addr = buffer_auto_out_aw_bits_addr;
  assign _T_39_aw_bits_len = buffer_auto_out_aw_bits_len;
  assign _T_39_aw_bits_size = buffer_auto_out_aw_bits_size;
  assign _T_39_aw_bits_burst = buffer_auto_out_aw_bits_burst;
  assign _T_39_aw_bits_lock = buffer_auto_out_aw_bits_lock;
  assign _T_39_aw_bits_cache = buffer_auto_out_aw_bits_cache;
  assign _T_39_aw_bits_prot = buffer_auto_out_aw_bits_prot;
  assign _T_39_aw_bits_qos = buffer_auto_out_aw_bits_qos;
  assign _T_39_w_ready = mem_axi4_0_w_ready;
  assign _T_39_w_valid = buffer_auto_out_w_valid;
  assign _T_39_w_bits_data = buffer_auto_out_w_bits_data;
  assign _T_39_w_bits_strb = buffer_auto_out_w_bits_strb;
  assign _T_39_w_bits_last = buffer_auto_out_w_bits_last;
  assign _T_39_b_ready = buffer_auto_out_b_ready;
  assign _T_39_b_valid = mem_axi4_0_b_valid;
  assign _T_39_b_bits_id = mem_axi4_0_b_bits_id;
  assign _T_39_b_bits_resp = mem_axi4_0_b_bits_resp;
  assign _T_39_ar_ready = mem_axi4_0_ar_ready;
  assign _T_39_ar_valid = buffer_auto_out_ar_valid;
  assign _T_39_ar_bits_id = buffer_auto_out_ar_bits_id;
  assign _T_39_ar_bits_addr = buffer_auto_out_ar_bits_addr;
  assign _T_39_ar_bits_len = buffer_auto_out_ar_bits_len;
  assign _T_39_ar_bits_size = buffer_auto_out_ar_bits_size;
  assign _T_39_ar_bits_burst = buffer_auto_out_ar_bits_burst;
  assign _T_39_ar_bits_lock = buffer_auto_out_ar_bits_lock;
  assign _T_39_ar_bits_cache = buffer_auto_out_ar_bits_cache;
  assign _T_39_ar_bits_prot = buffer_auto_out_ar_bits_prot;
  assign _T_39_ar_bits_qos = buffer_auto_out_ar_bits_qos;
  assign _T_39_r_ready = buffer_auto_out_r_ready;
  assign _T_39_r_valid = mem_axi4_0_r_valid;
  assign _T_39_r_bits_id = mem_axi4_0_r_bits_id;
  assign _T_39_r_bits_data = mem_axi4_0_r_bits_data;
  assign _T_39_r_bits_resp = mem_axi4_0_r_bits_resp;
  assign _T_39_r_bits_last = mem_axi4_0_r_bits_last;
  assign _T_97_aw_ready = mmio_axi4_0_aw_ready;
  assign _T_97_aw_valid = AXI4Buffer_auto_out_aw_valid;
  assign _T_97_aw_bits_id = AXI4Buffer_auto_out_aw_bits_id;
  assign _T_97_aw_bits_addr = AXI4Buffer_auto_out_aw_bits_addr;
  assign _T_97_aw_bits_len = AXI4Buffer_auto_out_aw_bits_len;
  assign _T_97_aw_bits_size = AXI4Buffer_auto_out_aw_bits_size;
  assign _T_97_aw_bits_burst = AXI4Buffer_auto_out_aw_bits_burst;
  assign _T_97_aw_bits_lock = AXI4Buffer_auto_out_aw_bits_lock;
  assign _T_97_aw_bits_cache = AXI4Buffer_auto_out_aw_bits_cache;
  assign _T_97_aw_bits_prot = AXI4Buffer_auto_out_aw_bits_prot;
  assign _T_97_aw_bits_qos = AXI4Buffer_auto_out_aw_bits_qos;
  assign _T_97_w_ready = mmio_axi4_0_w_ready;
  assign _T_97_w_valid = AXI4Buffer_auto_out_w_valid;
  assign _T_97_w_bits_data = AXI4Buffer_auto_out_w_bits_data;
  assign _T_97_w_bits_strb = AXI4Buffer_auto_out_w_bits_strb;
  assign _T_97_w_bits_last = AXI4Buffer_auto_out_w_bits_last;
  assign _T_97_b_ready = AXI4Buffer_auto_out_b_ready;
  assign _T_97_b_valid = mmio_axi4_0_b_valid;
  assign _T_97_b_bits_id = mmio_axi4_0_b_bits_id;
  assign _T_97_b_bits_resp = mmio_axi4_0_b_bits_resp;
  assign _T_97_ar_ready = mmio_axi4_0_ar_ready;
  assign _T_97_ar_valid = AXI4Buffer_auto_out_ar_valid;
  assign _T_97_ar_bits_id = AXI4Buffer_auto_out_ar_bits_id;
  assign _T_97_ar_bits_addr = AXI4Buffer_auto_out_ar_bits_addr;
  assign _T_97_ar_bits_len = AXI4Buffer_auto_out_ar_bits_len;
  assign _T_97_ar_bits_size = AXI4Buffer_auto_out_ar_bits_size;
  assign _T_97_ar_bits_burst = AXI4Buffer_auto_out_ar_bits_burst;
  assign _T_97_ar_bits_lock = AXI4Buffer_auto_out_ar_bits_lock;
  assign _T_97_ar_bits_cache = AXI4Buffer_auto_out_ar_bits_cache;
  assign _T_97_ar_bits_prot = AXI4Buffer_auto_out_ar_bits_prot;
  assign _T_97_ar_bits_qos = AXI4Buffer_auto_out_ar_bits_qos;
  assign _T_97_r_ready = AXI4Buffer_auto_out_r_ready;
  assign _T_97_r_valid = mmio_axi4_0_r_valid;
  assign _T_97_r_bits_id = mmio_axi4_0_r_bits_id;
  assign _T_97_r_bits_data = mmio_axi4_0_r_bits_data;
  assign _T_97_r_bits_resp = mmio_axi4_0_r_bits_resp;
  assign _T_97_r_bits_last = mmio_axi4_0_r_bits_last;
  assign _T_155_aw_ready = AXI4IdIndexer_1_auto_in_aw_ready;
  assign _T_155_aw_valid = l2_frontend_bus_axi4_0_aw_valid;
  assign _T_155_aw_bits_id = l2_frontend_bus_axi4_0_aw_bits_id;
  assign _T_155_aw_bits_addr = l2_frontend_bus_axi4_0_aw_bits_addr;
  assign _T_155_aw_bits_len = l2_frontend_bus_axi4_0_aw_bits_len;
  assign _T_155_aw_bits_size = l2_frontend_bus_axi4_0_aw_bits_size;
  assign _T_155_aw_bits_burst = l2_frontend_bus_axi4_0_aw_bits_burst;
  assign _T_155_w_ready = AXI4IdIndexer_1_auto_in_w_ready;
  assign _T_155_w_valid = l2_frontend_bus_axi4_0_w_valid;
  assign _T_155_w_bits_data = l2_frontend_bus_axi4_0_w_bits_data;
  assign _T_155_w_bits_strb = l2_frontend_bus_axi4_0_w_bits_strb;
  assign _T_155_w_bits_last = l2_frontend_bus_axi4_0_w_bits_last;
  assign _T_155_b_ready = l2_frontend_bus_axi4_0_b_ready;
  assign _T_155_b_valid = AXI4IdIndexer_1_auto_in_b_valid;
  assign _T_155_b_bits_id = AXI4IdIndexer_1_auto_in_b_bits_id;
  assign _T_155_b_bits_resp = AXI4IdIndexer_1_auto_in_b_bits_resp;
  assign _T_155_ar_ready = AXI4IdIndexer_1_auto_in_ar_ready;
  assign _T_155_ar_valid = l2_frontend_bus_axi4_0_ar_valid;
  assign _T_155_ar_bits_id = l2_frontend_bus_axi4_0_ar_bits_id;
  assign _T_155_ar_bits_addr = l2_frontend_bus_axi4_0_ar_bits_addr;
  assign _T_155_ar_bits_len = l2_frontend_bus_axi4_0_ar_bits_len;
  assign _T_155_ar_bits_size = l2_frontend_bus_axi4_0_ar_bits_size;
  assign _T_155_ar_bits_burst = l2_frontend_bus_axi4_0_ar_bits_burst;
  assign _T_155_r_ready = l2_frontend_bus_axi4_0_r_ready;
  assign _T_155_r_valid = AXI4IdIndexer_1_auto_in_r_valid;
  assign _T_155_r_bits_id = AXI4IdIndexer_1_auto_in_r_bits_id;
  assign _T_155_r_bits_data = AXI4IdIndexer_1_auto_in_r_bits_data;
  assign _T_155_r_bits_resp = AXI4IdIndexer_1_auto_in_r_bits_resp;
  assign _T_155_r_bits_last = AXI4IdIndexer_1_auto_in_r_bits_last;
  assign tile_inputs_0_clock = clock;
  assign tile_inputs_0_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (int_rtc_tick) begin
        value <= 7'h0;
      end else begin
        value <= _T_245;
      end
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [27:0] auto_in_aw_bits_addr,
  input         auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [27:0] auto_in_ar_bits_addr,
  input         auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_user
);
  wire  in_aw_ready;
  wire  in_aw_valid;
  wire [3:0] in_aw_bits_id;
  wire [27:0] in_aw_bits_addr;
  wire  in_aw_bits_user;
  wire  in_w_ready;
  wire  in_w_valid;
  wire [63:0] in_w_bits_data;
  wire [7:0] in_w_bits_strb;
  wire  in_b_ready;
  wire  in_b_valid;
  wire [3:0] in_b_bits_id;
  wire [1:0] in_b_bits_resp;
  wire  in_b_bits_user;
  wire  in_ar_ready;
  wire  in_ar_valid;
  wire [3:0] in_ar_bits_id;
  wire [27:0] in_ar_bits_addr;
  wire  in_ar_bits_user;
  wire  in_r_ready;
  wire  in_r_valid;
  wire [3:0] in_r_bits_id;
  wire [63:0] in_r_bits_data;
  wire [1:0] in_r_bits_resp;
  wire  in_r_bits_user;
  reg [7:0] mem_0 [0:33554431];
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_326_data;
  wire [24:0] mem_0__T_326_addr;
  wire [7:0] mem_0__T_281_data;
  wire [24:0] mem_0__T_281_addr;
  wire  mem_0__T_281_mask;
  wire  mem_0__T_281_en;
  wire  _GEN_57;
  reg [24:0] mem_0__T_326_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] mem_1 [0:33554431];
  reg [31:0] _RAND_2;
  wire [7:0] mem_1__T_326_data;
  wire [24:0] mem_1__T_326_addr;
  wire [7:0] mem_1__T_281_data;
  wire [24:0] mem_1__T_281_addr;
  wire  mem_1__T_281_mask;
  wire  mem_1__T_281_en;
  reg [24:0] mem_1__T_326_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [7:0] mem_2 [0:33554431];
  reg [31:0] _RAND_4;
  wire [7:0] mem_2__T_326_data;
  wire [24:0] mem_2__T_326_addr;
  wire [7:0] mem_2__T_281_data;
  wire [24:0] mem_2__T_281_addr;
  wire  mem_2__T_281_mask;
  wire  mem_2__T_281_en;
  reg [24:0] mem_2__T_326_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] mem_3 [0:33554431];
  reg [31:0] _RAND_6;
  wire [7:0] mem_3__T_326_data;
  wire [24:0] mem_3__T_326_addr;
  wire [7:0] mem_3__T_281_data;
  wire [24:0] mem_3__T_281_addr;
  wire  mem_3__T_281_mask;
  wire  mem_3__T_281_en;
  reg [24:0] mem_3__T_326_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [7:0] mem_4 [0:33554431];
  reg [31:0] _RAND_8;
  wire [7:0] mem_4__T_326_data;
  wire [24:0] mem_4__T_326_addr;
  wire [7:0] mem_4__T_281_data;
  wire [24:0] mem_4__T_281_addr;
  wire  mem_4__T_281_mask;
  wire  mem_4__T_281_en;
  reg [24:0] mem_4__T_326_addr_pipe_0;
  reg [31:0] _RAND_9;
  reg [7:0] mem_5 [0:33554431];
  reg [31:0] _RAND_10;
  wire [7:0] mem_5__T_326_data;
  wire [24:0] mem_5__T_326_addr;
  wire [7:0] mem_5__T_281_data;
  wire [24:0] mem_5__T_281_addr;
  wire  mem_5__T_281_mask;
  wire  mem_5__T_281_en;
  reg [24:0] mem_5__T_326_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] mem_6 [0:33554431];
  reg [31:0] _RAND_12;
  wire [7:0] mem_6__T_326_data;
  wire [24:0] mem_6__T_326_addr;
  wire [7:0] mem_6__T_281_data;
  wire [24:0] mem_6__T_281_addr;
  wire  mem_6__T_281_mask;
  wire  mem_6__T_281_en;
  reg [24:0] mem_6__T_326_addr_pipe_0;
  reg [31:0] _RAND_13;
  reg [7:0] mem_7 [0:33554431];
  reg [31:0] _RAND_14;
  wire [7:0] mem_7__T_326_data;
  wire [24:0] mem_7__T_326_addr;
  wire [7:0] mem_7__T_281_data;
  wire [24:0] mem_7__T_281_addr;
  wire  mem_7__T_281_mask;
  wire  mem_7__T_281_en;
  reg [24:0] mem_7__T_326_addr_pipe_0;
  reg [31:0] _RAND_15;
  wire [24:0] _T_130;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  _T_134;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_138;
  wire  _T_139;
  wire  _T_140;
  wire  _T_141;
  wire  _T_142;
  wire  _T_143;
  wire  _T_144;
  wire  _T_145;
  wire  _T_146;
  wire  _T_147;
  wire  _T_148;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire [1:0] _T_156;
  wire [2:0] _T_157;
  wire [1:0] _T_158;
  wire [2:0] _T_159;
  wire [5:0] _T_160;
  wire [1:0] _T_161;
  wire [2:0] _T_162;
  wire [1:0] _T_163;
  wire [2:0] _T_164;
  wire [5:0] _T_165;
  wire [11:0] _T_166;
  wire [1:0] _T_167;
  wire [2:0] _T_168;
  wire [1:0] _T_169;
  wire [2:0] _T_170;
  wire [5:0] _T_171;
  wire [1:0] _T_172;
  wire [2:0] _T_173;
  wire [1:0] _T_174;
  wire [1:0] _T_175;
  wire [3:0] _T_176;
  wire [6:0] _T_177;
  wire [12:0] _T_178;
  wire [24:0] r_addr;
  wire [24:0] _T_179;
  wire  _T_180;
  wire  _T_181;
  wire  _T_182;
  wire  _T_183;
  wire  _T_184;
  wire  _T_185;
  wire  _T_186;
  wire  _T_187;
  wire  _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire  _T_193;
  wire  _T_194;
  wire  _T_195;
  wire  _T_196;
  wire  _T_197;
  wire  _T_198;
  wire  _T_199;
  wire  _T_200;
  wire  _T_201;
  wire  _T_202;
  wire  _T_203;
  wire  _T_204;
  wire [1:0] _T_205;
  wire [2:0] _T_206;
  wire [1:0] _T_207;
  wire [2:0] _T_208;
  wire [5:0] _T_209;
  wire [1:0] _T_210;
  wire [2:0] _T_211;
  wire [1:0] _T_212;
  wire [2:0] _T_213;
  wire [5:0] _T_214;
  wire [11:0] _T_215;
  wire [1:0] _T_216;
  wire [2:0] _T_217;
  wire [1:0] _T_218;
  wire [2:0] _T_219;
  wire [5:0] _T_220;
  wire [1:0] _T_221;
  wire [2:0] _T_222;
  wire [1:0] _T_223;
  wire [1:0] _T_224;
  wire [3:0] _T_225;
  wire [6:0] _T_226;
  wire [12:0] _T_227;
  wire [24:0] w_addr;
  wire [28:0] _T_230;
  wire [28:0] _T_232;
  wire [28:0] _T_233;
  wire  r_sel0;
  wire [28:0] _T_237;
  wire [28:0] _T_239;
  wire [28:0] _T_240;
  wire  w_sel0;
  reg  w_full;
  reg [31:0] _RAND_16;
  reg [3:0] w_id;
  reg [31:0] _RAND_17;
  reg  w_user;
  reg [31:0] _RAND_18;
  reg  r_sel1;
  reg [31:0] _RAND_19;
  reg  w_sel1;
  reg [31:0] _RAND_20;
  wire  _T_246;
  wire  _GEN_0;
  wire  _T_248;
  wire  _GEN_1;
  wire [3:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [7:0] _T_251;
  wire [7:0] _T_252;
  wire [7:0] _T_253;
  wire [7:0] _T_254;
  wire [7:0] _T_255;
  wire [7:0] _T_256;
  wire [7:0] _T_257;
  wire [7:0] _T_258;
  wire [7:0] wdata_0;
  wire [7:0] wdata_1;
  wire [7:0] wdata_2;
  wire [7:0] wdata_3;
  wire [7:0] wdata_4;
  wire [7:0] wdata_5;
  wire [7:0] wdata_6;
  wire [7:0] wdata_7;
  wire  _T_272;
  wire  _T_273;
  wire  _T_274;
  wire  _T_275;
  wire  _T_276;
  wire  _T_277;
  wire  _T_278;
  wire  _T_279;
  wire  _T_280;
  wire  _GEN_25;
  wire  _GEN_27;
  wire  _GEN_29;
  wire  _GEN_31;
  wire  _GEN_33;
  wire  _GEN_35;
  wire  _GEN_37;
  wire  _GEN_39;
  wire  _T_302;
  wire  _T_303;
  wire  _T_304;
  wire  _T_308;
  wire [1:0] _T_311;
  reg  r_full;
  reg [31:0] _RAND_21;
  reg [3:0] r_id;
  reg [31:0] _RAND_22;
  reg  r_user;
  reg [31:0] _RAND_23;
  wire  _T_316;
  wire  _GEN_40;
  wire  _T_318;
  wire  _GEN_41;
  wire [3:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  ren;
  wire [24:0] _T_322;
  reg  _T_347;
  reg [31:0] _RAND_24;
  reg [7:0] _T_377_0;
  reg [31:0] _RAND_25;
  reg [7:0] _T_377_1;
  reg [31:0] _RAND_26;
  reg [7:0] _T_377_2;
  reg [31:0] _RAND_27;
  reg [7:0] _T_377_3;
  reg [31:0] _RAND_28;
  reg [7:0] _T_377_4;
  reg [31:0] _RAND_29;
  reg [7:0] _T_377_5;
  reg [31:0] _RAND_30;
  reg [7:0] _T_377_6;
  reg [31:0] _RAND_31;
  reg [7:0] _T_377_7;
  reg [31:0] _RAND_32;
  wire [7:0] _GEN_49;
  wire [7:0] _GEN_50;
  wire [7:0] _GEN_51;
  wire [7:0] _GEN_52;
  wire [7:0] _GEN_53;
  wire [7:0] _GEN_54;
  wire [7:0] _GEN_55;
  wire [7:0] _GEN_56;
  wire  _T_444;
  wire  _T_445;
  wire [1:0] _T_448;
  wire [15:0] _T_449;
  wire [15:0] _T_450;
  wire [31:0] _T_451;
  wire [15:0] _T_452;
  wire [15:0] _T_453;
  wire [31:0] _T_454;
  wire [63:0] _T_455;
  assign mem_0__T_326_addr = mem_0__T_326_addr_pipe_0;
  assign mem_0__T_326_data = mem_0[mem_0__T_326_addr];
  assign mem_0__T_281_data = wdata_0;
  assign mem_0__T_281_addr = w_addr;
  assign mem_0__T_281_mask = _GEN_25;
  assign mem_0__T_281_en = _T_272;
  assign _GEN_57 = ren;
  assign mem_1__T_326_addr = mem_1__T_326_addr_pipe_0;
  assign mem_1__T_326_data = mem_1[mem_1__T_326_addr];
  assign mem_1__T_281_data = wdata_1;
  assign mem_1__T_281_addr = w_addr;
  assign mem_1__T_281_mask = _GEN_27;
  assign mem_1__T_281_en = _T_272;
  assign mem_2__T_326_addr = mem_2__T_326_addr_pipe_0;
  assign mem_2__T_326_data = mem_2[mem_2__T_326_addr];
  assign mem_2__T_281_data = wdata_2;
  assign mem_2__T_281_addr = w_addr;
  assign mem_2__T_281_mask = _GEN_29;
  assign mem_2__T_281_en = _T_272;
  assign mem_3__T_326_addr = mem_3__T_326_addr_pipe_0;
  assign mem_3__T_326_data = mem_3[mem_3__T_326_addr];
  assign mem_3__T_281_data = wdata_3;
  assign mem_3__T_281_addr = w_addr;
  assign mem_3__T_281_mask = _GEN_31;
  assign mem_3__T_281_en = _T_272;
  assign mem_4__T_326_addr = mem_4__T_326_addr_pipe_0;
  assign mem_4__T_326_data = mem_4[mem_4__T_326_addr];
  assign mem_4__T_281_data = wdata_4;
  assign mem_4__T_281_addr = w_addr;
  assign mem_4__T_281_mask = _GEN_33;
  assign mem_4__T_281_en = _T_272;
  assign mem_5__T_326_addr = mem_5__T_326_addr_pipe_0;
  assign mem_5__T_326_data = mem_5[mem_5__T_326_addr];
  assign mem_5__T_281_data = wdata_5;
  assign mem_5__T_281_addr = w_addr;
  assign mem_5__T_281_mask = _GEN_35;
  assign mem_5__T_281_en = _T_272;
  assign mem_6__T_326_addr = mem_6__T_326_addr_pipe_0;
  assign mem_6__T_326_data = mem_6[mem_6__T_326_addr];
  assign mem_6__T_281_data = wdata_6;
  assign mem_6__T_281_addr = w_addr;
  assign mem_6__T_281_mask = _GEN_37;
  assign mem_6__T_281_en = _T_272;
  assign mem_7__T_326_addr = mem_7__T_326_addr_pipe_0;
  assign mem_7__T_326_data = mem_7[mem_7__T_326_addr];
  assign mem_7__T_281_data = wdata_7;
  assign mem_7__T_281_addr = w_addr;
  assign mem_7__T_281_mask = _GEN_39;
  assign mem_7__T_281_en = _T_272;
  assign _T_130 = in_ar_bits_addr[27:3];
  assign _T_131 = _T_130[0];
  assign _T_132 = _T_130[1];
  assign _T_133 = _T_130[2];
  assign _T_134 = _T_130[3];
  assign _T_135 = _T_130[4];
  assign _T_136 = _T_130[5];
  assign _T_137 = _T_130[6];
  assign _T_138 = _T_130[7];
  assign _T_139 = _T_130[8];
  assign _T_140 = _T_130[9];
  assign _T_141 = _T_130[10];
  assign _T_142 = _T_130[11];
  assign _T_143 = _T_130[12];
  assign _T_144 = _T_130[13];
  assign _T_145 = _T_130[14];
  assign _T_146 = _T_130[15];
  assign _T_147 = _T_130[16];
  assign _T_148 = _T_130[17];
  assign _T_149 = _T_130[18];
  assign _T_150 = _T_130[19];
  assign _T_151 = _T_130[20];
  assign _T_152 = _T_130[21];
  assign _T_153 = _T_130[22];
  assign _T_154 = _T_130[23];
  assign _T_155 = _T_130[24];
  assign _T_156 = {_T_133,_T_132};
  assign _T_157 = {_T_156,_T_131};
  assign _T_158 = {_T_136,_T_135};
  assign _T_159 = {_T_158,_T_134};
  assign _T_160 = {_T_159,_T_157};
  assign _T_161 = {_T_139,_T_138};
  assign _T_162 = {_T_161,_T_137};
  assign _T_163 = {_T_142,_T_141};
  assign _T_164 = {_T_163,_T_140};
  assign _T_165 = {_T_164,_T_162};
  assign _T_166 = {_T_165,_T_160};
  assign _T_167 = {_T_145,_T_144};
  assign _T_168 = {_T_167,_T_143};
  assign _T_169 = {_T_148,_T_147};
  assign _T_170 = {_T_169,_T_146};
  assign _T_171 = {_T_170,_T_168};
  assign _T_172 = {_T_151,_T_150};
  assign _T_173 = {_T_172,_T_149};
  assign _T_174 = {_T_153,_T_152};
  assign _T_175 = {_T_155,_T_154};
  assign _T_176 = {_T_175,_T_174};
  assign _T_177 = {_T_176,_T_173};
  assign _T_178 = {_T_177,_T_171};
  assign r_addr = {_T_178,_T_166};
  assign _T_179 = in_aw_bits_addr[27:3];
  assign _T_180 = _T_179[0];
  assign _T_181 = _T_179[1];
  assign _T_182 = _T_179[2];
  assign _T_183 = _T_179[3];
  assign _T_184 = _T_179[4];
  assign _T_185 = _T_179[5];
  assign _T_186 = _T_179[6];
  assign _T_187 = _T_179[7];
  assign _T_188 = _T_179[8];
  assign _T_189 = _T_179[9];
  assign _T_190 = _T_179[10];
  assign _T_191 = _T_179[11];
  assign _T_192 = _T_179[12];
  assign _T_193 = _T_179[13];
  assign _T_194 = _T_179[14];
  assign _T_195 = _T_179[15];
  assign _T_196 = _T_179[16];
  assign _T_197 = _T_179[17];
  assign _T_198 = _T_179[18];
  assign _T_199 = _T_179[19];
  assign _T_200 = _T_179[20];
  assign _T_201 = _T_179[21];
  assign _T_202 = _T_179[22];
  assign _T_203 = _T_179[23];
  assign _T_204 = _T_179[24];
  assign _T_205 = {_T_182,_T_181};
  assign _T_206 = {_T_205,_T_180};
  assign _T_207 = {_T_185,_T_184};
  assign _T_208 = {_T_207,_T_183};
  assign _T_209 = {_T_208,_T_206};
  assign _T_210 = {_T_188,_T_187};
  assign _T_211 = {_T_210,_T_186};
  assign _T_212 = {_T_191,_T_190};
  assign _T_213 = {_T_212,_T_189};
  assign _T_214 = {_T_213,_T_211};
  assign _T_215 = {_T_214,_T_209};
  assign _T_216 = {_T_194,_T_193};
  assign _T_217 = {_T_216,_T_192};
  assign _T_218 = {_T_197,_T_196};
  assign _T_219 = {_T_218,_T_195};
  assign _T_220 = {_T_219,_T_217};
  assign _T_221 = {_T_200,_T_199};
  assign _T_222 = {_T_221,_T_198};
  assign _T_223 = {_T_202,_T_201};
  assign _T_224 = {_T_204,_T_203};
  assign _T_225 = {_T_224,_T_223};
  assign _T_226 = {_T_225,_T_222};
  assign _T_227 = {_T_226,_T_220};
  assign w_addr = {_T_227,_T_215};
  assign _T_230 = {1'b0,$signed(in_ar_bits_addr)};
  assign _T_232 = $signed(_T_230) & $signed(-29'sh10000000);
  assign _T_233 = $signed(_T_232);
  assign r_sel0 = $signed(_T_233) == $signed(29'sh0);
  assign _T_237 = {1'b0,$signed(in_aw_bits_addr)};
  assign _T_239 = $signed(_T_237) & $signed(-29'sh10000000);
  assign _T_240 = $signed(_T_239);
  assign w_sel0 = $signed(_T_240) == $signed(29'sh0);
  assign _T_246 = in_b_ready & in_b_valid;
  assign _GEN_0 = _T_246 ? 1'h0 : w_full;
  assign _T_248 = in_aw_ready & in_aw_valid;
  assign _GEN_1 = _T_248 ? 1'h1 : _GEN_0;
  assign _GEN_2 = _T_248 ? in_aw_bits_id : w_id;
  assign _GEN_3 = _T_248 ? w_sel0 : w_sel1;
  assign _GEN_4 = _T_248 ? in_aw_bits_user : w_user;
  assign _T_251 = in_w_bits_data[7:0];
  assign _T_252 = in_w_bits_data[15:8];
  assign _T_253 = in_w_bits_data[23:16];
  assign _T_254 = in_w_bits_data[31:24];
  assign _T_255 = in_w_bits_data[39:32];
  assign _T_256 = in_w_bits_data[47:40];
  assign _T_257 = in_w_bits_data[55:48];
  assign _T_258 = in_w_bits_data[63:56];
  assign _T_272 = _T_248 & w_sel0;
  assign _T_273 = in_w_bits_strb[0];
  assign _T_274 = in_w_bits_strb[1];
  assign _T_275 = in_w_bits_strb[2];
  assign _T_276 = in_w_bits_strb[3];
  assign _T_277 = in_w_bits_strb[4];
  assign _T_278 = in_w_bits_strb[5];
  assign _T_279 = in_w_bits_strb[6];
  assign _T_280 = in_w_bits_strb[7];
  assign _GEN_25 = _T_272 ? _T_273 : 1'h0;
  assign _GEN_27 = _T_272 ? _T_274 : 1'h0;
  assign _GEN_29 = _T_272 ? _T_275 : 1'h0;
  assign _GEN_31 = _T_272 ? _T_276 : 1'h0;
  assign _GEN_33 = _T_272 ? _T_277 : 1'h0;
  assign _GEN_35 = _T_272 ? _T_278 : 1'h0;
  assign _GEN_37 = _T_272 ? _T_279 : 1'h0;
  assign _GEN_39 = _T_272 ? _T_280 : 1'h0;
  assign _T_302 = w_full == 1'h0;
  assign _T_303 = in_b_ready | _T_302;
  assign _T_304 = in_w_valid & _T_303;
  assign _T_308 = in_aw_valid & _T_303;
  assign _T_311 = w_sel1 ? 2'h0 : 2'h3;
  assign _T_316 = in_r_ready & in_r_valid;
  assign _GEN_40 = _T_316 ? 1'h0 : r_full;
  assign _T_318 = in_ar_ready & in_ar_valid;
  assign _GEN_41 = _T_318 ? 1'h1 : _GEN_40;
  assign _GEN_42 = _T_318 ? in_ar_bits_id : r_id;
  assign _GEN_43 = _T_318 ? r_sel0 : r_sel1;
  assign _GEN_44 = _T_318 ? in_ar_bits_user : r_user;
  assign ren = in_ar_ready & in_ar_valid;
  assign _GEN_49 = _T_347 ? mem_0__T_326_data : _T_377_0;
  assign _GEN_50 = _T_347 ? mem_1__T_326_data : _T_377_1;
  assign _GEN_51 = _T_347 ? mem_2__T_326_data : _T_377_2;
  assign _GEN_52 = _T_347 ? mem_3__T_326_data : _T_377_3;
  assign _GEN_53 = _T_347 ? mem_4__T_326_data : _T_377_4;
  assign _GEN_54 = _T_347 ? mem_5__T_326_data : _T_377_5;
  assign _GEN_55 = _T_347 ? mem_6__T_326_data : _T_377_6;
  assign _GEN_56 = _T_347 ? mem_7__T_326_data : _T_377_7;
  assign _T_444 = r_full == 1'h0;
  assign _T_445 = in_r_ready | _T_444;
  assign _T_448 = r_sel1 ? 2'h0 : 2'h3;
  assign _T_449 = {_GEN_50,_GEN_49};
  assign _T_450 = {_GEN_52,_GEN_51};
  assign _T_451 = {_T_450,_T_449};
  assign _T_452 = {_GEN_54,_GEN_53};
  assign _T_453 = {_GEN_56,_GEN_55};
  assign _T_454 = {_T_453,_T_452};
  assign _T_455 = {_T_454,_T_451};
  assign auto_in_aw_ready = in_aw_ready;
  assign auto_in_w_ready = in_w_ready;
  assign auto_in_b_valid = in_b_valid;
  assign auto_in_b_bits_id = in_b_bits_id;
  assign auto_in_b_bits_resp = in_b_bits_resp;
  assign auto_in_b_bits_user = in_b_bits_user;
  assign auto_in_ar_ready = in_ar_ready;
  assign auto_in_r_valid = in_r_valid;
  assign auto_in_r_bits_id = in_r_bits_id;
  assign auto_in_r_bits_data = in_r_bits_data;
  assign auto_in_r_bits_resp = in_r_bits_resp;
  assign auto_in_r_bits_user = in_r_bits_user;
  assign in_aw_ready = _T_304;
  assign in_aw_valid = auto_in_aw_valid;
  assign in_aw_bits_id = auto_in_aw_bits_id;
  assign in_aw_bits_addr = auto_in_aw_bits_addr;
  assign in_aw_bits_user = auto_in_aw_bits_user;
  assign in_w_ready = _T_308;
  assign in_w_valid = auto_in_w_valid;
  assign in_w_bits_data = auto_in_w_bits_data;
  assign in_w_bits_strb = auto_in_w_bits_strb;
  assign in_b_ready = auto_in_b_ready;
  assign in_b_valid = w_full;
  assign in_b_bits_id = w_id;
  assign in_b_bits_resp = _T_311;
  assign in_b_bits_user = w_user;
  assign in_ar_ready = _T_445;
  assign in_ar_valid = auto_in_ar_valid;
  assign in_ar_bits_id = auto_in_ar_bits_id;
  assign in_ar_bits_addr = auto_in_ar_bits_addr;
  assign in_ar_bits_user = auto_in_ar_bits_user;
  assign in_r_ready = auto_in_r_ready;
  assign in_r_valid = r_full;
  assign in_r_bits_id = r_id;
  assign in_r_bits_data = _T_455;
  assign in_r_bits_resp = _T_448;
  assign in_r_bits_user = r_user;
  assign wdata_0 = _T_251;
  assign wdata_1 = _T_252;
  assign wdata_2 = _T_253;
  assign wdata_3 = _T_254;
  assign wdata_4 = _T_255;
  assign wdata_5 = _T_256;
  assign wdata_6 = _T_257;
  assign wdata_7 = _T_258;
  assign _T_322 = r_addr;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0__T_326_addr_pipe_0 = _RAND_1[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_1[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_1__T_326_addr_pipe_0 = _RAND_3[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_2[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_2__T_326_addr_pipe_0 = _RAND_5[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_3[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_3__T_326_addr_pipe_0 = _RAND_7[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_4[initvar] = _RAND_8[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_4__T_326_addr_pipe_0 = _RAND_9[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_5[initvar] = _RAND_10[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_5__T_326_addr_pipe_0 = _RAND_11[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_6[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_6__T_326_addr_pipe_0 = _RAND_13[24:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 33554432; initvar = initvar+1)
    mem_7[initvar] = _RAND_14[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_7__T_326_addr_pipe_0 = _RAND_15[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  w_full = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  w_id = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  w_user = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  r_sel1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  w_sel1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  r_full = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  r_id = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  r_user = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_347 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_377_0 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_377_1 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_377_2 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_377_3 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_377_4 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_377_5 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_377_6 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_377_7 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_281_en & mem_0__T_281_mask) begin
      mem_0[mem_0__T_281_addr] <= mem_0__T_281_data;
    end
    if (_GEN_57) begin
      mem_0__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_1__T_281_en & mem_1__T_281_mask) begin
      mem_1[mem_1__T_281_addr] <= mem_1__T_281_data;
    end
    if (_GEN_57) begin
      mem_1__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_2__T_281_en & mem_2__T_281_mask) begin
      mem_2[mem_2__T_281_addr] <= mem_2__T_281_data;
    end
    if (_GEN_57) begin
      mem_2__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_3__T_281_en & mem_3__T_281_mask) begin
      mem_3[mem_3__T_281_addr] <= mem_3__T_281_data;
    end
    if (_GEN_57) begin
      mem_3__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_4__T_281_en & mem_4__T_281_mask) begin
      mem_4[mem_4__T_281_addr] <= mem_4__T_281_data;
    end
    if (_GEN_57) begin
      mem_4__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_5__T_281_en & mem_5__T_281_mask) begin
      mem_5[mem_5__T_281_addr] <= mem_5__T_281_data;
    end
    if (_GEN_57) begin
      mem_5__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_6__T_281_en & mem_6__T_281_mask) begin
      mem_6[mem_6__T_281_addr] <= mem_6__T_281_data;
    end
    if (_GEN_57) begin
      mem_6__T_326_addr_pipe_0 <= _T_322;
    end
    if(mem_7__T_281_en & mem_7__T_281_mask) begin
      mem_7[mem_7__T_281_addr] <= mem_7__T_281_data;
    end
    if (_GEN_57) begin
      mem_7__T_326_addr_pipe_0 <= _T_322;
    end
    if (reset) begin
      w_full <= 1'h0;
    end else begin
      if (_T_248) begin
        w_full <= 1'h1;
      end else begin
        if (_T_246) begin
          w_full <= 1'h0;
        end
      end
    end
    if (_T_248) begin
      w_id <= in_aw_bits_id;
    end
    if (_T_248) begin
      w_user <= in_aw_bits_user;
    end
    if (_T_318) begin
      r_sel1 <= r_sel0;
    end
    if (_T_248) begin
      w_sel1 <= w_sel0;
    end
    if (reset) begin
      r_full <= 1'h0;
    end else begin
      if (_T_318) begin
        r_full <= 1'h1;
      end else begin
        if (_T_316) begin
          r_full <= 1'h0;
        end
      end
    end
    if (_T_318) begin
      r_id <= in_ar_bits_id;
    end
    if (_T_318) begin
      r_user <= in_ar_bits_user;
    end
    _T_347 <= _T_318;
    if (_T_347) begin
      _T_377_0 <= mem_0__T_326_data;
    end
    if (_T_347) begin
      _T_377_1 <= mem_1__T_326_data;
    end
    if (_T_347) begin
      _T_377_2 <= mem_2__T_326_data;
    end
    if (_T_347) begin
      _T_377_3 <= mem_3__T_326_data;
    end
    if (_T_347) begin
      _T_377_4 <= mem_4__T_326_data;
    end
    if (_T_347) begin
      _T_377_5 <= mem_5__T_326_data;
    end
    if (_T_347) begin
      _T_377_6 <= mem_6__T_326_data;
    end
    if (_T_347) begin
      _T_377_7 <= mem_7__T_326_data;
    end
  end
endmodule
module Queue_115(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [27:0] io_enq_bits_addr,
  input         io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [27:0] io_deq_bits_addr,
  output        io_deq_bits_user
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [27:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [27:0] ram_addr__T_50_data;
  wire  ram_addr__T_50_addr;
  wire [27:0] ram_addr__T_36_data;
  wire  ram_addr__T_36_addr;
  wire  ram_addr__T_36_mask;
  wire  ram_addr__T_36_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_2;
  wire  ram_user__T_50_data;
  wire  ram_user__T_50_addr;
  wire  ram_user__T_36_data;
  wire  ram_user__T_36_addr;
  wire  ram_user__T_36_mask;
  wire  ram_user__T_36_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_13;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_14;
  wire  _T_45;
  wire  _GEN_15;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_addr__T_50_addr = value_1;
  assign ram_addr__T_50_data = ram_addr[ram_addr__T_50_addr];
  assign ram_addr__T_36_data = io_enq_bits_addr;
  assign ram_addr__T_36_addr = value;
  assign ram_addr__T_36_mask = do_enq;
  assign ram_addr__T_36_en = do_enq;
  assign ram_user__T_50_addr = value_1;
  assign ram_user__T_50_data = ram_user[ram_user__T_50_addr];
  assign ram_user__T_36_data = io_enq_bits_user;
  assign ram_user__T_36_addr = value;
  assign ram_user__T_36_mask = do_enq;
  assign ram_user__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_13 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_14 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_15 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_addr = ram_addr__T_50_data;
  assign io_deq_bits_user = ram_user__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[27:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_addr__T_36_en & ram_addr__T_36_mask) begin
      ram_addr[ram_addr__T_36_addr] <= ram_addr__T_36_data;
    end
    if(ram_user__T_36_en & ram_user__T_36_mask) begin
      ram_user[ram_user__T_36_addr] <= ram_user__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_117(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_enq_bits_user,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp,
  output       io_deq_bits_user
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_resp__T_50_data;
  wire  ram_resp__T_50_addr;
  wire [1:0] ram_resp__T_36_data;
  wire  ram_resp__T_36_addr;
  wire  ram_resp__T_36_mask;
  wire  ram_resp__T_36_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_2;
  wire  ram_user__T_50_data;
  wire  ram_user__T_50_addr;
  wire  ram_user__T_36_data;
  wire  ram_user__T_36_addr;
  wire  ram_user__T_36_mask;
  wire  ram_user__T_36_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_6;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_7;
  wire  _T_45;
  wire  _GEN_8;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_resp__T_50_addr = value_1;
  assign ram_resp__T_50_data = ram_resp[ram_resp__T_50_addr];
  assign ram_resp__T_36_data = io_enq_bits_resp;
  assign ram_resp__T_36_addr = value;
  assign ram_resp__T_36_mask = do_enq;
  assign ram_resp__T_36_en = do_enq;
  assign ram_user__T_50_addr = value_1;
  assign ram_user__T_50_data = ram_user[ram_user__T_50_addr];
  assign ram_user__T_36_data = io_enq_bits_user;
  assign ram_user__T_36_addr = value;
  assign ram_user__T_36_mask = do_enq;
  assign ram_user__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_6 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_7 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_8 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_resp = ram_resp__T_50_data;
  assign io_deq_bits_user = ram_user__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_resp__T_36_en & ram_resp__T_36_mask) begin
      ram_resp[ram_resp__T_36_addr] <= ram_resp__T_36_data;
    end
    if(ram_user__T_36_en & ram_user__T_36_mask) begin
      ram_user[ram_user__T_36_addr] <= ram_user__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_119(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_user,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_50_data;
  wire  ram_data__T_50_addr;
  wire [63:0] ram_data__T_36_data;
  wire  ram_data__T_36_addr;
  wire  ram_data__T_36_mask;
  wire  ram_data__T_36_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_50_data;
  wire  ram_resp__T_50_addr;
  wire [1:0] ram_resp__T_36_data;
  wire  ram_resp__T_36_addr;
  wire  ram_resp__T_36_mask;
  wire  ram_resp__T_36_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_3;
  wire  ram_user__T_50_data;
  wire  ram_user__T_50_addr;
  wire  ram_user__T_36_data;
  wire  ram_user__T_36_addr;
  wire  ram_user__T_36_mask;
  wire  ram_user__T_36_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_4;
  wire  ram_last__T_50_data;
  wire  ram_last__T_50_addr;
  wire  ram_last__T_36_data;
  wire  ram_last__T_36_addr;
  wire  ram_last__T_36_mask;
  wire  ram_last__T_36_en;
  reg  value;
  reg [31:0] _RAND_5;
  reg  value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_8;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_9;
  wire  _T_45;
  wire  _GEN_10;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_data__T_50_addr = value_1;
  assign ram_data__T_50_data = ram_data[ram_data__T_50_addr];
  assign ram_data__T_36_data = io_enq_bits_data;
  assign ram_data__T_36_addr = value;
  assign ram_data__T_36_mask = do_enq;
  assign ram_data__T_36_en = do_enq;
  assign ram_resp__T_50_addr = value_1;
  assign ram_resp__T_50_data = ram_resp[ram_resp__T_50_addr];
  assign ram_resp__T_36_data = io_enq_bits_resp;
  assign ram_resp__T_36_addr = value;
  assign ram_resp__T_36_mask = do_enq;
  assign ram_resp__T_36_en = do_enq;
  assign ram_user__T_50_addr = value_1;
  assign ram_user__T_50_data = ram_user[ram_user__T_50_addr];
  assign ram_user__T_36_data = io_enq_bits_user;
  assign ram_user__T_36_addr = value;
  assign ram_user__T_36_mask = do_enq;
  assign ram_user__T_36_en = do_enq;
  assign ram_last__T_50_addr = value_1;
  assign ram_last__T_50_data = ram_last[ram_last__T_50_addr];
  assign ram_last__T_36_data = 1'h1;
  assign ram_last__T_36_addr = value;
  assign ram_last__T_36_mask = do_enq;
  assign ram_last__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_8 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_9 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_10 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_data = ram_data__T_50_data;
  assign io_deq_bits_resp = ram_resp__T_50_data;
  assign io_deq_bits_user = ram_user__T_50_data;
  assign io_deq_bits_last = ram_last__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_data__T_36_en & ram_data__T_36_mask) begin
      ram_data[ram_data__T_36_addr] <= ram_data__T_36_data;
    end
    if(ram_resp__T_36_en & ram_resp__T_36_mask) begin
      ram_resp[ram_resp__T_36_addr] <= ram_resp__T_36_data;
    end
    if(ram_user__T_36_en & ram_user__T_36_mask) begin
      ram_user[ram_user__T_36_addr] <= ram_user__T_36_data;
    end
    if(ram_last__T_36_en & ram_last__T_36_mask) begin
      ram_last[ram_last__T_36_addr] <= ram_last__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Buffer_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [27:0] auto_in_aw_bits_addr,
  input         auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [27:0] auto_in_ar_bits_addr,
  input         auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [27:0] auto_out_aw_bits_addr,
  output        auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [27:0] auto_out_ar_bits_addr,
  output        auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_user
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [27:0] _T_31_aw_bits_addr;
  wire  _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [27:0] _T_31_ar_bits_addr;
  wire  _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [27:0] _T_89_aw_bits_addr;
  wire  _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [27:0] _T_89_ar_bits_addr;
  wire  _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_user;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [27:0] Queue_io_enq_bits_addr;
  wire  Queue_io_enq_bits_user;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [27:0] Queue_io_deq_bits_addr;
  wire  Queue_io_deq_bits_user;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [27:0] _T_207_bits_addr;
  wire  _T_207_bits_user;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_215_ready;
  wire  _T_215_valid;
  wire [63:0] _T_215_bits_data;
  wire [7:0] _T_215_bits_strb;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_enq_bits_user;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  Queue_2_io_deq_bits_user;
  wire  _T_223_ready;
  wire  _T_223_valid;
  wire [3:0] _T_223_bits_id;
  wire [1:0] _T_223_bits_resp;
  wire  _T_223_bits_user;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [27:0] Queue_3_io_enq_bits_addr;
  wire  Queue_3_io_enq_bits_user;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [27:0] Queue_3_io_deq_bits_addr;
  wire  Queue_3_io_deq_bits_user;
  wire  _T_231_ready;
  wire  _T_231_valid;
  wire [3:0] _T_231_bits_id;
  wire [27:0] _T_231_bits_addr;
  wire  _T_231_bits_user;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_user;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_user;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_239_ready;
  wire  _T_239_valid;
  wire [3:0] _T_239_bits_id;
  wire [63:0] _T_239_bits_data;
  wire [1:0] _T_239_bits_resp;
  wire  _T_239_bits_user;
  wire  _T_239_bits_last;
  Queue_115 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  Queue_67 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_117 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user)
  );
  Queue_115 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_user(Queue_3_io_deq_bits_user)
  );
  Queue_119 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_user(Queue_4_io_enq_bits_user),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_user(Queue_4_io_deq_bits_user),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = Queue_1_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_223_valid;
  assign _T_31_b_bits_id = _T_223_bits_id;
  assign _T_31_b_bits_resp = _T_223_bits_resp;
  assign _T_31_b_bits_user = _T_223_bits_user;
  assign _T_31_ar_ready = Queue_3_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_239_valid;
  assign _T_31_r_bits_id = _T_239_bits_id;
  assign _T_31_r_bits_data = _T_239_bits_data;
  assign _T_31_r_bits_resp = _T_239_bits_resp;
  assign _T_31_r_bits_user = _T_239_bits_user;
  assign _T_31_r_bits_last = _T_239_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_207_valid;
  assign _T_89_aw_bits_id = _T_207_bits_id;
  assign _T_89_aw_bits_addr = _T_207_bits_addr;
  assign _T_89_aw_bits_user = _T_207_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_215_valid;
  assign _T_89_w_bits_data = _T_215_bits_data;
  assign _T_89_w_bits_strb = _T_215_bits_strb;
  assign _T_89_b_ready = Queue_2_io_enq_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_231_valid;
  assign _T_89_ar_bits_id = _T_231_bits_id;
  assign _T_89_ar_bits_addr = _T_231_bits_addr;
  assign _T_89_ar_bits_user = _T_231_bits_user;
  assign _T_89_r_ready = Queue_4_io_enq_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign Queue_io_enq_valid = _T_31_aw_valid;
  assign Queue_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_io_enq_bits_user = _T_31_aw_bits_user;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_89_aw_ready;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_user = Queue_io_deq_bits_user;
  assign Queue_1_io_enq_valid = _T_31_w_valid;
  assign Queue_1_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_1_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_1_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_1_io_deq_ready = _T_215_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_215_ready = _T_89_w_ready;
  assign _T_215_valid = Queue_1_io_deq_valid;
  assign _T_215_bits_data = Queue_1_io_deq_bits_data;
  assign _T_215_bits_strb = Queue_1_io_deq_bits_strb;
  assign Queue_2_io_enq_valid = _T_89_b_valid;
  assign Queue_2_io_enq_bits_id = _T_89_b_bits_id;
  assign Queue_2_io_enq_bits_resp = _T_89_b_bits_resp;
  assign Queue_2_io_enq_bits_user = _T_89_b_bits_user;
  assign Queue_2_io_deq_ready = _T_223_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_223_ready = _T_31_b_ready;
  assign _T_223_valid = Queue_2_io_deq_valid;
  assign _T_223_bits_id = Queue_2_io_deq_bits_id;
  assign _T_223_bits_resp = Queue_2_io_deq_bits_resp;
  assign _T_223_bits_user = Queue_2_io_deq_bits_user;
  assign Queue_3_io_enq_valid = _T_31_ar_valid;
  assign Queue_3_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_3_io_enq_bits_user = _T_31_ar_bits_user;
  assign Queue_3_io_deq_ready = _T_231_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign _T_231_ready = _T_89_ar_ready;
  assign _T_231_valid = Queue_3_io_deq_valid;
  assign _T_231_bits_id = Queue_3_io_deq_bits_id;
  assign _T_231_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_231_bits_user = Queue_3_io_deq_bits_user;
  assign Queue_4_io_enq_valid = _T_89_r_valid;
  assign Queue_4_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_4_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_4_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_4_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_4_io_deq_ready = _T_239_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign _T_239_ready = _T_31_r_ready;
  assign _T_239_valid = Queue_4_io_deq_valid;
  assign _T_239_bits_id = Queue_4_io_deq_bits_id;
  assign _T_239_bits_data = Queue_4_io_deq_bits_data;
  assign _T_239_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_239_bits_user = Queue_4_io_deq_bits_user;
  assign _T_239_bits_last = Queue_4_io_deq_bits_last;
endmodule
module Queue_120(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [27:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [27:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst
);
  reg [3:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire [3:0] ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [27:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [27:0] ram_addr__T_42_data;
  wire  ram_addr__T_42_addr;
  wire [27:0] ram_addr__T_33_data;
  wire  ram_addr__T_33_addr;
  wire  ram_addr__T_33_mask;
  wire  ram_addr__T_33_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_42_data;
  wire  ram_len__T_42_addr;
  wire [7:0] ram_len__T_33_data;
  wire  ram_len__T_33_addr;
  wire  ram_len__T_33_mask;
  wire  ram_len__T_33_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [2:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_42_data;
  wire  ram_burst__T_42_addr;
  wire [1:0] ram_burst__T_33_data;
  wire  ram_burst__T_33_addr;
  wire  ram_burst__T_33_mask;
  wire  ram_burst__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_12;
  wire  _T_38;
  wire  _GEN_13;
  wire  _GEN_14;
  wire [1:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [7:0] _GEN_21;
  wire [27:0] _GEN_22;
  wire [3:0] _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_addr__T_42_addr = 1'h0;
  assign ram_addr__T_42_data = ram_addr[ram_addr__T_42_addr];
  assign ram_addr__T_33_data = io_enq_bits_addr;
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_mask = do_enq;
  assign ram_addr__T_33_en = do_enq;
  assign ram_len__T_42_addr = 1'h0;
  assign ram_len__T_42_data = ram_len[ram_len__T_42_addr];
  assign ram_len__T_33_data = io_enq_bits_len;
  assign ram_len__T_33_addr = 1'h0;
  assign ram_len__T_33_mask = do_enq;
  assign ram_len__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_burst__T_42_addr = 1'h0;
  assign ram_burst__T_42_data = ram_burst[ram_burst__T_42_addr];
  assign ram_burst__T_33_data = io_enq_bits_burst;
  assign ram_burst__T_33_addr = 1'h0;
  assign ram_burst__T_33_mask = do_enq;
  assign ram_burst__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_12 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_13 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_14 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_19 = empty ? io_enq_bits_burst : ram_burst__T_42_data;
  assign _GEN_20 = empty ? io_enq_bits_size : ram_size__T_42_data;
  assign _GEN_21 = empty ? io_enq_bits_len : ram_len__T_42_data;
  assign _GEN_22 = empty ? io_enq_bits_addr : ram_addr__T_42_data;
  assign _GEN_23 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_24 = empty ? 1'h0 : _T_30;
  assign _GEN_25 = empty ? _GEN_14 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_13;
  assign io_deq_bits_id = _GEN_23;
  assign io_deq_bits_addr = _GEN_22;
  assign io_deq_bits_len = _GEN_21;
  assign io_deq_bits_size = _GEN_20;
  assign io_deq_bits_burst = _GEN_19;
  assign do_enq = _GEN_25;
  assign do_deq = _GEN_24;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[27:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_addr__T_33_en & ram_addr__T_33_mask) begin
      ram_addr[ram_addr__T_33_addr] <= ram_addr__T_33_data;
    end
    if(ram_len__T_33_en & ram_len__T_33_mask) begin
      ram_len[ram_len__T_33_addr] <= ram_len__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_burst__T_33_en & ram_burst__T_33_mask) begin
      ram_burst[ram_burst__T_33_addr] <= ram_burst__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Fragmenter_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [27:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [27:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [27:0] auto_out_aw_bits_addr,
  output        auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [27:0] auto_out_ar_bits_addr,
  output        auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [27:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [27:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [27:0] _T_89_aw_bits_addr;
  wire  _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [27:0] _T_89_ar_bits_addr;
  wire  _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [27:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [27:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [27:0] _T_207_bits_addr;
  wire [7:0] _T_207_bits_len;
  wire [2:0] _T_207_bits_size;
  wire [1:0] _T_207_bits_burst;
  wire  _T_211_ready;
  wire  _T_211_valid;
  wire [3:0] _T_211_bits_id;
  wire [27:0] _T_211_bits_addr;
  reg  _T_217;
  reg [31:0] _RAND_0;
  reg [27:0] _T_219;
  reg [31:0] _RAND_1;
  reg [7:0] _T_221;
  reg [31:0] _RAND_2;
  wire [7:0] _T_222;
  wire [27:0] _T_223;
  wire  _T_271;
  wire [8:0] _T_277;
  wire [8:0] _T_279;
  wire [15:0] _GEN_54;
  wire [15:0] _T_284;
  wire [27:0] _GEN_55;
  wire [28:0] _T_285;
  wire [27:0] _T_286;
  wire [15:0] _T_288;
  wire [22:0] _GEN_56;
  wire [22:0] _T_289;
  wire [14:0] _T_290;
  wire [27:0] _T_292;
  wire  _T_294;
  wire [27:0] _GEN_57;
  wire [27:0] _T_295;
  wire [27:0] _T_296;
  wire [27:0] _T_297;
  wire [27:0] _T_298;
  wire [27:0] _T_299;
  wire [27:0] _GEN_1;
  wire [27:0] _GEN_2;
  wire  _T_302;
  wire  _T_303;
  wire [27:0] _T_304;
  wire [9:0] _T_307;
  wire [2:0] _T_308;
  wire [2:0] _T_309;
  wire [27:0] _GEN_59;
  wire [27:0] _T_310;
  wire [27:0] _T_311;
  wire  _T_312;
  wire  _T_314;
  wire [8:0] _GEN_60;
  wire [9:0] _T_315;
  wire [9:0] _T_316;
  wire [8:0] _T_317;
  wire  _GEN_3;
  wire [27:0] _GEN_4;
  wire [8:0] _GEN_5;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_id;
  wire [27:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_id;
  wire [27:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire  _T_322_ready;
  wire  _T_322_valid;
  wire [3:0] _T_322_bits_id;
  wire [27:0] _T_322_bits_addr;
  wire [7:0] _T_322_bits_len;
  wire [2:0] _T_322_bits_size;
  wire [1:0] _T_322_bits_burst;
  wire  _T_326_ready;
  wire  _T_326_valid;
  wire [3:0] _T_326_bits_id;
  wire [27:0] _T_326_bits_addr;
  reg  _T_332;
  reg [31:0] _RAND_3;
  reg [27:0] _T_334;
  reg [31:0] _RAND_4;
  reg [7:0] _T_336;
  reg [31:0] _RAND_5;
  wire [7:0] _T_337;
  wire [27:0] _T_338;
  wire  _T_386;
  wire [15:0] _T_399;
  wire [27:0] _GEN_72;
  wire [28:0] _T_400;
  wire [27:0] _T_401;
  wire [15:0] _T_403;
  wire [22:0] _GEN_73;
  wire [22:0] _T_404;
  wire [14:0] _T_405;
  wire [27:0] _T_407;
  wire  _T_409;
  wire [27:0] _GEN_74;
  wire [27:0] _T_410;
  wire [27:0] _T_411;
  wire [27:0] _T_412;
  wire [27:0] _T_413;
  wire [27:0] _T_414;
  wire [27:0] _GEN_6;
  wire [27:0] _GEN_7;
  wire  _T_417;
  wire  _T_418;
  wire [27:0] _T_419;
  wire [9:0] _T_422;
  wire [2:0] _T_423;
  wire [2:0] _T_424;
  wire [27:0] _GEN_76;
  wire [27:0] _T_425;
  wire [27:0] _T_426;
  wire  _T_427;
  wire  _T_429;
  wire [8:0] _GEN_77;
  wire [9:0] _T_430;
  wire [9:0] _T_431;
  wire [8:0] _T_432;
  wire  _GEN_8;
  wire [27:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [7:0] Queue_2_io_enq_bits_strb;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [7:0] Queue_2_io_deq_bits_strb;
  wire  Queue_2_io_deq_bits_last;
  wire  _T_437_ready;
  wire  _T_437_valid;
  wire [63:0] _T_437_bits_data;
  wire [7:0] _T_437_bits_strb;
  wire  _T_437_bits_last;
  reg  _T_443;
  reg [31:0] _RAND_6;
  wire  _T_445;
  wire  _T_447;
  wire  _T_448;
  wire  _GEN_11;
  wire  _T_450;
  wire  _GEN_12;
  wire  _T_452;
  wire  _T_453;
  wire  _T_455;
  wire  _T_457;
  wire  _T_458;
  reg [8:0] _T_461;
  reg [31:0] _RAND_7;
  wire  _T_463;
  wire [8:0] _T_465;
  wire [8:0] _T_466;
  wire  _T_468;
  wire  _T_469;
  wire [8:0] _GEN_78;
  wire [9:0] _T_470;
  wire [9:0] _T_471;
  wire [8:0] _T_472;
  wire  _T_475;
  wire  _T_477;
  wire  _T_478;
  wire  _T_480;
  wire  _T_482;
  wire  _T_484;
  wire  _T_485;
  wire  _T_486;
  wire  _T_490;
  wire  _T_492;
  wire  _T_494;
  wire  _T_495;
  wire  _T_496;
  wire  _T_498;
  wire  _T_500;
  wire  _T_502;
  wire  _T_504;
  wire  _T_506;
  wire  _T_507;
  reg [1:0] _T_581_0;
  reg [31:0] _RAND_8;
  reg [1:0] _T_581_1;
  reg [31:0] _RAND_9;
  reg [1:0] _T_581_2;
  reg [31:0] _RAND_10;
  reg [1:0] _T_581_3;
  reg [31:0] _RAND_11;
  reg [1:0] _T_581_4;
  reg [31:0] _RAND_12;
  reg [1:0] _T_581_5;
  reg [31:0] _RAND_13;
  reg [1:0] _T_581_6;
  reg [31:0] _RAND_14;
  reg [1:0] _T_581_7;
  reg [31:0] _RAND_15;
  reg [1:0] _T_581_8;
  reg [31:0] _RAND_16;
  reg [1:0] _T_581_9;
  reg [31:0] _RAND_17;
  reg [1:0] _T_581_10;
  reg [31:0] _RAND_18;
  reg [1:0] _T_581_11;
  reg [31:0] _RAND_19;
  reg [1:0] _T_581_12;
  reg [31:0] _RAND_20;
  reg [1:0] _T_581_13;
  reg [31:0] _RAND_21;
  reg [1:0] _T_581_14;
  reg [31:0] _RAND_22;
  reg [1:0] _T_581_15;
  reg [31:0] _RAND_23;
  wire [1:0] _GEN_0;
  wire [1:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire [1:0] _GEN_17;
  wire [1:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [1:0] _GEN_22;
  wire [1:0] _GEN_23;
  wire [1:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [1:0] _GEN_26;
  wire [1:0] _GEN_27;
  wire [1:0] _T_637;
  wire [15:0] _T_640;
  wire  _T_642;
  wire  _T_643;
  wire  _T_644;
  wire  _T_645;
  wire  _T_646;
  wire  _T_647;
  wire  _T_648;
  wire  _T_649;
  wire  _T_650;
  wire  _T_651;
  wire  _T_652;
  wire  _T_653;
  wire  _T_654;
  wire  _T_655;
  wire  _T_656;
  wire  _T_657;
  wire  _T_658;
  wire  _T_659;
  wire [1:0] _T_661;
  wire [1:0] _T_662;
  wire [1:0] _GEN_28;
  wire  _T_664;
  wire [1:0] _T_666;
  wire [1:0] _T_667;
  wire [1:0] _GEN_29;
  wire  _T_669;
  wire [1:0] _T_671;
  wire [1:0] _T_672;
  wire [1:0] _GEN_30;
  wire  _T_674;
  wire [1:0] _T_676;
  wire [1:0] _T_677;
  wire [1:0] _GEN_31;
  wire  _T_679;
  wire [1:0] _T_681;
  wire [1:0] _T_682;
  wire [1:0] _GEN_32;
  wire  _T_684;
  wire [1:0] _T_686;
  wire [1:0] _T_687;
  wire [1:0] _GEN_33;
  wire  _T_689;
  wire [1:0] _T_691;
  wire [1:0] _T_692;
  wire [1:0] _GEN_34;
  wire  _T_694;
  wire [1:0] _T_696;
  wire [1:0] _T_697;
  wire [1:0] _GEN_35;
  wire  _T_699;
  wire [1:0] _T_701;
  wire [1:0] _T_702;
  wire [1:0] _GEN_36;
  wire  _T_704;
  wire [1:0] _T_706;
  wire [1:0] _T_707;
  wire [1:0] _GEN_37;
  wire  _T_709;
  wire [1:0] _T_711;
  wire [1:0] _T_712;
  wire [1:0] _GEN_38;
  wire  _T_714;
  wire [1:0] _T_716;
  wire [1:0] _T_717;
  wire [1:0] _GEN_39;
  wire  _T_719;
  wire [1:0] _T_721;
  wire [1:0] _T_722;
  wire [1:0] _GEN_40;
  wire  _T_724;
  wire [1:0] _T_726;
  wire [1:0] _T_727;
  wire [1:0] _GEN_41;
  wire  _T_729;
  wire [1:0] _T_731;
  wire [1:0] _T_732;
  wire [1:0] _GEN_42;
  wire  _T_734;
  wire [1:0] _T_736;
  wire [1:0] _T_737;
  wire [1:0] _GEN_43;
  Queue_120 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst)
  );
  Queue_120 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst)
  );
  Queue_32 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign _T_222 = _T_217 ? _T_221 : _T_207_bits_len;
  assign _T_223 = _T_217 ? _T_219 : _T_207_bits_addr;
  assign _T_271 = _T_207_bits_burst == 2'h0;
  assign _T_277 = 9'h0 << 1;
  assign _T_279 = _T_277 | 9'h1;
  assign _GEN_54 = {{7'd0}, _T_279};
  assign _T_284 = _GEN_54 << _T_207_bits_size;
  assign _GEN_55 = {{12'd0}, _T_284};
  assign _T_285 = _T_223 + _GEN_55;
  assign _T_286 = _T_285[27:0];
  assign _T_288 = {_T_207_bits_len,8'hff};
  assign _GEN_56 = {{7'd0}, _T_288};
  assign _T_289 = _GEN_56 << _T_207_bits_size;
  assign _T_290 = _T_289[22:8];
  assign _T_294 = _T_207_bits_burst == 2'h2;
  assign _GEN_57 = {{13'd0}, _T_290};
  assign _T_295 = _T_286 & _GEN_57;
  assign _T_296 = ~ _T_207_bits_addr;
  assign _T_297 = _T_296 | _GEN_57;
  assign _T_298 = ~ _T_297;
  assign _T_299 = _T_295 | _T_298;
  assign _GEN_1 = _T_294 ? _T_299 : _T_286;
  assign _GEN_2 = _T_271 ? _T_207_bits_addr : _GEN_1;
  assign _T_302 = 8'h0 == _T_222;
  assign _T_303 = _T_211_ready & _T_302;
  assign _T_304 = ~ _T_223;
  assign _T_307 = 10'h7 << _T_207_bits_size;
  assign _T_308 = _T_307[2:0];
  assign _T_309 = ~ _T_308;
  assign _GEN_59 = {{25'd0}, _T_309};
  assign _T_310 = _T_304 | _GEN_59;
  assign _T_311 = ~ _T_310;
  assign _T_312 = _T_211_ready & _T_211_valid;
  assign _T_314 = _T_302 == 1'h0;
  assign _GEN_60 = {{1'd0}, _T_222};
  assign _T_315 = _GEN_60 - _T_279;
  assign _T_316 = $unsigned(_T_315);
  assign _T_317 = _T_316[8:0];
  assign _GEN_3 = _T_312 ? _T_314 : _T_217;
  assign _GEN_4 = _T_312 ? _T_292 : _T_219;
  assign _GEN_5 = _T_312 ? _T_317 : {{1'd0}, _T_221};
  assign _T_337 = _T_332 ? _T_336 : _T_322_bits_len;
  assign _T_338 = _T_332 ? _T_334 : _T_322_bits_addr;
  assign _T_386 = _T_322_bits_burst == 2'h0;
  assign _T_399 = _GEN_54 << _T_322_bits_size;
  assign _GEN_72 = {{12'd0}, _T_399};
  assign _T_400 = _T_338 + _GEN_72;
  assign _T_401 = _T_400[27:0];
  assign _T_403 = {_T_322_bits_len,8'hff};
  assign _GEN_73 = {{7'd0}, _T_403};
  assign _T_404 = _GEN_73 << _T_322_bits_size;
  assign _T_405 = _T_404[22:8];
  assign _T_409 = _T_322_bits_burst == 2'h2;
  assign _GEN_74 = {{13'd0}, _T_405};
  assign _T_410 = _T_401 & _GEN_74;
  assign _T_411 = ~ _T_322_bits_addr;
  assign _T_412 = _T_411 | _GEN_74;
  assign _T_413 = ~ _T_412;
  assign _T_414 = _T_410 | _T_413;
  assign _GEN_6 = _T_409 ? _T_414 : _T_401;
  assign _GEN_7 = _T_386 ? _T_322_bits_addr : _GEN_6;
  assign _T_417 = 8'h0 == _T_337;
  assign _T_418 = _T_326_ready & _T_417;
  assign _T_419 = ~ _T_338;
  assign _T_422 = 10'h7 << _T_322_bits_size;
  assign _T_423 = _T_422[2:0];
  assign _T_424 = ~ _T_423;
  assign _GEN_76 = {{25'd0}, _T_424};
  assign _T_425 = _T_419 | _GEN_76;
  assign _T_426 = ~ _T_425;
  assign _T_427 = _T_326_ready & _T_326_valid;
  assign _T_429 = _T_417 == 1'h0;
  assign _GEN_77 = {{1'd0}, _T_337};
  assign _T_430 = _GEN_77 - _T_279;
  assign _T_431 = $unsigned(_T_430);
  assign _T_432 = _T_431[8:0];
  assign _GEN_8 = _T_427 ? _T_429 : _T_332;
  assign _GEN_9 = _T_427 ? _T_407 : _T_334;
  assign _GEN_10 = _T_427 ? _T_432 : {{1'd0}, _T_336};
  assign _T_448 = _T_447 & _T_445;
  assign _GEN_11 = _T_448 ? 1'h1 : _T_443;
  assign _T_450 = _T_89_aw_ready & _T_89_aw_valid;
  assign _GEN_12 = _T_450 ? 1'h0 : _GEN_11;
  assign _T_452 = _T_445 | _T_443;
  assign _T_453 = _T_326_valid & _T_452;
  assign _T_455 = _T_89_aw_ready & _T_452;
  assign _T_457 = _T_443 == 1'h0;
  assign _T_458 = _T_326_valid & _T_457;
  assign _T_463 = _T_461 == 9'h0;
  assign _T_465 = _T_447 ? _T_279 : 9'h0;
  assign _T_466 = _T_463 ? _T_465 : _T_461;
  assign _T_468 = _T_466 == 9'h1;
  assign _T_469 = _T_89_w_ready & _T_89_w_valid;
  assign _GEN_78 = {{8'd0}, _T_469};
  assign _T_470 = _T_466 - _GEN_78;
  assign _T_471 = $unsigned(_T_470);
  assign _T_472 = _T_471[8:0];
  assign _T_475 = _T_469 == 1'h0;
  assign _T_477 = _T_466 != 9'h0;
  assign _T_478 = _T_475 | _T_477;
  assign _T_480 = _T_478 | reset;
  assign _T_482 = _T_480 == 1'h0;
  assign _T_484 = _T_445 == 1'h0;
  assign _T_485 = _T_484 | _T_447;
  assign _T_486 = _T_437_valid & _T_485;
  assign _T_490 = _T_89_w_ready & _T_485;
  assign _T_492 = _T_89_w_valid == 1'h0;
  assign _T_494 = _T_437_bits_last == 1'h0;
  assign _T_495 = _T_492 | _T_494;
  assign _T_496 = _T_495 | _T_468;
  assign _T_498 = _T_496 | reset;
  assign _T_500 = _T_498 == 1'h0;
  assign _T_502 = _T_89_r_bits_last & _T_89_r_bits_user;
  assign _T_504 = _T_89_b_valid & _T_89_b_bits_user;
  assign _T_506 = _T_89_b_bits_user == 1'h0;
  assign _T_507 = _T_31_b_ready | _T_506;
  assign _GEN_13 = 4'h1 == _T_89_b_bits_id ? _T_581_1 : _T_581_0;
  assign _GEN_14 = 4'h2 == _T_89_b_bits_id ? _T_581_2 : _GEN_13;
  assign _GEN_15 = 4'h3 == _T_89_b_bits_id ? _T_581_3 : _GEN_14;
  assign _GEN_16 = 4'h4 == _T_89_b_bits_id ? _T_581_4 : _GEN_15;
  assign _GEN_17 = 4'h5 == _T_89_b_bits_id ? _T_581_5 : _GEN_16;
  assign _GEN_18 = 4'h6 == _T_89_b_bits_id ? _T_581_6 : _GEN_17;
  assign _GEN_19 = 4'h7 == _T_89_b_bits_id ? _T_581_7 : _GEN_18;
  assign _GEN_20 = 4'h8 == _T_89_b_bits_id ? _T_581_8 : _GEN_19;
  assign _GEN_21 = 4'h9 == _T_89_b_bits_id ? _T_581_9 : _GEN_20;
  assign _GEN_22 = 4'ha == _T_89_b_bits_id ? _T_581_10 : _GEN_21;
  assign _GEN_23 = 4'hb == _T_89_b_bits_id ? _T_581_11 : _GEN_22;
  assign _GEN_24 = 4'hc == _T_89_b_bits_id ? _T_581_12 : _GEN_23;
  assign _GEN_25 = 4'hd == _T_89_b_bits_id ? _T_581_13 : _GEN_24;
  assign _GEN_26 = 4'he == _T_89_b_bits_id ? _T_581_14 : _GEN_25;
  assign _GEN_27 = 4'hf == _T_89_b_bits_id ? _T_581_15 : _GEN_26;
  assign _T_637 = _T_89_b_bits_resp | _GEN_0;
  assign _T_640 = 16'h1 << _T_89_b_bits_id;
  assign _T_642 = _T_640[0];
  assign _T_643 = _T_640[1];
  assign _T_644 = _T_640[2];
  assign _T_645 = _T_640[3];
  assign _T_646 = _T_640[4];
  assign _T_647 = _T_640[5];
  assign _T_648 = _T_640[6];
  assign _T_649 = _T_640[7];
  assign _T_650 = _T_640[8];
  assign _T_651 = _T_640[9];
  assign _T_652 = _T_640[10];
  assign _T_653 = _T_640[11];
  assign _T_654 = _T_640[12];
  assign _T_655 = _T_640[13];
  assign _T_656 = _T_640[14];
  assign _T_657 = _T_640[15];
  assign _T_658 = _T_89_b_ready & _T_89_b_valid;
  assign _T_659 = _T_642 & _T_658;
  assign _T_661 = _T_581_0 | _T_89_b_bits_resp;
  assign _T_662 = _T_89_b_bits_user ? 2'h0 : _T_661;
  assign _GEN_28 = _T_659 ? _T_662 : _T_581_0;
  assign _T_664 = _T_643 & _T_658;
  assign _T_666 = _T_581_1 | _T_89_b_bits_resp;
  assign _T_667 = _T_89_b_bits_user ? 2'h0 : _T_666;
  assign _GEN_29 = _T_664 ? _T_667 : _T_581_1;
  assign _T_669 = _T_644 & _T_658;
  assign _T_671 = _T_581_2 | _T_89_b_bits_resp;
  assign _T_672 = _T_89_b_bits_user ? 2'h0 : _T_671;
  assign _GEN_30 = _T_669 ? _T_672 : _T_581_2;
  assign _T_674 = _T_645 & _T_658;
  assign _T_676 = _T_581_3 | _T_89_b_bits_resp;
  assign _T_677 = _T_89_b_bits_user ? 2'h0 : _T_676;
  assign _GEN_31 = _T_674 ? _T_677 : _T_581_3;
  assign _T_679 = _T_646 & _T_658;
  assign _T_681 = _T_581_4 | _T_89_b_bits_resp;
  assign _T_682 = _T_89_b_bits_user ? 2'h0 : _T_681;
  assign _GEN_32 = _T_679 ? _T_682 : _T_581_4;
  assign _T_684 = _T_647 & _T_658;
  assign _T_686 = _T_581_5 | _T_89_b_bits_resp;
  assign _T_687 = _T_89_b_bits_user ? 2'h0 : _T_686;
  assign _GEN_33 = _T_684 ? _T_687 : _T_581_5;
  assign _T_689 = _T_648 & _T_658;
  assign _T_691 = _T_581_6 | _T_89_b_bits_resp;
  assign _T_692 = _T_89_b_bits_user ? 2'h0 : _T_691;
  assign _GEN_34 = _T_689 ? _T_692 : _T_581_6;
  assign _T_694 = _T_649 & _T_658;
  assign _T_696 = _T_581_7 | _T_89_b_bits_resp;
  assign _T_697 = _T_89_b_bits_user ? 2'h0 : _T_696;
  assign _GEN_35 = _T_694 ? _T_697 : _T_581_7;
  assign _T_699 = _T_650 & _T_658;
  assign _T_701 = _T_581_8 | _T_89_b_bits_resp;
  assign _T_702 = _T_89_b_bits_user ? 2'h0 : _T_701;
  assign _GEN_36 = _T_699 ? _T_702 : _T_581_8;
  assign _T_704 = _T_651 & _T_658;
  assign _T_706 = _T_581_9 | _T_89_b_bits_resp;
  assign _T_707 = _T_89_b_bits_user ? 2'h0 : _T_706;
  assign _GEN_37 = _T_704 ? _T_707 : _T_581_9;
  assign _T_709 = _T_652 & _T_658;
  assign _T_711 = _T_581_10 | _T_89_b_bits_resp;
  assign _T_712 = _T_89_b_bits_user ? 2'h0 : _T_711;
  assign _GEN_38 = _T_709 ? _T_712 : _T_581_10;
  assign _T_714 = _T_653 & _T_658;
  assign _T_716 = _T_581_11 | _T_89_b_bits_resp;
  assign _T_717 = _T_89_b_bits_user ? 2'h0 : _T_716;
  assign _GEN_39 = _T_714 ? _T_717 : _T_581_11;
  assign _T_719 = _T_654 & _T_658;
  assign _T_721 = _T_581_12 | _T_89_b_bits_resp;
  assign _T_722 = _T_89_b_bits_user ? 2'h0 : _T_721;
  assign _GEN_40 = _T_719 ? _T_722 : _T_581_12;
  assign _T_724 = _T_655 & _T_658;
  assign _T_726 = _T_581_13 | _T_89_b_bits_resp;
  assign _T_727 = _T_89_b_bits_user ? 2'h0 : _T_726;
  assign _GEN_41 = _T_724 ? _T_727 : _T_581_13;
  assign _T_729 = _T_656 & _T_658;
  assign _T_731 = _T_581_14 | _T_89_b_bits_resp;
  assign _T_732 = _T_89_b_bits_user ? 2'h0 : _T_731;
  assign _GEN_42 = _T_729 ? _T_732 : _T_581_14;
  assign _T_734 = _T_657 & _T_658;
  assign _T_736 = _T_581_15 | _T_89_b_bits_resp;
  assign _T_737 = _T_89_b_bits_user ? 2'h0 : _T_736;
  assign _GEN_43 = _T_734 ? _T_737 : _T_581_15;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_1_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_w_ready = Queue_2_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_504;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_637;
  assign _T_31_ar_ready = Queue_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_last = _T_502;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_453;
  assign _T_89_aw_bits_id = _T_326_bits_id;
  assign _T_89_aw_bits_addr = _T_326_bits_addr;
  assign _T_89_aw_bits_user = _T_417;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_486;
  assign _T_89_w_bits_data = _T_437_bits_data;
  assign _T_89_w_bits_strb = _T_437_bits_strb;
  assign _T_89_w_bits_last = _T_468;
  assign _T_89_b_ready = _T_507;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_211_valid;
  assign _T_89_ar_bits_id = _T_211_bits_id;
  assign _T_89_ar_bits_addr = _T_211_bits_addr;
  assign _T_89_ar_bits_user = _T_302;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_31_ar_valid;
  assign Queue_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_io_enq_bits_len = _T_31_ar_bits_len;
  assign Queue_io_enq_bits_size = _T_31_ar_bits_size;
  assign Queue_io_enq_bits_burst = _T_31_ar_bits_burst;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_303;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_len = Queue_io_deq_bits_len;
  assign _T_207_bits_size = Queue_io_deq_bits_size;
  assign _T_207_bits_burst = Queue_io_deq_bits_burst;
  assign _T_211_ready = _T_89_ar_ready;
  assign _T_211_valid = _T_207_valid;
  assign _T_211_bits_id = _T_207_bits_id;
  assign _T_211_bits_addr = _T_311;
  assign _T_292 = _GEN_2;
  assign Queue_1_io_enq_valid = _T_31_aw_valid;
  assign Queue_1_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_1_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_1_io_enq_bits_len = _T_31_aw_bits_len;
  assign Queue_1_io_enq_bits_size = _T_31_aw_bits_size;
  assign Queue_1_io_enq_bits_burst = _T_31_aw_bits_burst;
  assign Queue_1_io_deq_ready = _T_322_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_322_ready = _T_418;
  assign _T_322_valid = Queue_1_io_deq_valid;
  assign _T_322_bits_id = Queue_1_io_deq_bits_id;
  assign _T_322_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_322_bits_len = Queue_1_io_deq_bits_len;
  assign _T_322_bits_size = Queue_1_io_deq_bits_size;
  assign _T_322_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_326_ready = _T_455;
  assign _T_326_valid = _T_322_valid;
  assign _T_326_bits_id = _T_322_bits_id;
  assign _T_326_bits_addr = _T_426;
  assign _T_407 = _GEN_7;
  assign Queue_2_io_enq_valid = _T_31_w_valid;
  assign Queue_2_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_2_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_2_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_2_io_deq_ready = _T_437_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_437_ready = _T_490;
  assign _T_437_valid = Queue_2_io_deq_valid;
  assign _T_437_bits_data = Queue_2_io_deq_bits_data;
  assign _T_437_bits_strb = Queue_2_io_deq_bits_strb;
  assign _T_437_bits_last = Queue_2_io_deq_bits_last;
  assign _T_445 = _T_463;
  assign _T_447 = _T_458;
  assign _GEN_0 = _GEN_27;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_217 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_219 = _RAND_1[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_221 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_332 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_334 = _RAND_4[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_336 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_443 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_461 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_581_0 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_581_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_581_2 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_581_3 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_581_4 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_581_5 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_581_6 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_581_7 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_581_8 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_581_9 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_581_10 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_581_11 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_581_12 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_581_13 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_581_14 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_581_15 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_217 <= 1'h0;
    end else begin
      if (_T_312) begin
        _T_217 <= _T_314;
      end
    end
    if (_T_312) begin
      _T_219 <= _T_292;
    end
    _T_221 <= _GEN_5[7:0];
    if (reset) begin
      _T_332 <= 1'h0;
    end else begin
      if (_T_427) begin
        _T_332 <= _T_429;
      end
    end
    if (_T_427) begin
      _T_334 <= _T_407;
    end
    _T_336 <= _GEN_10[7:0];
    if (reset) begin
      _T_443 <= 1'h0;
    end else begin
      if (_T_450) begin
        _T_443 <= 1'h0;
      end else begin
        if (_T_448) begin
          _T_443 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_461 <= 9'h0;
    end else begin
      _T_461 <= _T_472;
    end
    if (reset) begin
      _T_581_0 <= 2'h0;
    end else begin
      if (_T_659) begin
        if (_T_89_b_bits_user) begin
          _T_581_0 <= 2'h0;
        end else begin
          _T_581_0 <= _T_661;
        end
      end
    end
    if (reset) begin
      _T_581_1 <= 2'h0;
    end else begin
      if (_T_664) begin
        if (_T_89_b_bits_user) begin
          _T_581_1 <= 2'h0;
        end else begin
          _T_581_1 <= _T_666;
        end
      end
    end
    if (reset) begin
      _T_581_2 <= 2'h0;
    end else begin
      if (_T_669) begin
        if (_T_89_b_bits_user) begin
          _T_581_2 <= 2'h0;
        end else begin
          _T_581_2 <= _T_671;
        end
      end
    end
    if (reset) begin
      _T_581_3 <= 2'h0;
    end else begin
      if (_T_674) begin
        if (_T_89_b_bits_user) begin
          _T_581_3 <= 2'h0;
        end else begin
          _T_581_3 <= _T_676;
        end
      end
    end
    if (reset) begin
      _T_581_4 <= 2'h0;
    end else begin
      if (_T_679) begin
        if (_T_89_b_bits_user) begin
          _T_581_4 <= 2'h0;
        end else begin
          _T_581_4 <= _T_681;
        end
      end
    end
    if (reset) begin
      _T_581_5 <= 2'h0;
    end else begin
      if (_T_684) begin
        if (_T_89_b_bits_user) begin
          _T_581_5 <= 2'h0;
        end else begin
          _T_581_5 <= _T_686;
        end
      end
    end
    if (reset) begin
      _T_581_6 <= 2'h0;
    end else begin
      if (_T_689) begin
        if (_T_89_b_bits_user) begin
          _T_581_6 <= 2'h0;
        end else begin
          _T_581_6 <= _T_691;
        end
      end
    end
    if (reset) begin
      _T_581_7 <= 2'h0;
    end else begin
      if (_T_694) begin
        if (_T_89_b_bits_user) begin
          _T_581_7 <= 2'h0;
        end else begin
          _T_581_7 <= _T_696;
        end
      end
    end
    if (reset) begin
      _T_581_8 <= 2'h0;
    end else begin
      if (_T_699) begin
        if (_T_89_b_bits_user) begin
          _T_581_8 <= 2'h0;
        end else begin
          _T_581_8 <= _T_701;
        end
      end
    end
    if (reset) begin
      _T_581_9 <= 2'h0;
    end else begin
      if (_T_704) begin
        if (_T_89_b_bits_user) begin
          _T_581_9 <= 2'h0;
        end else begin
          _T_581_9 <= _T_706;
        end
      end
    end
    if (reset) begin
      _T_581_10 <= 2'h0;
    end else begin
      if (_T_709) begin
        if (_T_89_b_bits_user) begin
          _T_581_10 <= 2'h0;
        end else begin
          _T_581_10 <= _T_711;
        end
      end
    end
    if (reset) begin
      _T_581_11 <= 2'h0;
    end else begin
      if (_T_714) begin
        if (_T_89_b_bits_user) begin
          _T_581_11 <= 2'h0;
        end else begin
          _T_581_11 <= _T_716;
        end
      end
    end
    if (reset) begin
      _T_581_12 <= 2'h0;
    end else begin
      if (_T_719) begin
        if (_T_89_b_bits_user) begin
          _T_581_12 <= 2'h0;
        end else begin
          _T_581_12 <= _T_721;
        end
      end
    end
    if (reset) begin
      _T_581_13 <= 2'h0;
    end else begin
      if (_T_724) begin
        if (_T_89_b_bits_user) begin
          _T_581_13 <= 2'h0;
        end else begin
          _T_581_13 <= _T_726;
        end
      end
    end
    if (reset) begin
      _T_581_14 <= 2'h0;
    end else begin
      if (_T_729) begin
        if (_T_89_b_bits_user) begin
          _T_581_14 <= 2'h0;
        end else begin
          _T_581_14 <= _T_731;
        end
      end
    end
    if (reset) begin
      _T_581_15 <= 2'h0;
    end else begin
      if (_T_734) begin
        if (_T_89_b_bits_user) begin
          _T_581_15 <= 2'h0;
        end else begin
          _T_581_15 <= _T_736;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_482) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:166 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_482) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_500) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:175 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_500) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimAXIMem(
  input         clock,
  input         reset,
  output        io_axi4_0_aw_ready,
  input         io_axi4_0_aw_valid,
  input  [3:0]  io_axi4_0_aw_bits_id,
  input  [27:0] io_axi4_0_aw_bits_addr,
  input  [7:0]  io_axi4_0_aw_bits_len,
  input  [2:0]  io_axi4_0_aw_bits_size,
  input  [1:0]  io_axi4_0_aw_bits_burst,
  output        io_axi4_0_w_ready,
  input         io_axi4_0_w_valid,
  input  [63:0] io_axi4_0_w_bits_data,
  input  [7:0]  io_axi4_0_w_bits_strb,
  input         io_axi4_0_w_bits_last,
  input         io_axi4_0_b_ready,
  output        io_axi4_0_b_valid,
  output [3:0]  io_axi4_0_b_bits_id,
  output [1:0]  io_axi4_0_b_bits_resp,
  output        io_axi4_0_ar_ready,
  input         io_axi4_0_ar_valid,
  input  [3:0]  io_axi4_0_ar_bits_id,
  input  [27:0] io_axi4_0_ar_bits_addr,
  input  [7:0]  io_axi4_0_ar_bits_len,
  input  [2:0]  io_axi4_0_ar_bits_size,
  input  [1:0]  io_axi4_0_ar_bits_burst,
  input         io_axi4_0_r_ready,
  output        io_axi4_0_r_valid,
  output [3:0]  io_axi4_0_r_bits_id,
  output [63:0] io_axi4_0_r_bits_data,
  output [1:0]  io_axi4_0_r_bits_resp,
  output        io_axi4_0_r_bits_last
);
  wire  AXI4RAM_clock;
  wire  AXI4RAM_reset;
  wire  AXI4RAM_auto_in_aw_ready;
  wire  AXI4RAM_auto_in_aw_valid;
  wire [3:0] AXI4RAM_auto_in_aw_bits_id;
  wire [27:0] AXI4RAM_auto_in_aw_bits_addr;
  wire  AXI4RAM_auto_in_aw_bits_user;
  wire  AXI4RAM_auto_in_w_ready;
  wire  AXI4RAM_auto_in_w_valid;
  wire [63:0] AXI4RAM_auto_in_w_bits_data;
  wire [7:0] AXI4RAM_auto_in_w_bits_strb;
  wire  AXI4RAM_auto_in_b_ready;
  wire  AXI4RAM_auto_in_b_valid;
  wire [3:0] AXI4RAM_auto_in_b_bits_id;
  wire [1:0] AXI4RAM_auto_in_b_bits_resp;
  wire  AXI4RAM_auto_in_b_bits_user;
  wire  AXI4RAM_auto_in_ar_ready;
  wire  AXI4RAM_auto_in_ar_valid;
  wire [3:0] AXI4RAM_auto_in_ar_bits_id;
  wire [27:0] AXI4RAM_auto_in_ar_bits_addr;
  wire  AXI4RAM_auto_in_ar_bits_user;
  wire  AXI4RAM_auto_in_r_ready;
  wire  AXI4RAM_auto_in_r_valid;
  wire [3:0] AXI4RAM_auto_in_r_bits_id;
  wire [63:0] AXI4RAM_auto_in_r_bits_data;
  wire [1:0] AXI4RAM_auto_in_r_bits_resp;
  wire  AXI4RAM_auto_in_r_bits_user;
  wire  AXI4Buffer_clock;
  wire  AXI4Buffer_reset;
  wire  AXI4Buffer_auto_in_aw_ready;
  wire  AXI4Buffer_auto_in_aw_valid;
  wire [3:0] AXI4Buffer_auto_in_aw_bits_id;
  wire [27:0] AXI4Buffer_auto_in_aw_bits_addr;
  wire  AXI4Buffer_auto_in_aw_bits_user;
  wire  AXI4Buffer_auto_in_w_ready;
  wire  AXI4Buffer_auto_in_w_valid;
  wire [63:0] AXI4Buffer_auto_in_w_bits_data;
  wire [7:0] AXI4Buffer_auto_in_w_bits_strb;
  wire  AXI4Buffer_auto_in_w_bits_last;
  wire  AXI4Buffer_auto_in_b_ready;
  wire  AXI4Buffer_auto_in_b_valid;
  wire [3:0] AXI4Buffer_auto_in_b_bits_id;
  wire [1:0] AXI4Buffer_auto_in_b_bits_resp;
  wire  AXI4Buffer_auto_in_b_bits_user;
  wire  AXI4Buffer_auto_in_ar_ready;
  wire  AXI4Buffer_auto_in_ar_valid;
  wire [3:0] AXI4Buffer_auto_in_ar_bits_id;
  wire [27:0] AXI4Buffer_auto_in_ar_bits_addr;
  wire  AXI4Buffer_auto_in_ar_bits_user;
  wire  AXI4Buffer_auto_in_r_ready;
  wire  AXI4Buffer_auto_in_r_valid;
  wire [3:0] AXI4Buffer_auto_in_r_bits_id;
  wire [63:0] AXI4Buffer_auto_in_r_bits_data;
  wire [1:0] AXI4Buffer_auto_in_r_bits_resp;
  wire  AXI4Buffer_auto_in_r_bits_user;
  wire  AXI4Buffer_auto_in_r_bits_last;
  wire  AXI4Buffer_auto_out_aw_ready;
  wire  AXI4Buffer_auto_out_aw_valid;
  wire [3:0] AXI4Buffer_auto_out_aw_bits_id;
  wire [27:0] AXI4Buffer_auto_out_aw_bits_addr;
  wire  AXI4Buffer_auto_out_aw_bits_user;
  wire  AXI4Buffer_auto_out_w_ready;
  wire  AXI4Buffer_auto_out_w_valid;
  wire [63:0] AXI4Buffer_auto_out_w_bits_data;
  wire [7:0] AXI4Buffer_auto_out_w_bits_strb;
  wire  AXI4Buffer_auto_out_b_ready;
  wire  AXI4Buffer_auto_out_b_valid;
  wire [3:0] AXI4Buffer_auto_out_b_bits_id;
  wire [1:0] AXI4Buffer_auto_out_b_bits_resp;
  wire  AXI4Buffer_auto_out_b_bits_user;
  wire  AXI4Buffer_auto_out_ar_ready;
  wire  AXI4Buffer_auto_out_ar_valid;
  wire [3:0] AXI4Buffer_auto_out_ar_bits_id;
  wire [27:0] AXI4Buffer_auto_out_ar_bits_addr;
  wire  AXI4Buffer_auto_out_ar_bits_user;
  wire  AXI4Buffer_auto_out_r_ready;
  wire  AXI4Buffer_auto_out_r_valid;
  wire [3:0] AXI4Buffer_auto_out_r_bits_id;
  wire [63:0] AXI4Buffer_auto_out_r_bits_data;
  wire [1:0] AXI4Buffer_auto_out_r_bits_resp;
  wire  AXI4Buffer_auto_out_r_bits_user;
  wire  AXI4Fragmenter_clock;
  wire  AXI4Fragmenter_reset;
  wire  AXI4Fragmenter_auto_in_aw_ready;
  wire  AXI4Fragmenter_auto_in_aw_valid;
  wire [3:0] AXI4Fragmenter_auto_in_aw_bits_id;
  wire [27:0] AXI4Fragmenter_auto_in_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_aw_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_aw_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_aw_bits_burst;
  wire  AXI4Fragmenter_auto_in_w_ready;
  wire  AXI4Fragmenter_auto_in_w_valid;
  wire [63:0] AXI4Fragmenter_auto_in_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_in_w_bits_strb;
  wire  AXI4Fragmenter_auto_in_w_bits_last;
  wire  AXI4Fragmenter_auto_in_b_ready;
  wire  AXI4Fragmenter_auto_in_b_valid;
  wire [3:0] AXI4Fragmenter_auto_in_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_in_b_bits_resp;
  wire  AXI4Fragmenter_auto_in_ar_ready;
  wire  AXI4Fragmenter_auto_in_ar_valid;
  wire [3:0] AXI4Fragmenter_auto_in_ar_bits_id;
  wire [27:0] AXI4Fragmenter_auto_in_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_ar_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_ar_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_ar_bits_burst;
  wire  AXI4Fragmenter_auto_in_r_ready;
  wire  AXI4Fragmenter_auto_in_r_valid;
  wire [3:0] AXI4Fragmenter_auto_in_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_in_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_in_r_bits_resp;
  wire  AXI4Fragmenter_auto_in_r_bits_last;
  wire  AXI4Fragmenter_auto_out_aw_ready;
  wire  AXI4Fragmenter_auto_out_aw_valid;
  wire [3:0] AXI4Fragmenter_auto_out_aw_bits_id;
  wire [27:0] AXI4Fragmenter_auto_out_aw_bits_addr;
  wire  AXI4Fragmenter_auto_out_aw_bits_user;
  wire  AXI4Fragmenter_auto_out_w_ready;
  wire  AXI4Fragmenter_auto_out_w_valid;
  wire [63:0] AXI4Fragmenter_auto_out_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_out_w_bits_strb;
  wire  AXI4Fragmenter_auto_out_w_bits_last;
  wire  AXI4Fragmenter_auto_out_b_ready;
  wire  AXI4Fragmenter_auto_out_b_valid;
  wire [3:0] AXI4Fragmenter_auto_out_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_out_b_bits_resp;
  wire  AXI4Fragmenter_auto_out_b_bits_user;
  wire  AXI4Fragmenter_auto_out_ar_ready;
  wire  AXI4Fragmenter_auto_out_ar_valid;
  wire [3:0] AXI4Fragmenter_auto_out_ar_bits_id;
  wire [27:0] AXI4Fragmenter_auto_out_ar_bits_addr;
  wire  AXI4Fragmenter_auto_out_ar_bits_user;
  wire  AXI4Fragmenter_auto_out_r_ready;
  wire  AXI4Fragmenter_auto_out_r_valid;
  wire [3:0] AXI4Fragmenter_auto_out_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_out_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_out_r_bits_resp;
  wire  AXI4Fragmenter_auto_out_r_bits_user;
  wire  AXI4Fragmenter_auto_out_r_bits_last;
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [27:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [27:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  AXI4RAM AXI4RAM (
    .clock(AXI4RAM_clock),
    .reset(AXI4RAM_reset),
    .auto_in_aw_ready(AXI4RAM_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4RAM_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4RAM_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4RAM_auto_in_aw_bits_addr),
    .auto_in_aw_bits_user(AXI4RAM_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4RAM_auto_in_w_ready),
    .auto_in_w_valid(AXI4RAM_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4RAM_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4RAM_auto_in_w_bits_strb),
    .auto_in_b_ready(AXI4RAM_auto_in_b_ready),
    .auto_in_b_valid(AXI4RAM_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4RAM_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4RAM_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4RAM_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4RAM_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4RAM_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4RAM_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4RAM_auto_in_ar_bits_addr),
    .auto_in_ar_bits_user(AXI4RAM_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4RAM_auto_in_r_ready),
    .auto_in_r_valid(AXI4RAM_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4RAM_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4RAM_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4RAM_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4RAM_auto_in_r_bits_user)
  );
  AXI4Buffer_1 AXI4Buffer (
    .clock(AXI4Buffer_clock),
    .reset(AXI4Buffer_reset),
    .auto_in_aw_ready(AXI4Buffer_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Buffer_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Buffer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Buffer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_user(AXI4Buffer_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4Buffer_auto_in_w_ready),
    .auto_in_w_valid(AXI4Buffer_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Buffer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Buffer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Buffer_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Buffer_auto_in_b_ready),
    .auto_in_b_valid(AXI4Buffer_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Buffer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Buffer_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4Buffer_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4Buffer_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Buffer_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Buffer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Buffer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_user(AXI4Buffer_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4Buffer_auto_in_r_ready),
    .auto_in_r_valid(AXI4Buffer_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Buffer_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Buffer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Buffer_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4Buffer_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4Buffer_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Buffer_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Buffer_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Buffer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Buffer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_user(AXI4Buffer_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Buffer_auto_out_w_ready),
    .auto_out_w_valid(AXI4Buffer_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Buffer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Buffer_auto_out_w_bits_strb),
    .auto_out_b_ready(AXI4Buffer_auto_out_b_ready),
    .auto_out_b_valid(AXI4Buffer_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Buffer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Buffer_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Buffer_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Buffer_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Buffer_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Buffer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Buffer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_user(AXI4Buffer_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Buffer_auto_out_r_ready),
    .auto_out_r_valid(AXI4Buffer_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Buffer_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Buffer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Buffer_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Buffer_auto_out_r_bits_user)
  );
  AXI4Fragmenter_1 AXI4Fragmenter (
    .clock(AXI4Fragmenter_clock),
    .reset(AXI4Fragmenter_reset),
    .auto_in_aw_ready(AXI4Fragmenter_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Fragmenter_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Fragmenter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Fragmenter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4Fragmenter_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4Fragmenter_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4Fragmenter_auto_in_aw_bits_burst),
    .auto_in_w_ready(AXI4Fragmenter_auto_in_w_ready),
    .auto_in_w_valid(AXI4Fragmenter_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Fragmenter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Fragmenter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Fragmenter_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Fragmenter_auto_in_b_ready),
    .auto_in_b_valid(AXI4Fragmenter_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Fragmenter_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Fragmenter_auto_in_b_bits_resp),
    .auto_in_ar_ready(AXI4Fragmenter_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Fragmenter_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Fragmenter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Fragmenter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4Fragmenter_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4Fragmenter_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4Fragmenter_auto_in_ar_bits_burst),
    .auto_in_r_ready(AXI4Fragmenter_auto_in_r_ready),
    .auto_in_r_valid(AXI4Fragmenter_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Fragmenter_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Fragmenter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Fragmenter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(AXI4Fragmenter_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Fragmenter_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Fragmenter_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Fragmenter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Fragmenter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_user(AXI4Fragmenter_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Fragmenter_auto_out_w_ready),
    .auto_out_w_valid(AXI4Fragmenter_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Fragmenter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Fragmenter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4Fragmenter_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4Fragmenter_auto_out_b_ready),
    .auto_out_b_valid(AXI4Fragmenter_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Fragmenter_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Fragmenter_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Fragmenter_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Fragmenter_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Fragmenter_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Fragmenter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Fragmenter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_user(AXI4Fragmenter_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Fragmenter_auto_out_r_ready),
    .auto_out_r_valid(AXI4Fragmenter_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Fragmenter_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Fragmenter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Fragmenter_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Fragmenter_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4Fragmenter_auto_out_r_bits_last)
  );
  assign io_axi4_0_aw_ready = _T_31_aw_ready;
  assign io_axi4_0_w_ready = _T_31_w_ready;
  assign io_axi4_0_b_valid = _T_31_b_valid;
  assign io_axi4_0_b_bits_id = _T_31_b_bits_id;
  assign io_axi4_0_b_bits_resp = _T_31_b_bits_resp;
  assign io_axi4_0_ar_ready = _T_31_ar_ready;
  assign io_axi4_0_r_valid = _T_31_r_valid;
  assign io_axi4_0_r_bits_id = _T_31_r_bits_id;
  assign io_axi4_0_r_bits_data = _T_31_r_bits_data;
  assign io_axi4_0_r_bits_resp = _T_31_r_bits_resp;
  assign io_axi4_0_r_bits_last = _T_31_r_bits_last;
  assign AXI4RAM_clock = clock;
  assign AXI4RAM_reset = reset;
  assign AXI4RAM_auto_in_aw_valid = AXI4Buffer_auto_out_aw_valid;
  assign AXI4RAM_auto_in_aw_bits_id = AXI4Buffer_auto_out_aw_bits_id;
  assign AXI4RAM_auto_in_aw_bits_addr = AXI4Buffer_auto_out_aw_bits_addr;
  assign AXI4RAM_auto_in_aw_bits_user = AXI4Buffer_auto_out_aw_bits_user;
  assign AXI4RAM_auto_in_w_valid = AXI4Buffer_auto_out_w_valid;
  assign AXI4RAM_auto_in_w_bits_data = AXI4Buffer_auto_out_w_bits_data;
  assign AXI4RAM_auto_in_w_bits_strb = AXI4Buffer_auto_out_w_bits_strb;
  assign AXI4RAM_auto_in_b_ready = AXI4Buffer_auto_out_b_ready;
  assign AXI4RAM_auto_in_ar_valid = AXI4Buffer_auto_out_ar_valid;
  assign AXI4RAM_auto_in_ar_bits_id = AXI4Buffer_auto_out_ar_bits_id;
  assign AXI4RAM_auto_in_ar_bits_addr = AXI4Buffer_auto_out_ar_bits_addr;
  assign AXI4RAM_auto_in_ar_bits_user = AXI4Buffer_auto_out_ar_bits_user;
  assign AXI4RAM_auto_in_r_ready = AXI4Buffer_auto_out_r_ready;
  assign AXI4Buffer_clock = clock;
  assign AXI4Buffer_reset = reset;
  assign AXI4Buffer_auto_in_aw_valid = AXI4Fragmenter_auto_out_aw_valid;
  assign AXI4Buffer_auto_in_aw_bits_id = AXI4Fragmenter_auto_out_aw_bits_id;
  assign AXI4Buffer_auto_in_aw_bits_addr = AXI4Fragmenter_auto_out_aw_bits_addr;
  assign AXI4Buffer_auto_in_aw_bits_user = AXI4Fragmenter_auto_out_aw_bits_user;
  assign AXI4Buffer_auto_in_w_valid = AXI4Fragmenter_auto_out_w_valid;
  assign AXI4Buffer_auto_in_w_bits_data = AXI4Fragmenter_auto_out_w_bits_data;
  assign AXI4Buffer_auto_in_w_bits_strb = AXI4Fragmenter_auto_out_w_bits_strb;
  assign AXI4Buffer_auto_in_w_bits_last = AXI4Fragmenter_auto_out_w_bits_last;
  assign AXI4Buffer_auto_in_b_ready = AXI4Fragmenter_auto_out_b_ready;
  assign AXI4Buffer_auto_in_ar_valid = AXI4Fragmenter_auto_out_ar_valid;
  assign AXI4Buffer_auto_in_ar_bits_id = AXI4Fragmenter_auto_out_ar_bits_id;
  assign AXI4Buffer_auto_in_ar_bits_addr = AXI4Fragmenter_auto_out_ar_bits_addr;
  assign AXI4Buffer_auto_in_ar_bits_user = AXI4Fragmenter_auto_out_ar_bits_user;
  assign AXI4Buffer_auto_in_r_ready = AXI4Fragmenter_auto_out_r_ready;
  assign AXI4Buffer_auto_out_aw_ready = AXI4RAM_auto_in_aw_ready;
  assign AXI4Buffer_auto_out_w_ready = AXI4RAM_auto_in_w_ready;
  assign AXI4Buffer_auto_out_b_valid = AXI4RAM_auto_in_b_valid;
  assign AXI4Buffer_auto_out_b_bits_id = AXI4RAM_auto_in_b_bits_id;
  assign AXI4Buffer_auto_out_b_bits_resp = AXI4RAM_auto_in_b_bits_resp;
  assign AXI4Buffer_auto_out_b_bits_user = AXI4RAM_auto_in_b_bits_user;
  assign AXI4Buffer_auto_out_ar_ready = AXI4RAM_auto_in_ar_ready;
  assign AXI4Buffer_auto_out_r_valid = AXI4RAM_auto_in_r_valid;
  assign AXI4Buffer_auto_out_r_bits_id = AXI4RAM_auto_in_r_bits_id;
  assign AXI4Buffer_auto_out_r_bits_data = AXI4RAM_auto_in_r_bits_data;
  assign AXI4Buffer_auto_out_r_bits_resp = AXI4RAM_auto_in_r_bits_resp;
  assign AXI4Buffer_auto_out_r_bits_user = AXI4RAM_auto_in_r_bits_user;
  assign AXI4Fragmenter_clock = clock;
  assign AXI4Fragmenter_reset = reset;
  assign AXI4Fragmenter_auto_in_aw_valid = _T_31_aw_valid;
  assign AXI4Fragmenter_auto_in_aw_bits_id = _T_31_aw_bits_id;
  assign AXI4Fragmenter_auto_in_aw_bits_addr = _T_31_aw_bits_addr;
  assign AXI4Fragmenter_auto_in_aw_bits_len = _T_31_aw_bits_len;
  assign AXI4Fragmenter_auto_in_aw_bits_size = _T_31_aw_bits_size;
  assign AXI4Fragmenter_auto_in_aw_bits_burst = _T_31_aw_bits_burst;
  assign AXI4Fragmenter_auto_in_w_valid = _T_31_w_valid;
  assign AXI4Fragmenter_auto_in_w_bits_data = _T_31_w_bits_data;
  assign AXI4Fragmenter_auto_in_w_bits_strb = _T_31_w_bits_strb;
  assign AXI4Fragmenter_auto_in_w_bits_last = _T_31_w_bits_last;
  assign AXI4Fragmenter_auto_in_b_ready = _T_31_b_ready;
  assign AXI4Fragmenter_auto_in_ar_valid = _T_31_ar_valid;
  assign AXI4Fragmenter_auto_in_ar_bits_id = _T_31_ar_bits_id;
  assign AXI4Fragmenter_auto_in_ar_bits_addr = _T_31_ar_bits_addr;
  assign AXI4Fragmenter_auto_in_ar_bits_len = _T_31_ar_bits_len;
  assign AXI4Fragmenter_auto_in_ar_bits_size = _T_31_ar_bits_size;
  assign AXI4Fragmenter_auto_in_ar_bits_burst = _T_31_ar_bits_burst;
  assign AXI4Fragmenter_auto_in_r_ready = _T_31_r_ready;
  assign AXI4Fragmenter_auto_out_aw_ready = AXI4Buffer_auto_in_aw_ready;
  assign AXI4Fragmenter_auto_out_w_ready = AXI4Buffer_auto_in_w_ready;
  assign AXI4Fragmenter_auto_out_b_valid = AXI4Buffer_auto_in_b_valid;
  assign AXI4Fragmenter_auto_out_b_bits_id = AXI4Buffer_auto_in_b_bits_id;
  assign AXI4Fragmenter_auto_out_b_bits_resp = AXI4Buffer_auto_in_b_bits_resp;
  assign AXI4Fragmenter_auto_out_b_bits_user = AXI4Buffer_auto_in_b_bits_user;
  assign AXI4Fragmenter_auto_out_ar_ready = AXI4Buffer_auto_in_ar_ready;
  assign AXI4Fragmenter_auto_out_r_valid = AXI4Buffer_auto_in_r_valid;
  assign AXI4Fragmenter_auto_out_r_bits_id = AXI4Buffer_auto_in_r_bits_id;
  assign AXI4Fragmenter_auto_out_r_bits_data = AXI4Buffer_auto_in_r_bits_data;
  assign AXI4Fragmenter_auto_out_r_bits_resp = AXI4Buffer_auto_in_r_bits_resp;
  assign AXI4Fragmenter_auto_out_r_bits_user = AXI4Buffer_auto_in_r_bits_user;
  assign AXI4Fragmenter_auto_out_r_bits_last = AXI4Buffer_auto_in_r_bits_last;
  assign _T_31_aw_ready = AXI4Fragmenter_auto_in_aw_ready;
  assign _T_31_aw_valid = io_axi4_0_aw_valid;
  assign _T_31_aw_bits_id = io_axi4_0_aw_bits_id;
  assign _T_31_aw_bits_addr = io_axi4_0_aw_bits_addr;
  assign _T_31_aw_bits_len = io_axi4_0_aw_bits_len;
  assign _T_31_aw_bits_size = io_axi4_0_aw_bits_size;
  assign _T_31_aw_bits_burst = io_axi4_0_aw_bits_burst;
  assign _T_31_w_ready = AXI4Fragmenter_auto_in_w_ready;
  assign _T_31_w_valid = io_axi4_0_w_valid;
  assign _T_31_w_bits_data = io_axi4_0_w_bits_data;
  assign _T_31_w_bits_strb = io_axi4_0_w_bits_strb;
  assign _T_31_w_bits_last = io_axi4_0_w_bits_last;
  assign _T_31_b_ready = io_axi4_0_b_ready;
  assign _T_31_b_valid = AXI4Fragmenter_auto_in_b_valid;
  assign _T_31_b_bits_id = AXI4Fragmenter_auto_in_b_bits_id;
  assign _T_31_b_bits_resp = AXI4Fragmenter_auto_in_b_bits_resp;
  assign _T_31_ar_ready = AXI4Fragmenter_auto_in_ar_ready;
  assign _T_31_ar_valid = io_axi4_0_ar_valid;
  assign _T_31_ar_bits_id = io_axi4_0_ar_bits_id;
  assign _T_31_ar_bits_addr = io_axi4_0_ar_bits_addr;
  assign _T_31_ar_bits_len = io_axi4_0_ar_bits_len;
  assign _T_31_ar_bits_size = io_axi4_0_ar_bits_size;
  assign _T_31_ar_bits_burst = io_axi4_0_ar_bits_burst;
  assign _T_31_r_ready = io_axi4_0_r_ready;
  assign _T_31_r_valid = AXI4Fragmenter_auto_in_r_valid;
  assign _T_31_r_bits_id = AXI4Fragmenter_auto_in_r_bits_id;
  assign _T_31_r_bits_data = AXI4Fragmenter_auto_in_r_bits_data;
  assign _T_31_r_bits_resp = AXI4Fragmenter_auto_in_r_bits_resp;
  assign _T_31_r_bits_last = AXI4Fragmenter_auto_in_r_bits_last;
endmodule
module AXI4RAM_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [11:0] auto_in_aw_bits_addr,
  input         auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [11:0] auto_in_ar_bits_addr,
  input         auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_user
);
  wire  in_aw_ready;
  wire  in_aw_valid;
  wire [3:0] in_aw_bits_id;
  wire [11:0] in_aw_bits_addr;
  wire  in_aw_bits_user;
  wire  in_w_ready;
  wire  in_w_valid;
  wire [63:0] in_w_bits_data;
  wire [7:0] in_w_bits_strb;
  wire  in_b_ready;
  wire  in_b_valid;
  wire [3:0] in_b_bits_id;
  wire [1:0] in_b_bits_resp;
  wire  in_b_bits_user;
  wire  in_ar_ready;
  wire  in_ar_valid;
  wire [3:0] in_ar_bits_id;
  wire [11:0] in_ar_bits_addr;
  wire  in_ar_bits_user;
  wire  in_r_ready;
  wire  in_r_valid;
  wire [3:0] in_r_bits_id;
  wire [63:0] in_r_bits_data;
  wire [1:0] in_r_bits_resp;
  wire  in_r_bits_user;
  reg [7:0] mem_0 [0:511];
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_262_data;
  wire [8:0] mem_0__T_262_addr;
  wire [7:0] mem_0__T_217_data;
  wire [8:0] mem_0__T_217_addr;
  wire  mem_0__T_217_mask;
  wire  mem_0__T_217_en;
  wire  _GEN_57;
  reg [8:0] mem_0__T_262_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] mem_1 [0:511];
  reg [31:0] _RAND_2;
  wire [7:0] mem_1__T_262_data;
  wire [8:0] mem_1__T_262_addr;
  wire [7:0] mem_1__T_217_data;
  wire [8:0] mem_1__T_217_addr;
  wire  mem_1__T_217_mask;
  wire  mem_1__T_217_en;
  reg [8:0] mem_1__T_262_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [7:0] mem_2 [0:511];
  reg [31:0] _RAND_4;
  wire [7:0] mem_2__T_262_data;
  wire [8:0] mem_2__T_262_addr;
  wire [7:0] mem_2__T_217_data;
  wire [8:0] mem_2__T_217_addr;
  wire  mem_2__T_217_mask;
  wire  mem_2__T_217_en;
  reg [8:0] mem_2__T_262_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] mem_3 [0:511];
  reg [31:0] _RAND_6;
  wire [7:0] mem_3__T_262_data;
  wire [8:0] mem_3__T_262_addr;
  wire [7:0] mem_3__T_217_data;
  wire [8:0] mem_3__T_217_addr;
  wire  mem_3__T_217_mask;
  wire  mem_3__T_217_en;
  reg [8:0] mem_3__T_262_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [7:0] mem_4 [0:511];
  reg [31:0] _RAND_8;
  wire [7:0] mem_4__T_262_data;
  wire [8:0] mem_4__T_262_addr;
  wire [7:0] mem_4__T_217_data;
  wire [8:0] mem_4__T_217_addr;
  wire  mem_4__T_217_mask;
  wire  mem_4__T_217_en;
  reg [8:0] mem_4__T_262_addr_pipe_0;
  reg [31:0] _RAND_9;
  reg [7:0] mem_5 [0:511];
  reg [31:0] _RAND_10;
  wire [7:0] mem_5__T_262_data;
  wire [8:0] mem_5__T_262_addr;
  wire [7:0] mem_5__T_217_data;
  wire [8:0] mem_5__T_217_addr;
  wire  mem_5__T_217_mask;
  wire  mem_5__T_217_en;
  reg [8:0] mem_5__T_262_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] mem_6 [0:511];
  reg [31:0] _RAND_12;
  wire [7:0] mem_6__T_262_data;
  wire [8:0] mem_6__T_262_addr;
  wire [7:0] mem_6__T_217_data;
  wire [8:0] mem_6__T_217_addr;
  wire  mem_6__T_217_mask;
  wire  mem_6__T_217_en;
  reg [8:0] mem_6__T_262_addr_pipe_0;
  reg [31:0] _RAND_13;
  reg [7:0] mem_7 [0:511];
  reg [31:0] _RAND_14;
  wire [7:0] mem_7__T_262_data;
  wire [8:0] mem_7__T_262_addr;
  wire [7:0] mem_7__T_217_data;
  wire [8:0] mem_7__T_217_addr;
  wire  mem_7__T_217_mask;
  wire  mem_7__T_217_en;
  reg [8:0] mem_7__T_262_addr_pipe_0;
  reg [31:0] _RAND_15;
  wire [8:0] _T_130;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  _T_134;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_138;
  wire  _T_139;
  wire [1:0] _T_140;
  wire [1:0] _T_141;
  wire [3:0] _T_142;
  wire [1:0] _T_143;
  wire [1:0] _T_144;
  wire [2:0] _T_145;
  wire [4:0] _T_146;
  wire [8:0] r_addr;
  wire [8:0] _T_147;
  wire  _T_148;
  wire  _T_149;
  wire  _T_150;
  wire  _T_151;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire  _T_156;
  wire [1:0] _T_157;
  wire [1:0] _T_158;
  wire [3:0] _T_159;
  wire [1:0] _T_160;
  wire [1:0] _T_161;
  wire [2:0] _T_162;
  wire [4:0] _T_163;
  wire [8:0] w_addr;
  wire [12:0] _T_166;
  wire [12:0] _T_168;
  wire [12:0] _T_169;
  wire  r_sel0;
  wire [12:0] _T_173;
  wire [12:0] _T_175;
  wire [12:0] _T_176;
  wire  w_sel0;
  reg  w_full;
  reg [31:0] _RAND_16;
  reg [3:0] w_id;
  reg [31:0] _RAND_17;
  reg  w_user;
  reg [31:0] _RAND_18;
  reg  r_sel1;
  reg [31:0] _RAND_19;
  reg  w_sel1;
  reg [31:0] _RAND_20;
  wire  _T_182;
  wire  _GEN_0;
  wire  _T_184;
  wire  _GEN_1;
  wire [3:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [7:0] _T_187;
  wire [7:0] _T_188;
  wire [7:0] _T_189;
  wire [7:0] _T_190;
  wire [7:0] _T_191;
  wire [7:0] _T_192;
  wire [7:0] _T_193;
  wire [7:0] _T_194;
  wire [7:0] wdata_0;
  wire [7:0] wdata_1;
  wire [7:0] wdata_2;
  wire [7:0] wdata_3;
  wire [7:0] wdata_4;
  wire [7:0] wdata_5;
  wire [7:0] wdata_6;
  wire [7:0] wdata_7;
  wire  _T_208;
  wire  _T_209;
  wire  _T_210;
  wire  _T_211;
  wire  _T_212;
  wire  _T_213;
  wire  _T_214;
  wire  _T_215;
  wire  _T_216;
  wire  _GEN_25;
  wire  _GEN_27;
  wire  _GEN_29;
  wire  _GEN_31;
  wire  _GEN_33;
  wire  _GEN_35;
  wire  _GEN_37;
  wire  _GEN_39;
  wire  _T_238;
  wire  _T_239;
  wire  _T_240;
  wire  _T_244;
  wire [1:0] _T_247;
  reg  r_full;
  reg [31:0] _RAND_21;
  reg [3:0] r_id;
  reg [31:0] _RAND_22;
  reg  r_user;
  reg [31:0] _RAND_23;
  wire  _T_252;
  wire  _GEN_40;
  wire  _T_254;
  wire  _GEN_41;
  wire [3:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  ren;
  wire [8:0] _T_258;
  reg  _T_283;
  reg [31:0] _RAND_24;
  reg [7:0] _T_313_0;
  reg [31:0] _RAND_25;
  reg [7:0] _T_313_1;
  reg [31:0] _RAND_26;
  reg [7:0] _T_313_2;
  reg [31:0] _RAND_27;
  reg [7:0] _T_313_3;
  reg [31:0] _RAND_28;
  reg [7:0] _T_313_4;
  reg [31:0] _RAND_29;
  reg [7:0] _T_313_5;
  reg [31:0] _RAND_30;
  reg [7:0] _T_313_6;
  reg [31:0] _RAND_31;
  reg [7:0] _T_313_7;
  reg [31:0] _RAND_32;
  wire [7:0] _GEN_49;
  wire [7:0] _GEN_50;
  wire [7:0] _GEN_51;
  wire [7:0] _GEN_52;
  wire [7:0] _GEN_53;
  wire [7:0] _GEN_54;
  wire [7:0] _GEN_55;
  wire [7:0] _GEN_56;
  wire  _T_380;
  wire  _T_381;
  wire [1:0] _T_384;
  wire [15:0] _T_385;
  wire [15:0] _T_386;
  wire [31:0] _T_387;
  wire [15:0] _T_388;
  wire [15:0] _T_389;
  wire [31:0] _T_390;
  wire [63:0] _T_391;
  assign mem_0__T_262_addr = mem_0__T_262_addr_pipe_0;
  assign mem_0__T_262_data = mem_0[mem_0__T_262_addr];
  assign mem_0__T_217_data = wdata_0;
  assign mem_0__T_217_addr = w_addr;
  assign mem_0__T_217_mask = _GEN_25;
  assign mem_0__T_217_en = _T_208;
  assign _GEN_57 = ren;
  assign mem_1__T_262_addr = mem_1__T_262_addr_pipe_0;
  assign mem_1__T_262_data = mem_1[mem_1__T_262_addr];
  assign mem_1__T_217_data = wdata_1;
  assign mem_1__T_217_addr = w_addr;
  assign mem_1__T_217_mask = _GEN_27;
  assign mem_1__T_217_en = _T_208;
  assign mem_2__T_262_addr = mem_2__T_262_addr_pipe_0;
  assign mem_2__T_262_data = mem_2[mem_2__T_262_addr];
  assign mem_2__T_217_data = wdata_2;
  assign mem_2__T_217_addr = w_addr;
  assign mem_2__T_217_mask = _GEN_29;
  assign mem_2__T_217_en = _T_208;
  assign mem_3__T_262_addr = mem_3__T_262_addr_pipe_0;
  assign mem_3__T_262_data = mem_3[mem_3__T_262_addr];
  assign mem_3__T_217_data = wdata_3;
  assign mem_3__T_217_addr = w_addr;
  assign mem_3__T_217_mask = _GEN_31;
  assign mem_3__T_217_en = _T_208;
  assign mem_4__T_262_addr = mem_4__T_262_addr_pipe_0;
  assign mem_4__T_262_data = mem_4[mem_4__T_262_addr];
  assign mem_4__T_217_data = wdata_4;
  assign mem_4__T_217_addr = w_addr;
  assign mem_4__T_217_mask = _GEN_33;
  assign mem_4__T_217_en = _T_208;
  assign mem_5__T_262_addr = mem_5__T_262_addr_pipe_0;
  assign mem_5__T_262_data = mem_5[mem_5__T_262_addr];
  assign mem_5__T_217_data = wdata_5;
  assign mem_5__T_217_addr = w_addr;
  assign mem_5__T_217_mask = _GEN_35;
  assign mem_5__T_217_en = _T_208;
  assign mem_6__T_262_addr = mem_6__T_262_addr_pipe_0;
  assign mem_6__T_262_data = mem_6[mem_6__T_262_addr];
  assign mem_6__T_217_data = wdata_6;
  assign mem_6__T_217_addr = w_addr;
  assign mem_6__T_217_mask = _GEN_37;
  assign mem_6__T_217_en = _T_208;
  assign mem_7__T_262_addr = mem_7__T_262_addr_pipe_0;
  assign mem_7__T_262_data = mem_7[mem_7__T_262_addr];
  assign mem_7__T_217_data = wdata_7;
  assign mem_7__T_217_addr = w_addr;
  assign mem_7__T_217_mask = _GEN_39;
  assign mem_7__T_217_en = _T_208;
  assign _T_130 = in_ar_bits_addr[11:3];
  assign _T_131 = _T_130[0];
  assign _T_132 = _T_130[1];
  assign _T_133 = _T_130[2];
  assign _T_134 = _T_130[3];
  assign _T_135 = _T_130[4];
  assign _T_136 = _T_130[5];
  assign _T_137 = _T_130[6];
  assign _T_138 = _T_130[7];
  assign _T_139 = _T_130[8];
  assign _T_140 = {_T_132,_T_131};
  assign _T_141 = {_T_134,_T_133};
  assign _T_142 = {_T_141,_T_140};
  assign _T_143 = {_T_136,_T_135};
  assign _T_144 = {_T_139,_T_138};
  assign _T_145 = {_T_144,_T_137};
  assign _T_146 = {_T_145,_T_143};
  assign r_addr = {_T_146,_T_142};
  assign _T_147 = in_aw_bits_addr[11:3];
  assign _T_148 = _T_147[0];
  assign _T_149 = _T_147[1];
  assign _T_150 = _T_147[2];
  assign _T_151 = _T_147[3];
  assign _T_152 = _T_147[4];
  assign _T_153 = _T_147[5];
  assign _T_154 = _T_147[6];
  assign _T_155 = _T_147[7];
  assign _T_156 = _T_147[8];
  assign _T_157 = {_T_149,_T_148};
  assign _T_158 = {_T_151,_T_150};
  assign _T_159 = {_T_158,_T_157};
  assign _T_160 = {_T_153,_T_152};
  assign _T_161 = {_T_156,_T_155};
  assign _T_162 = {_T_161,_T_154};
  assign _T_163 = {_T_162,_T_160};
  assign w_addr = {_T_163,_T_159};
  assign _T_166 = {1'b0,$signed(in_ar_bits_addr)};
  assign _T_168 = $signed(_T_166) & $signed(-13'sh1000);
  assign _T_169 = $signed(_T_168);
  assign r_sel0 = $signed(_T_169) == $signed(13'sh0);
  assign _T_173 = {1'b0,$signed(in_aw_bits_addr)};
  assign _T_175 = $signed(_T_173) & $signed(-13'sh1000);
  assign _T_176 = $signed(_T_175);
  assign w_sel0 = $signed(_T_176) == $signed(13'sh0);
  assign _T_182 = in_b_ready & in_b_valid;
  assign _GEN_0 = _T_182 ? 1'h0 : w_full;
  assign _T_184 = in_aw_ready & in_aw_valid;
  assign _GEN_1 = _T_184 ? 1'h1 : _GEN_0;
  assign _GEN_2 = _T_184 ? in_aw_bits_id : w_id;
  assign _GEN_3 = _T_184 ? w_sel0 : w_sel1;
  assign _GEN_4 = _T_184 ? in_aw_bits_user : w_user;
  assign _T_187 = in_w_bits_data[7:0];
  assign _T_188 = in_w_bits_data[15:8];
  assign _T_189 = in_w_bits_data[23:16];
  assign _T_190 = in_w_bits_data[31:24];
  assign _T_191 = in_w_bits_data[39:32];
  assign _T_192 = in_w_bits_data[47:40];
  assign _T_193 = in_w_bits_data[55:48];
  assign _T_194 = in_w_bits_data[63:56];
  assign _T_208 = _T_184 & w_sel0;
  assign _T_209 = in_w_bits_strb[0];
  assign _T_210 = in_w_bits_strb[1];
  assign _T_211 = in_w_bits_strb[2];
  assign _T_212 = in_w_bits_strb[3];
  assign _T_213 = in_w_bits_strb[4];
  assign _T_214 = in_w_bits_strb[5];
  assign _T_215 = in_w_bits_strb[6];
  assign _T_216 = in_w_bits_strb[7];
  assign _GEN_25 = _T_208 ? _T_209 : 1'h0;
  assign _GEN_27 = _T_208 ? _T_210 : 1'h0;
  assign _GEN_29 = _T_208 ? _T_211 : 1'h0;
  assign _GEN_31 = _T_208 ? _T_212 : 1'h0;
  assign _GEN_33 = _T_208 ? _T_213 : 1'h0;
  assign _GEN_35 = _T_208 ? _T_214 : 1'h0;
  assign _GEN_37 = _T_208 ? _T_215 : 1'h0;
  assign _GEN_39 = _T_208 ? _T_216 : 1'h0;
  assign _T_238 = w_full == 1'h0;
  assign _T_239 = in_b_ready | _T_238;
  assign _T_240 = in_w_valid & _T_239;
  assign _T_244 = in_aw_valid & _T_239;
  assign _T_247 = w_sel1 ? 2'h0 : 2'h3;
  assign _T_252 = in_r_ready & in_r_valid;
  assign _GEN_40 = _T_252 ? 1'h0 : r_full;
  assign _T_254 = in_ar_ready & in_ar_valid;
  assign _GEN_41 = _T_254 ? 1'h1 : _GEN_40;
  assign _GEN_42 = _T_254 ? in_ar_bits_id : r_id;
  assign _GEN_43 = _T_254 ? r_sel0 : r_sel1;
  assign _GEN_44 = _T_254 ? in_ar_bits_user : r_user;
  assign ren = in_ar_ready & in_ar_valid;
  assign _GEN_49 = _T_283 ? mem_0__T_262_data : _T_313_0;
  assign _GEN_50 = _T_283 ? mem_1__T_262_data : _T_313_1;
  assign _GEN_51 = _T_283 ? mem_2__T_262_data : _T_313_2;
  assign _GEN_52 = _T_283 ? mem_3__T_262_data : _T_313_3;
  assign _GEN_53 = _T_283 ? mem_4__T_262_data : _T_313_4;
  assign _GEN_54 = _T_283 ? mem_5__T_262_data : _T_313_5;
  assign _GEN_55 = _T_283 ? mem_6__T_262_data : _T_313_6;
  assign _GEN_56 = _T_283 ? mem_7__T_262_data : _T_313_7;
  assign _T_380 = r_full == 1'h0;
  assign _T_381 = in_r_ready | _T_380;
  assign _T_384 = r_sel1 ? 2'h0 : 2'h3;
  assign _T_385 = {_GEN_50,_GEN_49};
  assign _T_386 = {_GEN_52,_GEN_51};
  assign _T_387 = {_T_386,_T_385};
  assign _T_388 = {_GEN_54,_GEN_53};
  assign _T_389 = {_GEN_56,_GEN_55};
  assign _T_390 = {_T_389,_T_388};
  assign _T_391 = {_T_390,_T_387};
  assign auto_in_aw_ready = in_aw_ready;
  assign auto_in_w_ready = in_w_ready;
  assign auto_in_b_valid = in_b_valid;
  assign auto_in_b_bits_id = in_b_bits_id;
  assign auto_in_b_bits_resp = in_b_bits_resp;
  assign auto_in_b_bits_user = in_b_bits_user;
  assign auto_in_ar_ready = in_ar_ready;
  assign auto_in_r_valid = in_r_valid;
  assign auto_in_r_bits_id = in_r_bits_id;
  assign auto_in_r_bits_data = in_r_bits_data;
  assign auto_in_r_bits_resp = in_r_bits_resp;
  assign auto_in_r_bits_user = in_r_bits_user;
  assign in_aw_ready = _T_240;
  assign in_aw_valid = auto_in_aw_valid;
  assign in_aw_bits_id = auto_in_aw_bits_id;
  assign in_aw_bits_addr = auto_in_aw_bits_addr;
  assign in_aw_bits_user = auto_in_aw_bits_user;
  assign in_w_ready = _T_244;
  assign in_w_valid = auto_in_w_valid;
  assign in_w_bits_data = auto_in_w_bits_data;
  assign in_w_bits_strb = auto_in_w_bits_strb;
  assign in_b_ready = auto_in_b_ready;
  assign in_b_valid = w_full;
  assign in_b_bits_id = w_id;
  assign in_b_bits_resp = _T_247;
  assign in_b_bits_user = w_user;
  assign in_ar_ready = _T_381;
  assign in_ar_valid = auto_in_ar_valid;
  assign in_ar_bits_id = auto_in_ar_bits_id;
  assign in_ar_bits_addr = auto_in_ar_bits_addr;
  assign in_ar_bits_user = auto_in_ar_bits_user;
  assign in_r_ready = auto_in_r_ready;
  assign in_r_valid = r_full;
  assign in_r_bits_id = r_id;
  assign in_r_bits_data = _T_391;
  assign in_r_bits_resp = _T_384;
  assign in_r_bits_user = r_user;
  assign wdata_0 = _T_187;
  assign wdata_1 = _T_188;
  assign wdata_2 = _T_189;
  assign wdata_3 = _T_190;
  assign wdata_4 = _T_191;
  assign wdata_5 = _T_192;
  assign wdata_6 = _T_193;
  assign wdata_7 = _T_194;
  assign _T_258 = r_addr;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0__T_262_addr_pipe_0 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_1[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_1__T_262_addr_pipe_0 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_2[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_2__T_262_addr_pipe_0 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_3[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_3__T_262_addr_pipe_0 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_4[initvar] = _RAND_8[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_4__T_262_addr_pipe_0 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_5[initvar] = _RAND_10[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_5__T_262_addr_pipe_0 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_6[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_6__T_262_addr_pipe_0 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_7[initvar] = _RAND_14[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_7__T_262_addr_pipe_0 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  w_full = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  w_id = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  w_user = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  r_sel1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  w_sel1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  r_full = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  r_id = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  r_user = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_283 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_313_0 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_313_1 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_313_2 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_313_3 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_313_4 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_313_5 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_313_6 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_313_7 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_217_en & mem_0__T_217_mask) begin
      mem_0[mem_0__T_217_addr] <= mem_0__T_217_data;
    end
    if (_GEN_57) begin
      mem_0__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_1__T_217_en & mem_1__T_217_mask) begin
      mem_1[mem_1__T_217_addr] <= mem_1__T_217_data;
    end
    if (_GEN_57) begin
      mem_1__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_2__T_217_en & mem_2__T_217_mask) begin
      mem_2[mem_2__T_217_addr] <= mem_2__T_217_data;
    end
    if (_GEN_57) begin
      mem_2__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_3__T_217_en & mem_3__T_217_mask) begin
      mem_3[mem_3__T_217_addr] <= mem_3__T_217_data;
    end
    if (_GEN_57) begin
      mem_3__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_4__T_217_en & mem_4__T_217_mask) begin
      mem_4[mem_4__T_217_addr] <= mem_4__T_217_data;
    end
    if (_GEN_57) begin
      mem_4__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_5__T_217_en & mem_5__T_217_mask) begin
      mem_5[mem_5__T_217_addr] <= mem_5__T_217_data;
    end
    if (_GEN_57) begin
      mem_5__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_6__T_217_en & mem_6__T_217_mask) begin
      mem_6[mem_6__T_217_addr] <= mem_6__T_217_data;
    end
    if (_GEN_57) begin
      mem_6__T_262_addr_pipe_0 <= _T_258;
    end
    if(mem_7__T_217_en & mem_7__T_217_mask) begin
      mem_7[mem_7__T_217_addr] <= mem_7__T_217_data;
    end
    if (_GEN_57) begin
      mem_7__T_262_addr_pipe_0 <= _T_258;
    end
    if (reset) begin
      w_full <= 1'h0;
    end else begin
      if (_T_184) begin
        w_full <= 1'h1;
      end else begin
        if (_T_182) begin
          w_full <= 1'h0;
        end
      end
    end
    if (_T_184) begin
      w_id <= in_aw_bits_id;
    end
    if (_T_184) begin
      w_user <= in_aw_bits_user;
    end
    if (_T_254) begin
      r_sel1 <= r_sel0;
    end
    if (_T_184) begin
      w_sel1 <= w_sel0;
    end
    if (reset) begin
      r_full <= 1'h0;
    end else begin
      if (_T_254) begin
        r_full <= 1'h1;
      end else begin
        if (_T_252) begin
          r_full <= 1'h0;
        end
      end
    end
    if (_T_254) begin
      r_id <= in_ar_bits_id;
    end
    if (_T_254) begin
      r_user <= in_ar_bits_user;
    end
    _T_283 <= _T_254;
    if (_T_283) begin
      _T_313_0 <= mem_0__T_262_data;
    end
    if (_T_283) begin
      _T_313_1 <= mem_1__T_262_data;
    end
    if (_T_283) begin
      _T_313_2 <= mem_2__T_262_data;
    end
    if (_T_283) begin
      _T_313_3 <= mem_3__T_262_data;
    end
    if (_T_283) begin
      _T_313_4 <= mem_4__T_262_data;
    end
    if (_T_283) begin
      _T_313_5 <= mem_5__T_262_data;
    end
    if (_T_283) begin
      _T_313_6 <= mem_6__T_262_data;
    end
    if (_T_283) begin
      _T_313_7 <= mem_7__T_262_data;
    end
  end
endmodule
module Queue_123(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [11:0] io_enq_bits_addr,
  input         io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [11:0] io_deq_bits_addr,
  output        io_deq_bits_user
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_50_data;
  wire  ram_id__T_50_addr;
  wire [3:0] ram_id__T_36_data;
  wire  ram_id__T_36_addr;
  wire  ram_id__T_36_mask;
  wire  ram_id__T_36_en;
  reg [11:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [11:0] ram_addr__T_50_data;
  wire  ram_addr__T_50_addr;
  wire [11:0] ram_addr__T_36_data;
  wire  ram_addr__T_36_addr;
  wire  ram_addr__T_36_mask;
  wire  ram_addr__T_36_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_2;
  wire  ram_user__T_50_data;
  wire  ram_user__T_50_addr;
  wire  ram_user__T_36_data;
  wire  ram_user__T_36_addr;
  wire  ram_user__T_36_mask;
  wire  ram_user__T_36_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_28;
  wire  _T_30;
  wire  empty;
  wire  _T_31;
  wire  _T_32;
  wire  do_enq;
  wire  _T_34;
  wire  do_deq;
  wire [1:0] _T_39;
  wire  _T_40;
  wire  _GEN_13;
  wire [1:0] _T_43;
  wire  _T_44;
  wire  _GEN_14;
  wire  _T_45;
  wire  _GEN_15;
  wire  _T_47;
  wire  _T_49;
  assign ram_id__T_50_addr = value_1;
  assign ram_id__T_50_data = ram_id[ram_id__T_50_addr];
  assign ram_id__T_36_data = io_enq_bits_id;
  assign ram_id__T_36_addr = value;
  assign ram_id__T_36_mask = do_enq;
  assign ram_id__T_36_en = do_enq;
  assign ram_addr__T_50_addr = value_1;
  assign ram_addr__T_50_data = ram_addr[ram_addr__T_50_addr];
  assign ram_addr__T_36_data = io_enq_bits_addr;
  assign ram_addr__T_36_addr = value;
  assign ram_addr__T_36_mask = do_enq;
  assign ram_addr__T_36_en = do_enq;
  assign ram_user__T_50_addr = value_1;
  assign ram_user__T_50_data = ram_user[ram_user__T_50_addr];
  assign ram_user__T_36_data = io_enq_bits_user;
  assign ram_user__T_36_addr = value;
  assign ram_user__T_36_mask = do_enq;
  assign ram_user__T_36_en = do_enq;
  assign _T_28 = value == value_1;
  assign _T_30 = maybe_full == 1'h0;
  assign empty = _T_28 & _T_30;
  assign _T_31 = _T_28 & maybe_full;
  assign _T_32 = io_enq_ready & io_enq_valid;
  assign _T_34 = io_deq_ready & io_deq_valid;
  assign _T_39 = value + 1'h1;
  assign _T_40 = _T_39[0:0];
  assign _GEN_13 = do_enq ? _T_40 : value;
  assign _T_43 = value_1 + 1'h1;
  assign _T_44 = _T_43[0:0];
  assign _GEN_14 = do_deq ? _T_44 : value_1;
  assign _T_45 = do_enq != do_deq;
  assign _GEN_15 = _T_45 ? do_enq : maybe_full;
  assign _T_47 = empty == 1'h0;
  assign _T_49 = _T_31 == 1'h0;
  assign io_enq_ready = _T_49;
  assign io_deq_valid = _T_47;
  assign io_deq_bits_id = ram_id__T_50_data;
  assign io_deq_bits_addr = ram_addr__T_50_data;
  assign io_deq_bits_user = ram_user__T_50_data;
  assign do_enq = _T_32;
  assign do_deq = _T_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_36_en & ram_id__T_36_mask) begin
      ram_id[ram_id__T_36_addr] <= ram_id__T_36_data;
    end
    if(ram_addr__T_36_en & ram_addr__T_36_mask) begin
      ram_addr[ram_addr__T_36_addr] <= ram_addr__T_36_data;
    end
    if(ram_user__T_36_en & ram_user__T_36_mask) begin
      ram_user[ram_user__T_36_addr] <= ram_user__T_36_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (do_enq) begin
        value <= _T_40;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_44;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_45) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Buffer_2(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [11:0] auto_in_aw_bits_addr,
  input         auto_in_aw_bits_user,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_b_bits_user,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [11:0] auto_in_ar_bits_addr,
  input         auto_in_ar_bits_user,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_user,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [11:0] auto_out_aw_bits_addr,
  output        auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [11:0] auto_out_ar_bits_addr,
  output        auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_user
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [11:0] _T_31_aw_bits_addr;
  wire  _T_31_aw_bits_user;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_b_bits_user;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [11:0] _T_31_ar_bits_addr;
  wire  _T_31_ar_bits_user;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_user;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [11:0] _T_89_aw_bits_addr;
  wire  _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [11:0] _T_89_ar_bits_addr;
  wire  _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_user;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [11:0] Queue_io_enq_bits_addr;
  wire  Queue_io_enq_bits_user;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [11:0] Queue_io_deq_bits_addr;
  wire  Queue_io_deq_bits_user;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [11:0] _T_207_bits_addr;
  wire  _T_207_bits_user;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_215_ready;
  wire  _T_215_valid;
  wire [63:0] _T_215_bits_data;
  wire [7:0] _T_215_bits_strb;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_enq_bits_user;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  Queue_2_io_deq_bits_user;
  wire  _T_223_ready;
  wire  _T_223_valid;
  wire [3:0] _T_223_bits_id;
  wire [1:0] _T_223_bits_resp;
  wire  _T_223_bits_user;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [11:0] Queue_3_io_enq_bits_addr;
  wire  Queue_3_io_enq_bits_user;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [11:0] Queue_3_io_deq_bits_addr;
  wire  Queue_3_io_deq_bits_user;
  wire  _T_231_ready;
  wire  _T_231_valid;
  wire [3:0] _T_231_bits_id;
  wire [11:0] _T_231_bits_addr;
  wire  _T_231_bits_user;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_user;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_user;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_239_ready;
  wire  _T_239_valid;
  wire [3:0] _T_239_bits_id;
  wire [63:0] _T_239_bits_data;
  wire [1:0] _T_239_bits_resp;
  wire  _T_239_bits_user;
  wire  _T_239_bits_last;
  Queue_123 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  Queue_67 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_117 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user)
  );
  Queue_123 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_user(Queue_3_io_deq_bits_user)
  );
  Queue_119 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_user(Queue_4_io_enq_bits_user),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_user(Queue_4_io_deq_bits_user),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_b_bits_user = _T_31_b_bits_user;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_user = _T_31_r_bits_user;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_user = auto_in_aw_bits_user;
  assign _T_31_w_ready = Queue_1_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_223_valid;
  assign _T_31_b_bits_id = _T_223_bits_id;
  assign _T_31_b_bits_resp = _T_223_bits_resp;
  assign _T_31_b_bits_user = _T_223_bits_user;
  assign _T_31_ar_ready = Queue_3_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_user = auto_in_ar_bits_user;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_239_valid;
  assign _T_31_r_bits_id = _T_239_bits_id;
  assign _T_31_r_bits_data = _T_239_bits_data;
  assign _T_31_r_bits_resp = _T_239_bits_resp;
  assign _T_31_r_bits_user = _T_239_bits_user;
  assign _T_31_r_bits_last = _T_239_bits_last;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_207_valid;
  assign _T_89_aw_bits_id = _T_207_bits_id;
  assign _T_89_aw_bits_addr = _T_207_bits_addr;
  assign _T_89_aw_bits_user = _T_207_bits_user;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_215_valid;
  assign _T_89_w_bits_data = _T_215_bits_data;
  assign _T_89_w_bits_strb = _T_215_bits_strb;
  assign _T_89_b_ready = Queue_2_io_enq_ready;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_231_valid;
  assign _T_89_ar_bits_id = _T_231_bits_id;
  assign _T_89_ar_bits_addr = _T_231_bits_addr;
  assign _T_89_ar_bits_user = _T_231_bits_user;
  assign _T_89_r_ready = Queue_4_io_enq_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign Queue_io_enq_valid = _T_31_aw_valid;
  assign Queue_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_io_enq_bits_user = _T_31_aw_bits_user;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_89_aw_ready;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_user = Queue_io_deq_bits_user;
  assign Queue_1_io_enq_valid = _T_31_w_valid;
  assign Queue_1_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_1_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_1_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_1_io_deq_ready = _T_215_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_215_ready = _T_89_w_ready;
  assign _T_215_valid = Queue_1_io_deq_valid;
  assign _T_215_bits_data = Queue_1_io_deq_bits_data;
  assign _T_215_bits_strb = Queue_1_io_deq_bits_strb;
  assign Queue_2_io_enq_valid = _T_89_b_valid;
  assign Queue_2_io_enq_bits_id = _T_89_b_bits_id;
  assign Queue_2_io_enq_bits_resp = _T_89_b_bits_resp;
  assign Queue_2_io_enq_bits_user = _T_89_b_bits_user;
  assign Queue_2_io_deq_ready = _T_223_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_223_ready = _T_31_b_ready;
  assign _T_223_valid = Queue_2_io_deq_valid;
  assign _T_223_bits_id = Queue_2_io_deq_bits_id;
  assign _T_223_bits_resp = Queue_2_io_deq_bits_resp;
  assign _T_223_bits_user = Queue_2_io_deq_bits_user;
  assign Queue_3_io_enq_valid = _T_31_ar_valid;
  assign Queue_3_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_3_io_enq_bits_user = _T_31_ar_bits_user;
  assign Queue_3_io_deq_ready = _T_231_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign _T_231_ready = _T_89_ar_ready;
  assign _T_231_valid = Queue_3_io_deq_valid;
  assign _T_231_bits_id = Queue_3_io_deq_bits_id;
  assign _T_231_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_231_bits_user = Queue_3_io_deq_bits_user;
  assign Queue_4_io_enq_valid = _T_89_r_valid;
  assign Queue_4_io_enq_bits_id = _T_89_r_bits_id;
  assign Queue_4_io_enq_bits_data = _T_89_r_bits_data;
  assign Queue_4_io_enq_bits_resp = _T_89_r_bits_resp;
  assign Queue_4_io_enq_bits_user = _T_89_r_bits_user;
  assign Queue_4_io_deq_ready = _T_239_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign _T_239_ready = _T_31_r_ready;
  assign _T_239_valid = Queue_4_io_deq_valid;
  assign _T_239_bits_id = Queue_4_io_deq_bits_id;
  assign _T_239_bits_data = Queue_4_io_deq_bits_data;
  assign _T_239_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_239_bits_user = Queue_4_io_deq_bits_user;
  assign _T_239_bits_last = Queue_4_io_deq_bits_last;
endmodule
module Queue_128(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [11:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [11:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst
);
  reg [3:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_42_data;
  wire  ram_id__T_42_addr;
  wire [3:0] ram_id__T_33_data;
  wire  ram_id__T_33_addr;
  wire  ram_id__T_33_mask;
  wire  ram_id__T_33_en;
  reg [11:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [11:0] ram_addr__T_42_data;
  wire  ram_addr__T_42_addr;
  wire [11:0] ram_addr__T_33_data;
  wire  ram_addr__T_33_addr;
  wire  ram_addr__T_33_mask;
  wire  ram_addr__T_33_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_42_data;
  wire  ram_len__T_42_addr;
  wire [7:0] ram_len__T_33_data;
  wire  ram_len__T_33_addr;
  wire  ram_len__T_33_mask;
  wire  ram_len__T_33_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_42_data;
  wire  ram_size__T_42_addr;
  wire [2:0] ram_size__T_33_data;
  wire  ram_size__T_33_addr;
  wire  ram_size__T_33_mask;
  wire  ram_size__T_33_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_42_data;
  wire  ram_burst__T_42_addr;
  wire [1:0] ram_burst__T_33_data;
  wire  ram_burst__T_33_addr;
  wire  ram_burst__T_33_mask;
  wire  ram_burst__T_33_en;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  empty;
  wire  _T_28;
  wire  do_enq;
  wire  _T_30;
  wire  do_deq;
  wire  _T_36;
  wire  _GEN_12;
  wire  _T_38;
  wire  _GEN_13;
  wire  _GEN_14;
  wire [1:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [7:0] _GEN_21;
  wire [11:0] _GEN_22;
  wire [3:0] _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  assign ram_id__T_42_addr = 1'h0;
  assign ram_id__T_42_data = ram_id[ram_id__T_42_addr];
  assign ram_id__T_33_data = io_enq_bits_id;
  assign ram_id__T_33_addr = 1'h0;
  assign ram_id__T_33_mask = do_enq;
  assign ram_id__T_33_en = do_enq;
  assign ram_addr__T_42_addr = 1'h0;
  assign ram_addr__T_42_data = ram_addr[ram_addr__T_42_addr];
  assign ram_addr__T_33_data = io_enq_bits_addr;
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_mask = do_enq;
  assign ram_addr__T_33_en = do_enq;
  assign ram_len__T_42_addr = 1'h0;
  assign ram_len__T_42_data = ram_len[ram_len__T_42_addr];
  assign ram_len__T_33_data = io_enq_bits_len;
  assign ram_len__T_33_addr = 1'h0;
  assign ram_len__T_33_mask = do_enq;
  assign ram_len__T_33_en = do_enq;
  assign ram_size__T_42_addr = 1'h0;
  assign ram_size__T_42_data = ram_size[ram_size__T_42_addr];
  assign ram_size__T_33_data = io_enq_bits_size;
  assign ram_size__T_33_addr = 1'h0;
  assign ram_size__T_33_mask = do_enq;
  assign ram_size__T_33_en = do_enq;
  assign ram_burst__T_42_addr = 1'h0;
  assign ram_burst__T_42_data = ram_burst[ram_burst__T_42_addr];
  assign ram_burst__T_33_data = io_enq_bits_burst;
  assign ram_burst__T_33_addr = 1'h0;
  assign ram_burst__T_33_mask = do_enq;
  assign ram_burst__T_33_en = do_enq;
  assign empty = maybe_full == 1'h0;
  assign _T_28 = io_enq_ready & io_enq_valid;
  assign _T_30 = io_deq_ready & io_deq_valid;
  assign _T_36 = do_enq != do_deq;
  assign _GEN_12 = _T_36 ? do_enq : maybe_full;
  assign _T_38 = empty == 1'h0;
  assign _GEN_13 = io_enq_valid ? 1'h1 : _T_38;
  assign _GEN_14 = io_deq_ready ? 1'h0 : _T_28;
  assign _GEN_19 = empty ? io_enq_bits_burst : ram_burst__T_42_data;
  assign _GEN_20 = empty ? io_enq_bits_size : ram_size__T_42_data;
  assign _GEN_21 = empty ? io_enq_bits_len : ram_len__T_42_data;
  assign _GEN_22 = empty ? io_enq_bits_addr : ram_addr__T_42_data;
  assign _GEN_23 = empty ? io_enq_bits_id : ram_id__T_42_data;
  assign _GEN_24 = empty ? 1'h0 : _T_30;
  assign _GEN_25 = empty ? _GEN_14 : _T_28;
  assign io_enq_ready = empty;
  assign io_deq_valid = _GEN_13;
  assign io_deq_bits_id = _GEN_23;
  assign io_deq_bits_addr = _GEN_22;
  assign io_deq_bits_len = _GEN_21;
  assign io_deq_bits_size = _GEN_20;
  assign io_deq_bits_burst = _GEN_19;
  assign do_enq = _GEN_25;
  assign do_deq = _GEN_24;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_33_en & ram_id__T_33_mask) begin
      ram_id[ram_id__T_33_addr] <= ram_id__T_33_data;
    end
    if(ram_addr__T_33_en & ram_addr__T_33_mask) begin
      ram_addr[ram_addr__T_33_addr] <= ram_addr__T_33_data;
    end
    if(ram_len__T_33_en & ram_len__T_33_mask) begin
      ram_len[ram_len__T_33_addr] <= ram_len__T_33_data;
    end
    if(ram_size__T_33_en & ram_size__T_33_mask) begin
      ram_size[ram_size__T_33_addr] <= ram_size__T_33_data;
    end
    if(ram_burst__T_33_en & ram_burst__T_33_mask) begin
      ram_burst[ram_burst__T_33_addr] <= ram_burst__T_33_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_36) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module AXI4Fragmenter_2(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [11:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [11:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [11:0] auto_out_aw_bits_addr,
  output        auto_out_aw_bits_user,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_b_bits_user,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [11:0] auto_out_ar_bits_addr,
  output        auto_out_ar_bits_user,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_user,
  input         auto_out_r_bits_last
);
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [11:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [11:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  wire  _T_89_aw_ready;
  wire  _T_89_aw_valid;
  wire [3:0] _T_89_aw_bits_id;
  wire [11:0] _T_89_aw_bits_addr;
  wire  _T_89_aw_bits_user;
  wire  _T_89_w_ready;
  wire  _T_89_w_valid;
  wire [63:0] _T_89_w_bits_data;
  wire [7:0] _T_89_w_bits_strb;
  wire  _T_89_w_bits_last;
  wire  _T_89_b_ready;
  wire  _T_89_b_valid;
  wire [3:0] _T_89_b_bits_id;
  wire [1:0] _T_89_b_bits_resp;
  wire  _T_89_b_bits_user;
  wire  _T_89_ar_ready;
  wire  _T_89_ar_valid;
  wire [3:0] _T_89_ar_bits_id;
  wire [11:0] _T_89_ar_bits_addr;
  wire  _T_89_ar_bits_user;
  wire  _T_89_r_ready;
  wire  _T_89_r_valid;
  wire [3:0] _T_89_r_bits_id;
  wire [63:0] _T_89_r_bits_data;
  wire [1:0] _T_89_r_bits_resp;
  wire  _T_89_r_bits_user;
  wire  _T_89_r_bits_last;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [11:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [11:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  _T_207_ready;
  wire  _T_207_valid;
  wire [3:0] _T_207_bits_id;
  wire [11:0] _T_207_bits_addr;
  wire [7:0] _T_207_bits_len;
  wire [2:0] _T_207_bits_size;
  wire [1:0] _T_207_bits_burst;
  wire  _T_211_ready;
  wire  _T_211_valid;
  wire [3:0] _T_211_bits_id;
  wire [11:0] _T_211_bits_addr;
  reg  _T_217;
  reg [31:0] _RAND_0;
  reg [11:0] _T_219;
  reg [31:0] _RAND_1;
  reg [7:0] _T_221;
  reg [31:0] _RAND_2;
  wire [7:0] _T_222;
  wire [11:0] _T_223;
  wire  _T_271;
  wire [8:0] _T_277;
  wire [8:0] _T_279;
  wire [15:0] _GEN_54;
  wire [15:0] _T_284;
  wire [15:0] _GEN_55;
  wire [16:0] _T_285;
  wire [15:0] _T_286;
  wire [15:0] _T_288;
  wire [22:0] _GEN_56;
  wire [22:0] _T_289;
  wire [14:0] _T_290;
  wire [15:0] _T_292;
  wire  _T_294;
  wire [15:0] _GEN_57;
  wire [15:0] _T_295;
  wire [11:0] _T_296;
  wire [14:0] _GEN_58;
  wire [14:0] _T_297;
  wire [14:0] _T_298;
  wire [15:0] _GEN_59;
  wire [15:0] _T_299;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire  _T_302;
  wire  _T_303;
  wire [11:0] _T_304;
  wire [9:0] _T_307;
  wire [2:0] _T_308;
  wire [2:0] _T_309;
  wire [11:0] _GEN_60;
  wire [11:0] _T_310;
  wire [11:0] _T_311;
  wire  _T_312;
  wire  _T_314;
  wire [8:0] _GEN_61;
  wire [9:0] _T_315;
  wire [9:0] _T_316;
  wire [8:0] _T_317;
  wire  _GEN_3;
  wire [15:0] _GEN_4;
  wire [8:0] _GEN_5;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_id;
  wire [11:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_id;
  wire [11:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire  _T_322_ready;
  wire  _T_322_valid;
  wire [3:0] _T_322_bits_id;
  wire [11:0] _T_322_bits_addr;
  wire [7:0] _T_322_bits_len;
  wire [2:0] _T_322_bits_size;
  wire [1:0] _T_322_bits_burst;
  wire  _T_326_ready;
  wire  _T_326_valid;
  wire [3:0] _T_326_bits_id;
  wire [11:0] _T_326_bits_addr;
  reg  _T_332;
  reg [31:0] _RAND_3;
  reg [11:0] _T_334;
  reg [31:0] _RAND_4;
  reg [7:0] _T_336;
  reg [31:0] _RAND_5;
  wire [7:0] _T_337;
  wire [11:0] _T_338;
  wire  _T_386;
  wire [15:0] _T_399;
  wire [15:0] _GEN_73;
  wire [16:0] _T_400;
  wire [15:0] _T_401;
  wire [15:0] _T_403;
  wire [22:0] _GEN_74;
  wire [22:0] _T_404;
  wire [14:0] _T_405;
  wire [15:0] _T_407;
  wire  _T_409;
  wire [15:0] _GEN_75;
  wire [15:0] _T_410;
  wire [11:0] _T_411;
  wire [14:0] _GEN_76;
  wire [14:0] _T_412;
  wire [14:0] _T_413;
  wire [15:0] _GEN_77;
  wire [15:0] _T_414;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire  _T_417;
  wire  _T_418;
  wire [11:0] _T_419;
  wire [9:0] _T_422;
  wire [2:0] _T_423;
  wire [2:0] _T_424;
  wire [11:0] _GEN_78;
  wire [11:0] _T_425;
  wire [11:0] _T_426;
  wire  _T_427;
  wire  _T_429;
  wire [8:0] _GEN_79;
  wire [9:0] _T_430;
  wire [9:0] _T_431;
  wire [8:0] _T_432;
  wire  _GEN_8;
  wire [15:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [7:0] Queue_2_io_enq_bits_strb;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [7:0] Queue_2_io_deq_bits_strb;
  wire  Queue_2_io_deq_bits_last;
  wire  _T_437_ready;
  wire  _T_437_valid;
  wire [63:0] _T_437_bits_data;
  wire [7:0] _T_437_bits_strb;
  wire  _T_437_bits_last;
  reg  _T_443;
  reg [31:0] _RAND_6;
  wire  _T_445;
  wire  _T_447;
  wire  _T_448;
  wire  _GEN_11;
  wire  _T_450;
  wire  _GEN_12;
  wire  _T_452;
  wire  _T_453;
  wire  _T_455;
  wire  _T_457;
  wire  _T_458;
  reg [8:0] _T_461;
  reg [31:0] _RAND_7;
  wire  _T_463;
  wire [8:0] _T_465;
  wire [8:0] _T_466;
  wire  _T_468;
  wire  _T_469;
  wire [8:0] _GEN_80;
  wire [9:0] _T_470;
  wire [9:0] _T_471;
  wire [8:0] _T_472;
  wire  _T_475;
  wire  _T_477;
  wire  _T_478;
  wire  _T_480;
  wire  _T_482;
  wire  _T_484;
  wire  _T_485;
  wire  _T_486;
  wire  _T_490;
  wire  _T_492;
  wire  _T_494;
  wire  _T_495;
  wire  _T_496;
  wire  _T_498;
  wire  _T_500;
  wire  _T_502;
  wire  _T_504;
  wire  _T_506;
  wire  _T_507;
  reg [1:0] _T_581_0;
  reg [31:0] _RAND_8;
  reg [1:0] _T_581_1;
  reg [31:0] _RAND_9;
  reg [1:0] _T_581_2;
  reg [31:0] _RAND_10;
  reg [1:0] _T_581_3;
  reg [31:0] _RAND_11;
  reg [1:0] _T_581_4;
  reg [31:0] _RAND_12;
  reg [1:0] _T_581_5;
  reg [31:0] _RAND_13;
  reg [1:0] _T_581_6;
  reg [31:0] _RAND_14;
  reg [1:0] _T_581_7;
  reg [31:0] _RAND_15;
  reg [1:0] _T_581_8;
  reg [31:0] _RAND_16;
  reg [1:0] _T_581_9;
  reg [31:0] _RAND_17;
  reg [1:0] _T_581_10;
  reg [31:0] _RAND_18;
  reg [1:0] _T_581_11;
  reg [31:0] _RAND_19;
  reg [1:0] _T_581_12;
  reg [31:0] _RAND_20;
  reg [1:0] _T_581_13;
  reg [31:0] _RAND_21;
  reg [1:0] _T_581_14;
  reg [31:0] _RAND_22;
  reg [1:0] _T_581_15;
  reg [31:0] _RAND_23;
  wire [1:0] _GEN_0;
  wire [1:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire [1:0] _GEN_17;
  wire [1:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [1:0] _GEN_22;
  wire [1:0] _GEN_23;
  wire [1:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [1:0] _GEN_26;
  wire [1:0] _GEN_27;
  wire [1:0] _T_637;
  wire [15:0] _T_640;
  wire  _T_642;
  wire  _T_643;
  wire  _T_644;
  wire  _T_645;
  wire  _T_646;
  wire  _T_647;
  wire  _T_648;
  wire  _T_649;
  wire  _T_650;
  wire  _T_651;
  wire  _T_652;
  wire  _T_653;
  wire  _T_654;
  wire  _T_655;
  wire  _T_656;
  wire  _T_657;
  wire  _T_658;
  wire  _T_659;
  wire [1:0] _T_661;
  wire [1:0] _T_662;
  wire [1:0] _GEN_28;
  wire  _T_664;
  wire [1:0] _T_666;
  wire [1:0] _T_667;
  wire [1:0] _GEN_29;
  wire  _T_669;
  wire [1:0] _T_671;
  wire [1:0] _T_672;
  wire [1:0] _GEN_30;
  wire  _T_674;
  wire [1:0] _T_676;
  wire [1:0] _T_677;
  wire [1:0] _GEN_31;
  wire  _T_679;
  wire [1:0] _T_681;
  wire [1:0] _T_682;
  wire [1:0] _GEN_32;
  wire  _T_684;
  wire [1:0] _T_686;
  wire [1:0] _T_687;
  wire [1:0] _GEN_33;
  wire  _T_689;
  wire [1:0] _T_691;
  wire [1:0] _T_692;
  wire [1:0] _GEN_34;
  wire  _T_694;
  wire [1:0] _T_696;
  wire [1:0] _T_697;
  wire [1:0] _GEN_35;
  wire  _T_699;
  wire [1:0] _T_701;
  wire [1:0] _T_702;
  wire [1:0] _GEN_36;
  wire  _T_704;
  wire [1:0] _T_706;
  wire [1:0] _T_707;
  wire [1:0] _GEN_37;
  wire  _T_709;
  wire [1:0] _T_711;
  wire [1:0] _T_712;
  wire [1:0] _GEN_38;
  wire  _T_714;
  wire [1:0] _T_716;
  wire [1:0] _T_717;
  wire [1:0] _GEN_39;
  wire  _T_719;
  wire [1:0] _T_721;
  wire [1:0] _T_722;
  wire [1:0] _GEN_40;
  wire  _T_724;
  wire [1:0] _T_726;
  wire [1:0] _T_727;
  wire [1:0] _GEN_41;
  wire  _T_729;
  wire [1:0] _T_731;
  wire [1:0] _T_732;
  wire [1:0] _GEN_42;
  wire  _T_734;
  wire [1:0] _T_736;
  wire [1:0] _T_737;
  wire [1:0] _GEN_43;
  Queue_128 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst)
  );
  Queue_128 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst)
  );
  Queue_32 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign _T_222 = _T_217 ? _T_221 : _T_207_bits_len;
  assign _T_223 = _T_217 ? _T_219 : _T_207_bits_addr;
  assign _T_271 = _T_207_bits_burst == 2'h0;
  assign _T_277 = 9'h0 << 1;
  assign _T_279 = _T_277 | 9'h1;
  assign _GEN_54 = {{7'd0}, _T_279};
  assign _T_284 = _GEN_54 << _T_207_bits_size;
  assign _GEN_55 = {{4'd0}, _T_223};
  assign _T_285 = _GEN_55 + _T_284;
  assign _T_286 = _T_285[15:0];
  assign _T_288 = {_T_207_bits_len,8'hff};
  assign _GEN_56 = {{7'd0}, _T_288};
  assign _T_289 = _GEN_56 << _T_207_bits_size;
  assign _T_290 = _T_289[22:8];
  assign _T_294 = _T_207_bits_burst == 2'h2;
  assign _GEN_57 = {{1'd0}, _T_290};
  assign _T_295 = _T_286 & _GEN_57;
  assign _T_296 = ~ _T_207_bits_addr;
  assign _GEN_58 = {{3'd0}, _T_296};
  assign _T_297 = _GEN_58 | _T_290;
  assign _T_298 = ~ _T_297;
  assign _GEN_59 = {{1'd0}, _T_298};
  assign _T_299 = _T_295 | _GEN_59;
  assign _GEN_1 = _T_294 ? _T_299 : _T_286;
  assign _GEN_2 = _T_271 ? {{4'd0}, _T_207_bits_addr} : _GEN_1;
  assign _T_302 = 8'h0 == _T_222;
  assign _T_303 = _T_211_ready & _T_302;
  assign _T_304 = ~ _T_223;
  assign _T_307 = 10'h7 << _T_207_bits_size;
  assign _T_308 = _T_307[2:0];
  assign _T_309 = ~ _T_308;
  assign _GEN_60 = {{9'd0}, _T_309};
  assign _T_310 = _T_304 | _GEN_60;
  assign _T_311 = ~ _T_310;
  assign _T_312 = _T_211_ready & _T_211_valid;
  assign _T_314 = _T_302 == 1'h0;
  assign _GEN_61 = {{1'd0}, _T_222};
  assign _T_315 = _GEN_61 - _T_279;
  assign _T_316 = $unsigned(_T_315);
  assign _T_317 = _T_316[8:0];
  assign _GEN_3 = _T_312 ? _T_314 : _T_217;
  assign _GEN_4 = _T_312 ? _T_292 : {{4'd0}, _T_219};
  assign _GEN_5 = _T_312 ? _T_317 : {{1'd0}, _T_221};
  assign _T_337 = _T_332 ? _T_336 : _T_322_bits_len;
  assign _T_338 = _T_332 ? _T_334 : _T_322_bits_addr;
  assign _T_386 = _T_322_bits_burst == 2'h0;
  assign _T_399 = _GEN_54 << _T_322_bits_size;
  assign _GEN_73 = {{4'd0}, _T_338};
  assign _T_400 = _GEN_73 + _T_399;
  assign _T_401 = _T_400[15:0];
  assign _T_403 = {_T_322_bits_len,8'hff};
  assign _GEN_74 = {{7'd0}, _T_403};
  assign _T_404 = _GEN_74 << _T_322_bits_size;
  assign _T_405 = _T_404[22:8];
  assign _T_409 = _T_322_bits_burst == 2'h2;
  assign _GEN_75 = {{1'd0}, _T_405};
  assign _T_410 = _T_401 & _GEN_75;
  assign _T_411 = ~ _T_322_bits_addr;
  assign _GEN_76 = {{3'd0}, _T_411};
  assign _T_412 = _GEN_76 | _T_405;
  assign _T_413 = ~ _T_412;
  assign _GEN_77 = {{1'd0}, _T_413};
  assign _T_414 = _T_410 | _GEN_77;
  assign _GEN_6 = _T_409 ? _T_414 : _T_401;
  assign _GEN_7 = _T_386 ? {{4'd0}, _T_322_bits_addr} : _GEN_6;
  assign _T_417 = 8'h0 == _T_337;
  assign _T_418 = _T_326_ready & _T_417;
  assign _T_419 = ~ _T_338;
  assign _T_422 = 10'h7 << _T_322_bits_size;
  assign _T_423 = _T_422[2:0];
  assign _T_424 = ~ _T_423;
  assign _GEN_78 = {{9'd0}, _T_424};
  assign _T_425 = _T_419 | _GEN_78;
  assign _T_426 = ~ _T_425;
  assign _T_427 = _T_326_ready & _T_326_valid;
  assign _T_429 = _T_417 == 1'h0;
  assign _GEN_79 = {{1'd0}, _T_337};
  assign _T_430 = _GEN_79 - _T_279;
  assign _T_431 = $unsigned(_T_430);
  assign _T_432 = _T_431[8:0];
  assign _GEN_8 = _T_427 ? _T_429 : _T_332;
  assign _GEN_9 = _T_427 ? _T_407 : {{4'd0}, _T_334};
  assign _GEN_10 = _T_427 ? _T_432 : {{1'd0}, _T_336};
  assign _T_448 = _T_447 & _T_445;
  assign _GEN_11 = _T_448 ? 1'h1 : _T_443;
  assign _T_450 = _T_89_aw_ready & _T_89_aw_valid;
  assign _GEN_12 = _T_450 ? 1'h0 : _GEN_11;
  assign _T_452 = _T_445 | _T_443;
  assign _T_453 = _T_326_valid & _T_452;
  assign _T_455 = _T_89_aw_ready & _T_452;
  assign _T_457 = _T_443 == 1'h0;
  assign _T_458 = _T_326_valid & _T_457;
  assign _T_463 = _T_461 == 9'h0;
  assign _T_465 = _T_447 ? _T_279 : 9'h0;
  assign _T_466 = _T_463 ? _T_465 : _T_461;
  assign _T_468 = _T_466 == 9'h1;
  assign _T_469 = _T_89_w_ready & _T_89_w_valid;
  assign _GEN_80 = {{8'd0}, _T_469};
  assign _T_470 = _T_466 - _GEN_80;
  assign _T_471 = $unsigned(_T_470);
  assign _T_472 = _T_471[8:0];
  assign _T_475 = _T_469 == 1'h0;
  assign _T_477 = _T_466 != 9'h0;
  assign _T_478 = _T_475 | _T_477;
  assign _T_480 = _T_478 | reset;
  assign _T_482 = _T_480 == 1'h0;
  assign _T_484 = _T_445 == 1'h0;
  assign _T_485 = _T_484 | _T_447;
  assign _T_486 = _T_437_valid & _T_485;
  assign _T_490 = _T_89_w_ready & _T_485;
  assign _T_492 = _T_89_w_valid == 1'h0;
  assign _T_494 = _T_437_bits_last == 1'h0;
  assign _T_495 = _T_492 | _T_494;
  assign _T_496 = _T_495 | _T_468;
  assign _T_498 = _T_496 | reset;
  assign _T_500 = _T_498 == 1'h0;
  assign _T_502 = _T_89_r_bits_last & _T_89_r_bits_user;
  assign _T_504 = _T_89_b_valid & _T_89_b_bits_user;
  assign _T_506 = _T_89_b_bits_user == 1'h0;
  assign _T_507 = _T_31_b_ready | _T_506;
  assign _GEN_13 = 4'h1 == _T_89_b_bits_id ? _T_581_1 : _T_581_0;
  assign _GEN_14 = 4'h2 == _T_89_b_bits_id ? _T_581_2 : _GEN_13;
  assign _GEN_15 = 4'h3 == _T_89_b_bits_id ? _T_581_3 : _GEN_14;
  assign _GEN_16 = 4'h4 == _T_89_b_bits_id ? _T_581_4 : _GEN_15;
  assign _GEN_17 = 4'h5 == _T_89_b_bits_id ? _T_581_5 : _GEN_16;
  assign _GEN_18 = 4'h6 == _T_89_b_bits_id ? _T_581_6 : _GEN_17;
  assign _GEN_19 = 4'h7 == _T_89_b_bits_id ? _T_581_7 : _GEN_18;
  assign _GEN_20 = 4'h8 == _T_89_b_bits_id ? _T_581_8 : _GEN_19;
  assign _GEN_21 = 4'h9 == _T_89_b_bits_id ? _T_581_9 : _GEN_20;
  assign _GEN_22 = 4'ha == _T_89_b_bits_id ? _T_581_10 : _GEN_21;
  assign _GEN_23 = 4'hb == _T_89_b_bits_id ? _T_581_11 : _GEN_22;
  assign _GEN_24 = 4'hc == _T_89_b_bits_id ? _T_581_12 : _GEN_23;
  assign _GEN_25 = 4'hd == _T_89_b_bits_id ? _T_581_13 : _GEN_24;
  assign _GEN_26 = 4'he == _T_89_b_bits_id ? _T_581_14 : _GEN_25;
  assign _GEN_27 = 4'hf == _T_89_b_bits_id ? _T_581_15 : _GEN_26;
  assign _T_637 = _T_89_b_bits_resp | _GEN_0;
  assign _T_640 = 16'h1 << _T_89_b_bits_id;
  assign _T_642 = _T_640[0];
  assign _T_643 = _T_640[1];
  assign _T_644 = _T_640[2];
  assign _T_645 = _T_640[3];
  assign _T_646 = _T_640[4];
  assign _T_647 = _T_640[5];
  assign _T_648 = _T_640[6];
  assign _T_649 = _T_640[7];
  assign _T_650 = _T_640[8];
  assign _T_651 = _T_640[9];
  assign _T_652 = _T_640[10];
  assign _T_653 = _T_640[11];
  assign _T_654 = _T_640[12];
  assign _T_655 = _T_640[13];
  assign _T_656 = _T_640[14];
  assign _T_657 = _T_640[15];
  assign _T_658 = _T_89_b_ready & _T_89_b_valid;
  assign _T_659 = _T_642 & _T_658;
  assign _T_661 = _T_581_0 | _T_89_b_bits_resp;
  assign _T_662 = _T_89_b_bits_user ? 2'h0 : _T_661;
  assign _GEN_28 = _T_659 ? _T_662 : _T_581_0;
  assign _T_664 = _T_643 & _T_658;
  assign _T_666 = _T_581_1 | _T_89_b_bits_resp;
  assign _T_667 = _T_89_b_bits_user ? 2'h0 : _T_666;
  assign _GEN_29 = _T_664 ? _T_667 : _T_581_1;
  assign _T_669 = _T_644 & _T_658;
  assign _T_671 = _T_581_2 | _T_89_b_bits_resp;
  assign _T_672 = _T_89_b_bits_user ? 2'h0 : _T_671;
  assign _GEN_30 = _T_669 ? _T_672 : _T_581_2;
  assign _T_674 = _T_645 & _T_658;
  assign _T_676 = _T_581_3 | _T_89_b_bits_resp;
  assign _T_677 = _T_89_b_bits_user ? 2'h0 : _T_676;
  assign _GEN_31 = _T_674 ? _T_677 : _T_581_3;
  assign _T_679 = _T_646 & _T_658;
  assign _T_681 = _T_581_4 | _T_89_b_bits_resp;
  assign _T_682 = _T_89_b_bits_user ? 2'h0 : _T_681;
  assign _GEN_32 = _T_679 ? _T_682 : _T_581_4;
  assign _T_684 = _T_647 & _T_658;
  assign _T_686 = _T_581_5 | _T_89_b_bits_resp;
  assign _T_687 = _T_89_b_bits_user ? 2'h0 : _T_686;
  assign _GEN_33 = _T_684 ? _T_687 : _T_581_5;
  assign _T_689 = _T_648 & _T_658;
  assign _T_691 = _T_581_6 | _T_89_b_bits_resp;
  assign _T_692 = _T_89_b_bits_user ? 2'h0 : _T_691;
  assign _GEN_34 = _T_689 ? _T_692 : _T_581_6;
  assign _T_694 = _T_649 & _T_658;
  assign _T_696 = _T_581_7 | _T_89_b_bits_resp;
  assign _T_697 = _T_89_b_bits_user ? 2'h0 : _T_696;
  assign _GEN_35 = _T_694 ? _T_697 : _T_581_7;
  assign _T_699 = _T_650 & _T_658;
  assign _T_701 = _T_581_8 | _T_89_b_bits_resp;
  assign _T_702 = _T_89_b_bits_user ? 2'h0 : _T_701;
  assign _GEN_36 = _T_699 ? _T_702 : _T_581_8;
  assign _T_704 = _T_651 & _T_658;
  assign _T_706 = _T_581_9 | _T_89_b_bits_resp;
  assign _T_707 = _T_89_b_bits_user ? 2'h0 : _T_706;
  assign _GEN_37 = _T_704 ? _T_707 : _T_581_9;
  assign _T_709 = _T_652 & _T_658;
  assign _T_711 = _T_581_10 | _T_89_b_bits_resp;
  assign _T_712 = _T_89_b_bits_user ? 2'h0 : _T_711;
  assign _GEN_38 = _T_709 ? _T_712 : _T_581_10;
  assign _T_714 = _T_653 & _T_658;
  assign _T_716 = _T_581_11 | _T_89_b_bits_resp;
  assign _T_717 = _T_89_b_bits_user ? 2'h0 : _T_716;
  assign _GEN_39 = _T_714 ? _T_717 : _T_581_11;
  assign _T_719 = _T_654 & _T_658;
  assign _T_721 = _T_581_12 | _T_89_b_bits_resp;
  assign _T_722 = _T_89_b_bits_user ? 2'h0 : _T_721;
  assign _GEN_40 = _T_719 ? _T_722 : _T_581_12;
  assign _T_724 = _T_655 & _T_658;
  assign _T_726 = _T_581_13 | _T_89_b_bits_resp;
  assign _T_727 = _T_89_b_bits_user ? 2'h0 : _T_726;
  assign _GEN_41 = _T_724 ? _T_727 : _T_581_13;
  assign _T_729 = _T_656 & _T_658;
  assign _T_731 = _T_581_14 | _T_89_b_bits_resp;
  assign _T_732 = _T_89_b_bits_user ? 2'h0 : _T_731;
  assign _GEN_42 = _T_729 ? _T_732 : _T_581_14;
  assign _T_734 = _T_657 & _T_658;
  assign _T_736 = _T_581_15 | _T_89_b_bits_resp;
  assign _T_737 = _T_89_b_bits_user ? 2'h0 : _T_736;
  assign _GEN_43 = _T_734 ? _T_737 : _T_581_15;
  assign auto_in_aw_ready = _T_31_aw_ready;
  assign auto_in_w_ready = _T_31_w_ready;
  assign auto_in_b_valid = _T_31_b_valid;
  assign auto_in_b_bits_id = _T_31_b_bits_id;
  assign auto_in_b_bits_resp = _T_31_b_bits_resp;
  assign auto_in_ar_ready = _T_31_ar_ready;
  assign auto_in_r_valid = _T_31_r_valid;
  assign auto_in_r_bits_id = _T_31_r_bits_id;
  assign auto_in_r_bits_data = _T_31_r_bits_data;
  assign auto_in_r_bits_resp = _T_31_r_bits_resp;
  assign auto_in_r_bits_last = _T_31_r_bits_last;
  assign auto_out_aw_valid = _T_89_aw_valid;
  assign auto_out_aw_bits_id = _T_89_aw_bits_id;
  assign auto_out_aw_bits_addr = _T_89_aw_bits_addr;
  assign auto_out_aw_bits_user = _T_89_aw_bits_user;
  assign auto_out_w_valid = _T_89_w_valid;
  assign auto_out_w_bits_data = _T_89_w_bits_data;
  assign auto_out_w_bits_strb = _T_89_w_bits_strb;
  assign auto_out_w_bits_last = _T_89_w_bits_last;
  assign auto_out_b_ready = _T_89_b_ready;
  assign auto_out_ar_valid = _T_89_ar_valid;
  assign auto_out_ar_bits_id = _T_89_ar_bits_id;
  assign auto_out_ar_bits_addr = _T_89_ar_bits_addr;
  assign auto_out_ar_bits_user = _T_89_ar_bits_user;
  assign auto_out_r_ready = _T_89_r_ready;
  assign _T_31_aw_ready = Queue_1_io_enq_ready;
  assign _T_31_aw_valid = auto_in_aw_valid;
  assign _T_31_aw_bits_id = auto_in_aw_bits_id;
  assign _T_31_aw_bits_addr = auto_in_aw_bits_addr;
  assign _T_31_aw_bits_len = auto_in_aw_bits_len;
  assign _T_31_aw_bits_size = auto_in_aw_bits_size;
  assign _T_31_aw_bits_burst = auto_in_aw_bits_burst;
  assign _T_31_w_ready = Queue_2_io_enq_ready;
  assign _T_31_w_valid = auto_in_w_valid;
  assign _T_31_w_bits_data = auto_in_w_bits_data;
  assign _T_31_w_bits_strb = auto_in_w_bits_strb;
  assign _T_31_w_bits_last = auto_in_w_bits_last;
  assign _T_31_b_ready = auto_in_b_ready;
  assign _T_31_b_valid = _T_504;
  assign _T_31_b_bits_id = _T_89_b_bits_id;
  assign _T_31_b_bits_resp = _T_637;
  assign _T_31_ar_ready = Queue_io_enq_ready;
  assign _T_31_ar_valid = auto_in_ar_valid;
  assign _T_31_ar_bits_id = auto_in_ar_bits_id;
  assign _T_31_ar_bits_addr = auto_in_ar_bits_addr;
  assign _T_31_ar_bits_len = auto_in_ar_bits_len;
  assign _T_31_ar_bits_size = auto_in_ar_bits_size;
  assign _T_31_ar_bits_burst = auto_in_ar_bits_burst;
  assign _T_31_r_ready = auto_in_r_ready;
  assign _T_31_r_valid = _T_89_r_valid;
  assign _T_31_r_bits_id = _T_89_r_bits_id;
  assign _T_31_r_bits_data = _T_89_r_bits_data;
  assign _T_31_r_bits_resp = _T_89_r_bits_resp;
  assign _T_31_r_bits_last = _T_502;
  assign _T_89_aw_ready = auto_out_aw_ready;
  assign _T_89_aw_valid = _T_453;
  assign _T_89_aw_bits_id = _T_326_bits_id;
  assign _T_89_aw_bits_addr = _T_326_bits_addr;
  assign _T_89_aw_bits_user = _T_417;
  assign _T_89_w_ready = auto_out_w_ready;
  assign _T_89_w_valid = _T_486;
  assign _T_89_w_bits_data = _T_437_bits_data;
  assign _T_89_w_bits_strb = _T_437_bits_strb;
  assign _T_89_w_bits_last = _T_468;
  assign _T_89_b_ready = _T_507;
  assign _T_89_b_valid = auto_out_b_valid;
  assign _T_89_b_bits_id = auto_out_b_bits_id;
  assign _T_89_b_bits_resp = auto_out_b_bits_resp;
  assign _T_89_b_bits_user = auto_out_b_bits_user;
  assign _T_89_ar_ready = auto_out_ar_ready;
  assign _T_89_ar_valid = _T_211_valid;
  assign _T_89_ar_bits_id = _T_211_bits_id;
  assign _T_89_ar_bits_addr = _T_211_bits_addr;
  assign _T_89_ar_bits_user = _T_302;
  assign _T_89_r_ready = _T_31_r_ready;
  assign _T_89_r_valid = auto_out_r_valid;
  assign _T_89_r_bits_id = auto_out_r_bits_id;
  assign _T_89_r_bits_data = auto_out_r_bits_data;
  assign _T_89_r_bits_resp = auto_out_r_bits_resp;
  assign _T_89_r_bits_user = auto_out_r_bits_user;
  assign _T_89_r_bits_last = auto_out_r_bits_last;
  assign Queue_io_enq_valid = _T_31_ar_valid;
  assign Queue_io_enq_bits_id = _T_31_ar_bits_id;
  assign Queue_io_enq_bits_addr = _T_31_ar_bits_addr;
  assign Queue_io_enq_bits_len = _T_31_ar_bits_len;
  assign Queue_io_enq_bits_size = _T_31_ar_bits_size;
  assign Queue_io_enq_bits_burst = _T_31_ar_bits_burst;
  assign Queue_io_deq_ready = _T_207_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign _T_207_ready = _T_303;
  assign _T_207_valid = Queue_io_deq_valid;
  assign _T_207_bits_id = Queue_io_deq_bits_id;
  assign _T_207_bits_addr = Queue_io_deq_bits_addr;
  assign _T_207_bits_len = Queue_io_deq_bits_len;
  assign _T_207_bits_size = Queue_io_deq_bits_size;
  assign _T_207_bits_burst = Queue_io_deq_bits_burst;
  assign _T_211_ready = _T_89_ar_ready;
  assign _T_211_valid = _T_207_valid;
  assign _T_211_bits_id = _T_207_bits_id;
  assign _T_211_bits_addr = _T_311;
  assign _T_292 = _GEN_2;
  assign Queue_1_io_enq_valid = _T_31_aw_valid;
  assign Queue_1_io_enq_bits_id = _T_31_aw_bits_id;
  assign Queue_1_io_enq_bits_addr = _T_31_aw_bits_addr;
  assign Queue_1_io_enq_bits_len = _T_31_aw_bits_len;
  assign Queue_1_io_enq_bits_size = _T_31_aw_bits_size;
  assign Queue_1_io_enq_bits_burst = _T_31_aw_bits_burst;
  assign Queue_1_io_deq_ready = _T_322_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign _T_322_ready = _T_418;
  assign _T_322_valid = Queue_1_io_deq_valid;
  assign _T_322_bits_id = Queue_1_io_deq_bits_id;
  assign _T_322_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_322_bits_len = Queue_1_io_deq_bits_len;
  assign _T_322_bits_size = Queue_1_io_deq_bits_size;
  assign _T_322_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_326_ready = _T_455;
  assign _T_326_valid = _T_322_valid;
  assign _T_326_bits_id = _T_322_bits_id;
  assign _T_326_bits_addr = _T_426;
  assign _T_407 = _GEN_7;
  assign Queue_2_io_enq_valid = _T_31_w_valid;
  assign Queue_2_io_enq_bits_data = _T_31_w_bits_data;
  assign Queue_2_io_enq_bits_strb = _T_31_w_bits_strb;
  assign Queue_2_io_enq_bits_last = _T_31_w_bits_last;
  assign Queue_2_io_deq_ready = _T_437_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign _T_437_ready = _T_490;
  assign _T_437_valid = Queue_2_io_deq_valid;
  assign _T_437_bits_data = Queue_2_io_deq_bits_data;
  assign _T_437_bits_strb = Queue_2_io_deq_bits_strb;
  assign _T_437_bits_last = Queue_2_io_deq_bits_last;
  assign _T_445 = _T_463;
  assign _T_447 = _T_458;
  assign _GEN_0 = _GEN_27;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_217 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_219 = _RAND_1[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_221 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_332 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_334 = _RAND_4[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_336 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_443 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_461 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_581_0 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_581_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_581_2 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_581_3 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_581_4 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_581_5 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_581_6 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_581_7 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_581_8 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_581_9 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_581_10 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_581_11 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_581_12 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_581_13 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_581_14 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_581_15 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_217 <= 1'h0;
    end else begin
      if (_T_312) begin
        _T_217 <= _T_314;
      end
    end
    _T_219 <= _GEN_4[11:0];
    _T_221 <= _GEN_5[7:0];
    if (reset) begin
      _T_332 <= 1'h0;
    end else begin
      if (_T_427) begin
        _T_332 <= _T_429;
      end
    end
    _T_334 <= _GEN_9[11:0];
    _T_336 <= _GEN_10[7:0];
    if (reset) begin
      _T_443 <= 1'h0;
    end else begin
      if (_T_450) begin
        _T_443 <= 1'h0;
      end else begin
        if (_T_448) begin
          _T_443 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_461 <= 9'h0;
    end else begin
      _T_461 <= _T_472;
    end
    if (reset) begin
      _T_581_0 <= 2'h0;
    end else begin
      if (_T_659) begin
        if (_T_89_b_bits_user) begin
          _T_581_0 <= 2'h0;
        end else begin
          _T_581_0 <= _T_661;
        end
      end
    end
    if (reset) begin
      _T_581_1 <= 2'h0;
    end else begin
      if (_T_664) begin
        if (_T_89_b_bits_user) begin
          _T_581_1 <= 2'h0;
        end else begin
          _T_581_1 <= _T_666;
        end
      end
    end
    if (reset) begin
      _T_581_2 <= 2'h0;
    end else begin
      if (_T_669) begin
        if (_T_89_b_bits_user) begin
          _T_581_2 <= 2'h0;
        end else begin
          _T_581_2 <= _T_671;
        end
      end
    end
    if (reset) begin
      _T_581_3 <= 2'h0;
    end else begin
      if (_T_674) begin
        if (_T_89_b_bits_user) begin
          _T_581_3 <= 2'h0;
        end else begin
          _T_581_3 <= _T_676;
        end
      end
    end
    if (reset) begin
      _T_581_4 <= 2'h0;
    end else begin
      if (_T_679) begin
        if (_T_89_b_bits_user) begin
          _T_581_4 <= 2'h0;
        end else begin
          _T_581_4 <= _T_681;
        end
      end
    end
    if (reset) begin
      _T_581_5 <= 2'h0;
    end else begin
      if (_T_684) begin
        if (_T_89_b_bits_user) begin
          _T_581_5 <= 2'h0;
        end else begin
          _T_581_5 <= _T_686;
        end
      end
    end
    if (reset) begin
      _T_581_6 <= 2'h0;
    end else begin
      if (_T_689) begin
        if (_T_89_b_bits_user) begin
          _T_581_6 <= 2'h0;
        end else begin
          _T_581_6 <= _T_691;
        end
      end
    end
    if (reset) begin
      _T_581_7 <= 2'h0;
    end else begin
      if (_T_694) begin
        if (_T_89_b_bits_user) begin
          _T_581_7 <= 2'h0;
        end else begin
          _T_581_7 <= _T_696;
        end
      end
    end
    if (reset) begin
      _T_581_8 <= 2'h0;
    end else begin
      if (_T_699) begin
        if (_T_89_b_bits_user) begin
          _T_581_8 <= 2'h0;
        end else begin
          _T_581_8 <= _T_701;
        end
      end
    end
    if (reset) begin
      _T_581_9 <= 2'h0;
    end else begin
      if (_T_704) begin
        if (_T_89_b_bits_user) begin
          _T_581_9 <= 2'h0;
        end else begin
          _T_581_9 <= _T_706;
        end
      end
    end
    if (reset) begin
      _T_581_10 <= 2'h0;
    end else begin
      if (_T_709) begin
        if (_T_89_b_bits_user) begin
          _T_581_10 <= 2'h0;
        end else begin
          _T_581_10 <= _T_711;
        end
      end
    end
    if (reset) begin
      _T_581_11 <= 2'h0;
    end else begin
      if (_T_714) begin
        if (_T_89_b_bits_user) begin
          _T_581_11 <= 2'h0;
        end else begin
          _T_581_11 <= _T_716;
        end
      end
    end
    if (reset) begin
      _T_581_12 <= 2'h0;
    end else begin
      if (_T_719) begin
        if (_T_89_b_bits_user) begin
          _T_581_12 <= 2'h0;
        end else begin
          _T_581_12 <= _T_721;
        end
      end
    end
    if (reset) begin
      _T_581_13 <= 2'h0;
    end else begin
      if (_T_724) begin
        if (_T_89_b_bits_user) begin
          _T_581_13 <= 2'h0;
        end else begin
          _T_581_13 <= _T_726;
        end
      end
    end
    if (reset) begin
      _T_581_14 <= 2'h0;
    end else begin
      if (_T_729) begin
        if (_T_89_b_bits_user) begin
          _T_581_14 <= 2'h0;
        end else begin
          _T_581_14 <= _T_731;
        end
      end
    end
    if (reset) begin
      _T_581_15 <= 2'h0;
    end else begin
      if (_T_734) begin
        if (_T_89_b_bits_user) begin
          _T_581_15 <= 2'h0;
        end else begin
          _T_581_15 <= _T_736;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_482) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:166 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_482) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_500) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:175 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_500) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimAXIMem_1(
  input         clock,
  input         reset,
  output        io_axi4_0_aw_ready,
  input         io_axi4_0_aw_valid,
  input  [3:0]  io_axi4_0_aw_bits_id,
  input  [11:0] io_axi4_0_aw_bits_addr,
  input  [7:0]  io_axi4_0_aw_bits_len,
  input  [2:0]  io_axi4_0_aw_bits_size,
  input  [1:0]  io_axi4_0_aw_bits_burst,
  output        io_axi4_0_w_ready,
  input         io_axi4_0_w_valid,
  input  [63:0] io_axi4_0_w_bits_data,
  input  [7:0]  io_axi4_0_w_bits_strb,
  input         io_axi4_0_w_bits_last,
  input         io_axi4_0_b_ready,
  output        io_axi4_0_b_valid,
  output [3:0]  io_axi4_0_b_bits_id,
  output [1:0]  io_axi4_0_b_bits_resp,
  output        io_axi4_0_ar_ready,
  input         io_axi4_0_ar_valid,
  input  [3:0]  io_axi4_0_ar_bits_id,
  input  [11:0] io_axi4_0_ar_bits_addr,
  input  [7:0]  io_axi4_0_ar_bits_len,
  input  [2:0]  io_axi4_0_ar_bits_size,
  input  [1:0]  io_axi4_0_ar_bits_burst,
  input         io_axi4_0_r_ready,
  output        io_axi4_0_r_valid,
  output [3:0]  io_axi4_0_r_bits_id,
  output [63:0] io_axi4_0_r_bits_data,
  output [1:0]  io_axi4_0_r_bits_resp,
  output        io_axi4_0_r_bits_last
);
  wire  AXI4RAM_clock;
  wire  AXI4RAM_reset;
  wire  AXI4RAM_auto_in_aw_ready;
  wire  AXI4RAM_auto_in_aw_valid;
  wire [3:0] AXI4RAM_auto_in_aw_bits_id;
  wire [11:0] AXI4RAM_auto_in_aw_bits_addr;
  wire  AXI4RAM_auto_in_aw_bits_user;
  wire  AXI4RAM_auto_in_w_ready;
  wire  AXI4RAM_auto_in_w_valid;
  wire [63:0] AXI4RAM_auto_in_w_bits_data;
  wire [7:0] AXI4RAM_auto_in_w_bits_strb;
  wire  AXI4RAM_auto_in_b_ready;
  wire  AXI4RAM_auto_in_b_valid;
  wire [3:0] AXI4RAM_auto_in_b_bits_id;
  wire [1:0] AXI4RAM_auto_in_b_bits_resp;
  wire  AXI4RAM_auto_in_b_bits_user;
  wire  AXI4RAM_auto_in_ar_ready;
  wire  AXI4RAM_auto_in_ar_valid;
  wire [3:0] AXI4RAM_auto_in_ar_bits_id;
  wire [11:0] AXI4RAM_auto_in_ar_bits_addr;
  wire  AXI4RAM_auto_in_ar_bits_user;
  wire  AXI4RAM_auto_in_r_ready;
  wire  AXI4RAM_auto_in_r_valid;
  wire [3:0] AXI4RAM_auto_in_r_bits_id;
  wire [63:0] AXI4RAM_auto_in_r_bits_data;
  wire [1:0] AXI4RAM_auto_in_r_bits_resp;
  wire  AXI4RAM_auto_in_r_bits_user;
  wire  AXI4Buffer_clock;
  wire  AXI4Buffer_reset;
  wire  AXI4Buffer_auto_in_aw_ready;
  wire  AXI4Buffer_auto_in_aw_valid;
  wire [3:0] AXI4Buffer_auto_in_aw_bits_id;
  wire [11:0] AXI4Buffer_auto_in_aw_bits_addr;
  wire  AXI4Buffer_auto_in_aw_bits_user;
  wire  AXI4Buffer_auto_in_w_ready;
  wire  AXI4Buffer_auto_in_w_valid;
  wire [63:0] AXI4Buffer_auto_in_w_bits_data;
  wire [7:0] AXI4Buffer_auto_in_w_bits_strb;
  wire  AXI4Buffer_auto_in_w_bits_last;
  wire  AXI4Buffer_auto_in_b_ready;
  wire  AXI4Buffer_auto_in_b_valid;
  wire [3:0] AXI4Buffer_auto_in_b_bits_id;
  wire [1:0] AXI4Buffer_auto_in_b_bits_resp;
  wire  AXI4Buffer_auto_in_b_bits_user;
  wire  AXI4Buffer_auto_in_ar_ready;
  wire  AXI4Buffer_auto_in_ar_valid;
  wire [3:0] AXI4Buffer_auto_in_ar_bits_id;
  wire [11:0] AXI4Buffer_auto_in_ar_bits_addr;
  wire  AXI4Buffer_auto_in_ar_bits_user;
  wire  AXI4Buffer_auto_in_r_ready;
  wire  AXI4Buffer_auto_in_r_valid;
  wire [3:0] AXI4Buffer_auto_in_r_bits_id;
  wire [63:0] AXI4Buffer_auto_in_r_bits_data;
  wire [1:0] AXI4Buffer_auto_in_r_bits_resp;
  wire  AXI4Buffer_auto_in_r_bits_user;
  wire  AXI4Buffer_auto_in_r_bits_last;
  wire  AXI4Buffer_auto_out_aw_ready;
  wire  AXI4Buffer_auto_out_aw_valid;
  wire [3:0] AXI4Buffer_auto_out_aw_bits_id;
  wire [11:0] AXI4Buffer_auto_out_aw_bits_addr;
  wire  AXI4Buffer_auto_out_aw_bits_user;
  wire  AXI4Buffer_auto_out_w_ready;
  wire  AXI4Buffer_auto_out_w_valid;
  wire [63:0] AXI4Buffer_auto_out_w_bits_data;
  wire [7:0] AXI4Buffer_auto_out_w_bits_strb;
  wire  AXI4Buffer_auto_out_b_ready;
  wire  AXI4Buffer_auto_out_b_valid;
  wire [3:0] AXI4Buffer_auto_out_b_bits_id;
  wire [1:0] AXI4Buffer_auto_out_b_bits_resp;
  wire  AXI4Buffer_auto_out_b_bits_user;
  wire  AXI4Buffer_auto_out_ar_ready;
  wire  AXI4Buffer_auto_out_ar_valid;
  wire [3:0] AXI4Buffer_auto_out_ar_bits_id;
  wire [11:0] AXI4Buffer_auto_out_ar_bits_addr;
  wire  AXI4Buffer_auto_out_ar_bits_user;
  wire  AXI4Buffer_auto_out_r_ready;
  wire  AXI4Buffer_auto_out_r_valid;
  wire [3:0] AXI4Buffer_auto_out_r_bits_id;
  wire [63:0] AXI4Buffer_auto_out_r_bits_data;
  wire [1:0] AXI4Buffer_auto_out_r_bits_resp;
  wire  AXI4Buffer_auto_out_r_bits_user;
  wire  AXI4Fragmenter_clock;
  wire  AXI4Fragmenter_reset;
  wire  AXI4Fragmenter_auto_in_aw_ready;
  wire  AXI4Fragmenter_auto_in_aw_valid;
  wire [3:0] AXI4Fragmenter_auto_in_aw_bits_id;
  wire [11:0] AXI4Fragmenter_auto_in_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_aw_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_aw_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_aw_bits_burst;
  wire  AXI4Fragmenter_auto_in_w_ready;
  wire  AXI4Fragmenter_auto_in_w_valid;
  wire [63:0] AXI4Fragmenter_auto_in_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_in_w_bits_strb;
  wire  AXI4Fragmenter_auto_in_w_bits_last;
  wire  AXI4Fragmenter_auto_in_b_ready;
  wire  AXI4Fragmenter_auto_in_b_valid;
  wire [3:0] AXI4Fragmenter_auto_in_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_in_b_bits_resp;
  wire  AXI4Fragmenter_auto_in_ar_ready;
  wire  AXI4Fragmenter_auto_in_ar_valid;
  wire [3:0] AXI4Fragmenter_auto_in_ar_bits_id;
  wire [11:0] AXI4Fragmenter_auto_in_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_auto_in_ar_bits_len;
  wire [2:0] AXI4Fragmenter_auto_in_ar_bits_size;
  wire [1:0] AXI4Fragmenter_auto_in_ar_bits_burst;
  wire  AXI4Fragmenter_auto_in_r_ready;
  wire  AXI4Fragmenter_auto_in_r_valid;
  wire [3:0] AXI4Fragmenter_auto_in_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_in_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_in_r_bits_resp;
  wire  AXI4Fragmenter_auto_in_r_bits_last;
  wire  AXI4Fragmenter_auto_out_aw_ready;
  wire  AXI4Fragmenter_auto_out_aw_valid;
  wire [3:0] AXI4Fragmenter_auto_out_aw_bits_id;
  wire [11:0] AXI4Fragmenter_auto_out_aw_bits_addr;
  wire  AXI4Fragmenter_auto_out_aw_bits_user;
  wire  AXI4Fragmenter_auto_out_w_ready;
  wire  AXI4Fragmenter_auto_out_w_valid;
  wire [63:0] AXI4Fragmenter_auto_out_w_bits_data;
  wire [7:0] AXI4Fragmenter_auto_out_w_bits_strb;
  wire  AXI4Fragmenter_auto_out_w_bits_last;
  wire  AXI4Fragmenter_auto_out_b_ready;
  wire  AXI4Fragmenter_auto_out_b_valid;
  wire [3:0] AXI4Fragmenter_auto_out_b_bits_id;
  wire [1:0] AXI4Fragmenter_auto_out_b_bits_resp;
  wire  AXI4Fragmenter_auto_out_b_bits_user;
  wire  AXI4Fragmenter_auto_out_ar_ready;
  wire  AXI4Fragmenter_auto_out_ar_valid;
  wire [3:0] AXI4Fragmenter_auto_out_ar_bits_id;
  wire [11:0] AXI4Fragmenter_auto_out_ar_bits_addr;
  wire  AXI4Fragmenter_auto_out_ar_bits_user;
  wire  AXI4Fragmenter_auto_out_r_ready;
  wire  AXI4Fragmenter_auto_out_r_valid;
  wire [3:0] AXI4Fragmenter_auto_out_r_bits_id;
  wire [63:0] AXI4Fragmenter_auto_out_r_bits_data;
  wire [1:0] AXI4Fragmenter_auto_out_r_bits_resp;
  wire  AXI4Fragmenter_auto_out_r_bits_user;
  wire  AXI4Fragmenter_auto_out_r_bits_last;
  wire  _T_31_aw_ready;
  wire  _T_31_aw_valid;
  wire [3:0] _T_31_aw_bits_id;
  wire [11:0] _T_31_aw_bits_addr;
  wire [7:0] _T_31_aw_bits_len;
  wire [2:0] _T_31_aw_bits_size;
  wire [1:0] _T_31_aw_bits_burst;
  wire  _T_31_w_ready;
  wire  _T_31_w_valid;
  wire [63:0] _T_31_w_bits_data;
  wire [7:0] _T_31_w_bits_strb;
  wire  _T_31_w_bits_last;
  wire  _T_31_b_ready;
  wire  _T_31_b_valid;
  wire [3:0] _T_31_b_bits_id;
  wire [1:0] _T_31_b_bits_resp;
  wire  _T_31_ar_ready;
  wire  _T_31_ar_valid;
  wire [3:0] _T_31_ar_bits_id;
  wire [11:0] _T_31_ar_bits_addr;
  wire [7:0] _T_31_ar_bits_len;
  wire [2:0] _T_31_ar_bits_size;
  wire [1:0] _T_31_ar_bits_burst;
  wire  _T_31_r_ready;
  wire  _T_31_r_valid;
  wire [3:0] _T_31_r_bits_id;
  wire [63:0] _T_31_r_bits_data;
  wire [1:0] _T_31_r_bits_resp;
  wire  _T_31_r_bits_last;
  AXI4RAM_1 AXI4RAM (
    .clock(AXI4RAM_clock),
    .reset(AXI4RAM_reset),
    .auto_in_aw_ready(AXI4RAM_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4RAM_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4RAM_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4RAM_auto_in_aw_bits_addr),
    .auto_in_aw_bits_user(AXI4RAM_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4RAM_auto_in_w_ready),
    .auto_in_w_valid(AXI4RAM_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4RAM_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4RAM_auto_in_w_bits_strb),
    .auto_in_b_ready(AXI4RAM_auto_in_b_ready),
    .auto_in_b_valid(AXI4RAM_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4RAM_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4RAM_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4RAM_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4RAM_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4RAM_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4RAM_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4RAM_auto_in_ar_bits_addr),
    .auto_in_ar_bits_user(AXI4RAM_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4RAM_auto_in_r_ready),
    .auto_in_r_valid(AXI4RAM_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4RAM_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4RAM_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4RAM_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4RAM_auto_in_r_bits_user)
  );
  AXI4Buffer_2 AXI4Buffer (
    .clock(AXI4Buffer_clock),
    .reset(AXI4Buffer_reset),
    .auto_in_aw_ready(AXI4Buffer_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Buffer_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Buffer_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Buffer_auto_in_aw_bits_addr),
    .auto_in_aw_bits_user(AXI4Buffer_auto_in_aw_bits_user),
    .auto_in_w_ready(AXI4Buffer_auto_in_w_ready),
    .auto_in_w_valid(AXI4Buffer_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Buffer_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Buffer_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Buffer_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Buffer_auto_in_b_ready),
    .auto_in_b_valid(AXI4Buffer_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Buffer_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Buffer_auto_in_b_bits_resp),
    .auto_in_b_bits_user(AXI4Buffer_auto_in_b_bits_user),
    .auto_in_ar_ready(AXI4Buffer_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Buffer_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Buffer_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Buffer_auto_in_ar_bits_addr),
    .auto_in_ar_bits_user(AXI4Buffer_auto_in_ar_bits_user),
    .auto_in_r_ready(AXI4Buffer_auto_in_r_ready),
    .auto_in_r_valid(AXI4Buffer_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Buffer_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Buffer_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Buffer_auto_in_r_bits_resp),
    .auto_in_r_bits_user(AXI4Buffer_auto_in_r_bits_user),
    .auto_in_r_bits_last(AXI4Buffer_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Buffer_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Buffer_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Buffer_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Buffer_auto_out_aw_bits_addr),
    .auto_out_aw_bits_user(AXI4Buffer_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Buffer_auto_out_w_ready),
    .auto_out_w_valid(AXI4Buffer_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Buffer_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Buffer_auto_out_w_bits_strb),
    .auto_out_b_ready(AXI4Buffer_auto_out_b_ready),
    .auto_out_b_valid(AXI4Buffer_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Buffer_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Buffer_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Buffer_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Buffer_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Buffer_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Buffer_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Buffer_auto_out_ar_bits_addr),
    .auto_out_ar_bits_user(AXI4Buffer_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Buffer_auto_out_r_ready),
    .auto_out_r_valid(AXI4Buffer_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Buffer_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Buffer_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Buffer_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Buffer_auto_out_r_bits_user)
  );
  AXI4Fragmenter_2 AXI4Fragmenter (
    .clock(AXI4Fragmenter_clock),
    .reset(AXI4Fragmenter_reset),
    .auto_in_aw_ready(AXI4Fragmenter_auto_in_aw_ready),
    .auto_in_aw_valid(AXI4Fragmenter_auto_in_aw_valid),
    .auto_in_aw_bits_id(AXI4Fragmenter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(AXI4Fragmenter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(AXI4Fragmenter_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(AXI4Fragmenter_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(AXI4Fragmenter_auto_in_aw_bits_burst),
    .auto_in_w_ready(AXI4Fragmenter_auto_in_w_ready),
    .auto_in_w_valid(AXI4Fragmenter_auto_in_w_valid),
    .auto_in_w_bits_data(AXI4Fragmenter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(AXI4Fragmenter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(AXI4Fragmenter_auto_in_w_bits_last),
    .auto_in_b_ready(AXI4Fragmenter_auto_in_b_ready),
    .auto_in_b_valid(AXI4Fragmenter_auto_in_b_valid),
    .auto_in_b_bits_id(AXI4Fragmenter_auto_in_b_bits_id),
    .auto_in_b_bits_resp(AXI4Fragmenter_auto_in_b_bits_resp),
    .auto_in_ar_ready(AXI4Fragmenter_auto_in_ar_ready),
    .auto_in_ar_valid(AXI4Fragmenter_auto_in_ar_valid),
    .auto_in_ar_bits_id(AXI4Fragmenter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(AXI4Fragmenter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(AXI4Fragmenter_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(AXI4Fragmenter_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(AXI4Fragmenter_auto_in_ar_bits_burst),
    .auto_in_r_ready(AXI4Fragmenter_auto_in_r_ready),
    .auto_in_r_valid(AXI4Fragmenter_auto_in_r_valid),
    .auto_in_r_bits_id(AXI4Fragmenter_auto_in_r_bits_id),
    .auto_in_r_bits_data(AXI4Fragmenter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(AXI4Fragmenter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(AXI4Fragmenter_auto_in_r_bits_last),
    .auto_out_aw_ready(AXI4Fragmenter_auto_out_aw_ready),
    .auto_out_aw_valid(AXI4Fragmenter_auto_out_aw_valid),
    .auto_out_aw_bits_id(AXI4Fragmenter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(AXI4Fragmenter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_user(AXI4Fragmenter_auto_out_aw_bits_user),
    .auto_out_w_ready(AXI4Fragmenter_auto_out_w_ready),
    .auto_out_w_valid(AXI4Fragmenter_auto_out_w_valid),
    .auto_out_w_bits_data(AXI4Fragmenter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(AXI4Fragmenter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(AXI4Fragmenter_auto_out_w_bits_last),
    .auto_out_b_ready(AXI4Fragmenter_auto_out_b_ready),
    .auto_out_b_valid(AXI4Fragmenter_auto_out_b_valid),
    .auto_out_b_bits_id(AXI4Fragmenter_auto_out_b_bits_id),
    .auto_out_b_bits_resp(AXI4Fragmenter_auto_out_b_bits_resp),
    .auto_out_b_bits_user(AXI4Fragmenter_auto_out_b_bits_user),
    .auto_out_ar_ready(AXI4Fragmenter_auto_out_ar_ready),
    .auto_out_ar_valid(AXI4Fragmenter_auto_out_ar_valid),
    .auto_out_ar_bits_id(AXI4Fragmenter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(AXI4Fragmenter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_user(AXI4Fragmenter_auto_out_ar_bits_user),
    .auto_out_r_ready(AXI4Fragmenter_auto_out_r_ready),
    .auto_out_r_valid(AXI4Fragmenter_auto_out_r_valid),
    .auto_out_r_bits_id(AXI4Fragmenter_auto_out_r_bits_id),
    .auto_out_r_bits_data(AXI4Fragmenter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(AXI4Fragmenter_auto_out_r_bits_resp),
    .auto_out_r_bits_user(AXI4Fragmenter_auto_out_r_bits_user),
    .auto_out_r_bits_last(AXI4Fragmenter_auto_out_r_bits_last)
  );
  assign io_axi4_0_aw_ready = _T_31_aw_ready;
  assign io_axi4_0_w_ready = _T_31_w_ready;
  assign io_axi4_0_b_valid = _T_31_b_valid;
  assign io_axi4_0_b_bits_id = _T_31_b_bits_id;
  assign io_axi4_0_b_bits_resp = _T_31_b_bits_resp;
  assign io_axi4_0_ar_ready = _T_31_ar_ready;
  assign io_axi4_0_r_valid = _T_31_r_valid;
  assign io_axi4_0_r_bits_id = _T_31_r_bits_id;
  assign io_axi4_0_r_bits_data = _T_31_r_bits_data;
  assign io_axi4_0_r_bits_resp = _T_31_r_bits_resp;
  assign io_axi4_0_r_bits_last = _T_31_r_bits_last;
  assign AXI4RAM_clock = clock;
  assign AXI4RAM_reset = reset;
  assign AXI4RAM_auto_in_aw_valid = AXI4Buffer_auto_out_aw_valid;
  assign AXI4RAM_auto_in_aw_bits_id = AXI4Buffer_auto_out_aw_bits_id;
  assign AXI4RAM_auto_in_aw_bits_addr = AXI4Buffer_auto_out_aw_bits_addr;
  assign AXI4RAM_auto_in_aw_bits_user = AXI4Buffer_auto_out_aw_bits_user;
  assign AXI4RAM_auto_in_w_valid = AXI4Buffer_auto_out_w_valid;
  assign AXI4RAM_auto_in_w_bits_data = AXI4Buffer_auto_out_w_bits_data;
  assign AXI4RAM_auto_in_w_bits_strb = AXI4Buffer_auto_out_w_bits_strb;
  assign AXI4RAM_auto_in_b_ready = AXI4Buffer_auto_out_b_ready;
  assign AXI4RAM_auto_in_ar_valid = AXI4Buffer_auto_out_ar_valid;
  assign AXI4RAM_auto_in_ar_bits_id = AXI4Buffer_auto_out_ar_bits_id;
  assign AXI4RAM_auto_in_ar_bits_addr = AXI4Buffer_auto_out_ar_bits_addr;
  assign AXI4RAM_auto_in_ar_bits_user = AXI4Buffer_auto_out_ar_bits_user;
  assign AXI4RAM_auto_in_r_ready = AXI4Buffer_auto_out_r_ready;
  assign AXI4Buffer_clock = clock;
  assign AXI4Buffer_reset = reset;
  assign AXI4Buffer_auto_in_aw_valid = AXI4Fragmenter_auto_out_aw_valid;
  assign AXI4Buffer_auto_in_aw_bits_id = AXI4Fragmenter_auto_out_aw_bits_id;
  assign AXI4Buffer_auto_in_aw_bits_addr = AXI4Fragmenter_auto_out_aw_bits_addr;
  assign AXI4Buffer_auto_in_aw_bits_user = AXI4Fragmenter_auto_out_aw_bits_user;
  assign AXI4Buffer_auto_in_w_valid = AXI4Fragmenter_auto_out_w_valid;
  assign AXI4Buffer_auto_in_w_bits_data = AXI4Fragmenter_auto_out_w_bits_data;
  assign AXI4Buffer_auto_in_w_bits_strb = AXI4Fragmenter_auto_out_w_bits_strb;
  assign AXI4Buffer_auto_in_w_bits_last = AXI4Fragmenter_auto_out_w_bits_last;
  assign AXI4Buffer_auto_in_b_ready = AXI4Fragmenter_auto_out_b_ready;
  assign AXI4Buffer_auto_in_ar_valid = AXI4Fragmenter_auto_out_ar_valid;
  assign AXI4Buffer_auto_in_ar_bits_id = AXI4Fragmenter_auto_out_ar_bits_id;
  assign AXI4Buffer_auto_in_ar_bits_addr = AXI4Fragmenter_auto_out_ar_bits_addr;
  assign AXI4Buffer_auto_in_ar_bits_user = AXI4Fragmenter_auto_out_ar_bits_user;
  assign AXI4Buffer_auto_in_r_ready = AXI4Fragmenter_auto_out_r_ready;
  assign AXI4Buffer_auto_out_aw_ready = AXI4RAM_auto_in_aw_ready;
  assign AXI4Buffer_auto_out_w_ready = AXI4RAM_auto_in_w_ready;
  assign AXI4Buffer_auto_out_b_valid = AXI4RAM_auto_in_b_valid;
  assign AXI4Buffer_auto_out_b_bits_id = AXI4RAM_auto_in_b_bits_id;
  assign AXI4Buffer_auto_out_b_bits_resp = AXI4RAM_auto_in_b_bits_resp;
  assign AXI4Buffer_auto_out_b_bits_user = AXI4RAM_auto_in_b_bits_user;
  assign AXI4Buffer_auto_out_ar_ready = AXI4RAM_auto_in_ar_ready;
  assign AXI4Buffer_auto_out_r_valid = AXI4RAM_auto_in_r_valid;
  assign AXI4Buffer_auto_out_r_bits_id = AXI4RAM_auto_in_r_bits_id;
  assign AXI4Buffer_auto_out_r_bits_data = AXI4RAM_auto_in_r_bits_data;
  assign AXI4Buffer_auto_out_r_bits_resp = AXI4RAM_auto_in_r_bits_resp;
  assign AXI4Buffer_auto_out_r_bits_user = AXI4RAM_auto_in_r_bits_user;
  assign AXI4Fragmenter_clock = clock;
  assign AXI4Fragmenter_reset = reset;
  assign AXI4Fragmenter_auto_in_aw_valid = _T_31_aw_valid;
  assign AXI4Fragmenter_auto_in_aw_bits_id = _T_31_aw_bits_id;
  assign AXI4Fragmenter_auto_in_aw_bits_addr = _T_31_aw_bits_addr;
  assign AXI4Fragmenter_auto_in_aw_bits_len = _T_31_aw_bits_len;
  assign AXI4Fragmenter_auto_in_aw_bits_size = _T_31_aw_bits_size;
  assign AXI4Fragmenter_auto_in_aw_bits_burst = _T_31_aw_bits_burst;
  assign AXI4Fragmenter_auto_in_w_valid = _T_31_w_valid;
  assign AXI4Fragmenter_auto_in_w_bits_data = _T_31_w_bits_data;
  assign AXI4Fragmenter_auto_in_w_bits_strb = _T_31_w_bits_strb;
  assign AXI4Fragmenter_auto_in_w_bits_last = _T_31_w_bits_last;
  assign AXI4Fragmenter_auto_in_b_ready = _T_31_b_ready;
  assign AXI4Fragmenter_auto_in_ar_valid = _T_31_ar_valid;
  assign AXI4Fragmenter_auto_in_ar_bits_id = _T_31_ar_bits_id;
  assign AXI4Fragmenter_auto_in_ar_bits_addr = _T_31_ar_bits_addr;
  assign AXI4Fragmenter_auto_in_ar_bits_len = _T_31_ar_bits_len;
  assign AXI4Fragmenter_auto_in_ar_bits_size = _T_31_ar_bits_size;
  assign AXI4Fragmenter_auto_in_ar_bits_burst = _T_31_ar_bits_burst;
  assign AXI4Fragmenter_auto_in_r_ready = _T_31_r_ready;
  assign AXI4Fragmenter_auto_out_aw_ready = AXI4Buffer_auto_in_aw_ready;
  assign AXI4Fragmenter_auto_out_w_ready = AXI4Buffer_auto_in_w_ready;
  assign AXI4Fragmenter_auto_out_b_valid = AXI4Buffer_auto_in_b_valid;
  assign AXI4Fragmenter_auto_out_b_bits_id = AXI4Buffer_auto_in_b_bits_id;
  assign AXI4Fragmenter_auto_out_b_bits_resp = AXI4Buffer_auto_in_b_bits_resp;
  assign AXI4Fragmenter_auto_out_b_bits_user = AXI4Buffer_auto_in_b_bits_user;
  assign AXI4Fragmenter_auto_out_ar_ready = AXI4Buffer_auto_in_ar_ready;
  assign AXI4Fragmenter_auto_out_r_valid = AXI4Buffer_auto_in_r_valid;
  assign AXI4Fragmenter_auto_out_r_bits_id = AXI4Buffer_auto_in_r_bits_id;
  assign AXI4Fragmenter_auto_out_r_bits_data = AXI4Buffer_auto_in_r_bits_data;
  assign AXI4Fragmenter_auto_out_r_bits_resp = AXI4Buffer_auto_in_r_bits_resp;
  assign AXI4Fragmenter_auto_out_r_bits_user = AXI4Buffer_auto_in_r_bits_user;
  assign AXI4Fragmenter_auto_out_r_bits_last = AXI4Buffer_auto_in_r_bits_last;
  assign _T_31_aw_ready = AXI4Fragmenter_auto_in_aw_ready;
  assign _T_31_aw_valid = io_axi4_0_aw_valid;
  assign _T_31_aw_bits_id = io_axi4_0_aw_bits_id;
  assign _T_31_aw_bits_addr = io_axi4_0_aw_bits_addr;
  assign _T_31_aw_bits_len = io_axi4_0_aw_bits_len;
  assign _T_31_aw_bits_size = io_axi4_0_aw_bits_size;
  assign _T_31_aw_bits_burst = io_axi4_0_aw_bits_burst;
  assign _T_31_w_ready = AXI4Fragmenter_auto_in_w_ready;
  assign _T_31_w_valid = io_axi4_0_w_valid;
  assign _T_31_w_bits_data = io_axi4_0_w_bits_data;
  assign _T_31_w_bits_strb = io_axi4_0_w_bits_strb;
  assign _T_31_w_bits_last = io_axi4_0_w_bits_last;
  assign _T_31_b_ready = io_axi4_0_b_ready;
  assign _T_31_b_valid = AXI4Fragmenter_auto_in_b_valid;
  assign _T_31_b_bits_id = AXI4Fragmenter_auto_in_b_bits_id;
  assign _T_31_b_bits_resp = AXI4Fragmenter_auto_in_b_bits_resp;
  assign _T_31_ar_ready = AXI4Fragmenter_auto_in_ar_ready;
  assign _T_31_ar_valid = io_axi4_0_ar_valid;
  assign _T_31_ar_bits_id = io_axi4_0_ar_bits_id;
  assign _T_31_ar_bits_addr = io_axi4_0_ar_bits_addr;
  assign _T_31_ar_bits_len = io_axi4_0_ar_bits_len;
  assign _T_31_ar_bits_size = io_axi4_0_ar_bits_size;
  assign _T_31_ar_bits_burst = io_axi4_0_ar_bits_burst;
  assign _T_31_r_ready = io_axi4_0_r_ready;
  assign _T_31_r_valid = AXI4Fragmenter_auto_in_r_valid;
  assign _T_31_r_bits_id = AXI4Fragmenter_auto_in_r_bits_id;
  assign _T_31_r_bits_data = AXI4Fragmenter_auto_in_r_bits_data;
  assign _T_31_r_bits_resp = AXI4Fragmenter_auto_in_r_bits_resp;
  assign _T_31_r_bits_last = AXI4Fragmenter_auto_in_r_bits_last;
endmodule
module TestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  ExampleBoomSystem_clock;
  wire  ExampleBoomSystem_reset;
  wire  ExampleBoomSystem_debug_clockeddmi_dmi_req_ready;
  wire  ExampleBoomSystem_debug_clockeddmi_dmi_req_valid;
  wire [6:0] ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_addr;
  wire [31:0] ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_data;
  wire [1:0] ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_op;
  wire  ExampleBoomSystem_debug_clockeddmi_dmi_resp_ready;
  wire  ExampleBoomSystem_debug_clockeddmi_dmi_resp_valid;
  wire [31:0] ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_data;
  wire [1:0] ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_resp;
  wire  ExampleBoomSystem_debug_clockeddmi_dmiClock;
  wire  ExampleBoomSystem_debug_clockeddmi_dmiReset;
  wire  ExampleBoomSystem_debug_ndreset;
  wire  ExampleBoomSystem_debug_dmactive;
  wire [1:0] ExampleBoomSystem_interrupts;
  wire  ExampleBoomSystem_mem_axi4_0_aw_ready;
  wire  ExampleBoomSystem_mem_axi4_0_aw_valid;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_aw_bits_id;
  wire [31:0] ExampleBoomSystem_mem_axi4_0_aw_bits_addr;
  wire [7:0] ExampleBoomSystem_mem_axi4_0_aw_bits_len;
  wire [2:0] ExampleBoomSystem_mem_axi4_0_aw_bits_size;
  wire [1:0] ExampleBoomSystem_mem_axi4_0_aw_bits_burst;
  wire  ExampleBoomSystem_mem_axi4_0_aw_bits_lock;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_aw_bits_cache;
  wire [2:0] ExampleBoomSystem_mem_axi4_0_aw_bits_prot;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_aw_bits_qos;
  wire  ExampleBoomSystem_mem_axi4_0_w_ready;
  wire  ExampleBoomSystem_mem_axi4_0_w_valid;
  wire [63:0] ExampleBoomSystem_mem_axi4_0_w_bits_data;
  wire [7:0] ExampleBoomSystem_mem_axi4_0_w_bits_strb;
  wire  ExampleBoomSystem_mem_axi4_0_w_bits_last;
  wire  ExampleBoomSystem_mem_axi4_0_b_ready;
  wire  ExampleBoomSystem_mem_axi4_0_b_valid;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_b_bits_id;
  wire [1:0] ExampleBoomSystem_mem_axi4_0_b_bits_resp;
  wire  ExampleBoomSystem_mem_axi4_0_ar_ready;
  wire  ExampleBoomSystem_mem_axi4_0_ar_valid;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_ar_bits_id;
  wire [31:0] ExampleBoomSystem_mem_axi4_0_ar_bits_addr;
  wire [7:0] ExampleBoomSystem_mem_axi4_0_ar_bits_len;
  wire [2:0] ExampleBoomSystem_mem_axi4_0_ar_bits_size;
  wire [1:0] ExampleBoomSystem_mem_axi4_0_ar_bits_burst;
  wire  ExampleBoomSystem_mem_axi4_0_ar_bits_lock;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_ar_bits_cache;
  wire [2:0] ExampleBoomSystem_mem_axi4_0_ar_bits_prot;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_ar_bits_qos;
  wire  ExampleBoomSystem_mem_axi4_0_r_ready;
  wire  ExampleBoomSystem_mem_axi4_0_r_valid;
  wire [3:0] ExampleBoomSystem_mem_axi4_0_r_bits_id;
  wire [63:0] ExampleBoomSystem_mem_axi4_0_r_bits_data;
  wire [1:0] ExampleBoomSystem_mem_axi4_0_r_bits_resp;
  wire  ExampleBoomSystem_mem_axi4_0_r_bits_last;
  wire  ExampleBoomSystem_mmio_axi4_0_aw_ready;
  wire  ExampleBoomSystem_mmio_axi4_0_aw_valid;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_id;
  wire [30:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_addr;
  wire [7:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_len;
  wire [2:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_size;
  wire [1:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_burst;
  wire  ExampleBoomSystem_mmio_axi4_0_aw_bits_lock;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_cache;
  wire [2:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_prot;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_aw_bits_qos;
  wire  ExampleBoomSystem_mmio_axi4_0_w_ready;
  wire  ExampleBoomSystem_mmio_axi4_0_w_valid;
  wire [63:0] ExampleBoomSystem_mmio_axi4_0_w_bits_data;
  wire [7:0] ExampleBoomSystem_mmio_axi4_0_w_bits_strb;
  wire  ExampleBoomSystem_mmio_axi4_0_w_bits_last;
  wire  ExampleBoomSystem_mmio_axi4_0_b_ready;
  wire  ExampleBoomSystem_mmio_axi4_0_b_valid;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_b_bits_id;
  wire [1:0] ExampleBoomSystem_mmio_axi4_0_b_bits_resp;
  wire  ExampleBoomSystem_mmio_axi4_0_ar_ready;
  wire  ExampleBoomSystem_mmio_axi4_0_ar_valid;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_id;
  wire [30:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_addr;
  wire [7:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_len;
  wire [2:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_size;
  wire [1:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_burst;
  wire  ExampleBoomSystem_mmio_axi4_0_ar_bits_lock;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_cache;
  wire [2:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_prot;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_ar_bits_qos;
  wire  ExampleBoomSystem_mmio_axi4_0_r_ready;
  wire  ExampleBoomSystem_mmio_axi4_0_r_valid;
  wire [3:0] ExampleBoomSystem_mmio_axi4_0_r_bits_id;
  wire [63:0] ExampleBoomSystem_mmio_axi4_0_r_bits_data;
  wire [1:0] ExampleBoomSystem_mmio_axi4_0_r_bits_resp;
  wire  ExampleBoomSystem_mmio_axi4_0_r_bits_last;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_ready;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_valid;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_id;
  wire [31:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_addr;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_len;
  wire [2:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_size;
  wire [1:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_burst;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_lock;
  wire [3:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_cache;
  wire [2:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_prot;
  wire [3:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_qos;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_w_ready;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_w_valid;
  wire [63:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_data;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_strb;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_last;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_b_ready;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_b_valid;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_b_bits_id;
  wire [1:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_b_bits_resp;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_ready;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_valid;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_id;
  wire [31:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_addr;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_len;
  wire [2:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_size;
  wire [1:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_burst;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_lock;
  wire [3:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_cache;
  wire [2:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_prot;
  wire [3:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_qos;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_r_ready;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_r_valid;
  wire [7:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_id;
  wire [63:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_data;
  wire [1:0] ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_resp;
  wire  ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_last;
  wire  _T_180;
  wire  SimAXIMem_clock;
  wire  SimAXIMem_reset;
  wire  SimAXIMem_io_axi4_0_aw_ready;
  wire  SimAXIMem_io_axi4_0_aw_valid;
  wire [3:0] SimAXIMem_io_axi4_0_aw_bits_id;
  wire [27:0] SimAXIMem_io_axi4_0_aw_bits_addr;
  wire [7:0] SimAXIMem_io_axi4_0_aw_bits_len;
  wire [2:0] SimAXIMem_io_axi4_0_aw_bits_size;
  wire [1:0] SimAXIMem_io_axi4_0_aw_bits_burst;
  wire  SimAXIMem_io_axi4_0_w_ready;
  wire  SimAXIMem_io_axi4_0_w_valid;
  wire [63:0] SimAXIMem_io_axi4_0_w_bits_data;
  wire [7:0] SimAXIMem_io_axi4_0_w_bits_strb;
  wire  SimAXIMem_io_axi4_0_w_bits_last;
  wire  SimAXIMem_io_axi4_0_b_ready;
  wire  SimAXIMem_io_axi4_0_b_valid;
  wire [3:0] SimAXIMem_io_axi4_0_b_bits_id;
  wire [1:0] SimAXIMem_io_axi4_0_b_bits_resp;
  wire  SimAXIMem_io_axi4_0_ar_ready;
  wire  SimAXIMem_io_axi4_0_ar_valid;
  wire [3:0] SimAXIMem_io_axi4_0_ar_bits_id;
  wire [27:0] SimAXIMem_io_axi4_0_ar_bits_addr;
  wire [7:0] SimAXIMem_io_axi4_0_ar_bits_len;
  wire [2:0] SimAXIMem_io_axi4_0_ar_bits_size;
  wire [1:0] SimAXIMem_io_axi4_0_ar_bits_burst;
  wire  SimAXIMem_io_axi4_0_r_ready;
  wire  SimAXIMem_io_axi4_0_r_valid;
  wire [3:0] SimAXIMem_io_axi4_0_r_bits_id;
  wire [63:0] SimAXIMem_io_axi4_0_r_bits_data;
  wire [1:0] SimAXIMem_io_axi4_0_r_bits_resp;
  wire  SimAXIMem_io_axi4_0_r_bits_last;
  wire  SimAXIMem_1_clock;
  wire  SimAXIMem_1_reset;
  wire  SimAXIMem_1_io_axi4_0_aw_ready;
  wire  SimAXIMem_1_io_axi4_0_aw_valid;
  wire [3:0] SimAXIMem_1_io_axi4_0_aw_bits_id;
  wire [11:0] SimAXIMem_1_io_axi4_0_aw_bits_addr;
  wire [7:0] SimAXIMem_1_io_axi4_0_aw_bits_len;
  wire [2:0] SimAXIMem_1_io_axi4_0_aw_bits_size;
  wire [1:0] SimAXIMem_1_io_axi4_0_aw_bits_burst;
  wire  SimAXIMem_1_io_axi4_0_w_ready;
  wire  SimAXIMem_1_io_axi4_0_w_valid;
  wire [63:0] SimAXIMem_1_io_axi4_0_w_bits_data;
  wire [7:0] SimAXIMem_1_io_axi4_0_w_bits_strb;
  wire  SimAXIMem_1_io_axi4_0_w_bits_last;
  wire  SimAXIMem_1_io_axi4_0_b_ready;
  wire  SimAXIMem_1_io_axi4_0_b_valid;
  wire [3:0] SimAXIMem_1_io_axi4_0_b_bits_id;
  wire [1:0] SimAXIMem_1_io_axi4_0_b_bits_resp;
  wire  SimAXIMem_1_io_axi4_0_ar_ready;
  wire  SimAXIMem_1_io_axi4_0_ar_valid;
  wire [3:0] SimAXIMem_1_io_axi4_0_ar_bits_id;
  wire [11:0] SimAXIMem_1_io_axi4_0_ar_bits_addr;
  wire [7:0] SimAXIMem_1_io_axi4_0_ar_bits_len;
  wire [2:0] SimAXIMem_1_io_axi4_0_ar_bits_size;
  wire [1:0] SimAXIMem_1_io_axi4_0_ar_bits_burst;
  wire  SimAXIMem_1_io_axi4_0_r_ready;
  wire  SimAXIMem_1_io_axi4_0_r_valid;
  wire [3:0] SimAXIMem_1_io_axi4_0_r_bits_id;
  wire [63:0] SimAXIMem_1_io_axi4_0_r_bits_data;
  wire [1:0] SimAXIMem_1_io_axi4_0_r_bits_resp;
  wire  SimAXIMem_1_io_axi4_0_r_bits_last;
  wire [31:0] SimDTM_exit;
  wire  SimDTM_debug_req_ready;
  wire  SimDTM_debug_req_valid;
  wire [6:0] SimDTM_debug_req_bits_addr;
  wire [31:0] SimDTM_debug_req_bits_data;
  wire [1:0] SimDTM_debug_req_bits_op;
  wire  SimDTM_debug_resp_ready;
  wire  SimDTM_debug_resp_valid;
  wire [31:0] SimDTM_debug_resp_bits_data;
  wire [1:0] SimDTM_debug_resp_bits_resp;
  wire  SimDTM_reset;
  wire  SimDTM_clk;
  wire  _T_197;
  wire  _T_199;
  wire [31:0] _T_201;
  wire  _T_204;
  ExampleBoomSystem ExampleBoomSystem (
    .clock(ExampleBoomSystem_clock),
    .reset(ExampleBoomSystem_reset),
    .debug_clockeddmi_dmi_req_ready(ExampleBoomSystem_debug_clockeddmi_dmi_req_ready),
    .debug_clockeddmi_dmi_req_valid(ExampleBoomSystem_debug_clockeddmi_dmi_req_valid),
    .debug_clockeddmi_dmi_req_bits_addr(ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_addr),
    .debug_clockeddmi_dmi_req_bits_data(ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_data),
    .debug_clockeddmi_dmi_req_bits_op(ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_op),
    .debug_clockeddmi_dmi_resp_ready(ExampleBoomSystem_debug_clockeddmi_dmi_resp_ready),
    .debug_clockeddmi_dmi_resp_valid(ExampleBoomSystem_debug_clockeddmi_dmi_resp_valid),
    .debug_clockeddmi_dmi_resp_bits_data(ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_data),
    .debug_clockeddmi_dmi_resp_bits_resp(ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_resp),
    .debug_clockeddmi_dmiClock(ExampleBoomSystem_debug_clockeddmi_dmiClock),
    .debug_clockeddmi_dmiReset(ExampleBoomSystem_debug_clockeddmi_dmiReset),
    .debug_ndreset(ExampleBoomSystem_debug_ndreset),
    .debug_dmactive(ExampleBoomSystem_debug_dmactive),
    .interrupts(ExampleBoomSystem_interrupts),
    .mem_axi4_0_aw_ready(ExampleBoomSystem_mem_axi4_0_aw_ready),
    .mem_axi4_0_aw_valid(ExampleBoomSystem_mem_axi4_0_aw_valid),
    .mem_axi4_0_aw_bits_id(ExampleBoomSystem_mem_axi4_0_aw_bits_id),
    .mem_axi4_0_aw_bits_addr(ExampleBoomSystem_mem_axi4_0_aw_bits_addr),
    .mem_axi4_0_aw_bits_len(ExampleBoomSystem_mem_axi4_0_aw_bits_len),
    .mem_axi4_0_aw_bits_size(ExampleBoomSystem_mem_axi4_0_aw_bits_size),
    .mem_axi4_0_aw_bits_burst(ExampleBoomSystem_mem_axi4_0_aw_bits_burst),
    .mem_axi4_0_aw_bits_lock(ExampleBoomSystem_mem_axi4_0_aw_bits_lock),
    .mem_axi4_0_aw_bits_cache(ExampleBoomSystem_mem_axi4_0_aw_bits_cache),
    .mem_axi4_0_aw_bits_prot(ExampleBoomSystem_mem_axi4_0_aw_bits_prot),
    .mem_axi4_0_aw_bits_qos(ExampleBoomSystem_mem_axi4_0_aw_bits_qos),
    .mem_axi4_0_w_ready(ExampleBoomSystem_mem_axi4_0_w_ready),
    .mem_axi4_0_w_valid(ExampleBoomSystem_mem_axi4_0_w_valid),
    .mem_axi4_0_w_bits_data(ExampleBoomSystem_mem_axi4_0_w_bits_data),
    .mem_axi4_0_w_bits_strb(ExampleBoomSystem_mem_axi4_0_w_bits_strb),
    .mem_axi4_0_w_bits_last(ExampleBoomSystem_mem_axi4_0_w_bits_last),
    .mem_axi4_0_b_ready(ExampleBoomSystem_mem_axi4_0_b_ready),
    .mem_axi4_0_b_valid(ExampleBoomSystem_mem_axi4_0_b_valid),
    .mem_axi4_0_b_bits_id(ExampleBoomSystem_mem_axi4_0_b_bits_id),
    .mem_axi4_0_b_bits_resp(ExampleBoomSystem_mem_axi4_0_b_bits_resp),
    .mem_axi4_0_ar_ready(ExampleBoomSystem_mem_axi4_0_ar_ready),
    .mem_axi4_0_ar_valid(ExampleBoomSystem_mem_axi4_0_ar_valid),
    .mem_axi4_0_ar_bits_id(ExampleBoomSystem_mem_axi4_0_ar_bits_id),
    .mem_axi4_0_ar_bits_addr(ExampleBoomSystem_mem_axi4_0_ar_bits_addr),
    .mem_axi4_0_ar_bits_len(ExampleBoomSystem_mem_axi4_0_ar_bits_len),
    .mem_axi4_0_ar_bits_size(ExampleBoomSystem_mem_axi4_0_ar_bits_size),
    .mem_axi4_0_ar_bits_burst(ExampleBoomSystem_mem_axi4_0_ar_bits_burst),
    .mem_axi4_0_ar_bits_lock(ExampleBoomSystem_mem_axi4_0_ar_bits_lock),
    .mem_axi4_0_ar_bits_cache(ExampleBoomSystem_mem_axi4_0_ar_bits_cache),
    .mem_axi4_0_ar_bits_prot(ExampleBoomSystem_mem_axi4_0_ar_bits_prot),
    .mem_axi4_0_ar_bits_qos(ExampleBoomSystem_mem_axi4_0_ar_bits_qos),
    .mem_axi4_0_r_ready(ExampleBoomSystem_mem_axi4_0_r_ready),
    .mem_axi4_0_r_valid(ExampleBoomSystem_mem_axi4_0_r_valid),
    .mem_axi4_0_r_bits_id(ExampleBoomSystem_mem_axi4_0_r_bits_id),
    .mem_axi4_0_r_bits_data(ExampleBoomSystem_mem_axi4_0_r_bits_data),
    .mem_axi4_0_r_bits_resp(ExampleBoomSystem_mem_axi4_0_r_bits_resp),
    .mem_axi4_0_r_bits_last(ExampleBoomSystem_mem_axi4_0_r_bits_last),
    .mmio_axi4_0_aw_ready(ExampleBoomSystem_mmio_axi4_0_aw_ready),
    .mmio_axi4_0_aw_valid(ExampleBoomSystem_mmio_axi4_0_aw_valid),
    .mmio_axi4_0_aw_bits_id(ExampleBoomSystem_mmio_axi4_0_aw_bits_id),
    .mmio_axi4_0_aw_bits_addr(ExampleBoomSystem_mmio_axi4_0_aw_bits_addr),
    .mmio_axi4_0_aw_bits_len(ExampleBoomSystem_mmio_axi4_0_aw_bits_len),
    .mmio_axi4_0_aw_bits_size(ExampleBoomSystem_mmio_axi4_0_aw_bits_size),
    .mmio_axi4_0_aw_bits_burst(ExampleBoomSystem_mmio_axi4_0_aw_bits_burst),
    .mmio_axi4_0_aw_bits_lock(ExampleBoomSystem_mmio_axi4_0_aw_bits_lock),
    .mmio_axi4_0_aw_bits_cache(ExampleBoomSystem_mmio_axi4_0_aw_bits_cache),
    .mmio_axi4_0_aw_bits_prot(ExampleBoomSystem_mmio_axi4_0_aw_bits_prot),
    .mmio_axi4_0_aw_bits_qos(ExampleBoomSystem_mmio_axi4_0_aw_bits_qos),
    .mmio_axi4_0_w_ready(ExampleBoomSystem_mmio_axi4_0_w_ready),
    .mmio_axi4_0_w_valid(ExampleBoomSystem_mmio_axi4_0_w_valid),
    .mmio_axi4_0_w_bits_data(ExampleBoomSystem_mmio_axi4_0_w_bits_data),
    .mmio_axi4_0_w_bits_strb(ExampleBoomSystem_mmio_axi4_0_w_bits_strb),
    .mmio_axi4_0_w_bits_last(ExampleBoomSystem_mmio_axi4_0_w_bits_last),
    .mmio_axi4_0_b_ready(ExampleBoomSystem_mmio_axi4_0_b_ready),
    .mmio_axi4_0_b_valid(ExampleBoomSystem_mmio_axi4_0_b_valid),
    .mmio_axi4_0_b_bits_id(ExampleBoomSystem_mmio_axi4_0_b_bits_id),
    .mmio_axi4_0_b_bits_resp(ExampleBoomSystem_mmio_axi4_0_b_bits_resp),
    .mmio_axi4_0_ar_ready(ExampleBoomSystem_mmio_axi4_0_ar_ready),
    .mmio_axi4_0_ar_valid(ExampleBoomSystem_mmio_axi4_0_ar_valid),
    .mmio_axi4_0_ar_bits_id(ExampleBoomSystem_mmio_axi4_0_ar_bits_id),
    .mmio_axi4_0_ar_bits_addr(ExampleBoomSystem_mmio_axi4_0_ar_bits_addr),
    .mmio_axi4_0_ar_bits_len(ExampleBoomSystem_mmio_axi4_0_ar_bits_len),
    .mmio_axi4_0_ar_bits_size(ExampleBoomSystem_mmio_axi4_0_ar_bits_size),
    .mmio_axi4_0_ar_bits_burst(ExampleBoomSystem_mmio_axi4_0_ar_bits_burst),
    .mmio_axi4_0_ar_bits_lock(ExampleBoomSystem_mmio_axi4_0_ar_bits_lock),
    .mmio_axi4_0_ar_bits_cache(ExampleBoomSystem_mmio_axi4_0_ar_bits_cache),
    .mmio_axi4_0_ar_bits_prot(ExampleBoomSystem_mmio_axi4_0_ar_bits_prot),
    .mmio_axi4_0_ar_bits_qos(ExampleBoomSystem_mmio_axi4_0_ar_bits_qos),
    .mmio_axi4_0_r_ready(ExampleBoomSystem_mmio_axi4_0_r_ready),
    .mmio_axi4_0_r_valid(ExampleBoomSystem_mmio_axi4_0_r_valid),
    .mmio_axi4_0_r_bits_id(ExampleBoomSystem_mmio_axi4_0_r_bits_id),
    .mmio_axi4_0_r_bits_data(ExampleBoomSystem_mmio_axi4_0_r_bits_data),
    .mmio_axi4_0_r_bits_resp(ExampleBoomSystem_mmio_axi4_0_r_bits_resp),
    .mmio_axi4_0_r_bits_last(ExampleBoomSystem_mmio_axi4_0_r_bits_last),
    .l2_frontend_bus_axi4_0_aw_ready(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_ready),
    .l2_frontend_bus_axi4_0_aw_valid(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_valid),
    .l2_frontend_bus_axi4_0_aw_bits_id(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_id),
    .l2_frontend_bus_axi4_0_aw_bits_addr(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_addr),
    .l2_frontend_bus_axi4_0_aw_bits_len(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_len),
    .l2_frontend_bus_axi4_0_aw_bits_size(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_size),
    .l2_frontend_bus_axi4_0_aw_bits_burst(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_burst),
    .l2_frontend_bus_axi4_0_aw_bits_lock(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_lock),
    .l2_frontend_bus_axi4_0_aw_bits_cache(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_cache),
    .l2_frontend_bus_axi4_0_aw_bits_prot(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_prot),
    .l2_frontend_bus_axi4_0_aw_bits_qos(ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_qos),
    .l2_frontend_bus_axi4_0_w_ready(ExampleBoomSystem_l2_frontend_bus_axi4_0_w_ready),
    .l2_frontend_bus_axi4_0_w_valid(ExampleBoomSystem_l2_frontend_bus_axi4_0_w_valid),
    .l2_frontend_bus_axi4_0_w_bits_data(ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_data),
    .l2_frontend_bus_axi4_0_w_bits_strb(ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_strb),
    .l2_frontend_bus_axi4_0_w_bits_last(ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_last),
    .l2_frontend_bus_axi4_0_b_ready(ExampleBoomSystem_l2_frontend_bus_axi4_0_b_ready),
    .l2_frontend_bus_axi4_0_b_valid(ExampleBoomSystem_l2_frontend_bus_axi4_0_b_valid),
    .l2_frontend_bus_axi4_0_b_bits_id(ExampleBoomSystem_l2_frontend_bus_axi4_0_b_bits_id),
    .l2_frontend_bus_axi4_0_b_bits_resp(ExampleBoomSystem_l2_frontend_bus_axi4_0_b_bits_resp),
    .l2_frontend_bus_axi4_0_ar_ready(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_ready),
    .l2_frontend_bus_axi4_0_ar_valid(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_valid),
    .l2_frontend_bus_axi4_0_ar_bits_id(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_id),
    .l2_frontend_bus_axi4_0_ar_bits_addr(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_addr),
    .l2_frontend_bus_axi4_0_ar_bits_len(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_len),
    .l2_frontend_bus_axi4_0_ar_bits_size(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_size),
    .l2_frontend_bus_axi4_0_ar_bits_burst(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_burst),
    .l2_frontend_bus_axi4_0_ar_bits_lock(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_lock),
    .l2_frontend_bus_axi4_0_ar_bits_cache(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_cache),
    .l2_frontend_bus_axi4_0_ar_bits_prot(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_prot),
    .l2_frontend_bus_axi4_0_ar_bits_qos(ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_qos),
    .l2_frontend_bus_axi4_0_r_ready(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_ready),
    .l2_frontend_bus_axi4_0_r_valid(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_valid),
    .l2_frontend_bus_axi4_0_r_bits_id(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_id),
    .l2_frontend_bus_axi4_0_r_bits_data(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_data),
    .l2_frontend_bus_axi4_0_r_bits_resp(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_resp),
    .l2_frontend_bus_axi4_0_r_bits_last(ExampleBoomSystem_l2_frontend_bus_axi4_0_r_bits_last)
  );
  SimAXIMem SimAXIMem (
    .clock(SimAXIMem_clock),
    .reset(SimAXIMem_reset),
    .io_axi4_0_aw_ready(SimAXIMem_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(SimAXIMem_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(SimAXIMem_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(SimAXIMem_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(SimAXIMem_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(SimAXIMem_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(SimAXIMem_io_axi4_0_aw_bits_burst),
    .io_axi4_0_w_ready(SimAXIMem_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(SimAXIMem_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(SimAXIMem_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(SimAXIMem_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(SimAXIMem_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(SimAXIMem_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(SimAXIMem_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(SimAXIMem_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(SimAXIMem_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(SimAXIMem_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(SimAXIMem_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(SimAXIMem_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(SimAXIMem_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(SimAXIMem_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(SimAXIMem_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(SimAXIMem_io_axi4_0_ar_bits_burst),
    .io_axi4_0_r_ready(SimAXIMem_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(SimAXIMem_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(SimAXIMem_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(SimAXIMem_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(SimAXIMem_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(SimAXIMem_io_axi4_0_r_bits_last)
  );
  SimAXIMem_1 SimAXIMem_1 (
    .clock(SimAXIMem_1_clock),
    .reset(SimAXIMem_1_reset),
    .io_axi4_0_aw_ready(SimAXIMem_1_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(SimAXIMem_1_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(SimAXIMem_1_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(SimAXIMem_1_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(SimAXIMem_1_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(SimAXIMem_1_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(SimAXIMem_1_io_axi4_0_aw_bits_burst),
    .io_axi4_0_w_ready(SimAXIMem_1_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(SimAXIMem_1_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(SimAXIMem_1_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(SimAXIMem_1_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(SimAXIMem_1_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(SimAXIMem_1_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(SimAXIMem_1_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(SimAXIMem_1_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(SimAXIMem_1_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(SimAXIMem_1_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(SimAXIMem_1_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(SimAXIMem_1_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(SimAXIMem_1_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(SimAXIMem_1_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(SimAXIMem_1_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(SimAXIMem_1_io_axi4_0_ar_bits_burst),
    .io_axi4_0_r_ready(SimAXIMem_1_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(SimAXIMem_1_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(SimAXIMem_1_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(SimAXIMem_1_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(SimAXIMem_1_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(SimAXIMem_1_io_axi4_0_r_bits_last)
  );
  SimDTM SimDTM (
    .exit(SimDTM_exit),
    .debug_req_ready(SimDTM_debug_req_ready),
    .debug_req_valid(SimDTM_debug_req_valid),
    .debug_req_bits_addr(SimDTM_debug_req_bits_addr),
    .debug_req_bits_data(SimDTM_debug_req_bits_data),
    .debug_req_bits_op(SimDTM_debug_req_bits_op),
    .debug_resp_ready(SimDTM_debug_resp_ready),
    .debug_resp_valid(SimDTM_debug_resp_valid),
    .debug_resp_bits_data(SimDTM_debug_resp_bits_data),
    .debug_resp_bits_resp(SimDTM_debug_resp_bits_resp),
    .reset(SimDTM_reset),
    .clk(SimDTM_clk)
  );
  assign _T_180 = reset | ExampleBoomSystem_debug_ndreset;
  assign _T_197 = SimDTM_exit == 32'h1;
  assign _T_199 = SimDTM_exit >= 32'h2;
  assign _T_201 = SimDTM_exit >> 1'h1;
  assign _T_204 = reset == 1'h0;
  assign io_success = _T_197;
  assign ExampleBoomSystem_clock = clock;
  assign ExampleBoomSystem_reset = _T_180;
  assign ExampleBoomSystem_debug_clockeddmi_dmi_req_valid = SimDTM_debug_req_valid;
  assign ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_addr = SimDTM_debug_req_bits_addr;
  assign ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_data = SimDTM_debug_req_bits_data;
  assign ExampleBoomSystem_debug_clockeddmi_dmi_req_bits_op = SimDTM_debug_req_bits_op;
  assign ExampleBoomSystem_debug_clockeddmi_dmi_resp_ready = SimDTM_debug_resp_ready;
  assign ExampleBoomSystem_debug_clockeddmi_dmiClock = clock;
  assign ExampleBoomSystem_debug_clockeddmi_dmiReset = reset;
  assign ExampleBoomSystem_interrupts = 2'h0;
  assign ExampleBoomSystem_mem_axi4_0_aw_ready = SimAXIMem_io_axi4_0_aw_ready;
  assign ExampleBoomSystem_mem_axi4_0_w_ready = SimAXIMem_io_axi4_0_w_ready;
  assign ExampleBoomSystem_mem_axi4_0_b_valid = SimAXIMem_io_axi4_0_b_valid;
  assign ExampleBoomSystem_mem_axi4_0_b_bits_id = SimAXIMem_io_axi4_0_b_bits_id;
  assign ExampleBoomSystem_mem_axi4_0_b_bits_resp = SimAXIMem_io_axi4_0_b_bits_resp;
  assign ExampleBoomSystem_mem_axi4_0_ar_ready = SimAXIMem_io_axi4_0_ar_ready;
  assign ExampleBoomSystem_mem_axi4_0_r_valid = SimAXIMem_io_axi4_0_r_valid;
  assign ExampleBoomSystem_mem_axi4_0_r_bits_id = SimAXIMem_io_axi4_0_r_bits_id;
  assign ExampleBoomSystem_mem_axi4_0_r_bits_data = SimAXIMem_io_axi4_0_r_bits_data;
  assign ExampleBoomSystem_mem_axi4_0_r_bits_resp = SimAXIMem_io_axi4_0_r_bits_resp;
  assign ExampleBoomSystem_mem_axi4_0_r_bits_last = SimAXIMem_io_axi4_0_r_bits_last;
  assign ExampleBoomSystem_mmio_axi4_0_aw_ready = SimAXIMem_1_io_axi4_0_aw_ready;
  assign ExampleBoomSystem_mmio_axi4_0_w_ready = SimAXIMem_1_io_axi4_0_w_ready;
  assign ExampleBoomSystem_mmio_axi4_0_b_valid = SimAXIMem_1_io_axi4_0_b_valid;
  assign ExampleBoomSystem_mmio_axi4_0_b_bits_id = SimAXIMem_1_io_axi4_0_b_bits_id;
  assign ExampleBoomSystem_mmio_axi4_0_b_bits_resp = SimAXIMem_1_io_axi4_0_b_bits_resp;
  assign ExampleBoomSystem_mmio_axi4_0_ar_ready = SimAXIMem_1_io_axi4_0_ar_ready;
  assign ExampleBoomSystem_mmio_axi4_0_r_valid = SimAXIMem_1_io_axi4_0_r_valid;
  assign ExampleBoomSystem_mmio_axi4_0_r_bits_id = SimAXIMem_1_io_axi4_0_r_bits_id;
  assign ExampleBoomSystem_mmio_axi4_0_r_bits_data = SimAXIMem_1_io_axi4_0_r_bits_data;
  assign ExampleBoomSystem_mmio_axi4_0_r_bits_resp = SimAXIMem_1_io_axi4_0_r_bits_resp;
  assign ExampleBoomSystem_mmio_axi4_0_r_bits_last = SimAXIMem_1_io_axi4_0_r_bits_last;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_valid = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_id = 8'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_addr = 32'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_len = 8'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_size = 3'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_burst = 2'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_lock = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_cache = 4'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_prot = 3'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_aw_bits_qos = 4'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_w_valid = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_data = 64'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_strb = 8'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_w_bits_last = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_b_ready = 1'h1;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_valid = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_id = 8'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_addr = 32'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_len = 8'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_size = 3'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_burst = 2'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_lock = 1'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_cache = 4'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_prot = 3'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_ar_bits_qos = 4'h0;
  assign ExampleBoomSystem_l2_frontend_bus_axi4_0_r_ready = 1'h1;
  assign SimAXIMem_clock = clock;
  assign SimAXIMem_reset = reset;
  assign SimAXIMem_io_axi4_0_aw_valid = ExampleBoomSystem_mem_axi4_0_aw_valid;
  assign SimAXIMem_io_axi4_0_aw_bits_id = ExampleBoomSystem_mem_axi4_0_aw_bits_id;
  assign SimAXIMem_io_axi4_0_aw_bits_addr = ExampleBoomSystem_mem_axi4_0_aw_bits_addr[27:0];
  assign SimAXIMem_io_axi4_0_aw_bits_len = ExampleBoomSystem_mem_axi4_0_aw_bits_len;
  assign SimAXIMem_io_axi4_0_aw_bits_size = ExampleBoomSystem_mem_axi4_0_aw_bits_size;
  assign SimAXIMem_io_axi4_0_aw_bits_burst = ExampleBoomSystem_mem_axi4_0_aw_bits_burst;
  assign SimAXIMem_io_axi4_0_w_valid = ExampleBoomSystem_mem_axi4_0_w_valid;
  assign SimAXIMem_io_axi4_0_w_bits_data = ExampleBoomSystem_mem_axi4_0_w_bits_data;
  assign SimAXIMem_io_axi4_0_w_bits_strb = ExampleBoomSystem_mem_axi4_0_w_bits_strb;
  assign SimAXIMem_io_axi4_0_w_bits_last = ExampleBoomSystem_mem_axi4_0_w_bits_last;
  assign SimAXIMem_io_axi4_0_b_ready = ExampleBoomSystem_mem_axi4_0_b_ready;
  assign SimAXIMem_io_axi4_0_ar_valid = ExampleBoomSystem_mem_axi4_0_ar_valid;
  assign SimAXIMem_io_axi4_0_ar_bits_id = ExampleBoomSystem_mem_axi4_0_ar_bits_id;
  assign SimAXIMem_io_axi4_0_ar_bits_addr = ExampleBoomSystem_mem_axi4_0_ar_bits_addr[27:0];
  assign SimAXIMem_io_axi4_0_ar_bits_len = ExampleBoomSystem_mem_axi4_0_ar_bits_len;
  assign SimAXIMem_io_axi4_0_ar_bits_size = ExampleBoomSystem_mem_axi4_0_ar_bits_size;
  assign SimAXIMem_io_axi4_0_ar_bits_burst = ExampleBoomSystem_mem_axi4_0_ar_bits_burst;
  assign SimAXIMem_io_axi4_0_r_ready = ExampleBoomSystem_mem_axi4_0_r_ready;
  assign SimAXIMem_1_clock = clock;
  assign SimAXIMem_1_reset = reset;
  assign SimAXIMem_1_io_axi4_0_aw_valid = ExampleBoomSystem_mmio_axi4_0_aw_valid;
  assign SimAXIMem_1_io_axi4_0_aw_bits_id = ExampleBoomSystem_mmio_axi4_0_aw_bits_id;
  assign SimAXIMem_1_io_axi4_0_aw_bits_addr = ExampleBoomSystem_mmio_axi4_0_aw_bits_addr[11:0];
  assign SimAXIMem_1_io_axi4_0_aw_bits_len = ExampleBoomSystem_mmio_axi4_0_aw_bits_len;
  assign SimAXIMem_1_io_axi4_0_aw_bits_size = ExampleBoomSystem_mmio_axi4_0_aw_bits_size;
  assign SimAXIMem_1_io_axi4_0_aw_bits_burst = ExampleBoomSystem_mmio_axi4_0_aw_bits_burst;
  assign SimAXIMem_1_io_axi4_0_w_valid = ExampleBoomSystem_mmio_axi4_0_w_valid;
  assign SimAXIMem_1_io_axi4_0_w_bits_data = ExampleBoomSystem_mmio_axi4_0_w_bits_data;
  assign SimAXIMem_1_io_axi4_0_w_bits_strb = ExampleBoomSystem_mmio_axi4_0_w_bits_strb;
  assign SimAXIMem_1_io_axi4_0_w_bits_last = ExampleBoomSystem_mmio_axi4_0_w_bits_last;
  assign SimAXIMem_1_io_axi4_0_b_ready = ExampleBoomSystem_mmio_axi4_0_b_ready;
  assign SimAXIMem_1_io_axi4_0_ar_valid = ExampleBoomSystem_mmio_axi4_0_ar_valid;
  assign SimAXIMem_1_io_axi4_0_ar_bits_id = ExampleBoomSystem_mmio_axi4_0_ar_bits_id;
  assign SimAXIMem_1_io_axi4_0_ar_bits_addr = ExampleBoomSystem_mmio_axi4_0_ar_bits_addr[11:0];
  assign SimAXIMem_1_io_axi4_0_ar_bits_len = ExampleBoomSystem_mmio_axi4_0_ar_bits_len;
  assign SimAXIMem_1_io_axi4_0_ar_bits_size = ExampleBoomSystem_mmio_axi4_0_ar_bits_size;
  assign SimAXIMem_1_io_axi4_0_ar_bits_burst = ExampleBoomSystem_mmio_axi4_0_ar_bits_burst;
  assign SimAXIMem_1_io_axi4_0_r_ready = ExampleBoomSystem_mmio_axi4_0_r_ready;
  assign SimDTM_debug_req_ready = ExampleBoomSystem_debug_clockeddmi_dmi_req_ready;
  assign SimDTM_debug_resp_valid = ExampleBoomSystem_debug_clockeddmi_dmi_resp_valid;
  assign SimDTM_debug_resp_bits_data = ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_data;
  assign SimDTM_debug_resp_bits_resp = ExampleBoomSystem_debug_clockeddmi_dmi_resp_bits_resp;
  assign SimDTM_reset = reset;
  assign SimDTM_clk = clock;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_199 & _T_204) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_201);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_199 & _T_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
