module trivial2a( input a, output c, output d);
assign c = ~a;
assign d = a;
endmodule

