module tup_out1 (
  output [1:0] out_a
  output [2:0] out_b
);

  assign out_a = 2'h1;
  assign out_b = 3'h2;

endmodule
