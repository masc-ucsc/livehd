module PMPChecker_1(
  input         clock,
  input         reset,
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_res,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_res,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_res,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_res,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_res,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_res,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_res,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_res,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  input  [1:0]  io_size,
  output        io_r,
  output        io_w,
  output        io_x
);
  wire  default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  wire [5:0] _T_3 = 6'h7 << io_size; // @[package.scala 189:77]
  wire [2:0] _T_5 = ~_T_3[2:0]; // @[package.scala 189:46]
  wire [31:0] _GEN_0 = {{29'd0}, _T_5}; // @[PMP.scala 70:26]
  wire [31:0] _T_6 = io_pmp_7_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [31:0] _T_8 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_9 = ~_T_8; // @[PMP.scala 62:29]
  wire [31:0] _T_10 = _T_9 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_11 = ~_T_10; // @[PMP.scala 62:27]
  wire [28:0] _T_14 = io_addr[31:3] ^ _T_11[31:3]; // @[PMP.scala 65:47]
  wire [28:0] _T_15 = ~io_pmp_7_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_16 = _T_14 & _T_15; // @[PMP.scala 65:52]
  wire  _T_17 = _T_16 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_25 = io_addr[2:0] ^ _T_11[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_26 = ~_T_6[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_27 = _T_25 & _T_26; // @[PMP.scala 65:52]
  wire  _T_28 = _T_27 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_29 = _T_17 & _T_28; // @[PMP.scala 73:16]
  wire [31:0] _T_36 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_37 = ~_T_36; // @[PMP.scala 62:29]
  wire [31:0] _T_38 = _T_37 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_39 = ~_T_38; // @[PMP.scala 62:27]
  wire  _T_41 = io_addr[31:3] < _T_39[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_48 = io_addr[31:3] ^ _T_39[31:3]; // @[PMP.scala 83:41]
  wire  _T_49 = _T_48 == 29'h0; // @[PMP.scala 83:69]
  wire [2:0] _T_51 = io_addr[2:0] | _T_5; // @[PMP.scala 84:42]
  wire  _T_57 = _T_51 < _T_39[2:0]; // @[PMP.scala 84:53]
  wire  _T_59 = _T_41 | _T_49 & _T_57; // @[PMP.scala 85:16]
  wire  _T_60 = ~_T_59; // @[PMP.scala 90:5]
  wire  _T_67 = io_addr[31:3] < _T_11[31:3]; // @[PMP.scala 82:39]
  wire  _T_75 = _T_14 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_83 = io_addr[2:0] < _T_11[2:0]; // @[PMP.scala 84:53]
  wire  _T_85 = _T_67 | _T_75 & _T_83; // @[PMP.scala 85:16]
  wire  _T_86 = _T_60 & _T_85; // @[PMP.scala 96:48]
  wire  _T_88 = io_pmp_7_cfg_a[1] ? _T_29 : io_pmp_7_cfg_a[0] & _T_86; // @[PMP.scala 134:8]
  wire  _T_90 = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_109 = ~io_addr[2:0]; // @[PMP.scala 125:125]
  wire [2:0] _T_110 = _T_39[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_112 = _T_49 & _T_110 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_128 = _T_11[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_130 = _T_75 & _T_128 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_132 = ~(_T_112 | _T_130); // @[PMP.scala 127:24]
  wire [2:0] _T_134 = ~io_pmp_7_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_135 = _T_5 & _T_134; // @[PMP.scala 128:32]
  wire  _T_136 = _T_135 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_138 = io_pmp_7_cfg_a[1] ? _T_136 : _T_132; // @[PMP.scala 129:8]
  wire  _T_191 = _T_138 & (io_pmp_7_cfg_r | _T_90); // @[PMP.scala 183:26]
  wire  _T_193 = _T_138 & (io_pmp_7_cfg_w | _T_90); // @[PMP.scala 184:26]
  wire  _T_195 = _T_138 & (io_pmp_7_cfg_x | _T_90); // @[PMP.scala 185:26]
  wire  _T_196_cfg_x = _T_88 ? _T_195 : default_; // @[PMP.scala 186:8]
  wire  _T_196_cfg_w = _T_88 ? _T_193 : default_; // @[PMP.scala 186:8]
  wire  _T_196_cfg_r = _T_88 ? _T_191 : default_; // @[PMP.scala 186:8]
  wire [31:0] _T_202 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_211 = ~io_pmp_6_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_212 = _T_48 & _T_211; // @[PMP.scala 65:52]
  wire  _T_213 = _T_212 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_221 = io_addr[2:0] ^ _T_39[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_222 = ~_T_202[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_223 = _T_221 & _T_222; // @[PMP.scala 65:52]
  wire  _T_224 = _T_223 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_225 = _T_213 & _T_224; // @[PMP.scala 73:16]
  wire [31:0] _T_232 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_233 = ~_T_232; // @[PMP.scala 62:29]
  wire [31:0] _T_234 = _T_233 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_235 = ~_T_234; // @[PMP.scala 62:27]
  wire  _T_237 = io_addr[31:3] < _T_235[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_244 = io_addr[31:3] ^ _T_235[31:3]; // @[PMP.scala 83:41]
  wire  _T_245 = _T_244 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_253 = _T_51 < _T_235[2:0]; // @[PMP.scala 84:53]
  wire  _T_255 = _T_237 | _T_245 & _T_253; // @[PMP.scala 85:16]
  wire  _T_256 = ~_T_255; // @[PMP.scala 90:5]
  wire  _T_279 = io_addr[2:0] < _T_39[2:0]; // @[PMP.scala 84:53]
  wire  _T_281 = _T_41 | _T_49 & _T_279; // @[PMP.scala 85:16]
  wire  _T_282 = _T_256 & _T_281; // @[PMP.scala 96:48]
  wire  _T_284 = io_pmp_6_cfg_a[1] ? _T_225 : io_pmp_6_cfg_a[0] & _T_282; // @[PMP.scala 134:8]
  wire  _T_286 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_306 = _T_235[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_308 = _T_245 & _T_306 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_324 = _T_39[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_326 = _T_49 & _T_324 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_328 = ~(_T_308 | _T_326); // @[PMP.scala 127:24]
  wire [2:0] _T_330 = ~io_pmp_6_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_331 = _T_5 & _T_330; // @[PMP.scala 128:32]
  wire  _T_332 = _T_331 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_334 = io_pmp_6_cfg_a[1] ? _T_332 : _T_328; // @[PMP.scala 129:8]
  wire  _T_387 = _T_334 & (io_pmp_6_cfg_r | _T_286); // @[PMP.scala 183:26]
  wire  _T_389 = _T_334 & (io_pmp_6_cfg_w | _T_286); // @[PMP.scala 184:26]
  wire  _T_391 = _T_334 & (io_pmp_6_cfg_x | _T_286); // @[PMP.scala 185:26]
  wire  _T_392_cfg_x = _T_284 ? _T_391 : _T_196_cfg_x; // @[PMP.scala 186:8]
  wire  _T_392_cfg_w = _T_284 ? _T_389 : _T_196_cfg_w; // @[PMP.scala 186:8]
  wire  _T_392_cfg_r = _T_284 ? _T_387 : _T_196_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_398 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_407 = ~io_pmp_5_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_408 = _T_244 & _T_407; // @[PMP.scala 65:52]
  wire  _T_409 = _T_408 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_417 = io_addr[2:0] ^ _T_235[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_418 = ~_T_398[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_419 = _T_417 & _T_418; // @[PMP.scala 65:52]
  wire  _T_420 = _T_419 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_421 = _T_409 & _T_420; // @[PMP.scala 73:16]
  wire [31:0] _T_428 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_429 = ~_T_428; // @[PMP.scala 62:29]
  wire [31:0] _T_430 = _T_429 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_431 = ~_T_430; // @[PMP.scala 62:27]
  wire  _T_433 = io_addr[31:3] < _T_431[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_440 = io_addr[31:3] ^ _T_431[31:3]; // @[PMP.scala 83:41]
  wire  _T_441 = _T_440 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_449 = _T_51 < _T_431[2:0]; // @[PMP.scala 84:53]
  wire  _T_451 = _T_433 | _T_441 & _T_449; // @[PMP.scala 85:16]
  wire  _T_452 = ~_T_451; // @[PMP.scala 90:5]
  wire  _T_475 = io_addr[2:0] < _T_235[2:0]; // @[PMP.scala 84:53]
  wire  _T_477 = _T_237 | _T_245 & _T_475; // @[PMP.scala 85:16]
  wire  _T_478 = _T_452 & _T_477; // @[PMP.scala 96:48]
  wire  _T_480 = io_pmp_5_cfg_a[1] ? _T_421 : io_pmp_5_cfg_a[0] & _T_478; // @[PMP.scala 134:8]
  wire  _T_482 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_502 = _T_431[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_504 = _T_441 & _T_502 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_520 = _T_235[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_522 = _T_245 & _T_520 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_524 = ~(_T_504 | _T_522); // @[PMP.scala 127:24]
  wire [2:0] _T_526 = ~io_pmp_5_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_527 = _T_5 & _T_526; // @[PMP.scala 128:32]
  wire  _T_528 = _T_527 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_530 = io_pmp_5_cfg_a[1] ? _T_528 : _T_524; // @[PMP.scala 129:8]
  wire  _T_583 = _T_530 & (io_pmp_5_cfg_r | _T_482); // @[PMP.scala 183:26]
  wire  _T_585 = _T_530 & (io_pmp_5_cfg_w | _T_482); // @[PMP.scala 184:26]
  wire  _T_587 = _T_530 & (io_pmp_5_cfg_x | _T_482); // @[PMP.scala 185:26]
  wire  _T_588_cfg_x = _T_480 ? _T_587 : _T_392_cfg_x; // @[PMP.scala 186:8]
  wire  _T_588_cfg_w = _T_480 ? _T_585 : _T_392_cfg_w; // @[PMP.scala 186:8]
  wire  _T_588_cfg_r = _T_480 ? _T_583 : _T_392_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_594 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_603 = ~io_pmp_4_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_604 = _T_440 & _T_603; // @[PMP.scala 65:52]
  wire  _T_605 = _T_604 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_613 = io_addr[2:0] ^ _T_431[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_614 = ~_T_594[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_615 = _T_613 & _T_614; // @[PMP.scala 65:52]
  wire  _T_616 = _T_615 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_617 = _T_605 & _T_616; // @[PMP.scala 73:16]
  wire [31:0] _T_624 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_625 = ~_T_624; // @[PMP.scala 62:29]
  wire [31:0] _T_626 = _T_625 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_627 = ~_T_626; // @[PMP.scala 62:27]
  wire  _T_629 = io_addr[31:3] < _T_627[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_636 = io_addr[31:3] ^ _T_627[31:3]; // @[PMP.scala 83:41]
  wire  _T_637 = _T_636 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_645 = _T_51 < _T_627[2:0]; // @[PMP.scala 84:53]
  wire  _T_647 = _T_629 | _T_637 & _T_645; // @[PMP.scala 85:16]
  wire  _T_648 = ~_T_647; // @[PMP.scala 90:5]
  wire  _T_671 = io_addr[2:0] < _T_431[2:0]; // @[PMP.scala 84:53]
  wire  _T_673 = _T_433 | _T_441 & _T_671; // @[PMP.scala 85:16]
  wire  _T_674 = _T_648 & _T_673; // @[PMP.scala 96:48]
  wire  _T_676 = io_pmp_4_cfg_a[1] ? _T_617 : io_pmp_4_cfg_a[0] & _T_674; // @[PMP.scala 134:8]
  wire  _T_678 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_698 = _T_627[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_700 = _T_637 & _T_698 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_716 = _T_431[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_718 = _T_441 & _T_716 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_720 = ~(_T_700 | _T_718); // @[PMP.scala 127:24]
  wire [2:0] _T_722 = ~io_pmp_4_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_723 = _T_5 & _T_722; // @[PMP.scala 128:32]
  wire  _T_724 = _T_723 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_726 = io_pmp_4_cfg_a[1] ? _T_724 : _T_720; // @[PMP.scala 129:8]
  wire  _T_779 = _T_726 & (io_pmp_4_cfg_r | _T_678); // @[PMP.scala 183:26]
  wire  _T_781 = _T_726 & (io_pmp_4_cfg_w | _T_678); // @[PMP.scala 184:26]
  wire  _T_783 = _T_726 & (io_pmp_4_cfg_x | _T_678); // @[PMP.scala 185:26]
  wire  _T_784_cfg_x = _T_676 ? _T_783 : _T_588_cfg_x; // @[PMP.scala 186:8]
  wire  _T_784_cfg_w = _T_676 ? _T_781 : _T_588_cfg_w; // @[PMP.scala 186:8]
  wire  _T_784_cfg_r = _T_676 ? _T_779 : _T_588_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_790 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_799 = ~io_pmp_3_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_800 = _T_636 & _T_799; // @[PMP.scala 65:52]
  wire  _T_801 = _T_800 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_809 = io_addr[2:0] ^ _T_627[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_810 = ~_T_790[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_811 = _T_809 & _T_810; // @[PMP.scala 65:52]
  wire  _T_812 = _T_811 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_813 = _T_801 & _T_812; // @[PMP.scala 73:16]
  wire [31:0] _T_820 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_821 = ~_T_820; // @[PMP.scala 62:29]
  wire [31:0] _T_822 = _T_821 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_823 = ~_T_822; // @[PMP.scala 62:27]
  wire  _T_825 = io_addr[31:3] < _T_823[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_832 = io_addr[31:3] ^ _T_823[31:3]; // @[PMP.scala 83:41]
  wire  _T_833 = _T_832 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_841 = _T_51 < _T_823[2:0]; // @[PMP.scala 84:53]
  wire  _T_843 = _T_825 | _T_833 & _T_841; // @[PMP.scala 85:16]
  wire  _T_844 = ~_T_843; // @[PMP.scala 90:5]
  wire  _T_867 = io_addr[2:0] < _T_627[2:0]; // @[PMP.scala 84:53]
  wire  _T_869 = _T_629 | _T_637 & _T_867; // @[PMP.scala 85:16]
  wire  _T_870 = _T_844 & _T_869; // @[PMP.scala 96:48]
  wire  _T_872 = io_pmp_3_cfg_a[1] ? _T_813 : io_pmp_3_cfg_a[0] & _T_870; // @[PMP.scala 134:8]
  wire  _T_874 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_894 = _T_823[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_896 = _T_833 & _T_894 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_912 = _T_627[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_914 = _T_637 & _T_912 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_916 = ~(_T_896 | _T_914); // @[PMP.scala 127:24]
  wire [2:0] _T_918 = ~io_pmp_3_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_919 = _T_5 & _T_918; // @[PMP.scala 128:32]
  wire  _T_920 = _T_919 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_922 = io_pmp_3_cfg_a[1] ? _T_920 : _T_916; // @[PMP.scala 129:8]
  wire  _T_975 = _T_922 & (io_pmp_3_cfg_r | _T_874); // @[PMP.scala 183:26]
  wire  _T_977 = _T_922 & (io_pmp_3_cfg_w | _T_874); // @[PMP.scala 184:26]
  wire  _T_979 = _T_922 & (io_pmp_3_cfg_x | _T_874); // @[PMP.scala 185:26]
  wire  _T_980_cfg_x = _T_872 ? _T_979 : _T_784_cfg_x; // @[PMP.scala 186:8]
  wire  _T_980_cfg_w = _T_872 ? _T_977 : _T_784_cfg_w; // @[PMP.scala 186:8]
  wire  _T_980_cfg_r = _T_872 ? _T_975 : _T_784_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_986 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_995 = ~io_pmp_2_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_996 = _T_832 & _T_995; // @[PMP.scala 65:52]
  wire  _T_997 = _T_996 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1005 = io_addr[2:0] ^ _T_823[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1006 = ~_T_986[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1007 = _T_1005 & _T_1006; // @[PMP.scala 65:52]
  wire  _T_1008 = _T_1007 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1009 = _T_997 & _T_1008; // @[PMP.scala 73:16]
  wire [31:0] _T_1016 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_1017 = ~_T_1016; // @[PMP.scala 62:29]
  wire [31:0] _T_1018 = _T_1017 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_1019 = ~_T_1018; // @[PMP.scala 62:27]
  wire  _T_1021 = io_addr[31:3] < _T_1019[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_1028 = io_addr[31:3] ^ _T_1019[31:3]; // @[PMP.scala 83:41]
  wire  _T_1029 = _T_1028 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_1037 = _T_51 < _T_1019[2:0]; // @[PMP.scala 84:53]
  wire  _T_1039 = _T_1021 | _T_1029 & _T_1037; // @[PMP.scala 85:16]
  wire  _T_1040 = ~_T_1039; // @[PMP.scala 90:5]
  wire  _T_1063 = io_addr[2:0] < _T_823[2:0]; // @[PMP.scala 84:53]
  wire  _T_1065 = _T_825 | _T_833 & _T_1063; // @[PMP.scala 85:16]
  wire  _T_1066 = _T_1040 & _T_1065; // @[PMP.scala 96:48]
  wire  _T_1068 = io_pmp_2_cfg_a[1] ? _T_1009 : io_pmp_2_cfg_a[0] & _T_1066; // @[PMP.scala 134:8]
  wire  _T_1070 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1090 = _T_1019[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_1092 = _T_1029 & _T_1090 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_1108 = _T_823[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1110 = _T_833 & _T_1108 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1112 = ~(_T_1092 | _T_1110); // @[PMP.scala 127:24]
  wire [2:0] _T_1114 = ~io_pmp_2_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1115 = _T_5 & _T_1114; // @[PMP.scala 128:32]
  wire  _T_1116 = _T_1115 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1118 = io_pmp_2_cfg_a[1] ? _T_1116 : _T_1112; // @[PMP.scala 129:8]
  wire  _T_1171 = _T_1118 & (io_pmp_2_cfg_r | _T_1070); // @[PMP.scala 183:26]
  wire  _T_1173 = _T_1118 & (io_pmp_2_cfg_w | _T_1070); // @[PMP.scala 184:26]
  wire  _T_1175 = _T_1118 & (io_pmp_2_cfg_x | _T_1070); // @[PMP.scala 185:26]
  wire  _T_1176_cfg_x = _T_1068 ? _T_1175 : _T_980_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_w = _T_1068 ? _T_1173 : _T_980_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1176_cfg_r = _T_1068 ? _T_1171 : _T_980_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1182 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_1191 = ~io_pmp_1_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_1192 = _T_1028 & _T_1191; // @[PMP.scala 65:52]
  wire  _T_1193 = _T_1192 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1201 = io_addr[2:0] ^ _T_1019[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1202 = ~_T_1182[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1203 = _T_1201 & _T_1202; // @[PMP.scala 65:52]
  wire  _T_1204 = _T_1203 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1205 = _T_1193 & _T_1204; // @[PMP.scala 73:16]
  wire [31:0] _T_1212 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  wire [31:0] _T_1213 = ~_T_1212; // @[PMP.scala 62:29]
  wire [31:0] _T_1214 = _T_1213 | 32'h3; // @[PMP.scala 62:48]
  wire [31:0] _T_1215 = ~_T_1214; // @[PMP.scala 62:27]
  wire  _T_1217 = io_addr[31:3] < _T_1215[31:3]; // @[PMP.scala 82:39]
  wire [28:0] _T_1224 = io_addr[31:3] ^ _T_1215[31:3]; // @[PMP.scala 83:41]
  wire  _T_1225 = _T_1224 == 29'h0; // @[PMP.scala 83:69]
  wire  _T_1233 = _T_51 < _T_1215[2:0]; // @[PMP.scala 84:53]
  wire  _T_1235 = _T_1217 | _T_1225 & _T_1233; // @[PMP.scala 85:16]
  wire  _T_1236 = ~_T_1235; // @[PMP.scala 90:5]
  wire  _T_1259 = io_addr[2:0] < _T_1019[2:0]; // @[PMP.scala 84:53]
  wire  _T_1261 = _T_1021 | _T_1029 & _T_1259; // @[PMP.scala 85:16]
  wire  _T_1262 = _T_1236 & _T_1261; // @[PMP.scala 96:48]
  wire  _T_1264 = io_pmp_1_cfg_a[1] ? _T_1205 : io_pmp_1_cfg_a[0] & _T_1262; // @[PMP.scala 134:8]
  wire  _T_1266 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1286 = _T_1215[2:0] & _T_109; // @[PMP.scala 125:123]
  wire  _T_1288 = _T_1225 & _T_1286 != 3'h0; // @[PMP.scala 125:88]
  wire [2:0] _T_1304 = _T_1019[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1306 = _T_1029 & _T_1304 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1308 = ~(_T_1288 | _T_1306); // @[PMP.scala 127:24]
  wire [2:0] _T_1310 = ~io_pmp_1_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1311 = _T_5 & _T_1310; // @[PMP.scala 128:32]
  wire  _T_1312 = _T_1311 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1314 = io_pmp_1_cfg_a[1] ? _T_1312 : _T_1308; // @[PMP.scala 129:8]
  wire  _T_1367 = _T_1314 & (io_pmp_1_cfg_r | _T_1266); // @[PMP.scala 183:26]
  wire  _T_1369 = _T_1314 & (io_pmp_1_cfg_w | _T_1266); // @[PMP.scala 184:26]
  wire  _T_1371 = _T_1314 & (io_pmp_1_cfg_x | _T_1266); // @[PMP.scala 185:26]
  wire  _T_1372_cfg_x = _T_1264 ? _T_1371 : _T_1176_cfg_x; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_w = _T_1264 ? _T_1369 : _T_1176_cfg_w; // @[PMP.scala 186:8]
  wire  _T_1372_cfg_r = _T_1264 ? _T_1367 : _T_1176_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _T_1378 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 70:26]
  wire [28:0] _T_1387 = ~io_pmp_0_mask[31:3]; // @[PMP.scala 65:54]
  wire [28:0] _T_1388 = _T_1224 & _T_1387; // @[PMP.scala 65:52]
  wire  _T_1389 = _T_1388 == 29'h0; // @[PMP.scala 65:58]
  wire [2:0] _T_1397 = io_addr[2:0] ^ _T_1215[2:0]; // @[PMP.scala 65:47]
  wire [2:0] _T_1398 = ~_T_1378[2:0]; // @[PMP.scala 65:54]
  wire [2:0] _T_1399 = _T_1397 & _T_1398; // @[PMP.scala 65:52]
  wire  _T_1400 = _T_1399 == 3'h0; // @[PMP.scala 65:58]
  wire  _T_1401 = _T_1389 & _T_1400; // @[PMP.scala 73:16]
  wire  _T_1455 = io_addr[2:0] < _T_1215[2:0]; // @[PMP.scala 84:53]
  wire  _T_1457 = _T_1217 | _T_1225 & _T_1455; // @[PMP.scala 85:16]
  wire  _T_1460 = io_pmp_0_cfg_a[1] ? _T_1401 : io_pmp_0_cfg_a[0] & _T_1457; // @[PMP.scala 134:8]
  wire  _T_1462 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  wire [2:0] _T_1500 = _T_1215[2:0] & _T_51; // @[PMP.scala 126:113]
  wire  _T_1502 = _T_1225 & _T_1500 != 3'h0; // @[PMP.scala 126:83]
  wire  _T_1504 = ~_T_1502; // @[PMP.scala 127:24]
  wire [2:0] _T_1506 = ~io_pmp_0_mask[2:0]; // @[PMP.scala 128:34]
  wire [2:0] _T_1507 = _T_5 & _T_1506; // @[PMP.scala 128:32]
  wire  _T_1508 = _T_1507 == 3'h0; // @[PMP.scala 128:57]
  wire  _T_1510 = io_pmp_0_cfg_a[1] ? _T_1508 : _T_1504; // @[PMP.scala 129:8]
  wire  _T_1563 = _T_1510 & (io_pmp_0_cfg_r | _T_1462); // @[PMP.scala 183:26]
  wire  _T_1565 = _T_1510 & (io_pmp_0_cfg_w | _T_1462); // @[PMP.scala 184:26]
  wire  _T_1567 = _T_1510 & (io_pmp_0_cfg_x | _T_1462); // @[PMP.scala 185:26]
  assign io_r = _T_1460 ? _T_1563 : _T_1372_cfg_r; // @[PMP.scala 186:8]
  assign io_w = _T_1460 ? _T_1565 : _T_1372_cfg_w; // @[PMP.scala 186:8]
  assign io_x = _T_1460 ? _T_1567 : _T_1372_cfg_x; // @[PMP.scala 186:8]
endmodule
