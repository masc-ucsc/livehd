module SnxnLv4Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 83028:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 83029:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 83030:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 83031:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 83032:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 83033:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 83034:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 83035:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 83036:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 83037:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 83038:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 83039:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 83040:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 83041:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 83042:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 83043:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 83044:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 83045:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 83046:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 83047:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 83048:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 83049:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 83050:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 83051:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 83052:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 83053:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 83054:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 83055:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 83056:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 83057:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 83058:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 83059:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 83060:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 83061:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 83062:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 83063:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 83064:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 83065:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 83066:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 83067:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 83068:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 83069:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 83070:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 83071:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 83072:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 83073:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 83074:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 83075:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 83076:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 83077:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 83078:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 83079:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 83080:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 83081:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 83082:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 83083:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 83084:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 83085:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 83086:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 83087:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 83088:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 83089:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 83090:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 83091:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 83092:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 83093:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 83094:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 83095:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 83096:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 83097:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 83098:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 83099:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 83100:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 83101:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 83102:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 83103:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 83104:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 83105:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 83106:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 83107:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 83108:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 83109:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 83110:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 83111:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 83112:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 83113:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 83114:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 83115:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 83116:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 83117:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 83118:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 83119:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 83120:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 83121:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 83122:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 83123:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 83124:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 83125:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 83126:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 83127:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 83128:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 83129:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 83130:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 83131:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 83132:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 83133:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 83134:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 83135:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 83136:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 83137:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 83138:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 83139:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 83140:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 83141:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 83142:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 83143:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 83144:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 83145:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 83146:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 83147:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 83148:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 83149:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 83150:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 83151:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 83152:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 83153:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 83154:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 83155:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 83156:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 83157:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 83158:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 83159:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 83160:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 83161:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 83162:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 83163:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 83164:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 83165:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 83166:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 83167:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 83168:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 83169:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 83170:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 83171:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 83172:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 83173:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 83174:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 83175:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 83176:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 83177:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 83178:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 83179:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 83180:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 83181:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 83182:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 83183:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 83184:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 83185:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 83186:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 83187:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 83188:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 83189:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 83190:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 83191:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 83192:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 83193:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 83194:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 83195:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 83196:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 83197:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 83198:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 83199:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 83200:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 83201:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 83202:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 83203:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 83204:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 83205:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 83206:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 83207:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 83208:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 83209:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 83210:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 83211:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 83212:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 83213:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 83214:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 83215:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 83216:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 83217:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 83218:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 83219:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 83220:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 83221:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 83222:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 83223:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 83224:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 83225:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 83226:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 83227:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 83228:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 83229:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 83230:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 83231:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 83232:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 83233:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 83234:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 83235:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 83236:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 83237:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 83238:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 83239:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 83240:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 83241:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 83242:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 83243:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 83244:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 83245:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 83246:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 83247:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 83248:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 83249:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 83250:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 83251:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 83252:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 83253:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 83254:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 83255:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 83256:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 83257:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 83258:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 83259:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 83260:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 83261:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 83262:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 83263:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 83264:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 83265:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 83266:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 83267:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 83268:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 83269:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 83270:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 83271:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 83272:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 83273:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 83274:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 83275:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 83276:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 83277:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 83278:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 83279:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 83280:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 83281:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 83282:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 83283:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 83284:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 83285:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 83286:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 83287:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 83288:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 83289:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 83290:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 83291:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 83292:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 83293:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 83294:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 83295:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 83296:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 83297:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 83298:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 83299:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 83300:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 83301:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 83302:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 83303:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 83304:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 83305:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 83306:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 83307:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 83308:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 83309:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 83310:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 83311:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 83312:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 83313:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 83314:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 83315:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 83316:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 83317:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 83318:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 83319:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 83320:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 83321:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 83322:20]
  assign io_z = ~x73; // @[Snxn100k.scala 83323:16]
endmodule
module SnxnLv4Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 83672:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 83673:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 83674:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 83675:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 83676:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 83677:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 83678:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 83679:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 83680:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 83681:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 83682:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 83683:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 83684:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 83685:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 83686:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 83687:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 83688:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 83689:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 83690:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 83691:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 83692:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 83693:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 83694:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 83695:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 83696:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 83697:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 83698:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 83699:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 83700:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 83701:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 83702:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 83703:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 83704:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 83705:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 83706:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 83707:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 83708:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 83709:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 83710:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 83711:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 83712:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 83713:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 83714:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 83715:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 83716:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 83717:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 83718:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 83719:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 83720:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 83721:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 83722:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 83723:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 83724:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 83725:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 83726:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 83727:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 83728:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 83729:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 83730:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 83731:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 83732:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 83733:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 83734:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 83735:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 83736:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 83737:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 83738:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 83739:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 83740:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 83741:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 83742:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 83743:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 83744:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 83745:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 83746:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 83747:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 83748:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 83749:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 83750:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 83751:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 83752:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 83753:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 83754:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 83755:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 83756:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 83757:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 83758:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 83759:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 83760:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 83761:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 83762:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 83763:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 83764:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 83765:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 83766:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 83767:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 83768:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 83769:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 83770:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 83771:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 83772:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 83773:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 83774:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 83775:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 83776:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 83777:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 83778:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 83779:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 83780:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 83781:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 83782:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 83783:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 83784:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 83785:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 83786:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 83787:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 83788:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 83789:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 83790:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 83791:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 83792:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 83793:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 83794:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 83795:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 83796:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 83797:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 83798:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 83799:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 83800:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 83801:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 83802:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 83803:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 83804:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 83805:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 83806:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 83807:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 83808:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 83809:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 83810:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 83811:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 83812:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 83813:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 83814:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 83815:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 83816:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 83817:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 83818:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 83819:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 83820:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 83821:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 83822:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 83823:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 83824:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 83825:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 83826:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 83827:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 83828:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 83829:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 83830:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 83831:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 83832:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 83833:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 83834:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 83835:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 83836:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 83837:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 83838:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 83839:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 83840:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 83841:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 83842:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 83843:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 83844:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 83845:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 83846:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 83847:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 83848:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 83849:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 83850:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 83851:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 83852:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 83853:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 83854:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 83855:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 83856:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 83857:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 83858:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 83859:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 83860:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 83861:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 83862:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 83863:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 83864:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 83865:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 83866:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 83867:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 83868:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 83869:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 83870:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 83871:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 83872:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 83873:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 83874:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 83875:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 83876:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 83877:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 83878:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 83879:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 83880:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 83881:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 83882:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 83883:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 83884:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 83885:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 83886:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 83887:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 83888:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 83889:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 83890:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 83891:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 83892:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 83893:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 83894:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 83895:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 83896:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 83897:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 83898:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 83899:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 83900:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 83901:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 83902:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 83903:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 83904:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 83905:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 83906:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 83907:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 83908:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 83909:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 83910:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 83911:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 83912:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 83913:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 83914:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 83915:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 83916:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 83917:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 83918:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 83919:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 83920:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 83921:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 83922:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 83923:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 83924:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 83925:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 83926:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 83927:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 83928:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 83929:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 83930:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 83931:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 83932:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 83933:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 83934:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 83935:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 83936:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 83937:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 83938:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 83939:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 83940:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 83941:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 83942:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 83943:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 83944:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 83945:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 83946:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 83947:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 83948:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 83949:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 83950:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 83951:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 83952:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 83953:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 83954:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 83955:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 83956:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 83957:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 83958:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 83959:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 83960:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 83961:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 83962:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 83963:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 83964:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 83965:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 83966:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 83967:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 83968:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 83969:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 83970:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 83971:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 83972:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 83973:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 83974:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 83975:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 83976:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 83977:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 83978:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 83979:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 83980:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 83981:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 83982:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 83983:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 83984:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 83985:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 83986:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 83987:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 83988:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 83989:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 83990:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 83991:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 83992:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 83993:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 83994:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 83995:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 83996:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 83997:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 83998:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 83999:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 84000:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 84001:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 84002:20]
  assign io_z = ~x82; // @[Snxn100k.scala 84003:16]
endmodule
module SnxnLv4Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 84014:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 84015:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 84016:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 84017:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 84018:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 84019:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 84020:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 84021:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 84022:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 84023:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 84024:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 84025:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 84026:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 84027:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 84028:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 84029:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 84030:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 84031:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 84032:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 84033:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 84034:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 84035:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 84036:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 84037:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 84038:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 84039:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 84040:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 84041:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 84042:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 84043:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 84044:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 84045:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 84046:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 84047:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 84048:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 84049:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 84050:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 84051:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 84052:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 84053:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 84054:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 84055:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 84056:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 84057:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 84058:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 84059:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 84060:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 84061:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 84062:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 84063:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 84064:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 84065:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 84066:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 84067:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 84068:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 84069:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 84070:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 84071:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 84072:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 84073:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 84074:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 84075:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 84076:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 84077:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 84078:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 84079:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 84080:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 84081:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 84082:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 84083:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 84084:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 84085:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 84086:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 84087:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 84088:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 84089:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 84090:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 84091:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 84092:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 84093:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 84094:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 84095:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 84096:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 84097:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 84098:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 84099:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 84100:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 84101:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 84102:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 84103:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 84104:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 84105:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 84106:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 84107:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 84108:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 84109:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 84110:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 84111:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 84112:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 84113:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 84114:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 84115:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 84116:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 84117:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 84118:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 84119:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 84120:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 84121:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 84122:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 84123:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 84124:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 84125:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 84126:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 84127:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 84128:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 84129:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 84130:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 84131:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 84132:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 84133:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 84134:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 84135:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 84136:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 84137:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 84138:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 84139:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 84140:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 84141:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 84142:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 84143:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 84144:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 84145:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 84146:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 84147:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 84148:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 84149:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 84150:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 84151:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 84152:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 84153:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 84154:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 84155:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 84156:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 84157:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 84158:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 84159:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 84160:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 84161:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 84162:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 84163:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 84164:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 84165:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 84166:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 84167:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 84168:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 84169:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 84170:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 84171:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 84172:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 84173:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 84174:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 84175:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 84176:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 84177:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 84178:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 84179:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 84180:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 84181:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 84182:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 84183:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 84184:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 84185:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 84186:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 84187:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 84188:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 84189:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 84190:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 84191:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 84192:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 84193:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 84194:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 84195:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 84196:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 84197:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 84198:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 84199:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 84200:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 84201:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 84202:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 84203:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 84204:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 84205:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 84206:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 84207:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 84208:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 84209:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 84210:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 84211:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 84212:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 84213:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 84214:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 84215:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 84216:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 84217:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 84218:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 84219:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 84220:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 84221:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 84222:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 84223:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 84224:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 84225:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 84226:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 84227:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 84228:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 84229:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 84230:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 84231:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 84232:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 84233:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 84234:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 84235:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 84236:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 84237:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 84238:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 84239:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 84240:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 84241:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 84242:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 84243:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 84244:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 84245:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 84246:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 84247:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 84248:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 84249:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 84250:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 84251:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 84252:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 84253:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 84254:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 84255:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 84256:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 84257:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 84258:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 84259:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 84260:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 84261:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 84262:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 84263:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 84264:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 84265:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 84266:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 84267:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 84268:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 84269:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 84270:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 84271:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 84272:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 84273:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 84274:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 84275:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 84276:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 84277:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 84278:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 84279:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 84280:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 84281:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 84282:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 84283:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 84284:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 84285:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 84286:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 84287:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 84288:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 84289:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 84290:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 84291:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 84292:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 84293:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 84294:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 84295:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 84296:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 84297:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 84298:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 84299:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 84300:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 84301:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 84302:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 84303:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 84304:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 84305:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 84306:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 84307:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 84308:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 84309:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 84310:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 84311:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 84312:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 84313:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 84314:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 84315:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 84316:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 84317:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 84318:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 84319:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 84320:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 84321:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 84322:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 84323:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 84324:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 84325:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 84326:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 84327:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 84328:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 84329:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 84330:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 84331:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 84332:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 84333:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 84334:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 84335:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 84336:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 84337:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 84338:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 84339:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 84340:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 84341:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 84342:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 84343:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 84344:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 84345:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 84346:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 84347:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 84348:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 84349:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 84350:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 84351:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 84352:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 84353:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 84354:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 84355:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 84356:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 84357:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 84358:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 84359:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 84360:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 84361:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 84362:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 84363:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 84364:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 84365:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 84366:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 84367:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 84368:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 84369:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 84370:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 84371:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 84372:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 84373:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 84374:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 84375:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 84376:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 84377:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 84378:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 84379:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 84380:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 84381:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 84382:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 84383:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 84384:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 84385:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 84386:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 84387:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 84388:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 84389:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 84390:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 84391:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 84392:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 84393:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 84394:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 84395:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 84396:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 84397:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 84398:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 84399:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 84400:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 84401:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 84402:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 84403:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 84404:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 84405:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 84406:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 84407:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 84408:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 84409:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 84410:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 84411:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 84412:20]
  assign io_z = ~x99; // @[Snxn100k.scala 84413:16]
endmodule
module SnxnLv4Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 83334:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 83335:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 83336:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 83337:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 83338:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 83339:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 83340:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 83341:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 83342:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 83343:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 83344:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 83345:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 83346:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 83347:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 83348:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 83349:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 83350:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 83351:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 83352:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 83353:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 83354:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 83355:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 83356:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 83357:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 83358:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 83359:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 83360:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 83361:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 83362:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 83363:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 83364:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 83365:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 83366:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 83367:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 83368:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 83369:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 83370:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 83371:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 83372:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 83373:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 83374:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 83375:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 83376:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 83377:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 83378:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 83379:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 83380:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 83381:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 83382:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 83383:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 83384:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 83385:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 83386:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 83387:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 83388:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 83389:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 83390:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 83391:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 83392:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 83393:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 83394:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 83395:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 83396:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 83397:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 83398:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 83399:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 83400:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 83401:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 83402:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 83403:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 83404:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 83405:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 83406:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 83407:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 83408:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 83409:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 83410:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 83411:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 83412:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 83413:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 83414:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 83415:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 83416:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 83417:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 83418:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 83419:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 83420:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 83421:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 83422:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 83423:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 83424:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 83425:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 83426:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 83427:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 83428:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 83429:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 83430:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 83431:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 83432:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 83433:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 83434:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 83435:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 83436:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 83437:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 83438:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 83439:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 83440:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 83441:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 83442:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 83443:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 83444:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 83445:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 83446:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 83447:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 83448:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 83449:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 83450:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 83451:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 83452:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 83453:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 83454:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 83455:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 83456:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 83457:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 83458:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 83459:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 83460:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 83461:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 83462:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 83463:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 83464:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 83465:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 83466:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 83467:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 83468:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 83469:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 83470:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 83471:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 83472:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 83473:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 83474:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 83475:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 83476:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 83477:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 83478:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 83479:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 83480:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 83481:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 83482:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 83483:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 83484:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 83485:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 83486:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 83487:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 83488:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 83489:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 83490:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 83491:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 83492:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 83493:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 83494:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 83495:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 83496:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 83497:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 83498:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 83499:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 83500:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 83501:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 83502:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 83503:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 83504:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 83505:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 83506:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 83507:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 83508:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 83509:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 83510:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 83511:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 83512:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 83513:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 83514:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 83515:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 83516:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 83517:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 83518:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 83519:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 83520:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 83521:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 83522:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 83523:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 83524:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 83525:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 83526:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 83527:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 83528:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 83529:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 83530:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 83531:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 83532:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 83533:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 83534:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 83535:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 83536:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 83537:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 83538:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 83539:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 83540:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 83541:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 83542:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 83543:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 83544:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 83545:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 83546:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 83547:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 83548:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 83549:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 83550:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 83551:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 83552:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 83553:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 83554:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 83555:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 83556:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 83557:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 83558:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 83559:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 83560:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 83561:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 83562:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 83563:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 83564:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 83565:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 83566:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 83567:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 83568:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 83569:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 83570:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 83571:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 83572:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 83573:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 83574:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 83575:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 83576:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 83577:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 83578:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 83579:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 83580:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 83581:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 83582:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 83583:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 83584:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 83585:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 83586:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 83587:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 83588:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 83589:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 83590:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 83591:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 83592:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 83593:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 83594:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 83595:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 83596:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 83597:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 83598:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 83599:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 83600:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 83601:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 83602:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 83603:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 83604:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 83605:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 83606:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 83607:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 83608:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 83609:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 83610:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 83611:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 83612:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 83613:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 83614:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 83615:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 83616:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 83617:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 83618:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 83619:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 83620:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 83621:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 83622:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 83623:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 83624:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 83625:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 83626:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 83627:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 83628:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 83629:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 83630:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 83631:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 83632:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 83633:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 83634:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 83635:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 83636:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 83637:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 83638:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 83639:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 83640:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 83641:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 83642:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 83643:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 83644:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 83645:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 83646:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 83647:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 83648:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 83649:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 83650:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 83651:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 83652:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 83653:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 83654:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 83655:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 83656:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 83657:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 83658:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 83659:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 83660:20]
  assign io_z = ~x81; // @[Snxn100k.scala 83661:16]
endmodule
module SnxnLv3Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst0_io_a; // @[Snxn100k.scala 21805:33]
  wire  inst_SnxnLv4Inst0_io_b; // @[Snxn100k.scala 21805:33]
  wire  inst_SnxnLv4Inst0_io_z; // @[Snxn100k.scala 21805:33]
  wire  inst_SnxnLv4Inst1_io_a; // @[Snxn100k.scala 21809:33]
  wire  inst_SnxnLv4Inst1_io_b; // @[Snxn100k.scala 21809:33]
  wire  inst_SnxnLv4Inst1_io_z; // @[Snxn100k.scala 21809:33]
  wire  inst_SnxnLv4Inst2_io_a; // @[Snxn100k.scala 21813:33]
  wire  inst_SnxnLv4Inst2_io_b; // @[Snxn100k.scala 21813:33]
  wire  inst_SnxnLv4Inst2_io_z; // @[Snxn100k.scala 21813:33]
  wire  inst_SnxnLv4Inst3_io_a; // @[Snxn100k.scala 21817:33]
  wire  inst_SnxnLv4Inst3_io_b; // @[Snxn100k.scala 21817:33]
  wire  inst_SnxnLv4Inst3_io_z; // @[Snxn100k.scala 21817:33]
  wire  _sum_T_1 = inst_SnxnLv4Inst0_io_z + inst_SnxnLv4Inst1_io_z; // @[Snxn100k.scala 21821:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst2_io_z; // @[Snxn100k.scala 21821:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst3_io_z; // @[Snxn100k.scala 21821:86]
  SnxnLv4Inst0 inst_SnxnLv4Inst0 ( // @[Snxn100k.scala 21805:33]
    .io_a(inst_SnxnLv4Inst0_io_a),
    .io_b(inst_SnxnLv4Inst0_io_b),
    .io_z(inst_SnxnLv4Inst0_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst1 ( // @[Snxn100k.scala 21809:33]
    .io_a(inst_SnxnLv4Inst1_io_a),
    .io_b(inst_SnxnLv4Inst1_io_b),
    .io_z(inst_SnxnLv4Inst1_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst2 ( // @[Snxn100k.scala 21813:33]
    .io_a(inst_SnxnLv4Inst2_io_a),
    .io_b(inst_SnxnLv4Inst2_io_b),
    .io_z(inst_SnxnLv4Inst2_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst3 ( // @[Snxn100k.scala 21817:33]
    .io_a(inst_SnxnLv4Inst3_io_a),
    .io_b(inst_SnxnLv4Inst3_io_b),
    .io_z(inst_SnxnLv4Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21822:15]
  assign inst_SnxnLv4Inst0_io_a = io_a; // @[Snxn100k.scala 21806:26]
  assign inst_SnxnLv4Inst0_io_b = io_b; // @[Snxn100k.scala 21807:26]
  assign inst_SnxnLv4Inst1_io_a = io_a; // @[Snxn100k.scala 21810:26]
  assign inst_SnxnLv4Inst1_io_b = io_b; // @[Snxn100k.scala 21811:26]
  assign inst_SnxnLv4Inst2_io_a = io_a; // @[Snxn100k.scala 21814:26]
  assign inst_SnxnLv4Inst2_io_b = io_b; // @[Snxn100k.scala 21815:26]
  assign inst_SnxnLv4Inst3_io_a = io_a; // @[Snxn100k.scala 21818:26]
  assign inst_SnxnLv4Inst3_io_b = io_b; // @[Snxn100k.scala 21819:26]
endmodule
module SnxnLv4Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 80604:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 80605:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 80606:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 80607:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 80608:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 80609:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 80610:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 80611:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 80612:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 80613:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 80614:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 80615:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 80616:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 80617:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 80618:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 80619:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 80620:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 80621:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 80622:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 80623:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 80624:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 80625:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 80626:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 80627:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 80628:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 80629:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 80630:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 80631:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 80632:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 80633:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 80634:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 80635:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 80636:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 80637:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 80638:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 80639:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 80640:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 80641:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 80642:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 80643:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 80644:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 80645:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 80646:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 80647:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 80648:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 80649:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 80650:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 80651:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 80652:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 80653:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 80654:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 80655:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 80656:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 80657:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 80658:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 80659:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 80660:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 80661:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 80662:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 80663:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 80664:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 80665:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 80666:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 80667:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 80668:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 80669:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 80670:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 80671:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 80672:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 80673:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 80674:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 80675:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 80676:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 80677:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 80678:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 80679:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 80680:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 80681:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 80682:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 80683:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 80684:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 80685:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 80686:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 80687:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 80688:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 80689:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 80690:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 80691:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 80692:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 80693:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 80694:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 80695:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 80696:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 80697:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 80698:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 80699:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 80700:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 80701:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 80702:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 80703:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 80704:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 80705:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 80706:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 80707:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 80708:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 80709:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 80710:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 80711:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 80712:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 80713:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 80714:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 80715:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 80716:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 80717:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 80718:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 80719:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 80720:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 80721:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 80722:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 80723:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 80724:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 80725:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 80726:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 80727:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 80728:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 80729:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 80730:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 80731:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 80732:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 80733:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 80734:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 80735:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 80736:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 80737:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 80738:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 80739:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 80740:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 80741:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 80742:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 80743:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 80744:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 80745:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 80746:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 80747:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 80748:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 80749:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 80750:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 80751:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 80752:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 80753:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 80754:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 80755:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 80756:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 80757:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 80758:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 80759:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 80760:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 80761:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 80762:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 80763:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 80764:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 80765:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 80766:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 80767:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 80768:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 80769:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 80770:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 80771:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 80772:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 80773:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 80774:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 80775:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 80776:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 80777:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 80778:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 80779:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 80780:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 80781:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 80782:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 80783:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 80784:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 80785:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 80786:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 80787:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 80788:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 80789:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 80790:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 80791:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 80792:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 80793:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 80794:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 80795:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 80796:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 80797:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 80798:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 80799:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 80800:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 80801:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 80802:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 80803:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 80804:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 80805:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 80806:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 80807:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 80808:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 80809:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 80810:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 80811:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 80812:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 80813:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 80814:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 80815:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 80816:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 80817:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 80818:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 80819:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 80820:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 80821:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 80822:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 80823:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 80824:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 80825:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 80826:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 80827:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 80828:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 80829:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 80830:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 80831:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 80832:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 80833:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 80834:20]
  assign io_z = ~x57; // @[Snxn100k.scala 80835:16]
endmodule
module SnxnLv4Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81522:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81523:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81524:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81525:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81526:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81527:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81528:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81529:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81530:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81531:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81532:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81533:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81534:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81535:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81536:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81537:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81538:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81539:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81540:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81541:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81542:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81543:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81544:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81545:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81546:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81547:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81548:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81549:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81550:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81551:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81552:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81553:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81554:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81555:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81556:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81557:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81558:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81559:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81560:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81561:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81562:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81563:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81564:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81565:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81566:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81567:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81568:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81569:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81570:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81571:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81572:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81573:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81574:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81575:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81576:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81577:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81578:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81579:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81580:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81581:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81582:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81583:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81584:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81585:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81586:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81587:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81588:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81589:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81590:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81591:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81592:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81593:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81594:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81595:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81596:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81597:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81598:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81599:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81600:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81601:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 81602:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 81603:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 81604:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 81605:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 81606:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 81607:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 81608:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 81609:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 81610:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 81611:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 81612:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 81613:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 81614:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 81615:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 81616:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 81617:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 81618:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 81619:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 81620:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 81621:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 81622:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 81623:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 81624:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 81625:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 81626:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 81627:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 81628:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 81629:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 81630:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 81631:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 81632:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 81633:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 81634:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 81635:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 81636:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 81637:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 81638:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 81639:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 81640:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 81641:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 81642:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 81643:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 81644:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 81645:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 81646:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 81647:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 81648:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 81649:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 81650:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 81651:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 81652:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 81653:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 81654:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 81655:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 81656:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 81657:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 81658:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 81659:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 81660:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 81661:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 81662:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 81663:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 81664:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 81665:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 81666:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 81667:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 81668:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 81669:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 81670:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 81671:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 81672:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 81673:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 81674:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 81675:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81676:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 81677:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 81678:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 81679:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 81680:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 81681:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 81682:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 81683:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 81684:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 81685:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 81686:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 81687:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 81688:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 81689:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 81690:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 81691:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 81692:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 81693:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 81694:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 81695:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 81696:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 81697:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 81698:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 81699:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 81700:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 81701:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 81702:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 81703:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 81704:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 81705:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 81706:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 81707:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 81708:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 81709:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 81710:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 81711:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 81712:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 81713:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 81714:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 81715:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 81716:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 81717:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 81718:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 81719:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 81720:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 81721:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 81722:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 81723:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 81724:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 81725:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 81726:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 81727:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 81728:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 81729:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 81730:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 81731:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 81732:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 81733:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 81734:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 81735:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 81736:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 81737:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 81738:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 81739:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 81740:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 81741:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 81742:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 81743:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 81744:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 81745:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 81746:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 81747:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 81748:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 81749:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 81750:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 81751:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 81752:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 81753:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 81754:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 81755:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 81756:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 81757:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 81758:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 81759:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 81760:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 81761:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 81762:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 81763:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 81764:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 81765:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 81766:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 81767:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 81768:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 81769:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 81770:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 81771:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 81772:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 81773:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 81774:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 81775:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 81776:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 81777:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 81778:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 81779:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 81780:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 81781:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 81782:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 81783:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 81784:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 81785:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 81786:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 81787:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 81788:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 81789:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 81790:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 81791:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 81792:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 81793:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 81794:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 81795:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 81796:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 81797:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 81798:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 81799:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 81800:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 81801:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 81802:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 81803:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 81804:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 81805:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 81806:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 81807:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 81808:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 81809:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 81810:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 81811:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 81812:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 81813:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 81814:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 81815:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 81816:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 81817:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 81818:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 81819:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 81820:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 81821:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 81822:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 81823:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 81824:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 81825:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 81826:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 81827:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 81828:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 81829:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 81830:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 81831:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 81832:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 81833:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 81834:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 81835:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 81836:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 81837:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 81838:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 81839:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 81840:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 81841:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 81842:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 81843:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 81844:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 81845:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 81846:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 81847:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 81848:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 81849:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 81850:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 81851:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 81852:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 81853:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 81854:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 81855:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 81856:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 81857:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 81858:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 81859:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 81860:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 81861:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 81862:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 81863:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 81864:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 81865:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 81866:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 81867:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 81868:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 81869:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 81870:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 81871:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 81872:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 81873:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 81874:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 81875:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 81876:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 81877:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 81878:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 81879:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 81880:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 81881:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 81882:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 81883:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 81884:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 81885:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 81886:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 81887:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 81888:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 81889:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 81890:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 81891:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 81892:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 81893:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 81894:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 81895:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 81896:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 81897:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 81898:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 81899:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 81900:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 81901:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 81902:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 81903:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 81904:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 81905:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 81906:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 81907:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 81908:20]
  assign io_z = ~x96; // @[Snxn100k.scala 81909:16]
endmodule
module SnxnLv4Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 80846:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 80847:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 80848:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 80849:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 80850:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 80851:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 80852:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 80853:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 80854:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 80855:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 80856:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 80857:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 80858:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 80859:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 80860:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 80861:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 80862:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 80863:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 80864:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 80865:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 80866:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 80867:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 80868:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 80869:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 80870:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 80871:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 80872:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 80873:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 80874:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 80875:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 80876:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 80877:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 80878:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 80879:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 80880:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 80881:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 80882:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 80883:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 80884:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 80885:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 80886:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 80887:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 80888:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 80889:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 80890:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 80891:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 80892:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 80893:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 80894:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 80895:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 80896:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 80897:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 80898:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 80899:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 80900:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 80901:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 80902:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 80903:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 80904:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 80905:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 80906:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 80907:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 80908:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 80909:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 80910:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 80911:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 80912:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 80913:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 80914:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 80915:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 80916:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 80917:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 80918:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 80919:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 80920:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 80921:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 80922:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 80923:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 80924:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 80925:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 80926:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 80927:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 80928:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 80929:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 80930:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 80931:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 80932:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 80933:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 80934:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 80935:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 80936:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 80937:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 80938:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 80939:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 80940:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 80941:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 80942:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 80943:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 80944:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 80945:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 80946:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 80947:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 80948:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 80949:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 80950:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 80951:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 80952:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 80953:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 80954:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 80955:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 80956:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 80957:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 80958:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 80959:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 80960:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 80961:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 80962:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 80963:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 80964:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 80965:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 80966:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 80967:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 80968:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 80969:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 80970:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 80971:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 80972:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 80973:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 80974:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 80975:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 80976:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 80977:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 80978:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 80979:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 80980:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 80981:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 80982:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 80983:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 80984:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 80985:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 80986:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 80987:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 80988:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 80989:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 80990:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 80991:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 80992:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 80993:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 80994:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 80995:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 80996:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 80997:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 80998:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 80999:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81000:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 81001:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 81002:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 81003:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 81004:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 81005:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 81006:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 81007:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 81008:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 81009:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 81010:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 81011:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 81012:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 81013:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 81014:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 81015:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 81016:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 81017:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 81018:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 81019:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 81020:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 81021:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 81022:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 81023:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 81024:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 81025:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 81026:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 81027:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 81028:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 81029:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 81030:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 81031:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 81032:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 81033:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 81034:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 81035:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 81036:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 81037:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 81038:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 81039:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 81040:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 81041:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 81042:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 81043:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 81044:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 81045:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 81046:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 81047:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 81048:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 81049:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 81050:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 81051:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 81052:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 81053:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 81054:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 81055:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 81056:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 81057:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 81058:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 81059:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 81060:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 81061:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 81062:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 81063:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 81064:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 81065:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 81066:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 81067:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 81068:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 81069:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 81070:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 81071:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 81072:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 81073:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 81074:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 81075:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 81076:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 81077:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 81078:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 81079:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 81080:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 81081:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 81082:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 81083:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 81084:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 81085:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 81086:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 81087:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 81088:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 81089:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 81090:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 81091:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 81092:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 81093:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 81094:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 81095:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 81096:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 81097:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 81098:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 81099:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 81100:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 81101:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 81102:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 81103:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 81104:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 81105:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 81106:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 81107:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 81108:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 81109:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 81110:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 81111:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 81112:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 81113:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 81114:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 81115:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 81116:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 81117:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 81118:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 81119:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 81120:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 81121:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 81122:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 81123:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 81124:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 81125:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 81126:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 81127:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 81128:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 81129:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 81130:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 81131:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 81132:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 81133:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 81134:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 81135:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 81136:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 81137:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 81138:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 81139:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 81140:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 81141:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 81142:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 81143:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 81144:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 81145:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 81146:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 81147:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 81148:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 81149:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 81150:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 81151:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 81152:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 81153:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 81154:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 81155:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 81156:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 81157:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 81158:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 81159:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 81160:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 81161:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 81162:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 81163:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 81164:20]
  assign io_z = ~x79; // @[Snxn100k.scala 81165:16]
endmodule
module SnxnLv4Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81176:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81177:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81178:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81179:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81180:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81181:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81182:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81183:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81184:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81185:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81186:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81187:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81188:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81189:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81190:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81191:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81192:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81193:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81194:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81195:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81196:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81197:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81198:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81199:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81200:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81201:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81202:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81203:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81204:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81205:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81206:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81207:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81208:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81209:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81210:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81211:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81212:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81213:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81214:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81215:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81216:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81217:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81218:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81219:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81220:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81221:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81222:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81223:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81224:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81225:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81226:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81227:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81228:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81229:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81230:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81231:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81232:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81233:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81234:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81235:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81236:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81237:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81238:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81239:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81240:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81241:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81242:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81243:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81244:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81245:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81246:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81247:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81248:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81249:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81250:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81251:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81252:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81253:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81254:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81255:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 81256:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 81257:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 81258:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 81259:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 81260:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 81261:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 81262:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 81263:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 81264:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 81265:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 81266:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 81267:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 81268:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 81269:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 81270:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 81271:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 81272:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 81273:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 81274:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 81275:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 81276:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 81277:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 81278:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 81279:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 81280:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 81281:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 81282:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 81283:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 81284:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 81285:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 81286:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 81287:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 81288:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 81289:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 81290:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 81291:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 81292:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 81293:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 81294:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 81295:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 81296:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 81297:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 81298:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 81299:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 81300:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 81301:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 81302:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 81303:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 81304:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 81305:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 81306:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 81307:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 81308:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 81309:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 81310:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 81311:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 81312:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 81313:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 81314:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 81315:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 81316:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 81317:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 81318:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 81319:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 81320:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 81321:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 81322:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 81323:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 81324:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 81325:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 81326:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 81327:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 81328:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 81329:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81330:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 81331:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 81332:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 81333:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 81334:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 81335:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 81336:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 81337:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 81338:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 81339:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 81340:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 81341:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 81342:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 81343:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 81344:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 81345:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 81346:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 81347:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 81348:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 81349:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 81350:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 81351:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 81352:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 81353:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 81354:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 81355:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 81356:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 81357:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 81358:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 81359:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 81360:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 81361:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 81362:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 81363:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 81364:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 81365:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 81366:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 81367:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 81368:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 81369:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 81370:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 81371:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 81372:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 81373:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 81374:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 81375:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 81376:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 81377:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 81378:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 81379:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 81380:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 81381:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 81382:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 81383:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 81384:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 81385:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 81386:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 81387:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 81388:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 81389:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 81390:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 81391:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 81392:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 81393:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 81394:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 81395:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 81396:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 81397:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 81398:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 81399:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 81400:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 81401:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 81402:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 81403:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 81404:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 81405:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 81406:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 81407:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 81408:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 81409:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 81410:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 81411:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 81412:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 81413:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 81414:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 81415:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 81416:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 81417:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 81418:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 81419:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 81420:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 81421:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 81422:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 81423:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 81424:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 81425:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 81426:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 81427:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 81428:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 81429:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 81430:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 81431:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 81432:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 81433:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 81434:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 81435:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 81436:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 81437:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 81438:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 81439:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 81440:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 81441:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 81442:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 81443:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 81444:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 81445:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 81446:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 81447:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 81448:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 81449:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 81450:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 81451:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 81452:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 81453:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 81454:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 81455:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 81456:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 81457:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 81458:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 81459:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 81460:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 81461:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 81462:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 81463:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 81464:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 81465:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 81466:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 81467:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 81468:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 81469:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 81470:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 81471:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 81472:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 81473:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 81474:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 81475:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 81476:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 81477:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 81478:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 81479:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 81480:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 81481:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 81482:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 81483:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 81484:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 81485:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 81486:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 81487:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 81488:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 81489:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 81490:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 81491:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 81492:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 81493:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 81494:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 81495:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 81496:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 81497:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 81498:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 81499:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 81500:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 81501:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 81502:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 81503:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 81504:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 81505:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 81506:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 81507:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 81508:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 81509:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 81510:20]
  assign io_z = ~x83; // @[Snxn100k.scala 81511:16]
endmodule
module SnxnLv3Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst4_io_a; // @[Snxn100k.scala 21151:33]
  wire  inst_SnxnLv4Inst4_io_b; // @[Snxn100k.scala 21151:33]
  wire  inst_SnxnLv4Inst4_io_z; // @[Snxn100k.scala 21151:33]
  wire  inst_SnxnLv4Inst5_io_a; // @[Snxn100k.scala 21155:33]
  wire  inst_SnxnLv4Inst5_io_b; // @[Snxn100k.scala 21155:33]
  wire  inst_SnxnLv4Inst5_io_z; // @[Snxn100k.scala 21155:33]
  wire  inst_SnxnLv4Inst6_io_a; // @[Snxn100k.scala 21159:33]
  wire  inst_SnxnLv4Inst6_io_b; // @[Snxn100k.scala 21159:33]
  wire  inst_SnxnLv4Inst6_io_z; // @[Snxn100k.scala 21159:33]
  wire  inst_SnxnLv4Inst7_io_a; // @[Snxn100k.scala 21163:33]
  wire  inst_SnxnLv4Inst7_io_b; // @[Snxn100k.scala 21163:33]
  wire  inst_SnxnLv4Inst7_io_z; // @[Snxn100k.scala 21163:33]
  wire  _sum_T_1 = inst_SnxnLv4Inst4_io_z + inst_SnxnLv4Inst5_io_z; // @[Snxn100k.scala 21167:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst6_io_z; // @[Snxn100k.scala 21167:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst7_io_z; // @[Snxn100k.scala 21167:86]
  SnxnLv4Inst4 inst_SnxnLv4Inst4 ( // @[Snxn100k.scala 21151:33]
    .io_a(inst_SnxnLv4Inst4_io_a),
    .io_b(inst_SnxnLv4Inst4_io_b),
    .io_z(inst_SnxnLv4Inst4_io_z)
  );
  SnxnLv4Inst5 inst_SnxnLv4Inst5 ( // @[Snxn100k.scala 21155:33]
    .io_a(inst_SnxnLv4Inst5_io_a),
    .io_b(inst_SnxnLv4Inst5_io_b),
    .io_z(inst_SnxnLv4Inst5_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst6 ( // @[Snxn100k.scala 21159:33]
    .io_a(inst_SnxnLv4Inst6_io_a),
    .io_b(inst_SnxnLv4Inst6_io_b),
    .io_z(inst_SnxnLv4Inst6_io_z)
  );
  SnxnLv4Inst7 inst_SnxnLv4Inst7 ( // @[Snxn100k.scala 21163:33]
    .io_a(inst_SnxnLv4Inst7_io_a),
    .io_b(inst_SnxnLv4Inst7_io_b),
    .io_z(inst_SnxnLv4Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21168:15]
  assign inst_SnxnLv4Inst4_io_a = io_a; // @[Snxn100k.scala 21152:26]
  assign inst_SnxnLv4Inst4_io_b = io_b; // @[Snxn100k.scala 21153:26]
  assign inst_SnxnLv4Inst5_io_a = io_a; // @[Snxn100k.scala 21156:26]
  assign inst_SnxnLv4Inst5_io_b = io_b; // @[Snxn100k.scala 21157:26]
  assign inst_SnxnLv4Inst6_io_a = io_a; // @[Snxn100k.scala 21160:26]
  assign inst_SnxnLv4Inst6_io_b = io_b; // @[Snxn100k.scala 21161:26]
  assign inst_SnxnLv4Inst7_io_a = io_a; // @[Snxn100k.scala 21164:26]
  assign inst_SnxnLv4Inst7_io_b = io_b; // @[Snxn100k.scala 21165:26]
endmodule
module SnxnLv4Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 80070:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 80071:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 80072:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 80073:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 80074:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 80075:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 80076:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 80077:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 80078:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 80079:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 80080:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 80081:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 80082:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 80083:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 80084:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 80085:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 80086:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 80087:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 80088:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 80089:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 80090:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 80091:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 80092:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 80093:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 80094:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 80095:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 80096:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 80097:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 80098:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 80099:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 80100:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 80101:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 80102:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 80103:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 80104:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 80105:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 80106:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 80107:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 80108:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 80109:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 80110:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 80111:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 80112:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 80113:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 80114:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 80115:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 80116:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 80117:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 80118:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 80119:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 80120:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 80121:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 80122:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 80123:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 80124:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 80125:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 80126:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 80127:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 80128:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 80129:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 80130:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 80131:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 80132:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 80133:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 80134:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 80135:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 80136:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 80137:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 80138:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 80139:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 80140:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 80141:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 80142:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 80143:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 80144:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 80145:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 80146:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 80147:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 80148:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 80149:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 80150:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 80151:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 80152:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 80153:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 80154:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 80155:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 80156:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 80157:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 80158:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 80159:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 80160:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 80161:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 80162:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 80163:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 80164:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 80165:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 80166:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 80167:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 80168:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 80169:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 80170:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 80171:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 80172:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 80173:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 80174:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 80175:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 80176:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 80177:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 80178:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 80179:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 80180:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 80181:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 80182:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 80183:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 80184:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 80185:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 80186:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 80187:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 80188:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 80189:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 80190:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 80191:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 80192:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 80193:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 80194:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 80195:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 80196:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 80197:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 80198:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 80199:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 80200:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 80201:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 80202:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 80203:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 80204:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 80205:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 80206:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 80207:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 80208:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 80209:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 80210:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 80211:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 80212:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 80213:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 80214:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 80215:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 80216:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 80217:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 80218:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 80219:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 80220:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 80221:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 80222:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 80223:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 80224:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 80225:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 80226:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 80227:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 80228:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 80229:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 80230:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 80231:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 80232:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 80233:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 80234:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 80235:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 80236:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 80237:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 80238:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 80239:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 80240:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 80241:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 80242:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 80243:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 80244:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 80245:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 80246:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 80247:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 80248:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 80249:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 80250:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 80251:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 80252:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 80253:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 80254:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 80255:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 80256:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 80257:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 80258:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 80259:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 80260:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 80261:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 80262:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 80263:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 80264:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 80265:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 80266:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 80267:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 80268:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 80269:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 80270:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 80271:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 80272:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 80273:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 80274:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 80275:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 80276:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 80277:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 80278:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 80279:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 80280:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 80281:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 80282:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 80283:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 80284:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 80285:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 80286:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 80287:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 80288:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 80289:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 80290:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 80291:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 80292:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 80293:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 80294:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 80295:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 80296:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 80297:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 80298:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 80299:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 80300:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 80301:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 80302:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 80303:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 80304:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 80305:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 80306:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 80307:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 80308:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 80309:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 80310:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 80311:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 80312:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 80313:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 80314:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 80315:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 80316:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 80317:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 80318:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 80319:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 80320:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 80321:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 80322:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 80323:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 80324:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 80325:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 80326:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 80327:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 80328:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 80329:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 80330:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 80331:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 80332:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 80333:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 80334:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 80335:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 80336:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 80337:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 80338:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 80339:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 80340:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 80341:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 80342:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 80343:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 80344:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 80345:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 80346:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 80347:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 80348:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 80349:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 80350:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 80351:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 80352:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 80353:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 80354:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 80355:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 80356:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 80357:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 80358:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 80359:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 80360:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 80361:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 80362:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 80363:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 80364:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 80365:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 80366:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 80367:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 80368:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 80369:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 80370:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 80371:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 80372:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 80373:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 80374:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 80375:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 80376:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 80377:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 80378:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 80379:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 80380:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 80381:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 80382:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 80383:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 80384:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 80385:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 80386:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 80387:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 80388:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 80389:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 80390:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 80391:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 80392:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 80393:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 80394:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 80395:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 80396:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 80397:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 80398:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 80399:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 80400:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 80401:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 80402:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 80403:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 80404:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 80405:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 80406:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 80407:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 80408:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 80409:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 80410:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 80411:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 80412:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 80413:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 80414:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 80415:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 80416:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 80417:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 80418:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 80419:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 80420:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 80421:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 80422:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 80423:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 80424:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 80425:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 80426:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 80427:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 80428:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 80429:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 80430:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 80431:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 80432:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 80433:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 80434:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 80435:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 80436:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 80437:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 80438:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 80439:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 80440:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 80441:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 80442:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 80443:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 80444:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 80445:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 80446:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 80447:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 80448:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 80449:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 80450:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 80451:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 80452:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 80453:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 80454:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 80455:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 80456:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 80457:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 80458:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 80459:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 80460:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 80461:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 80462:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 80463:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 80464:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 80465:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 80466:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 80467:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 80468:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 80469:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 80470:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 80471:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 80472:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 80473:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 80474:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 80475:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 80476:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 80477:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 80478:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 80479:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 80480:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 80481:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 80482:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 80483:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 80484:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 80485:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 80486:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 80487:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 80488:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 80489:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 80490:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 80491:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 80492:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 80493:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 80494:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 80495:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 80496:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 80497:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 80498:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 80499:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 80500:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 80501:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 80502:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 80503:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 80504:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 80505:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 80506:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 80507:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 80508:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 80509:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 80510:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 80511:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 80512:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 80513:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 80514:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 80515:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 80516:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 80517:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 80518:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 80519:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 80520:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 80521:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 80522:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 80523:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 80524:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 80525:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 80526:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 80527:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 80528:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 80529:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 80530:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 80531:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 80532:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 80533:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 80534:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 80535:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 80536:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 80537:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 80538:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 80539:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 80540:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 80541:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 80542:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 80543:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 80544:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 80545:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 80546:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 80547:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 80548:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 80549:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 80550:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 80551:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 80552:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 80553:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 80554:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 80555:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 80556:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 80557:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 80558:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 80559:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 80560:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 80561:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 80562:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 80563:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 80564:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 80565:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 80566:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 80567:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 80568:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 80569:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 80570:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 80571:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 80572:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 80573:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 80574:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 80575:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 80576:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 80577:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 80578:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 80579:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 80580:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 80581:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 80582:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 80583:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 80584:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 80585:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 80586:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 80587:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 80588:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 80589:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 80590:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 80591:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 80592:22]
  assign io_z = ~x130; // @[Snxn100k.scala 80593:17]
endmodule
module SnxnLv4Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78936:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78937:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78938:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78939:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78940:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78941:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78942:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78943:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78944:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78945:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78946:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78947:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78948:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78949:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78950:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78951:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78952:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78953:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78954:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78955:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78956:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78957:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78958:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78959:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78960:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78961:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78962:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78963:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78964:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78965:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78966:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78967:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78968:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78969:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78970:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78971:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78972:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78973:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78974:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78975:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78976:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78977:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78978:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78979:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78980:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78981:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78982:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78983:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78984:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78985:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78986:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78987:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78988:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78989:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78990:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78991:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78992:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78993:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78994:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78995:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78996:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78997:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78998:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78999:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 79000:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 79001:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 79002:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 79003:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 79004:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 79005:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 79006:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 79007:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 79008:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 79009:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 79010:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 79011:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 79012:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 79013:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 79014:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 79015:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 79016:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 79017:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 79018:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 79019:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 79020:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 79021:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 79022:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 79023:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 79024:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 79025:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 79026:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 79027:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 79028:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 79029:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 79030:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 79031:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 79032:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 79033:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 79034:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 79035:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 79036:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 79037:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 79038:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 79039:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 79040:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 79041:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 79042:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 79043:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 79044:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 79045:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 79046:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 79047:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 79048:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 79049:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 79050:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 79051:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 79052:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 79053:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 79054:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 79055:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 79056:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 79057:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 79058:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 79059:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 79060:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 79061:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 79062:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79063:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79064:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79065:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79066:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79067:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79068:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79069:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79070:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79071:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79072:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79073:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79074:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79075:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79076:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79077:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79078:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79079:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79080:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79081:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79082:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79083:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79084:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79085:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79086:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79087:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79088:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79089:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79090:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79091:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79092:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79093:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79094:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79095:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79096:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79097:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79098:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79099:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79100:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79101:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79102:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79103:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79104:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79105:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79106:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79107:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79108:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79109:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79110:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79111:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79112:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79113:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79114:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79115:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79116:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79117:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79118:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79119:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79120:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79121:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79122:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79123:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79124:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79125:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79126:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79127:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79128:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79129:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79130:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79131:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79132:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79133:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79134:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 79135:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 79136:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 79137:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 79138:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 79139:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 79140:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 79141:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 79142:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 79143:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 79144:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 79145:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 79146:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 79147:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 79148:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 79149:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 79150:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 79151:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 79152:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 79153:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 79154:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 79155:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 79156:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 79157:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 79158:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 79159:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 79160:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 79161:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 79162:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 79163:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 79164:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 79165:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 79166:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 79167:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 79168:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 79169:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 79170:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 79171:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 79172:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 79173:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 79174:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 79175:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 79176:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 79177:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 79178:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 79179:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 79180:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 79181:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 79182:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 79183:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 79184:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 79185:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 79186:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 79187:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 79188:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 79189:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 79190:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 79191:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 79192:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 79193:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 79194:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 79195:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 79196:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 79197:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 79198:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 79199:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 79200:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 79201:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 79202:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 79203:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 79204:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 79205:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 79206:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 79207:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 79208:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 79209:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 79210:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 79211:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 79212:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 79213:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 79214:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 79215:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 79216:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 79217:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 79218:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 79219:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 79220:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 79221:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 79222:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 79223:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 79224:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 79225:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 79226:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 79227:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 79228:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 79229:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 79230:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 79231:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 79232:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 79233:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 79234:20]
  assign io_z = ~x74; // @[Snxn100k.scala 79235:16]
endmodule
module SnxnLv4Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 79616:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 79617:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 79618:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 79619:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 79620:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 79621:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 79622:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 79623:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 79624:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 79625:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 79626:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 79627:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 79628:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 79629:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 79630:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 79631:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 79632:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 79633:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 79634:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 79635:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 79636:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 79637:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 79638:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 79639:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 79640:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 79641:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 79642:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 79643:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 79644:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 79645:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 79646:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 79647:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 79648:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 79649:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 79650:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 79651:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 79652:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 79653:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 79654:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 79655:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 79656:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 79657:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 79658:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 79659:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 79660:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 79661:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 79662:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 79663:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 79664:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 79665:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 79666:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 79667:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 79668:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 79669:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 79670:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 79671:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 79672:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 79673:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 79674:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 79675:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 79676:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 79677:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 79678:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 79679:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 79680:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 79681:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 79682:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 79683:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 79684:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 79685:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 79686:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 79687:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 79688:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 79689:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 79690:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 79691:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 79692:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 79693:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 79694:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 79695:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 79696:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 79697:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 79698:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 79699:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 79700:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 79701:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 79702:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 79703:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 79704:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 79705:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 79706:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 79707:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 79708:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 79709:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 79710:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 79711:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 79712:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 79713:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 79714:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 79715:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 79716:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 79717:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 79718:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 79719:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 79720:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 79721:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 79722:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 79723:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 79724:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 79725:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 79726:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 79727:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 79728:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 79729:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 79730:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 79731:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 79732:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 79733:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 79734:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 79735:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 79736:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 79737:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 79738:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 79739:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 79740:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 79741:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 79742:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79743:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79744:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79745:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79746:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79747:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79748:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79749:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79750:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79751:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79752:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79753:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79754:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79755:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79756:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79757:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79758:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79759:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79760:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79761:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79762:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79763:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79764:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79765:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79766:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79767:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79768:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79769:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79770:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79771:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79772:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79773:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79774:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79775:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79776:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79777:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79778:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79779:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79780:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79781:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79782:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79783:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79784:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79785:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79786:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79787:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79788:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79789:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79790:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79791:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79792:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79793:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79794:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79795:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79796:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79797:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79798:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79799:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79800:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79801:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79802:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79803:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79804:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79805:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79806:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79807:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79808:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79809:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79810:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79811:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79812:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79813:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79814:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 79815:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 79816:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 79817:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 79818:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 79819:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 79820:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 79821:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 79822:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 79823:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 79824:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 79825:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 79826:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 79827:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 79828:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 79829:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 79830:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 79831:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 79832:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 79833:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 79834:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 79835:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 79836:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 79837:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 79838:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 79839:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 79840:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 79841:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 79842:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 79843:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 79844:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 79845:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 79846:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 79847:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 79848:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 79849:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 79850:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 79851:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 79852:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 79853:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 79854:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 79855:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 79856:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 79857:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 79858:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 79859:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 79860:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 79861:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 79862:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 79863:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 79864:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 79865:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 79866:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 79867:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 79868:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 79869:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 79870:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 79871:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 79872:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 79873:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 79874:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 79875:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 79876:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 79877:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 79878:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 79879:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 79880:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 79881:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 79882:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 79883:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 79884:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 79885:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 79886:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 79887:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 79888:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 79889:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 79890:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 79891:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 79892:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 79893:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 79894:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 79895:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 79896:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 79897:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 79898:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 79899:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 79900:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 79901:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 79902:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 79903:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 79904:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 79905:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 79906:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 79907:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 79908:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 79909:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 79910:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 79911:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 79912:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 79913:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 79914:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 79915:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 79916:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 79917:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 79918:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 79919:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 79920:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 79921:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 79922:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 79923:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 79924:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 79925:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 79926:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 79927:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 79928:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 79929:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 79930:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 79931:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 79932:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 79933:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 79934:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 79935:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 79936:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 79937:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 79938:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 79939:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 79940:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 79941:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 79942:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 79943:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 79944:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 79945:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 79946:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 79947:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 79948:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 79949:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 79950:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 79951:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 79952:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 79953:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 79954:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 79955:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 79956:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 79957:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 79958:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 79959:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 79960:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 79961:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 79962:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 79963:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 79964:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 79965:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 79966:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 79967:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 79968:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 79969:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 79970:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 79971:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 79972:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 79973:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 79974:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 79975:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 79976:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 79977:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 79978:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 79979:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 79980:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 79981:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 79982:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 79983:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 79984:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 79985:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 79986:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 79987:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 79988:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 79989:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 79990:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 79991:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 79992:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 79993:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 79994:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 79995:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 79996:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 79997:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 79998:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 79999:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 80000:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 80001:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 80002:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 80003:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 80004:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 80005:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 80006:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 80007:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 80008:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 80009:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 80010:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 80011:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 80012:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 80013:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 80014:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 80015:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 80016:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 80017:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 80018:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 80019:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 80020:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 80021:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 80022:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 80023:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 80024:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 80025:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 80026:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 80027:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 80028:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 80029:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 80030:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 80031:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 80032:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 80033:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 80034:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 80035:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 80036:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 80037:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 80038:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 80039:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 80040:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 80041:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 80042:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 80043:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 80044:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 80045:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 80046:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 80047:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 80048:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 80049:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 80050:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 80051:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 80052:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 80053:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 80054:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 80055:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 80056:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 80057:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 80058:22]
  assign io_z = ~x110; // @[Snxn100k.scala 80059:17]
endmodule
module SnxnLv4Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 79246:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 79247:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 79248:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 79249:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 79250:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 79251:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 79252:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 79253:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 79254:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 79255:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 79256:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 79257:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 79258:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 79259:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 79260:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 79261:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 79262:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 79263:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 79264:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 79265:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 79266:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 79267:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 79268:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 79269:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 79270:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 79271:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 79272:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 79273:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 79274:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 79275:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 79276:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 79277:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 79278:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 79279:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 79280:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 79281:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 79282:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 79283:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 79284:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 79285:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 79286:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 79287:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 79288:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 79289:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 79290:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 79291:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 79292:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 79293:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 79294:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 79295:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 79296:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 79297:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 79298:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 79299:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 79300:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 79301:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 79302:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 79303:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 79304:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 79305:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 79306:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 79307:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 79308:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 79309:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 79310:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 79311:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 79312:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 79313:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 79314:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 79315:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 79316:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 79317:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 79318:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 79319:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 79320:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 79321:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 79322:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 79323:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 79324:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 79325:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 79326:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 79327:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 79328:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 79329:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 79330:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 79331:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 79332:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 79333:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 79334:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 79335:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 79336:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 79337:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 79338:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 79339:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 79340:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 79341:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 79342:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 79343:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 79344:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 79345:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 79346:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 79347:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 79348:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 79349:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 79350:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 79351:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 79352:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 79353:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 79354:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 79355:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 79356:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 79357:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 79358:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 79359:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 79360:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 79361:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 79362:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 79363:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 79364:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 79365:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 79366:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 79367:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 79368:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 79369:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 79370:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 79371:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 79372:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79373:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79374:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79375:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79376:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79377:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79378:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79379:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79380:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79381:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79382:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79383:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79384:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79385:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79386:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79387:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79388:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79389:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79390:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79391:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79392:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79393:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79394:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79395:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79396:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79397:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79398:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79399:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79400:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79401:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79402:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79403:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79404:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79405:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79406:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79407:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79408:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79409:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79410:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79411:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79412:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79413:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79414:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79415:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79416:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79417:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79418:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79419:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79420:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79421:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79422:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79423:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79424:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79425:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79426:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79427:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79428:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79429:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79430:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79431:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79432:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79433:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79434:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79435:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79436:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79437:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79438:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79439:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79440:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79441:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79442:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79443:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79444:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 79445:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 79446:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 79447:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 79448:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 79449:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 79450:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 79451:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 79452:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 79453:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 79454:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 79455:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 79456:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 79457:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 79458:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 79459:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 79460:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 79461:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 79462:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 79463:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 79464:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 79465:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 79466:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 79467:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 79468:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 79469:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 79470:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 79471:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 79472:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 79473:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 79474:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 79475:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 79476:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 79477:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 79478:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 79479:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 79480:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 79481:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 79482:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 79483:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 79484:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 79485:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 79486:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 79487:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 79488:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 79489:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 79490:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 79491:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 79492:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 79493:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 79494:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 79495:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 79496:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 79497:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 79498:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 79499:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 79500:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 79501:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 79502:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 79503:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 79504:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 79505:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 79506:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 79507:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 79508:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 79509:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 79510:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 79511:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 79512:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 79513:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 79514:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 79515:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 79516:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 79517:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 79518:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 79519:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 79520:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 79521:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 79522:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 79523:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 79524:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 79525:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 79526:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 79527:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 79528:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 79529:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 79530:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 79531:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 79532:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 79533:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 79534:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 79535:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 79536:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 79537:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 79538:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 79539:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 79540:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 79541:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 79542:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 79543:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 79544:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 79545:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 79546:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 79547:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 79548:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 79549:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 79550:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 79551:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 79552:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 79553:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 79554:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 79555:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 79556:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 79557:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 79558:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 79559:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 79560:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 79561:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 79562:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 79563:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 79564:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 79565:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 79566:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 79567:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 79568:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 79569:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 79570:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 79571:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 79572:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 79573:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 79574:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 79575:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 79576:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 79577:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 79578:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 79579:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 79580:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 79581:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 79582:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 79583:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 79584:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 79585:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 79586:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 79587:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 79588:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 79589:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 79590:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 79591:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 79592:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 79593:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 79594:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 79595:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 79596:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 79597:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 79598:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 79599:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 79600:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 79601:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 79602:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 79603:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 79604:20]
  assign io_z = ~x89; // @[Snxn100k.scala 79605:16]
endmodule
module SnxnLv3Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst8_io_a; // @[Snxn100k.scala 20856:33]
  wire  inst_SnxnLv4Inst8_io_b; // @[Snxn100k.scala 20856:33]
  wire  inst_SnxnLv4Inst8_io_z; // @[Snxn100k.scala 20856:33]
  wire  inst_SnxnLv4Inst9_io_a; // @[Snxn100k.scala 20860:33]
  wire  inst_SnxnLv4Inst9_io_b; // @[Snxn100k.scala 20860:33]
  wire  inst_SnxnLv4Inst9_io_z; // @[Snxn100k.scala 20860:33]
  wire  inst_SnxnLv4Inst10_io_a; // @[Snxn100k.scala 20864:34]
  wire  inst_SnxnLv4Inst10_io_b; // @[Snxn100k.scala 20864:34]
  wire  inst_SnxnLv4Inst10_io_z; // @[Snxn100k.scala 20864:34]
  wire  inst_SnxnLv4Inst11_io_a; // @[Snxn100k.scala 20868:34]
  wire  inst_SnxnLv4Inst11_io_b; // @[Snxn100k.scala 20868:34]
  wire  inst_SnxnLv4Inst11_io_z; // @[Snxn100k.scala 20868:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst8_io_z + inst_SnxnLv4Inst9_io_z; // @[Snxn100k.scala 20872:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst10_io_z; // @[Snxn100k.scala 20872:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst11_io_z; // @[Snxn100k.scala 20872:87]
  SnxnLv4Inst8 inst_SnxnLv4Inst8 ( // @[Snxn100k.scala 20856:33]
    .io_a(inst_SnxnLv4Inst8_io_a),
    .io_b(inst_SnxnLv4Inst8_io_b),
    .io_z(inst_SnxnLv4Inst8_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst9 ( // @[Snxn100k.scala 20860:33]
    .io_a(inst_SnxnLv4Inst9_io_a),
    .io_b(inst_SnxnLv4Inst9_io_b),
    .io_z(inst_SnxnLv4Inst9_io_z)
  );
  SnxnLv4Inst10 inst_SnxnLv4Inst10 ( // @[Snxn100k.scala 20864:34]
    .io_a(inst_SnxnLv4Inst10_io_a),
    .io_b(inst_SnxnLv4Inst10_io_b),
    .io_z(inst_SnxnLv4Inst10_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst11 ( // @[Snxn100k.scala 20868:34]
    .io_a(inst_SnxnLv4Inst11_io_a),
    .io_b(inst_SnxnLv4Inst11_io_b),
    .io_z(inst_SnxnLv4Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 20873:15]
  assign inst_SnxnLv4Inst8_io_a = io_a; // @[Snxn100k.scala 20857:26]
  assign inst_SnxnLv4Inst8_io_b = io_b; // @[Snxn100k.scala 20858:26]
  assign inst_SnxnLv4Inst9_io_a = io_a; // @[Snxn100k.scala 20861:26]
  assign inst_SnxnLv4Inst9_io_b = io_b; // @[Snxn100k.scala 20862:26]
  assign inst_SnxnLv4Inst10_io_a = io_a; // @[Snxn100k.scala 20865:27]
  assign inst_SnxnLv4Inst10_io_b = io_b; // @[Snxn100k.scala 20866:27]
  assign inst_SnxnLv4Inst11_io_a = io_a; // @[Snxn100k.scala 20869:27]
  assign inst_SnxnLv4Inst11_io_b = io_b; // @[Snxn100k.scala 20870:27]
endmodule
module SnxnLv4Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82106:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82107:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82108:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82109:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82110:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82111:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82112:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82113:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82114:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82115:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82116:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82117:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82118:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82119:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82120:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82121:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82122:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82123:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82124:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 82125:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 82126:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 82127:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 82128:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 82129:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 82130:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 82131:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 82132:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 82133:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 82134:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 82135:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 82136:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 82137:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 82138:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 82139:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 82140:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 82141:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 82142:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 82143:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 82144:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 82145:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 82146:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 82147:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 82148:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 82149:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 82150:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 82151:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 82152:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 82153:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 82154:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 82155:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 82156:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 82157:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 82158:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 82159:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 82160:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 82161:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 82162:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 82163:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 82164:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 82165:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 82166:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 82167:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 82168:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 82169:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 82170:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 82171:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 82172:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 82173:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 82174:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 82175:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 82176:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 82177:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 82178:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 82179:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 82180:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 82181:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 82182:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 82183:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 82184:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 82185:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82186:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82187:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82188:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82189:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82190:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82191:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82192:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82193:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82194:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82195:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82196:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82197:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82198:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82199:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82200:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82201:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82202:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82203:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82204:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82205:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82206:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82207:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82208:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82209:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82210:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82211:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82212:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82213:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82214:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82215:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82216:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82217:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82218:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82219:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82220:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82221:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82222:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82223:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82224:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82225:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82226:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82227:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82228:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82229:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82230:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82231:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82232:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82233:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82234:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82235:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82236:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82237:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82238:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82239:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82240:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82241:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82242:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82243:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82244:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82245:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82246:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82247:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82248:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82249:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82250:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82251:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82252:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82253:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82254:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82255:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82256:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82257:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82258:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82259:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82260:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82261:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82262:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82263:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82264:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82265:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82266:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82267:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82268:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82269:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82270:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82271:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82272:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82273:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82274:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82275:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82276:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82277:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82278:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82279:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82280:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 82281:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 82282:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 82283:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 82284:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 82285:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 82286:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 82287:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 82288:20]
  assign io_z = ~x45; // @[Snxn100k.scala 82289:16]
endmodule
module SnxnLv4Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81920:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81921:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81922:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81923:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81924:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81925:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81926:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81927:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81928:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81929:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81930:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81931:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81932:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81933:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81934:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81935:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81936:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81937:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81938:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81939:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81940:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81941:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81942:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81943:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81944:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81945:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81946:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81947:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81948:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81949:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81950:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81951:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81952:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81953:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81954:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81955:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81956:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81957:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81958:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81959:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81960:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81961:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81962:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81963:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81964:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81965:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81966:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81967:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81968:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81969:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81970:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81971:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81972:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81973:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81974:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81975:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81976:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81977:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81978:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81979:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81980:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81981:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81982:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81983:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81984:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81985:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81986:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81987:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81988:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81989:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81990:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81991:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81992:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81993:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81994:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81995:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81996:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81997:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81998:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81999:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82000:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82001:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82002:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82003:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82004:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82005:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82006:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82007:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82008:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82009:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82010:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82011:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82012:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82013:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82014:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82015:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82016:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82017:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82018:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82019:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82020:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82021:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82022:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82023:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82024:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82025:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82026:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82027:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82028:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82029:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82030:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82031:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82032:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82033:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82034:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82035:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82036:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82037:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82038:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82039:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82040:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82041:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82042:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82043:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82044:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82045:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82046:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82047:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82048:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82049:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82050:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82051:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82052:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82053:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82054:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82055:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82056:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82057:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82058:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82059:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82060:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82061:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82062:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82063:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82064:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82065:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82066:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82067:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82068:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82069:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82070:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82071:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82072:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82073:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82074:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82075:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82076:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82077:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82078:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82079:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82080:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82081:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82082:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82083:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82084:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82085:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82086:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82087:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82088:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82089:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82090:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82091:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82092:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82093:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82094:20]
  assign io_z = ~x43; // @[Snxn100k.scala 82095:16]
endmodule
module SnxnLv4Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82300:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82301:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82302:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82303:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82304:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82305:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82306:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82307:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82308:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82309:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82310:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82311:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82312:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82313:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82314:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82315:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82316:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82317:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82318:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 82319:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 82320:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 82321:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 82322:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 82323:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 82324:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 82325:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 82326:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 82327:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 82328:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 82329:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 82330:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 82331:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 82332:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 82333:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 82334:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 82335:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 82336:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 82337:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 82338:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 82339:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 82340:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 82341:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 82342:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 82343:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 82344:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 82345:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 82346:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 82347:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 82348:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 82349:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 82350:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 82351:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 82352:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 82353:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 82354:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 82355:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 82356:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 82357:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 82358:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 82359:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 82360:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 82361:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 82362:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 82363:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 82364:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 82365:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 82366:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 82367:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 82368:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 82369:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 82370:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 82371:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 82372:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 82373:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 82374:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 82375:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 82376:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 82377:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 82378:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 82379:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82380:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82381:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82382:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82383:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82384:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82385:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82386:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82387:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82388:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82389:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82390:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82391:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82392:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82393:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82394:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82395:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82396:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82397:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82398:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82399:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82400:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82401:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82402:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82403:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82404:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82405:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82406:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82407:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82408:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82409:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82410:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82411:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82412:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82413:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82414:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82415:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82416:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82417:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82418:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82419:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82420:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82421:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82422:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82423:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82424:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82425:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82426:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82427:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82428:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82429:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82430:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82431:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82432:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82433:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82434:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82435:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82436:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82437:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82438:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82439:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82440:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82441:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82442:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82443:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82444:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82445:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82446:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82447:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82448:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82449:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82450:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82451:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82452:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82453:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82454:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82455:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82456:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82457:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82458:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82459:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82460:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82461:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82462:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82463:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82464:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82465:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82466:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82467:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82468:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82469:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82470:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82471:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82472:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82473:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82474:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 82475:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 82476:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 82477:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 82478:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 82479:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 82480:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 82481:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 82482:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 82483:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 82484:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 82485:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 82486:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 82487:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 82488:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 82489:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 82490:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 82491:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 82492:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 82493:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 82494:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 82495:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 82496:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 82497:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 82498:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 82499:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 82500:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 82501:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 82502:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 82503:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 82504:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 82505:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 82506:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 82507:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 82508:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 82509:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 82510:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 82511:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 82512:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 82513:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 82514:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 82515:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 82516:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 82517:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 82518:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 82519:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 82520:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 82521:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 82522:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 82523:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 82524:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 82525:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 82526:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 82527:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 82528:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 82529:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 82530:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 82531:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 82532:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 82533:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 82534:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 82535:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 82536:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 82537:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 82538:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 82539:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 82540:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 82541:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 82542:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 82543:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 82544:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 82545:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 82546:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 82547:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 82548:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 82549:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 82550:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 82551:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 82552:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 82553:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 82554:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 82555:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 82556:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 82557:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 82558:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 82559:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 82560:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 82561:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 82562:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 82563:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 82564:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 82565:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 82566:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 82567:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 82568:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 82569:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 82570:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 82571:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 82572:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 82573:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 82574:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 82575:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 82576:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 82577:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 82578:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 82579:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 82580:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 82581:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 82582:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 82583:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 82584:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 82585:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 82586:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 82587:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 82588:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 82589:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 82590:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 82591:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 82592:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 82593:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 82594:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 82595:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 82596:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 82597:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 82598:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 82599:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 82600:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 82601:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 82602:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 82603:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 82604:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 82605:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 82606:20]
  assign io_z = ~x76; // @[Snxn100k.scala 82607:16]
endmodule
module SnxnLv3Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst12_io_a; // @[Snxn100k.scala 21462:34]
  wire  inst_SnxnLv4Inst12_io_b; // @[Snxn100k.scala 21462:34]
  wire  inst_SnxnLv4Inst12_io_z; // @[Snxn100k.scala 21462:34]
  wire  inst_SnxnLv4Inst13_io_a; // @[Snxn100k.scala 21466:34]
  wire  inst_SnxnLv4Inst13_io_b; // @[Snxn100k.scala 21466:34]
  wire  inst_SnxnLv4Inst13_io_z; // @[Snxn100k.scala 21466:34]
  wire  inst_SnxnLv4Inst14_io_a; // @[Snxn100k.scala 21470:34]
  wire  inst_SnxnLv4Inst14_io_b; // @[Snxn100k.scala 21470:34]
  wire  inst_SnxnLv4Inst14_io_z; // @[Snxn100k.scala 21470:34]
  wire  inst_SnxnLv4Inst15_io_a; // @[Snxn100k.scala 21474:34]
  wire  inst_SnxnLv4Inst15_io_b; // @[Snxn100k.scala 21474:34]
  wire  inst_SnxnLv4Inst15_io_z; // @[Snxn100k.scala 21474:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst12_io_z + inst_SnxnLv4Inst13_io_z; // @[Snxn100k.scala 21478:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst14_io_z; // @[Snxn100k.scala 21478:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst15_io_z; // @[Snxn100k.scala 21478:89]
  SnxnLv4Inst12 inst_SnxnLv4Inst12 ( // @[Snxn100k.scala 21462:34]
    .io_a(inst_SnxnLv4Inst12_io_a),
    .io_b(inst_SnxnLv4Inst12_io_b),
    .io_z(inst_SnxnLv4Inst12_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst13 ( // @[Snxn100k.scala 21466:34]
    .io_a(inst_SnxnLv4Inst13_io_a),
    .io_b(inst_SnxnLv4Inst13_io_b),
    .io_z(inst_SnxnLv4Inst13_io_z)
  );
  SnxnLv4Inst14 inst_SnxnLv4Inst14 ( // @[Snxn100k.scala 21470:34]
    .io_a(inst_SnxnLv4Inst14_io_a),
    .io_b(inst_SnxnLv4Inst14_io_b),
    .io_z(inst_SnxnLv4Inst14_io_z)
  );
  SnxnLv4Inst15 inst_SnxnLv4Inst15 ( // @[Snxn100k.scala 21474:34]
    .io_a(inst_SnxnLv4Inst15_io_a),
    .io_b(inst_SnxnLv4Inst15_io_b),
    .io_z(inst_SnxnLv4Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21479:15]
  assign inst_SnxnLv4Inst12_io_a = io_a; // @[Snxn100k.scala 21463:27]
  assign inst_SnxnLv4Inst12_io_b = io_b; // @[Snxn100k.scala 21464:27]
  assign inst_SnxnLv4Inst13_io_a = io_a; // @[Snxn100k.scala 21467:27]
  assign inst_SnxnLv4Inst13_io_b = io_b; // @[Snxn100k.scala 21468:27]
  assign inst_SnxnLv4Inst14_io_a = io_a; // @[Snxn100k.scala 21471:27]
  assign inst_SnxnLv4Inst14_io_b = io_b; // @[Snxn100k.scala 21472:27]
  assign inst_SnxnLv4Inst15_io_a = io_a; // @[Snxn100k.scala 21475:27]
  assign inst_SnxnLv4Inst15_io_b = io_b; // @[Snxn100k.scala 21476:27]
endmodule
module SnxnLv2Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst0_io_a; // @[Snxn100k.scala 4862:33]
  wire  inst_SnxnLv3Inst0_io_b; // @[Snxn100k.scala 4862:33]
  wire  inst_SnxnLv3Inst0_io_z; // @[Snxn100k.scala 4862:33]
  wire  inst_SnxnLv3Inst1_io_a; // @[Snxn100k.scala 4866:33]
  wire  inst_SnxnLv3Inst1_io_b; // @[Snxn100k.scala 4866:33]
  wire  inst_SnxnLv3Inst1_io_z; // @[Snxn100k.scala 4866:33]
  wire  inst_SnxnLv3Inst2_io_a; // @[Snxn100k.scala 4870:33]
  wire  inst_SnxnLv3Inst2_io_b; // @[Snxn100k.scala 4870:33]
  wire  inst_SnxnLv3Inst2_io_z; // @[Snxn100k.scala 4870:33]
  wire  inst_SnxnLv3Inst3_io_a; // @[Snxn100k.scala 4874:33]
  wire  inst_SnxnLv3Inst3_io_b; // @[Snxn100k.scala 4874:33]
  wire  inst_SnxnLv3Inst3_io_z; // @[Snxn100k.scala 4874:33]
  wire  _sum_T_1 = inst_SnxnLv3Inst0_io_z + inst_SnxnLv3Inst1_io_z; // @[Snxn100k.scala 4878:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst2_io_z; // @[Snxn100k.scala 4878:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst3_io_z; // @[Snxn100k.scala 4878:86]
  SnxnLv3Inst0 inst_SnxnLv3Inst0 ( // @[Snxn100k.scala 4862:33]
    .io_a(inst_SnxnLv3Inst0_io_a),
    .io_b(inst_SnxnLv3Inst0_io_b),
    .io_z(inst_SnxnLv3Inst0_io_z)
  );
  SnxnLv3Inst1 inst_SnxnLv3Inst1 ( // @[Snxn100k.scala 4866:33]
    .io_a(inst_SnxnLv3Inst1_io_a),
    .io_b(inst_SnxnLv3Inst1_io_b),
    .io_z(inst_SnxnLv3Inst1_io_z)
  );
  SnxnLv3Inst2 inst_SnxnLv3Inst2 ( // @[Snxn100k.scala 4870:33]
    .io_a(inst_SnxnLv3Inst2_io_a),
    .io_b(inst_SnxnLv3Inst2_io_b),
    .io_z(inst_SnxnLv3Inst2_io_z)
  );
  SnxnLv3Inst3 inst_SnxnLv3Inst3 ( // @[Snxn100k.scala 4874:33]
    .io_a(inst_SnxnLv3Inst3_io_a),
    .io_b(inst_SnxnLv3Inst3_io_b),
    .io_z(inst_SnxnLv3Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 4879:15]
  assign inst_SnxnLv3Inst0_io_a = io_a; // @[Snxn100k.scala 4863:26]
  assign inst_SnxnLv3Inst0_io_b = io_b; // @[Snxn100k.scala 4864:26]
  assign inst_SnxnLv3Inst1_io_a = io_a; // @[Snxn100k.scala 4867:26]
  assign inst_SnxnLv3Inst1_io_b = io_b; // @[Snxn100k.scala 4868:26]
  assign inst_SnxnLv3Inst2_io_a = io_a; // @[Snxn100k.scala 4871:26]
  assign inst_SnxnLv3Inst2_io_b = io_b; // @[Snxn100k.scala 4872:26]
  assign inst_SnxnLv3Inst3_io_a = io_a; // @[Snxn100k.scala 4875:26]
  assign inst_SnxnLv3Inst3_io_b = io_b; // @[Snxn100k.scala 4876:26]
endmodule
module SnxnLv4Inst16(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 69084:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 69085:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 69086:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 69087:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 69088:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 69089:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 69090:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 69091:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 69092:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 69093:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 69094:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 69095:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 69096:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 69097:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 69098:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 69099:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 69100:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 69101:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 69102:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 69103:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 69104:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 69105:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 69106:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 69107:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 69108:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 69109:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 69110:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 69111:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 69112:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 69113:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 69114:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 69115:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 69116:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 69117:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 69118:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 69119:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 69120:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 69121:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 69122:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 69123:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 69124:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 69125:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 69126:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 69127:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 69128:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 69129:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 69130:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 69131:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 69132:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 69133:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 69134:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 69135:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 69136:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 69137:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 69138:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 69139:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 69140:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 69141:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 69142:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 69143:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 69144:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 69145:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 69146:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 69147:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 69148:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 69149:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 69150:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 69151:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 69152:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 69153:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 69154:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 69155:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 69156:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 69157:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 69158:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 69159:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 69160:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 69161:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 69162:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 69163:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 69164:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 69165:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 69166:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 69167:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 69168:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 69169:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 69170:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 69171:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 69172:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 69173:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 69174:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 69175:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 69176:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 69177:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 69178:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 69179:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 69180:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 69181:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 69182:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 69183:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 69184:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 69185:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 69186:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 69187:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 69188:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 69189:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 69190:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 69191:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 69192:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 69193:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 69194:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 69195:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 69196:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 69197:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 69198:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 69199:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 69200:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 69201:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69202:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69203:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69204:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69205:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69206:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69207:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69208:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69209:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69210:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69211:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69212:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69213:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69214:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69215:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69216:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69217:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69218:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69219:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69220:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69221:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69222:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69223:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69224:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69225:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69226:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69227:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69228:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69229:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69230:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69231:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69232:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69233:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69234:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69235:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69236:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69237:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69238:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69239:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69240:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69241:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69242:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69243:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69244:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69245:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69246:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69247:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69248:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69249:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69250:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69251:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69252:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69253:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69254:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69255:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69256:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69257:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69258:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69259:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69260:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69261:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69262:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69263:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69264:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69265:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69266:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69267:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69268:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69269:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69270:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69271:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69272:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69273:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69274:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 69275:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 69276:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 69277:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 69278:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 69279:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 69280:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 69281:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 69282:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 69283:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 69284:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 69285:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 69286:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 69287:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 69288:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 69289:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 69290:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 69291:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 69292:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 69293:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 69294:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 69295:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 69296:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 69297:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 69298:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 69299:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 69300:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 69301:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 69302:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 69303:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 69304:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 69305:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 69306:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 69307:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 69308:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 69309:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 69310:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 69311:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 69312:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 69313:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 69314:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 69315:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 69316:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 69317:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 69318:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 69319:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 69320:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 69321:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 69322:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 69323:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 69324:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 69325:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 69326:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 69327:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 69328:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 69329:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 69330:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 69331:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 69332:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 69333:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 69334:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 69335:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 69336:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 69337:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 69338:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 69339:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 69340:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 69341:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 69342:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 69343:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 69344:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 69345:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 69346:20]
  assign io_z = ~x65; // @[Snxn100k.scala 69347:16]
endmodule
module SnxnLv4Inst17(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 68882:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 68883:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 68884:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 68885:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 68886:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 68887:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 68888:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 68889:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 68890:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 68891:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 68892:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 68893:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 68894:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 68895:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 68896:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 68897:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 68898:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 68899:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 68900:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 68901:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 68902:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 68903:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 68904:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 68905:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 68906:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 68907:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 68908:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 68909:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 68910:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 68911:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 68912:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 68913:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 68914:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 68915:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 68916:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 68917:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 68918:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 68919:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 68920:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 68921:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 68922:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 68923:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 68924:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 68925:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 68926:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 68927:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 68928:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 68929:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 68930:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 68931:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 68932:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 68933:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 68934:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 68935:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 68936:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 68937:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 68938:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 68939:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 68940:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 68941:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 68942:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 68943:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 68944:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 68945:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 68946:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 68947:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 68948:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 68949:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 68950:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 68951:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 68952:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 68953:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 68954:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 68955:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 68956:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 68957:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 68958:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 68959:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 68960:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 68961:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 68962:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 68963:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 68964:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 68965:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 68966:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 68967:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 68968:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 68969:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 68970:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 68971:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 68972:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 68973:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 68974:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 68975:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 68976:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 68977:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 68978:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 68979:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 68980:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 68981:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 68982:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 68983:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 68984:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 68985:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 68986:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 68987:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 68988:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 68989:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 68990:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 68991:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 68992:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 68993:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 68994:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 68995:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 68996:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 68997:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 68998:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 68999:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69000:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69001:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69002:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69003:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69004:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69005:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69006:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69007:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69008:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69009:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69010:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69011:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69012:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69013:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69014:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69015:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69016:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69017:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69018:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69019:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69020:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69021:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69022:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69023:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69024:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69025:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69026:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69027:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69028:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69029:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69030:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69031:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69032:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69033:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69034:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69035:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69036:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69037:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69038:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69039:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69040:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69041:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69042:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69043:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69044:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69045:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69046:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69047:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69048:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69049:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69050:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69051:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69052:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69053:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69054:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69055:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69056:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69057:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69058:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69059:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69060:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69061:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69062:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69063:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69064:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69065:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69066:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69067:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69068:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69069:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69070:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69071:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69072:20]
  assign io_z = ~x47; // @[Snxn100k.scala 69073:16]
endmodule
module SnxnLv4Inst18(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 68768:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 68769:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 68770:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 68771:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 68772:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 68773:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 68774:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 68775:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 68776:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 68777:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 68778:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 68779:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 68780:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 68781:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 68782:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 68783:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 68784:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 68785:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 68786:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 68787:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 68788:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 68789:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 68790:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 68791:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 68792:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 68793:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 68794:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 68795:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 68796:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 68797:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 68798:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 68799:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 68800:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 68801:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 68802:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 68803:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 68804:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 68805:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 68806:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 68807:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 68808:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 68809:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 68810:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 68811:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 68812:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 68813:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 68814:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 68815:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 68816:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 68817:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 68818:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 68819:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 68820:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 68821:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 68822:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 68823:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 68824:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 68825:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 68826:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 68827:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 68828:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 68829:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 68830:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 68831:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 68832:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 68833:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 68834:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 68835:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 68836:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 68837:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 68838:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 68839:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 68840:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 68841:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 68842:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 68843:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 68844:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 68845:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 68846:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 68847:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 68848:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 68849:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 68850:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 68851:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 68852:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 68853:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 68854:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 68855:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 68856:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 68857:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 68858:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 68859:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 68860:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 68861:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 68862:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 68863:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 68864:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 68865:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 68866:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 68867:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 68868:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 68869:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 68870:20]
  assign io_z = ~x25; // @[Snxn100k.scala 68871:16]
endmodule
module SnxnLv4Inst19(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 69358:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 69359:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 69360:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 69361:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 69362:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 69363:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 69364:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 69365:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 69366:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 69367:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 69368:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 69369:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 69370:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 69371:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 69372:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 69373:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 69374:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 69375:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 69376:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 69377:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 69378:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 69379:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 69380:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 69381:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 69382:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 69383:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 69384:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 69385:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 69386:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 69387:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 69388:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 69389:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 69390:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 69391:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 69392:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 69393:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 69394:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 69395:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 69396:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 69397:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 69398:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 69399:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 69400:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 69401:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 69402:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 69403:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 69404:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 69405:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 69406:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 69407:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 69408:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 69409:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 69410:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 69411:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 69412:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 69413:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 69414:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 69415:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 69416:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 69417:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 69418:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 69419:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 69420:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 69421:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 69422:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 69423:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 69424:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 69425:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 69426:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 69427:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 69428:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 69429:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 69430:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 69431:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 69432:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 69433:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 69434:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 69435:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 69436:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 69437:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 69438:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 69439:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 69440:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 69441:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 69442:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 69443:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 69444:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 69445:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 69446:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 69447:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 69448:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 69449:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 69450:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 69451:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 69452:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 69453:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 69454:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 69455:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 69456:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 69457:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 69458:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 69459:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 69460:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 69461:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 69462:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 69463:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 69464:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 69465:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 69466:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 69467:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 69468:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 69469:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 69470:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 69471:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 69472:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 69473:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 69474:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 69475:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69476:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69477:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69478:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69479:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69480:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69481:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69482:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69483:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69484:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69485:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69486:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69487:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69488:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69489:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69490:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69491:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69492:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69493:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69494:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69495:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69496:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69497:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69498:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69499:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69500:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69501:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69502:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69503:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69504:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69505:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69506:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69507:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69508:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69509:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69510:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69511:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69512:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69513:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69514:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69515:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69516:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69517:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69518:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69519:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69520:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69521:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69522:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69523:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69524:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69525:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69526:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69527:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69528:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69529:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69530:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69531:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69532:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69533:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69534:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69535:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69536:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69537:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69538:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69539:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69540:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69541:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69542:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69543:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69544:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69545:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69546:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69547:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69548:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 69549:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 69550:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 69551:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 69552:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 69553:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 69554:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 69555:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 69556:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 69557:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 69558:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 69559:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 69560:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 69561:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 69562:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 69563:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 69564:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 69565:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 69566:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 69567:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 69568:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 69569:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 69570:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 69571:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 69572:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 69573:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 69574:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 69575:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 69576:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 69577:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 69578:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 69579:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 69580:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 69581:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 69582:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 69583:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 69584:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 69585:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 69586:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 69587:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 69588:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 69589:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 69590:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 69591:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 69592:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 69593:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 69594:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 69595:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 69596:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 69597:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 69598:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 69599:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 69600:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 69601:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 69602:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 69603:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 69604:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 69605:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 69606:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 69607:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 69608:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 69609:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 69610:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 69611:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 69612:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 69613:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 69614:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 69615:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 69616:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 69617:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 69618:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 69619:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 69620:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 69621:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 69622:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 69623:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 69624:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 69625:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 69626:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 69627:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 69628:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 69629:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 69630:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 69631:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 69632:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 69633:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 69634:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 69635:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 69636:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 69637:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 69638:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 69639:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 69640:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 69641:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 69642:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 69643:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 69644:20]
  assign io_z = ~x71; // @[Snxn100k.scala 69645:16]
endmodule
module SnxnLv3Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst16_io_a; // @[Snxn100k.scala 18252:34]
  wire  inst_SnxnLv4Inst16_io_b; // @[Snxn100k.scala 18252:34]
  wire  inst_SnxnLv4Inst16_io_z; // @[Snxn100k.scala 18252:34]
  wire  inst_SnxnLv4Inst17_io_a; // @[Snxn100k.scala 18256:34]
  wire  inst_SnxnLv4Inst17_io_b; // @[Snxn100k.scala 18256:34]
  wire  inst_SnxnLv4Inst17_io_z; // @[Snxn100k.scala 18256:34]
  wire  inst_SnxnLv4Inst18_io_a; // @[Snxn100k.scala 18260:34]
  wire  inst_SnxnLv4Inst18_io_b; // @[Snxn100k.scala 18260:34]
  wire  inst_SnxnLv4Inst18_io_z; // @[Snxn100k.scala 18260:34]
  wire  inst_SnxnLv4Inst19_io_a; // @[Snxn100k.scala 18264:34]
  wire  inst_SnxnLv4Inst19_io_b; // @[Snxn100k.scala 18264:34]
  wire  inst_SnxnLv4Inst19_io_z; // @[Snxn100k.scala 18264:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst16_io_z + inst_SnxnLv4Inst17_io_z; // @[Snxn100k.scala 18268:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst18_io_z; // @[Snxn100k.scala 18268:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst19_io_z; // @[Snxn100k.scala 18268:89]
  SnxnLv4Inst16 inst_SnxnLv4Inst16 ( // @[Snxn100k.scala 18252:34]
    .io_a(inst_SnxnLv4Inst16_io_a),
    .io_b(inst_SnxnLv4Inst16_io_b),
    .io_z(inst_SnxnLv4Inst16_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst17 ( // @[Snxn100k.scala 18256:34]
    .io_a(inst_SnxnLv4Inst17_io_a),
    .io_b(inst_SnxnLv4Inst17_io_b),
    .io_z(inst_SnxnLv4Inst17_io_z)
  );
  SnxnLv4Inst18 inst_SnxnLv4Inst18 ( // @[Snxn100k.scala 18260:34]
    .io_a(inst_SnxnLv4Inst18_io_a),
    .io_b(inst_SnxnLv4Inst18_io_b),
    .io_z(inst_SnxnLv4Inst18_io_z)
  );
  SnxnLv4Inst19 inst_SnxnLv4Inst19 ( // @[Snxn100k.scala 18264:34]
    .io_a(inst_SnxnLv4Inst19_io_a),
    .io_b(inst_SnxnLv4Inst19_io_b),
    .io_z(inst_SnxnLv4Inst19_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 18269:15]
  assign inst_SnxnLv4Inst16_io_a = io_a; // @[Snxn100k.scala 18253:27]
  assign inst_SnxnLv4Inst16_io_b = io_b; // @[Snxn100k.scala 18254:27]
  assign inst_SnxnLv4Inst17_io_a = io_a; // @[Snxn100k.scala 18257:27]
  assign inst_SnxnLv4Inst17_io_b = io_b; // @[Snxn100k.scala 18258:27]
  assign inst_SnxnLv4Inst18_io_a = io_a; // @[Snxn100k.scala 18261:27]
  assign inst_SnxnLv4Inst18_io_b = io_b; // @[Snxn100k.scala 18262:27]
  assign inst_SnxnLv4Inst19_io_a = io_a; // @[Snxn100k.scala 18265:27]
  assign inst_SnxnLv4Inst19_io_b = io_b; // @[Snxn100k.scala 18266:27]
endmodule
module SnxnLv4Inst20(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71412:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71413:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71414:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71415:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71416:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71417:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71418:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71419:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71420:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71421:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71422:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71423:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71424:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71425:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71426:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71427:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71428:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71429:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71430:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71431:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71432:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71433:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71434:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71435:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71436:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71437:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71438:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71439:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71440:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71441:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71442:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71443:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71444:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71445:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71446:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71447:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71448:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71449:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71450:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71451:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71452:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71453:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71454:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71455:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71456:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71457:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71458:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71459:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71460:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71461:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71462:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71463:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71464:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71465:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71466:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71467:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71468:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71469:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71470:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71471:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71472:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71473:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71474:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71475:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71476:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71477:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71478:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71479:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71480:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71481:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71482:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71483:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71484:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71485:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71486:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71487:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71488:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71489:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71490:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71491:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71492:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71493:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71494:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71495:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71496:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71497:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71498:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71499:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71500:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71501:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71502:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71503:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71504:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71505:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71506:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71507:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71508:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71509:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71510:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71511:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71512:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71513:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71514:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71515:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71516:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71517:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71518:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71519:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71520:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71521:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71522:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71523:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71524:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71525:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71526:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71527:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71528:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71529:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71530:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71531:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71532:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71533:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71534:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71535:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71536:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71537:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71538:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71539:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71540:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71541:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71542:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71543:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71544:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71545:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71546:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71547:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71548:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71549:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71550:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 71551:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 71552:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 71553:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 71554:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 71555:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 71556:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 71557:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 71558:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 71559:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 71560:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 71561:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 71562:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 71563:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 71564:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 71565:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 71566:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 71567:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 71568:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 71569:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 71570:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 71571:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 71572:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 71573:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 71574:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 71575:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 71576:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 71577:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 71578:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 71579:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 71580:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 71581:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 71582:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 71583:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 71584:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 71585:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 71586:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 71587:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 71588:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 71589:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 71590:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 71591:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 71592:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 71593:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 71594:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 71595:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 71596:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 71597:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 71598:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 71599:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 71600:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 71601:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 71602:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 71603:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 71604:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 71605:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 71606:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 71607:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 71608:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 71609:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 71610:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 71611:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 71612:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 71613:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 71614:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 71615:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 71616:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 71617:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 71618:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 71619:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 71620:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 71621:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 71622:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 71623:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 71624:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 71625:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 71626:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 71627:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 71628:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 71629:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 71630:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 71631:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 71632:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 71633:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 71634:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 71635:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 71636:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 71637:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 71638:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 71639:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 71640:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 71641:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 71642:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 71643:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 71644:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 71645:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 71646:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 71647:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 71648:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 71649:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 71650:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 71651:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 71652:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 71653:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 71654:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 71655:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 71656:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 71657:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 71658:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 71659:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 71660:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 71661:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 71662:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 71663:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 71664:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 71665:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 71666:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 71667:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 71668:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 71669:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 71670:20]
  assign io_z = ~x64; // @[Snxn100k.scala 71671:16]
endmodule
module SnxnLv4Inst22(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71150:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71151:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71152:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71153:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71154:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71155:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71156:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71157:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71158:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71159:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71160:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71161:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71162:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71163:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71164:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71165:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71166:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71167:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71168:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71169:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71170:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71171:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71172:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71173:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71174:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71175:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71176:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71177:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71178:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71179:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71180:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71181:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71182:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71183:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71184:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71185:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71186:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71187:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71188:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71189:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71190:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71191:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71192:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71193:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71194:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71195:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71196:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71197:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71198:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71199:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71200:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71201:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71202:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71203:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71204:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71205:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71206:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71207:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71208:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71209:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71210:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71211:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71212:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71213:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71214:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71215:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71216:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71217:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71218:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71219:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71220:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71221:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71222:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71223:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71224:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71225:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71226:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71227:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71228:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71229:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71230:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71231:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71232:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71233:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71234:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71235:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71236:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71237:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71238:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71239:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71240:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71241:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71242:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71243:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71244:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71245:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71246:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71247:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71248:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71249:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71250:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71251:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71252:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71253:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71254:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71255:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71256:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71257:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71258:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71259:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71260:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71261:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71262:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71263:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71264:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71265:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71266:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71267:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71268:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71269:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71270:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71271:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71272:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71273:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71274:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71275:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71276:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71277:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71278:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71279:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71280:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71281:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71282:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71283:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71284:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71285:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71286:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71287:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71288:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 71289:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 71290:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 71291:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 71292:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 71293:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 71294:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 71295:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 71296:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 71297:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 71298:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 71299:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 71300:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 71301:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 71302:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 71303:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 71304:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 71305:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 71306:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 71307:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 71308:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 71309:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 71310:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 71311:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 71312:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 71313:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 71314:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 71315:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 71316:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 71317:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 71318:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 71319:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 71320:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 71321:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 71322:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 71323:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 71324:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 71325:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 71326:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 71327:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 71328:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 71329:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 71330:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 71331:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 71332:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 71333:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 71334:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 71335:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 71336:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 71337:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 71338:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 71339:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 71340:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 71341:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 71342:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 71343:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 71344:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 71345:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 71346:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 71347:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 71348:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 71349:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 71350:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 71351:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 71352:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 71353:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 71354:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 71355:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 71356:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 71357:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 71358:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 71359:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 71360:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 71361:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 71362:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 71363:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 71364:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 71365:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 71366:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 71367:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 71368:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 71369:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 71370:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 71371:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 71372:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 71373:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 71374:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 71375:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 71376:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 71377:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 71378:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 71379:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 71380:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 71381:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 71382:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 71383:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 71384:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 71385:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 71386:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 71387:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 71388:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 71389:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 71390:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 71391:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 71392:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 71393:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 71394:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 71395:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 71396:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 71397:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 71398:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 71399:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 71400:20]
  assign io_z = ~x62; // @[Snxn100k.scala 71401:16]
endmodule
module SnxnLv4Inst23(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71682:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71683:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71684:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71685:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71686:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71687:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71688:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71689:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71690:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71691:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71692:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71693:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71694:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71695:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71696:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71697:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71698:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71699:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71700:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71701:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71702:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71703:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71704:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71705:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71706:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71707:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71708:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71709:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71710:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71711:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71712:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71713:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71714:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71715:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71716:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71717:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71718:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71719:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71720:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71721:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71722:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71723:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71724:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71725:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71726:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71727:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71728:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71729:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71730:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71731:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71732:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71733:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71734:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71735:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71736:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71737:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71738:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71739:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71740:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71741:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71742:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71743:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71744:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71745:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71746:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71747:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71748:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71749:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71750:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71751:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71752:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71753:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71754:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71755:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71756:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71757:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71758:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71759:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71760:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71761:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71762:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71763:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71764:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71765:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71766:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71767:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71768:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71769:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71770:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71771:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71772:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71773:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71774:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71775:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71776:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71777:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71778:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71779:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71780:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71781:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71782:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71783:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71784:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71785:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71786:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71787:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71788:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71789:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71790:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71791:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71792:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71793:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71794:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71795:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71796:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71797:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71798:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71799:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71800:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71801:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71802:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71803:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71804:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71805:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71806:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71807:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71808:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71809:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71810:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71811:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71812:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71813:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71814:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71815:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71816:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71817:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71818:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71819:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71820:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 71821:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 71822:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 71823:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 71824:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 71825:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 71826:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 71827:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 71828:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 71829:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 71830:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 71831:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 71832:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 71833:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 71834:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 71835:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 71836:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 71837:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 71838:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 71839:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 71840:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 71841:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 71842:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 71843:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 71844:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 71845:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 71846:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 71847:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 71848:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 71849:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 71850:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 71851:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 71852:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 71853:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 71854:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 71855:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 71856:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 71857:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 71858:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 71859:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 71860:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 71861:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 71862:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 71863:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 71864:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 71865:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 71866:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 71867:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 71868:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 71869:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 71870:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 71871:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 71872:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 71873:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 71874:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 71875:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 71876:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 71877:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 71878:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 71879:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 71880:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 71881:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 71882:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 71883:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 71884:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 71885:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 71886:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 71887:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 71888:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 71889:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 71890:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 71891:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 71892:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 71893:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 71894:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 71895:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 71896:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 71897:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 71898:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 71899:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 71900:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 71901:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 71902:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 71903:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 71904:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 71905:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 71906:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 71907:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 71908:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 71909:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 71910:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 71911:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 71912:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 71913:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 71914:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 71915:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 71916:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 71917:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 71918:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 71919:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 71920:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 71921:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 71922:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 71923:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 71924:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 71925:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 71926:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 71927:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 71928:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 71929:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 71930:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 71931:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 71932:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 71933:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 71934:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 71935:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 71936:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 71937:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 71938:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 71939:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 71940:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 71941:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 71942:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 71943:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 71944:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 71945:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 71946:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 71947:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 71948:20]
  assign io_z = ~x66; // @[Snxn100k.scala 71949:16]
endmodule
module SnxnLv3Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst20_io_a; // @[Snxn100k.scala 18950:34]
  wire  inst_SnxnLv4Inst20_io_b; // @[Snxn100k.scala 18950:34]
  wire  inst_SnxnLv4Inst20_io_z; // @[Snxn100k.scala 18950:34]
  wire  inst_SnxnLv4Inst21_io_a; // @[Snxn100k.scala 18954:34]
  wire  inst_SnxnLv4Inst21_io_b; // @[Snxn100k.scala 18954:34]
  wire  inst_SnxnLv4Inst21_io_z; // @[Snxn100k.scala 18954:34]
  wire  inst_SnxnLv4Inst22_io_a; // @[Snxn100k.scala 18958:34]
  wire  inst_SnxnLv4Inst22_io_b; // @[Snxn100k.scala 18958:34]
  wire  inst_SnxnLv4Inst22_io_z; // @[Snxn100k.scala 18958:34]
  wire  inst_SnxnLv4Inst23_io_a; // @[Snxn100k.scala 18962:34]
  wire  inst_SnxnLv4Inst23_io_b; // @[Snxn100k.scala 18962:34]
  wire  inst_SnxnLv4Inst23_io_z; // @[Snxn100k.scala 18962:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst20_io_z + inst_SnxnLv4Inst21_io_z; // @[Snxn100k.scala 18966:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst22_io_z; // @[Snxn100k.scala 18966:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst23_io_z; // @[Snxn100k.scala 18966:89]
  SnxnLv4Inst20 inst_SnxnLv4Inst20 ( // @[Snxn100k.scala 18950:34]
    .io_a(inst_SnxnLv4Inst20_io_a),
    .io_b(inst_SnxnLv4Inst20_io_b),
    .io_z(inst_SnxnLv4Inst20_io_z)
  );
  SnxnLv4Inst18 inst_SnxnLv4Inst21 ( // @[Snxn100k.scala 18954:34]
    .io_a(inst_SnxnLv4Inst21_io_a),
    .io_b(inst_SnxnLv4Inst21_io_b),
    .io_z(inst_SnxnLv4Inst21_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst22 ( // @[Snxn100k.scala 18958:34]
    .io_a(inst_SnxnLv4Inst22_io_a),
    .io_b(inst_SnxnLv4Inst22_io_b),
    .io_z(inst_SnxnLv4Inst22_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst23 ( // @[Snxn100k.scala 18962:34]
    .io_a(inst_SnxnLv4Inst23_io_a),
    .io_b(inst_SnxnLv4Inst23_io_b),
    .io_z(inst_SnxnLv4Inst23_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 18967:15]
  assign inst_SnxnLv4Inst20_io_a = io_a; // @[Snxn100k.scala 18951:27]
  assign inst_SnxnLv4Inst20_io_b = io_b; // @[Snxn100k.scala 18952:27]
  assign inst_SnxnLv4Inst21_io_a = io_a; // @[Snxn100k.scala 18955:27]
  assign inst_SnxnLv4Inst21_io_b = io_b; // @[Snxn100k.scala 18956:27]
  assign inst_SnxnLv4Inst22_io_a = io_a; // @[Snxn100k.scala 18959:27]
  assign inst_SnxnLv4Inst22_io_b = io_b; // @[Snxn100k.scala 18960:27]
  assign inst_SnxnLv4Inst23_io_a = io_a; // @[Snxn100k.scala 18963:27]
  assign inst_SnxnLv4Inst23_io_b = io_b; // @[Snxn100k.scala 18964:27]
endmodule
module SnxnLv4Inst24(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72142:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72143:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72144:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72145:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72146:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72147:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72148:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 72149:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 72150:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 72151:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 72152:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 72153:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 72154:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 72155:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 72156:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 72157:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 72158:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 72159:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 72160:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 72161:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 72162:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 72163:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 72164:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 72165:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 72166:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72167:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72168:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72169:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 72170:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 72171:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 72172:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 72173:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 72174:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 72175:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 72176:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 72177:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 72178:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 72179:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 72180:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 72181:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72182:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72183:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72184:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72185:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72186:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72187:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72188:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72189:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72190:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72191:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72192:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72193:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72194:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72195:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72196:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72197:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72198:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72199:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72200:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72201:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72202:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72203:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72204:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72205:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72206:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72207:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72208:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72209:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72210:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72211:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72212:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72213:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72214:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72215:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72216:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72217:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72218:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72219:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72220:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72221:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72222:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72223:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72224:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72225:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72226:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72227:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72228:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72229:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72230:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72231:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72232:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72233:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72234:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72235:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72236:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72237:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72238:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72239:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72240:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 72241:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 72242:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 72243:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 72244:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 72245:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 72246:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 72247:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 72248:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 72249:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 72250:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 72251:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 72252:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 72253:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 72254:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 72255:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 72256:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 72257:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 72258:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 72259:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 72260:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 72261:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 72262:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 72263:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 72264:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 72265:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 72266:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 72267:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 72268:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 72269:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 72270:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 72271:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 72272:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 72273:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 72274:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 72275:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 72276:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 72277:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 72278:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 72279:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 72280:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 72281:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 72282:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 72283:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 72284:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 72285:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 72286:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 72287:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 72288:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 72289:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 72290:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 72291:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 72292:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 72293:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 72294:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 72295:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 72296:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 72297:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 72298:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 72299:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 72300:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 72301:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 72302:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 72303:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 72304:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 72305:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 72306:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 72307:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 72308:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 72309:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 72310:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 72311:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 72312:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 72313:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 72314:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 72315:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 72316:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 72317:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 72318:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 72319:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 72320:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 72321:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 72322:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 72323:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 72324:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 72325:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 72326:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 72327:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 72328:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 72329:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 72330:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 72331:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 72332:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 72333:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 72334:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 72335:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 72336:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 72337:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 72338:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 72339:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 72340:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 72341:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 72342:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 72343:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 72344:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 72345:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 72346:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 72347:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 72348:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 72349:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 72350:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 72351:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 72352:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 72353:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 72354:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 72355:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 72356:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 72357:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 72358:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 72359:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 72360:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 72361:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 72362:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 72363:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 72364:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 72365:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 72366:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 72367:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 72368:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 72369:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 72370:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 72371:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 72372:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 72373:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 72374:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 72375:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 72376:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 72377:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 72378:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 72379:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 72380:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 72381:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 72382:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 72383:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 72384:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 72385:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 72386:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 72387:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 72388:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 72389:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 72390:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 72391:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 72392:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 72393:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 72394:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 72395:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 72396:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 72397:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 72398:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 72399:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 72400:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 72401:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 72402:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 72403:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 72404:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 72405:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 72406:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 72407:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 72408:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 72409:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 72410:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 72411:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 72412:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 72413:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 72414:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 72415:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 72416:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 72417:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 72418:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 72419:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 72420:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 72421:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 72422:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 72423:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 72424:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 72425:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 72426:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 72427:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 72428:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 72429:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 72430:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 72431:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 72432:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 72433:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 72434:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 72435:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 72436:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 72437:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 72438:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 72439:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 72440:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 72441:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 72442:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 72443:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 72444:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 72445:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 72446:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 72447:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 72448:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 72449:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 72450:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 72451:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 72452:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 72453:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 72454:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 72455:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 72456:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 72457:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 72458:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 72459:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 72460:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 72461:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 72462:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 72463:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 72464:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 72465:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 72466:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 72467:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 72468:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 72469:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 72470:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 72471:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 72472:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 72473:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 72474:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 72475:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 72476:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 72477:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 72478:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 72479:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 72480:20]
  assign io_z = ~x84; // @[Snxn100k.scala 72481:16]
endmodule
module SnxnLv4Inst25(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72862:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72863:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72864:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72865:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72866:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72867:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72868:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 72869:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 72870:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 72871:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 72872:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 72873:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 72874:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 72875:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 72876:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 72877:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 72878:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 72879:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 72880:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 72881:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 72882:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 72883:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 72884:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 72885:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 72886:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72887:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72888:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72889:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 72890:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 72891:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 72892:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 72893:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 72894:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 72895:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 72896:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 72897:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 72898:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 72899:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 72900:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 72901:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72902:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72903:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72904:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72905:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72906:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72907:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72908:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72909:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72910:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72911:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72912:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72913:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72914:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72915:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72916:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72917:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72918:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72919:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72920:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72921:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72922:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72923:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72924:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72925:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72926:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72927:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72928:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72929:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72930:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72931:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72932:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72933:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72934:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72935:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72936:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72937:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72938:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72939:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72940:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72941:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72942:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72943:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72944:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72945:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72946:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72947:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72948:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72949:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72950:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72951:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72952:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72953:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72954:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72955:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72956:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72957:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72958:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72959:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72960:20]
  assign io_z = ~x24; // @[Snxn100k.scala 72961:16]
endmodule
module SnxnLv4Inst26(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71960:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71961:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71962:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71963:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71964:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71965:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71966:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71967:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71968:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71969:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71970:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71971:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71972:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71973:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71974:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71975:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71976:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71977:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71978:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71979:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71980:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71981:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71982:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71983:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71984:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71985:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71986:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71987:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71988:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71989:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71990:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71991:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71992:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71993:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71994:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71995:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71996:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71997:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71998:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71999:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72000:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72001:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72002:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72003:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72004:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72005:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72006:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72007:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72008:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72009:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72010:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72011:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72012:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72013:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72014:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72015:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72016:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72017:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72018:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72019:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72020:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72021:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72022:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72023:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72024:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72025:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72026:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72027:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72028:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72029:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72030:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72031:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72032:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72033:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72034:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72035:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72036:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72037:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72038:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72039:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72040:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72041:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72042:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72043:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72044:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72045:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72046:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72047:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72048:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72049:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72050:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72051:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72052:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72053:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72054:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72055:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72056:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72057:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72058:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 72059:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 72060:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 72061:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 72062:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 72063:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 72064:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 72065:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 72066:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 72067:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 72068:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 72069:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 72070:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 72071:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 72072:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 72073:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 72074:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 72075:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 72076:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 72077:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 72078:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 72079:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 72080:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 72081:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 72082:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 72083:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 72084:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 72085:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 72086:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 72087:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 72088:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 72089:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 72090:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 72091:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 72092:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 72093:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 72094:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 72095:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 72096:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 72097:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 72098:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 72099:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 72100:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 72101:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 72102:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 72103:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 72104:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 72105:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 72106:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 72107:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 72108:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 72109:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 72110:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 72111:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 72112:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 72113:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 72114:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 72115:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 72116:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 72117:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 72118:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 72119:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 72120:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 72121:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 72122:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 72123:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 72124:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 72125:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 72126:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 72127:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 72128:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 72129:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 72130:20]
  assign io_z = ~x42; // @[Snxn100k.scala 72131:16]
endmodule
module SnxnLv3Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst24_io_a; // @[Snxn100k.scala 19405:34]
  wire  inst_SnxnLv4Inst24_io_b; // @[Snxn100k.scala 19405:34]
  wire  inst_SnxnLv4Inst24_io_z; // @[Snxn100k.scala 19405:34]
  wire  inst_SnxnLv4Inst25_io_a; // @[Snxn100k.scala 19409:34]
  wire  inst_SnxnLv4Inst25_io_b; // @[Snxn100k.scala 19409:34]
  wire  inst_SnxnLv4Inst25_io_z; // @[Snxn100k.scala 19409:34]
  wire  inst_SnxnLv4Inst26_io_a; // @[Snxn100k.scala 19413:34]
  wire  inst_SnxnLv4Inst26_io_b; // @[Snxn100k.scala 19413:34]
  wire  inst_SnxnLv4Inst26_io_z; // @[Snxn100k.scala 19413:34]
  wire  inst_SnxnLv4Inst27_io_a; // @[Snxn100k.scala 19417:34]
  wire  inst_SnxnLv4Inst27_io_b; // @[Snxn100k.scala 19417:34]
  wire  inst_SnxnLv4Inst27_io_z; // @[Snxn100k.scala 19417:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst24_io_z + inst_SnxnLv4Inst25_io_z; // @[Snxn100k.scala 19421:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst26_io_z; // @[Snxn100k.scala 19421:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst27_io_z; // @[Snxn100k.scala 19421:89]
  SnxnLv4Inst24 inst_SnxnLv4Inst24 ( // @[Snxn100k.scala 19405:34]
    .io_a(inst_SnxnLv4Inst24_io_a),
    .io_b(inst_SnxnLv4Inst24_io_b),
    .io_z(inst_SnxnLv4Inst24_io_z)
  );
  SnxnLv4Inst25 inst_SnxnLv4Inst25 ( // @[Snxn100k.scala 19409:34]
    .io_a(inst_SnxnLv4Inst25_io_a),
    .io_b(inst_SnxnLv4Inst25_io_b),
    .io_z(inst_SnxnLv4Inst25_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst26 ( // @[Snxn100k.scala 19413:34]
    .io_a(inst_SnxnLv4Inst26_io_a),
    .io_b(inst_SnxnLv4Inst26_io_b),
    .io_z(inst_SnxnLv4Inst26_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst27 ( // @[Snxn100k.scala 19417:34]
    .io_a(inst_SnxnLv4Inst27_io_a),
    .io_b(inst_SnxnLv4Inst27_io_b),
    .io_z(inst_SnxnLv4Inst27_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 19422:15]
  assign inst_SnxnLv4Inst24_io_a = io_a; // @[Snxn100k.scala 19406:27]
  assign inst_SnxnLv4Inst24_io_b = io_b; // @[Snxn100k.scala 19407:27]
  assign inst_SnxnLv4Inst25_io_a = io_a; // @[Snxn100k.scala 19410:27]
  assign inst_SnxnLv4Inst25_io_b = io_b; // @[Snxn100k.scala 19411:27]
  assign inst_SnxnLv4Inst26_io_a = io_a; // @[Snxn100k.scala 19414:27]
  assign inst_SnxnLv4Inst26_io_b = io_b; // @[Snxn100k.scala 19415:27]
  assign inst_SnxnLv4Inst27_io_a = io_a; // @[Snxn100k.scala 19418:27]
  assign inst_SnxnLv4Inst27_io_b = io_b; // @[Snxn100k.scala 19419:27]
endmodule
module SnxnLv4Inst28(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 70236:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 70237:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 70238:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 70239:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 70240:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 70241:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 70242:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 70243:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 70244:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 70245:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 70246:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 70247:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 70248:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 70249:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 70250:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 70251:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 70252:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 70253:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 70254:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 70255:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 70256:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 70257:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 70258:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 70259:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 70260:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 70261:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 70262:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 70263:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 70264:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 70265:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 70266:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 70267:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 70268:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 70269:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 70270:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 70271:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 70272:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 70273:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 70274:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 70275:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 70276:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 70277:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 70278:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 70279:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 70280:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 70281:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 70282:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 70283:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 70284:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 70285:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 70286:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 70287:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 70288:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 70289:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 70290:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 70291:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 70292:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 70293:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 70294:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 70295:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 70296:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 70297:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 70298:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 70299:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 70300:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 70301:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 70302:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 70303:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 70304:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 70305:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 70306:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 70307:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 70308:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 70309:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 70310:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 70311:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 70312:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 70313:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 70314:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 70315:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 70316:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 70317:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 70318:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 70319:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 70320:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 70321:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 70322:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 70323:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 70324:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 70325:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 70326:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 70327:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 70328:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 70329:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 70330:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 70331:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 70332:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 70333:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 70334:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 70335:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 70336:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 70337:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 70338:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 70339:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 70340:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 70341:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 70342:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 70343:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 70344:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 70345:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 70346:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 70347:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 70348:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 70349:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 70350:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 70351:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 70352:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 70353:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 70354:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 70355:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 70356:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 70357:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 70358:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 70359:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 70360:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 70361:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 70362:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 70363:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 70364:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 70365:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 70366:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 70367:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 70368:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 70369:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 70370:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 70371:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 70372:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 70373:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 70374:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 70375:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 70376:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 70377:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 70378:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 70379:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 70380:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 70381:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 70382:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 70383:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 70384:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 70385:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 70386:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 70387:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 70388:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 70389:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 70390:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 70391:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 70392:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 70393:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 70394:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 70395:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 70396:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 70397:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 70398:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 70399:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 70400:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 70401:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 70402:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 70403:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 70404:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 70405:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 70406:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 70407:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 70408:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 70409:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 70410:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 70411:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 70412:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 70413:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 70414:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 70415:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 70416:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 70417:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 70418:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 70419:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 70420:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 70421:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 70422:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 70423:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 70424:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 70425:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 70426:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 70427:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 70428:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 70429:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 70430:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 70431:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 70432:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 70433:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 70434:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 70435:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 70436:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 70437:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 70438:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 70439:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 70440:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 70441:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 70442:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 70443:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 70444:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 70445:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 70446:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 70447:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 70448:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 70449:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 70450:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 70451:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 70452:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 70453:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 70454:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 70455:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 70456:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 70457:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 70458:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 70459:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 70460:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 70461:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 70462:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 70463:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 70464:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 70465:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 70466:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 70467:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 70468:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 70469:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 70470:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 70471:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 70472:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 70473:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 70474:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 70475:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 70476:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 70477:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 70478:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 70479:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 70480:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 70481:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 70482:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 70483:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 70484:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 70485:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 70486:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 70487:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 70488:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 70489:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 70490:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 70491:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 70492:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 70493:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 70494:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 70495:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 70496:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 70497:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 70498:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 70499:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 70500:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 70501:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 70502:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 70503:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 70504:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 70505:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 70506:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 70507:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 70508:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 70509:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 70510:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 70511:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 70512:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 70513:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 70514:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 70515:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 70516:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 70517:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 70518:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 70519:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 70520:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 70521:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 70522:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 70523:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 70524:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 70525:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 70526:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 70527:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 70528:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 70529:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 70530:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 70531:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 70532:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 70533:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 70534:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 70535:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 70536:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 70537:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 70538:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 70539:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 70540:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 70541:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 70542:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 70543:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 70544:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 70545:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 70546:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 70547:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 70548:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 70549:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 70550:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 70551:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 70552:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 70553:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 70554:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 70555:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 70556:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 70557:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 70558:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 70559:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 70560:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 70561:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 70562:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 70563:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 70564:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 70565:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 70566:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 70567:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 70568:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 70569:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 70570:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 70571:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 70572:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 70573:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 70574:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 70575:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 70576:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 70577:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 70578:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 70579:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 70580:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 70581:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 70582:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 70583:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 70584:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 70585:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 70586:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 70587:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 70588:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 70589:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 70590:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 70591:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 70592:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 70593:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 70594:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 70595:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 70596:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 70597:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 70598:20]
  assign io_z = ~x90; // @[Snxn100k.scala 70599:16]
endmodule
module SnxnLv4Inst29(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 70610:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 70611:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 70612:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 70613:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 70614:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 70615:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 70616:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 70617:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 70618:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 70619:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 70620:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 70621:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 70622:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 70623:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 70624:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 70625:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 70626:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 70627:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 70628:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 70629:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 70630:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 70631:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 70632:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 70633:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 70634:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 70635:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 70636:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 70637:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 70638:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 70639:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 70640:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 70641:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 70642:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 70643:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 70644:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 70645:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 70646:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 70647:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 70648:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 70649:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 70650:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 70651:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 70652:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 70653:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 70654:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 70655:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 70656:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 70657:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 70658:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 70659:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 70660:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 70661:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 70662:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 70663:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 70664:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 70665:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 70666:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 70667:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 70668:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 70669:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 70670:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 70671:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 70672:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 70673:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 70674:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 70675:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 70676:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 70677:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 70678:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 70679:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 70680:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 70681:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 70682:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 70683:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 70684:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 70685:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 70686:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 70687:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 70688:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 70689:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 70690:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 70691:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 70692:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 70693:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 70694:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 70695:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 70696:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 70697:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 70698:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 70699:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 70700:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 70701:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 70702:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 70703:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 70704:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 70705:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 70706:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 70707:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 70708:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 70709:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 70710:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 70711:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 70712:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 70713:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 70714:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 70715:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 70716:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 70717:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 70718:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 70719:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 70720:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 70721:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 70722:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 70723:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 70724:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 70725:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 70726:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 70727:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 70728:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 70729:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 70730:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 70731:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 70732:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 70733:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 70734:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 70735:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 70736:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 70737:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 70738:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 70739:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 70740:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 70741:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 70742:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 70743:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 70744:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 70745:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 70746:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 70747:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 70748:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 70749:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 70750:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 70751:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 70752:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 70753:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 70754:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 70755:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 70756:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 70757:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 70758:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 70759:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 70760:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 70761:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 70762:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 70763:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 70764:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 70765:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 70766:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 70767:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 70768:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 70769:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 70770:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 70771:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 70772:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 70773:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 70774:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 70775:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 70776:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 70777:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 70778:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 70779:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 70780:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 70781:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 70782:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 70783:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 70784:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 70785:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 70786:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 70787:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 70788:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 70789:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 70790:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 70791:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 70792:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 70793:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 70794:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 70795:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 70796:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 70797:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 70798:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 70799:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 70800:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 70801:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 70802:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 70803:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 70804:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 70805:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 70806:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 70807:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 70808:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 70809:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 70810:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 70811:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 70812:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 70813:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 70814:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 70815:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 70816:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 70817:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 70818:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 70819:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 70820:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 70821:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 70822:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 70823:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 70824:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 70825:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 70826:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 70827:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 70828:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 70829:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 70830:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 70831:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 70832:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 70833:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 70834:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 70835:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 70836:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 70837:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 70838:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 70839:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 70840:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 70841:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 70842:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 70843:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 70844:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 70845:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 70846:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 70847:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 70848:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 70849:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 70850:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 70851:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 70852:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 70853:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 70854:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 70855:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 70856:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 70857:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 70858:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 70859:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 70860:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 70861:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 70862:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 70863:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 70864:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 70865:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 70866:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 70867:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 70868:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 70869:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 70870:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 70871:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 70872:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 70873:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 70874:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 70875:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 70876:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 70877:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 70878:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 70879:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 70880:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 70881:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 70882:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 70883:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 70884:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 70885:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 70886:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 70887:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 70888:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 70889:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 70890:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 70891:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 70892:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 70893:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 70894:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 70895:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 70896:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 70897:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 70898:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 70899:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 70900:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 70901:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 70902:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 70903:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 70904:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 70905:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 70906:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 70907:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 70908:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 70909:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 70910:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 70911:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 70912:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 70913:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 70914:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 70915:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 70916:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 70917:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 70918:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 70919:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 70920:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 70921:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 70922:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 70923:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 70924:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 70925:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 70926:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 70927:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 70928:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 70929:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 70930:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 70931:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 70932:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 70933:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 70934:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 70935:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 70936:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 70937:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 70938:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 70939:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 70940:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 70941:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 70942:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 70943:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 70944:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 70945:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 70946:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 70947:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 70948:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 70949:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 70950:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 70951:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 70952:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 70953:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 70954:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 70955:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 70956:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 70957:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 70958:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 70959:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 70960:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 70961:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 70962:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 70963:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 70964:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 70965:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 70966:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 70967:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 70968:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 70969:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 70970:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 70971:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 70972:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 70973:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 70974:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 70975:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 70976:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 70977:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 70978:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 70979:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 70980:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 70981:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 70982:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 70983:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 70984:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 70985:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 70986:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 70987:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 70988:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 70989:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 70990:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 70991:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 70992:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 70993:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 70994:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 70995:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 70996:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 70997:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 70998:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 70999:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 71000:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 71001:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 71002:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 71003:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 71004:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 71005:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 71006:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 71007:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 71008:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 71009:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 71010:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 71011:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 71012:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 71013:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 71014:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 71015:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 71016:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 71017:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 71018:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 71019:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 71020:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 71021:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 71022:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 71023:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 71024:22]
  assign io_z = ~x103; // @[Snxn100k.scala 71025:17]
endmodule
module SnxnLv3Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst28_io_a; // @[Snxn100k.scala 18527:34]
  wire  inst_SnxnLv4Inst28_io_b; // @[Snxn100k.scala 18527:34]
  wire  inst_SnxnLv4Inst28_io_z; // @[Snxn100k.scala 18527:34]
  wire  inst_SnxnLv4Inst29_io_a; // @[Snxn100k.scala 18531:34]
  wire  inst_SnxnLv4Inst29_io_b; // @[Snxn100k.scala 18531:34]
  wire  inst_SnxnLv4Inst29_io_z; // @[Snxn100k.scala 18531:34]
  wire  inst_SnxnLv4Inst30_io_a; // @[Snxn100k.scala 18535:34]
  wire  inst_SnxnLv4Inst30_io_b; // @[Snxn100k.scala 18535:34]
  wire  inst_SnxnLv4Inst30_io_z; // @[Snxn100k.scala 18535:34]
  wire  inst_SnxnLv4Inst31_io_a; // @[Snxn100k.scala 18539:34]
  wire  inst_SnxnLv4Inst31_io_b; // @[Snxn100k.scala 18539:34]
  wire  inst_SnxnLv4Inst31_io_z; // @[Snxn100k.scala 18539:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst28_io_z + inst_SnxnLv4Inst29_io_z; // @[Snxn100k.scala 18543:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst30_io_z; // @[Snxn100k.scala 18543:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst31_io_z; // @[Snxn100k.scala 18543:89]
  SnxnLv4Inst28 inst_SnxnLv4Inst28 ( // @[Snxn100k.scala 18527:34]
    .io_a(inst_SnxnLv4Inst28_io_a),
    .io_b(inst_SnxnLv4Inst28_io_b),
    .io_z(inst_SnxnLv4Inst28_io_z)
  );
  SnxnLv4Inst29 inst_SnxnLv4Inst29 ( // @[Snxn100k.scala 18531:34]
    .io_a(inst_SnxnLv4Inst29_io_a),
    .io_b(inst_SnxnLv4Inst29_io_b),
    .io_z(inst_SnxnLv4Inst29_io_z)
  );
  SnxnLv4Inst4 inst_SnxnLv4Inst30 ( // @[Snxn100k.scala 18535:34]
    .io_a(inst_SnxnLv4Inst30_io_a),
    .io_b(inst_SnxnLv4Inst30_io_b),
    .io_z(inst_SnxnLv4Inst30_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst31 ( // @[Snxn100k.scala 18539:34]
    .io_a(inst_SnxnLv4Inst31_io_a),
    .io_b(inst_SnxnLv4Inst31_io_b),
    .io_z(inst_SnxnLv4Inst31_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 18544:15]
  assign inst_SnxnLv4Inst28_io_a = io_a; // @[Snxn100k.scala 18528:27]
  assign inst_SnxnLv4Inst28_io_b = io_b; // @[Snxn100k.scala 18529:27]
  assign inst_SnxnLv4Inst29_io_a = io_a; // @[Snxn100k.scala 18532:27]
  assign inst_SnxnLv4Inst29_io_b = io_b; // @[Snxn100k.scala 18533:27]
  assign inst_SnxnLv4Inst30_io_a = io_a; // @[Snxn100k.scala 18536:27]
  assign inst_SnxnLv4Inst30_io_b = io_b; // @[Snxn100k.scala 18537:27]
  assign inst_SnxnLv4Inst31_io_a = io_a; // @[Snxn100k.scala 18540:27]
  assign inst_SnxnLv4Inst31_io_b = io_b; // @[Snxn100k.scala 18541:27]
endmodule
module SnxnLv2Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst4_io_a; // @[Snxn100k.scala 4164:33]
  wire  inst_SnxnLv3Inst4_io_b; // @[Snxn100k.scala 4164:33]
  wire  inst_SnxnLv3Inst4_io_z; // @[Snxn100k.scala 4164:33]
  wire  inst_SnxnLv3Inst5_io_a; // @[Snxn100k.scala 4168:33]
  wire  inst_SnxnLv3Inst5_io_b; // @[Snxn100k.scala 4168:33]
  wire  inst_SnxnLv3Inst5_io_z; // @[Snxn100k.scala 4168:33]
  wire  inst_SnxnLv3Inst6_io_a; // @[Snxn100k.scala 4172:33]
  wire  inst_SnxnLv3Inst6_io_b; // @[Snxn100k.scala 4172:33]
  wire  inst_SnxnLv3Inst6_io_z; // @[Snxn100k.scala 4172:33]
  wire  inst_SnxnLv3Inst7_io_a; // @[Snxn100k.scala 4176:33]
  wire  inst_SnxnLv3Inst7_io_b; // @[Snxn100k.scala 4176:33]
  wire  inst_SnxnLv3Inst7_io_z; // @[Snxn100k.scala 4176:33]
  wire  _sum_T_1 = inst_SnxnLv3Inst4_io_z + inst_SnxnLv3Inst5_io_z; // @[Snxn100k.scala 4180:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst6_io_z; // @[Snxn100k.scala 4180:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst7_io_z; // @[Snxn100k.scala 4180:86]
  SnxnLv3Inst4 inst_SnxnLv3Inst4 ( // @[Snxn100k.scala 4164:33]
    .io_a(inst_SnxnLv3Inst4_io_a),
    .io_b(inst_SnxnLv3Inst4_io_b),
    .io_z(inst_SnxnLv3Inst4_io_z)
  );
  SnxnLv3Inst5 inst_SnxnLv3Inst5 ( // @[Snxn100k.scala 4168:33]
    .io_a(inst_SnxnLv3Inst5_io_a),
    .io_b(inst_SnxnLv3Inst5_io_b),
    .io_z(inst_SnxnLv3Inst5_io_z)
  );
  SnxnLv3Inst6 inst_SnxnLv3Inst6 ( // @[Snxn100k.scala 4172:33]
    .io_a(inst_SnxnLv3Inst6_io_a),
    .io_b(inst_SnxnLv3Inst6_io_b),
    .io_z(inst_SnxnLv3Inst6_io_z)
  );
  SnxnLv3Inst7 inst_SnxnLv3Inst7 ( // @[Snxn100k.scala 4176:33]
    .io_a(inst_SnxnLv3Inst7_io_a),
    .io_b(inst_SnxnLv3Inst7_io_b),
    .io_z(inst_SnxnLv3Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 4181:15]
  assign inst_SnxnLv3Inst4_io_a = io_a; // @[Snxn100k.scala 4165:26]
  assign inst_SnxnLv3Inst4_io_b = io_b; // @[Snxn100k.scala 4166:26]
  assign inst_SnxnLv3Inst5_io_a = io_a; // @[Snxn100k.scala 4169:26]
  assign inst_SnxnLv3Inst5_io_b = io_b; // @[Snxn100k.scala 4170:26]
  assign inst_SnxnLv3Inst6_io_a = io_a; // @[Snxn100k.scala 4173:26]
  assign inst_SnxnLv3Inst6_io_b = io_b; // @[Snxn100k.scala 4174:26]
  assign inst_SnxnLv3Inst7_io_a = io_a; // @[Snxn100k.scala 4177:26]
  assign inst_SnxnLv3Inst7_io_b = io_b; // @[Snxn100k.scala 4178:26]
endmodule
module SnxnLv4Inst33(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 88298:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 88299:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 88300:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 88301:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 88302:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 88303:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 88304:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 88305:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 88306:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 88307:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 88308:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 88309:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 88310:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 88311:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 88312:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 88313:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 88314:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 88315:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 88316:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 88317:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 88318:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 88319:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 88320:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 88321:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 88322:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 88323:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 88324:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 88325:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 88326:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 88327:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 88328:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 88329:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 88330:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 88331:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 88332:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 88333:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 88334:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 88335:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 88336:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 88337:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 88338:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 88339:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 88340:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 88341:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 88342:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 88343:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 88344:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 88345:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 88346:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 88347:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 88348:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 88349:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 88350:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 88351:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 88352:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 88353:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 88354:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 88355:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 88356:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 88357:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 88358:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 88359:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 88360:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 88361:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 88362:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 88363:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 88364:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 88365:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 88366:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 88367:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 88368:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 88369:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 88370:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 88371:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 88372:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 88373:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 88374:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 88375:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 88376:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 88377:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 88378:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 88379:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 88380:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 88381:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 88382:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 88383:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 88384:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 88385:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 88386:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 88387:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 88388:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 88389:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 88390:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 88391:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 88392:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 88393:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 88394:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 88395:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 88396:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 88397:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 88398:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 88399:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 88400:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 88401:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 88402:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 88403:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 88404:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 88405:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 88406:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 88407:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 88408:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 88409:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 88410:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 88411:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 88412:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 88413:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 88414:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 88415:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 88416:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 88417:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 88418:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 88419:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 88420:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 88421:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 88422:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 88423:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 88424:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 88425:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 88426:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 88427:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 88428:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 88429:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 88430:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 88431:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 88432:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 88433:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 88434:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 88435:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 88436:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 88437:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 88438:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 88439:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 88440:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 88441:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 88442:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 88443:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 88444:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 88445:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 88446:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 88447:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 88448:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 88449:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 88450:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 88451:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 88452:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 88453:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 88454:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 88455:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 88456:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 88457:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 88458:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 88459:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 88460:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 88461:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 88462:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 88463:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 88464:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 88465:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 88466:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 88467:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 88468:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 88469:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 88470:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 88471:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 88472:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 88473:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 88474:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 88475:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 88476:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 88477:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 88478:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 88479:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 88480:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 88481:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 88482:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 88483:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 88484:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 88485:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 88486:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 88487:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 88488:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 88489:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 88490:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 88491:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 88492:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 88493:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 88494:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 88495:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 88496:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 88497:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 88498:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 88499:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 88500:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 88501:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 88502:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 88503:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 88504:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 88505:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 88506:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 88507:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 88508:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 88509:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 88510:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 88511:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 88512:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 88513:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 88514:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 88515:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 88516:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 88517:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 88518:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 88519:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 88520:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 88521:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 88522:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 88523:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 88524:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 88525:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 88526:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 88527:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 88528:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 88529:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 88530:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 88531:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 88532:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 88533:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 88534:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 88535:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 88536:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 88537:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 88538:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 88539:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 88540:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 88541:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 88542:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 88543:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 88544:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 88545:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 88546:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 88547:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 88548:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 88549:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 88550:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 88551:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 88552:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 88553:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 88554:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 88555:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 88556:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 88557:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 88558:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 88559:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 88560:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 88561:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 88562:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 88563:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 88564:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 88565:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 88566:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 88567:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 88568:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 88569:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 88570:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 88571:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 88572:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 88573:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 88574:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 88575:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 88576:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 88577:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 88578:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 88579:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 88580:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 88581:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 88582:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 88583:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 88584:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 88585:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 88586:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 88587:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 88588:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 88589:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 88590:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 88591:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 88592:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 88593:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 88594:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 88595:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 88596:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 88597:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 88598:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 88599:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 88600:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 88601:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 88602:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 88603:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 88604:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 88605:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 88606:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 88607:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 88608:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 88609:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 88610:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 88611:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 88612:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 88613:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 88614:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 88615:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 88616:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 88617:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 88618:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 88619:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 88620:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 88621:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 88622:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 88623:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 88624:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 88625:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 88626:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 88627:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 88628:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 88629:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 88630:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 88631:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 88632:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 88633:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 88634:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 88635:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 88636:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 88637:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 88638:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 88639:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 88640:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 88641:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 88642:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 88643:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 88644:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 88645:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 88646:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 88647:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 88648:20]
  assign io_z = ~x87; // @[Snxn100k.scala 88649:16]
endmodule
module SnxnLv4Inst34(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 89110:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 89111:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 89112:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 89113:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 89114:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 89115:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 89116:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 89117:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 89118:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 89119:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 89120:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 89121:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 89122:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 89123:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 89124:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 89125:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 89126:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 89127:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 89128:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 89129:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 89130:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 89131:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 89132:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 89133:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 89134:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 89135:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 89136:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 89137:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 89138:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 89139:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 89140:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 89141:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 89142:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 89143:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 89144:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 89145:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 89146:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 89147:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 89148:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 89149:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 89150:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 89151:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 89152:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 89153:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 89154:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 89155:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 89156:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 89157:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 89158:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 89159:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 89160:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 89161:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 89162:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 89163:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 89164:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 89165:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 89166:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 89167:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 89168:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 89169:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 89170:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 89171:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 89172:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 89173:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 89174:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 89175:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 89176:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 89177:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 89178:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 89179:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 89180:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 89181:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 89182:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 89183:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 89184:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 89185:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 89186:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 89187:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 89188:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 89189:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 89190:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 89191:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 89192:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 89193:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 89194:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 89195:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 89196:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 89197:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 89198:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 89199:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 89200:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 89201:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 89202:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 89203:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 89204:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 89205:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 89206:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 89207:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 89208:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 89209:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 89210:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 89211:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 89212:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 89213:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 89214:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 89215:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 89216:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 89217:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 89218:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 89219:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 89220:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 89221:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 89222:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 89223:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 89224:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 89225:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 89226:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 89227:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 89228:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 89229:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 89230:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 89231:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 89232:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 89233:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 89234:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 89235:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 89236:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 89237:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 89238:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 89239:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 89240:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 89241:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 89242:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 89243:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 89244:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 89245:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 89246:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 89247:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 89248:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 89249:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 89250:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 89251:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 89252:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 89253:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 89254:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 89255:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 89256:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 89257:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 89258:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 89259:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 89260:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 89261:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 89262:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 89263:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 89264:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 89265:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 89266:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 89267:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 89268:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 89269:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 89270:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 89271:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 89272:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 89273:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 89274:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 89275:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 89276:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 89277:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 89278:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 89279:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 89280:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 89281:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 89282:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 89283:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 89284:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 89285:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 89286:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 89287:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 89288:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 89289:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 89290:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 89291:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 89292:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 89293:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 89294:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 89295:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 89296:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 89297:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 89298:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 89299:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 89300:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 89301:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 89302:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 89303:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 89304:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 89305:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 89306:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 89307:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 89308:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 89309:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 89310:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 89311:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 89312:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 89313:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 89314:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 89315:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 89316:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 89317:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 89318:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 89319:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 89320:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 89321:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 89322:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 89323:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 89324:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 89325:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 89326:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 89327:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 89328:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 89329:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 89330:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 89331:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 89332:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 89333:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 89334:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 89335:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 89336:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 89337:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 89338:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 89339:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 89340:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 89341:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 89342:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 89343:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 89344:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 89345:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 89346:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 89347:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 89348:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 89349:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 89350:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 89351:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 89352:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 89353:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 89354:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 89355:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 89356:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 89357:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 89358:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 89359:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 89360:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 89361:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 89362:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 89363:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 89364:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 89365:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 89366:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 89367:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 89368:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 89369:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 89370:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 89371:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 89372:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 89373:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 89374:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 89375:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 89376:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 89377:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 89378:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 89379:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 89380:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 89381:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 89382:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 89383:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 89384:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 89385:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 89386:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 89387:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 89388:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 89389:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 89390:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 89391:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 89392:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 89393:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 89394:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 89395:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 89396:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 89397:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 89398:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 89399:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 89400:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 89401:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 89402:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 89403:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 89404:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 89405:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 89406:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 89407:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 89408:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 89409:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 89410:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 89411:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 89412:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 89413:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 89414:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 89415:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 89416:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 89417:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 89418:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 89419:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 89420:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 89421:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 89422:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 89423:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 89424:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 89425:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 89426:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 89427:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 89428:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 89429:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 89430:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 89431:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 89432:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 89433:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 89434:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 89435:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 89436:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 89437:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 89438:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 89439:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 89440:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 89441:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 89442:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 89443:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 89444:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 89445:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 89446:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 89447:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 89448:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 89449:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 89450:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 89451:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 89452:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 89453:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 89454:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 89455:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 89456:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 89457:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 89458:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 89459:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 89460:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 89461:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 89462:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 89463:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 89464:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 89465:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 89466:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 89467:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 89468:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 89469:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 89470:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 89471:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 89472:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 89473:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 89474:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 89475:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 89476:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 89477:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 89478:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 89479:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 89480:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 89481:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 89482:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 89483:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 89484:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 89485:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 89486:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 89487:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 89488:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 89489:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 89490:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 89491:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 89492:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 89493:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 89494:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 89495:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 89496:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 89497:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 89498:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 89499:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 89500:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 89501:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 89502:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 89503:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 89504:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 89505:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 89506:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 89507:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 89508:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 89509:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 89510:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 89511:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 89512:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 89513:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 89514:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 89515:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 89516:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 89517:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 89518:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 89519:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 89520:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 89521:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 89522:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 89523:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 89524:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 89525:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 89526:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 89527:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 89528:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 89529:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 89530:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 89531:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 89532:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 89533:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 89534:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 89535:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 89536:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 89537:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 89538:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 89539:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 89540:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 89541:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 89542:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 89543:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 89544:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 89545:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 89546:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 89547:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 89548:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 89549:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 89550:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 89551:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 89552:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 89553:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 89554:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 89555:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 89556:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 89557:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 89558:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 89559:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 89560:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 89561:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 89562:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 89563:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 89564:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 89565:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 89566:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 89567:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 89568:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 89569:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 89570:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 89571:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 89572:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 89573:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 89574:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 89575:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 89576:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 89577:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 89578:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 89579:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 89580:22]
  assign io_z = ~x117; // @[Snxn100k.scala 89581:17]
endmodule
module SnxnLv4Inst35(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 88660:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 88661:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 88662:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 88663:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 88664:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 88665:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 88666:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 88667:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 88668:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 88669:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 88670:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 88671:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 88672:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 88673:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 88674:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 88675:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 88676:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 88677:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 88678:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 88679:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 88680:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 88681:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 88682:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 88683:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 88684:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 88685:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 88686:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 88687:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 88688:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 88689:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 88690:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 88691:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 88692:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 88693:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 88694:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 88695:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 88696:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 88697:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 88698:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 88699:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 88700:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 88701:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 88702:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 88703:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 88704:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 88705:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 88706:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 88707:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 88708:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 88709:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 88710:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 88711:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 88712:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 88713:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 88714:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 88715:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 88716:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 88717:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 88718:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 88719:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 88720:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 88721:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 88722:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 88723:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 88724:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 88725:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 88726:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 88727:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 88728:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 88729:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 88730:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 88731:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 88732:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 88733:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 88734:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 88735:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 88736:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 88737:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 88738:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 88739:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 88740:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 88741:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 88742:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 88743:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 88744:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 88745:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 88746:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 88747:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 88748:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 88749:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 88750:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 88751:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 88752:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 88753:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 88754:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 88755:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 88756:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 88757:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 88758:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 88759:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 88760:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 88761:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 88762:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 88763:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 88764:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 88765:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 88766:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 88767:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 88768:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 88769:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 88770:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 88771:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 88772:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 88773:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 88774:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 88775:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 88776:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 88777:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 88778:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 88779:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 88780:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 88781:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 88782:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 88783:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 88784:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 88785:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 88786:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 88787:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 88788:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 88789:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 88790:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 88791:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 88792:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 88793:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 88794:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 88795:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 88796:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 88797:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 88798:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 88799:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 88800:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 88801:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 88802:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 88803:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 88804:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 88805:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 88806:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 88807:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 88808:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 88809:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 88810:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 88811:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 88812:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 88813:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 88814:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 88815:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 88816:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 88817:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 88818:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 88819:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 88820:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 88821:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 88822:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 88823:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 88824:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 88825:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 88826:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 88827:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 88828:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 88829:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 88830:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 88831:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 88832:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 88833:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 88834:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 88835:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 88836:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 88837:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 88838:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 88839:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 88840:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 88841:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 88842:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 88843:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 88844:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 88845:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 88846:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 88847:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 88848:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 88849:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 88850:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 88851:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 88852:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 88853:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 88854:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 88855:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 88856:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 88857:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 88858:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 88859:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 88860:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 88861:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 88862:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 88863:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 88864:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 88865:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 88866:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 88867:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 88868:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 88869:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 88870:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 88871:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 88872:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 88873:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 88874:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 88875:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 88876:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 88877:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 88878:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 88879:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 88880:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 88881:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 88882:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 88883:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 88884:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 88885:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 88886:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 88887:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 88888:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 88889:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 88890:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 88891:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 88892:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 88893:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 88894:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 88895:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 88896:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 88897:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 88898:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 88899:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 88900:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 88901:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 88902:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 88903:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 88904:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 88905:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 88906:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 88907:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 88908:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 88909:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 88910:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 88911:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 88912:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 88913:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 88914:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 88915:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 88916:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 88917:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 88918:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 88919:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 88920:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 88921:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 88922:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 88923:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 88924:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 88925:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 88926:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 88927:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 88928:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 88929:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 88930:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 88931:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 88932:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 88933:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 88934:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 88935:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 88936:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 88937:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 88938:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 88939:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 88940:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 88941:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 88942:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 88943:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 88944:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 88945:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 88946:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 88947:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 88948:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 88949:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 88950:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 88951:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 88952:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 88953:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 88954:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 88955:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 88956:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 88957:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 88958:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 88959:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 88960:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 88961:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 88962:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 88963:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 88964:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 88965:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 88966:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 88967:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 88968:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 88969:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 88970:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 88971:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 88972:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 88973:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 88974:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 88975:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 88976:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 88977:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 88978:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 88979:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 88980:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 88981:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 88982:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 88983:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 88984:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 88985:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 88986:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 88987:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 88988:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 88989:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 88990:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 88991:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 88992:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 88993:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 88994:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 88995:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 88996:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 88997:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 88998:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 88999:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 89000:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 89001:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 89002:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 89003:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 89004:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 89005:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 89006:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 89007:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 89008:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 89009:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 89010:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 89011:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 89012:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 89013:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 89014:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 89015:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 89016:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 89017:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 89018:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 89019:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 89020:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 89021:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 89022:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 89023:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 89024:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 89025:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 89026:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 89027:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 89028:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 89029:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 89030:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 89031:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 89032:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 89033:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 89034:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 89035:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 89036:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 89037:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 89038:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 89039:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 89040:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 89041:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 89042:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 89043:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 89044:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 89045:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 89046:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 89047:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 89048:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 89049:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 89050:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 89051:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 89052:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 89053:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 89054:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 89055:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 89056:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 89057:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 89058:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 89059:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 89060:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 89061:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 89062:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 89063:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 89064:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 89065:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 89066:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 89067:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 89068:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 89069:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 89070:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 89071:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 89072:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 89073:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 89074:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 89075:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 89076:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 89077:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 89078:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 89079:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 89080:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 89081:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 89082:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 89083:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 89084:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 89085:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 89086:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 89087:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 89088:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 89089:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 89090:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 89091:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 89092:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 89093:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 89094:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 89095:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 89096:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 89097:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 89098:22]
  assign io_z = ~x109; // @[Snxn100k.scala 89099:17]
endmodule
module SnxnLv3Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst32_io_a; // @[Snxn100k.scala 22809:34]
  wire  inst_SnxnLv4Inst32_io_b; // @[Snxn100k.scala 22809:34]
  wire  inst_SnxnLv4Inst32_io_z; // @[Snxn100k.scala 22809:34]
  wire  inst_SnxnLv4Inst33_io_a; // @[Snxn100k.scala 22813:34]
  wire  inst_SnxnLv4Inst33_io_b; // @[Snxn100k.scala 22813:34]
  wire  inst_SnxnLv4Inst33_io_z; // @[Snxn100k.scala 22813:34]
  wire  inst_SnxnLv4Inst34_io_a; // @[Snxn100k.scala 22817:34]
  wire  inst_SnxnLv4Inst34_io_b; // @[Snxn100k.scala 22817:34]
  wire  inst_SnxnLv4Inst34_io_z; // @[Snxn100k.scala 22817:34]
  wire  inst_SnxnLv4Inst35_io_a; // @[Snxn100k.scala 22821:34]
  wire  inst_SnxnLv4Inst35_io_b; // @[Snxn100k.scala 22821:34]
  wire  inst_SnxnLv4Inst35_io_z; // @[Snxn100k.scala 22821:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst32_io_z + inst_SnxnLv4Inst33_io_z; // @[Snxn100k.scala 22825:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst34_io_z; // @[Snxn100k.scala 22825:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst35_io_z; // @[Snxn100k.scala 22825:89]
  SnxnLv4Inst7 inst_SnxnLv4Inst32 ( // @[Snxn100k.scala 22809:34]
    .io_a(inst_SnxnLv4Inst32_io_a),
    .io_b(inst_SnxnLv4Inst32_io_b),
    .io_z(inst_SnxnLv4Inst32_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst33 ( // @[Snxn100k.scala 22813:34]
    .io_a(inst_SnxnLv4Inst33_io_a),
    .io_b(inst_SnxnLv4Inst33_io_b),
    .io_z(inst_SnxnLv4Inst33_io_z)
  );
  SnxnLv4Inst34 inst_SnxnLv4Inst34 ( // @[Snxn100k.scala 22817:34]
    .io_a(inst_SnxnLv4Inst34_io_a),
    .io_b(inst_SnxnLv4Inst34_io_b),
    .io_z(inst_SnxnLv4Inst34_io_z)
  );
  SnxnLv4Inst35 inst_SnxnLv4Inst35 ( // @[Snxn100k.scala 22821:34]
    .io_a(inst_SnxnLv4Inst35_io_a),
    .io_b(inst_SnxnLv4Inst35_io_b),
    .io_z(inst_SnxnLv4Inst35_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22826:15]
  assign inst_SnxnLv4Inst32_io_a = io_a; // @[Snxn100k.scala 22810:27]
  assign inst_SnxnLv4Inst32_io_b = io_b; // @[Snxn100k.scala 22811:27]
  assign inst_SnxnLv4Inst33_io_a = io_a; // @[Snxn100k.scala 22814:27]
  assign inst_SnxnLv4Inst33_io_b = io_b; // @[Snxn100k.scala 22815:27]
  assign inst_SnxnLv4Inst34_io_a = io_a; // @[Snxn100k.scala 22818:27]
  assign inst_SnxnLv4Inst34_io_b = io_b; // @[Snxn100k.scala 22819:27]
  assign inst_SnxnLv4Inst35_io_a = io_a; // @[Snxn100k.scala 22822:27]
  assign inst_SnxnLv4Inst35_io_b = io_b; // @[Snxn100k.scala 22823:27]
endmodule
module SnxnLv4Inst36(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 84424:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 84425:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 84426:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 84427:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 84428:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 84429:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 84430:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 84431:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 84432:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 84433:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 84434:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 84435:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 84436:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 84437:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 84438:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 84439:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 84440:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 84441:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 84442:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 84443:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 84444:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 84445:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 84446:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 84447:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 84448:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 84449:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 84450:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 84451:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 84452:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 84453:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 84454:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 84455:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 84456:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 84457:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 84458:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 84459:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 84460:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 84461:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 84462:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 84463:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 84464:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 84465:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 84466:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 84467:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 84468:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 84469:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 84470:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 84471:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 84472:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 84473:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 84474:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 84475:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 84476:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 84477:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 84478:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 84479:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 84480:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 84481:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 84482:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 84483:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 84484:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 84485:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 84486:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 84487:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 84488:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 84489:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 84490:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 84491:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 84492:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 84493:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 84494:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 84495:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 84496:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 84497:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 84498:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 84499:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 84500:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 84501:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 84502:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 84503:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 84504:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 84505:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 84506:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 84507:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 84508:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 84509:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 84510:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 84511:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 84512:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 84513:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 84514:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 84515:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 84516:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 84517:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 84518:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 84519:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 84520:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 84521:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 84522:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 84523:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 84524:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 84525:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 84526:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 84527:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 84528:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 84529:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 84530:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 84531:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 84532:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 84533:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 84534:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 84535:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 84536:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 84537:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 84538:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 84539:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 84540:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 84541:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 84542:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 84543:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 84544:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 84545:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 84546:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 84547:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 84548:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 84549:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 84550:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 84551:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 84552:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 84553:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 84554:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 84555:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 84556:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 84557:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 84558:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 84559:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 84560:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 84561:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 84562:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 84563:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 84564:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 84565:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 84566:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 84567:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 84568:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 84569:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 84570:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 84571:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 84572:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 84573:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 84574:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 84575:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 84576:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 84577:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 84578:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 84579:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 84580:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 84581:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 84582:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 84583:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 84584:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 84585:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 84586:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 84587:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 84588:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 84589:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 84590:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 84591:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 84592:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 84593:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 84594:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 84595:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 84596:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 84597:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 84598:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 84599:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 84600:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 84601:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 84602:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 84603:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 84604:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 84605:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 84606:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 84607:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 84608:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 84609:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 84610:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 84611:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 84612:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 84613:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 84614:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 84615:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 84616:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 84617:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 84618:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 84619:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 84620:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 84621:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 84622:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 84623:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 84624:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 84625:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 84626:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 84627:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 84628:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 84629:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 84630:20]
  assign io_z = ~x51; // @[Snxn100k.scala 84631:16]
endmodule
module SnxnLv4Inst38(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 85202:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 85203:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 85204:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 85205:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 85206:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 85207:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 85208:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 85209:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 85210:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 85211:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 85212:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 85213:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 85214:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 85215:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 85216:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 85217:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 85218:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 85219:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 85220:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 85221:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 85222:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 85223:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 85224:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 85225:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 85226:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 85227:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 85228:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 85229:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 85230:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 85231:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 85232:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 85233:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 85234:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 85235:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 85236:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 85237:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 85238:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 85239:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 85240:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 85241:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 85242:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 85243:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 85244:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 85245:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 85246:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 85247:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 85248:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 85249:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 85250:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 85251:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 85252:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 85253:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 85254:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 85255:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 85256:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 85257:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 85258:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 85259:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 85260:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 85261:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 85262:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 85263:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 85264:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 85265:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 85266:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 85267:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 85268:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 85269:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 85270:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 85271:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 85272:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 85273:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 85274:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 85275:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 85276:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 85277:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 85278:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 85279:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 85280:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 85281:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 85282:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 85283:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 85284:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 85285:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 85286:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 85287:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 85288:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 85289:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 85290:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 85291:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 85292:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 85293:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 85294:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 85295:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 85296:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 85297:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 85298:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 85299:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 85300:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 85301:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 85302:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 85303:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 85304:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 85305:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 85306:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 85307:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 85308:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 85309:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 85310:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 85311:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 85312:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 85313:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 85314:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 85315:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 85316:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 85317:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 85318:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 85319:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 85320:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 85321:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 85322:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 85323:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 85324:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 85325:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 85326:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 85327:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 85328:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 85329:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 85330:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 85331:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 85332:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 85333:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 85334:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 85335:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 85336:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 85337:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 85338:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 85339:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 85340:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 85341:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 85342:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 85343:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 85344:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 85345:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 85346:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 85347:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 85348:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 85349:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 85350:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 85351:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 85352:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 85353:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 85354:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 85355:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 85356:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 85357:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 85358:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 85359:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 85360:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 85361:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 85362:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 85363:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 85364:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 85365:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 85366:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 85367:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 85368:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 85369:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 85370:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 85371:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 85372:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 85373:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 85374:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 85375:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 85376:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 85377:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 85378:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 85379:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 85380:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 85381:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 85382:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 85383:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 85384:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 85385:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 85386:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 85387:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 85388:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 85389:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 85390:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 85391:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 85392:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 85393:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 85394:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 85395:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 85396:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 85397:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 85398:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 85399:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 85400:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 85401:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 85402:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 85403:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 85404:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 85405:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 85406:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 85407:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 85408:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 85409:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 85410:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 85411:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 85412:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 85413:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 85414:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 85415:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 85416:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 85417:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 85418:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 85419:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 85420:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 85421:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 85422:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 85423:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 85424:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 85425:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 85426:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 85427:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 85428:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 85429:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 85430:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 85431:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 85432:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 85433:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 85434:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 85435:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 85436:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 85437:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 85438:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 85439:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 85440:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 85441:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 85442:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 85443:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 85444:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 85445:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 85446:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 85447:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 85448:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 85449:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 85450:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 85451:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 85452:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 85453:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 85454:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 85455:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 85456:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 85457:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 85458:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 85459:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 85460:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 85461:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 85462:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 85463:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 85464:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 85465:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 85466:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 85467:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 85468:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 85469:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 85470:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 85471:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 85472:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 85473:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 85474:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 85475:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 85476:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 85477:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 85478:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 85479:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 85480:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 85481:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 85482:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 85483:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 85484:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 85485:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 85486:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 85487:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 85488:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 85489:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 85490:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 85491:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 85492:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 85493:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 85494:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 85495:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 85496:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 85497:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 85498:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 85499:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 85500:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 85501:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 85502:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 85503:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 85504:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 85505:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 85506:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 85507:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 85508:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 85509:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 85510:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 85511:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 85512:20]
  assign io_z = ~x77; // @[Snxn100k.scala 85513:16]
endmodule
module SnxnLv4Inst39(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 84642:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 84643:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 84644:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 84645:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 84646:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 84647:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 84648:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 84649:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 84650:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 84651:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 84652:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 84653:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 84654:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 84655:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 84656:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 84657:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 84658:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 84659:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 84660:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 84661:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 84662:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 84663:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 84664:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 84665:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 84666:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 84667:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 84668:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 84669:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 84670:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 84671:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 84672:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 84673:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 84674:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 84675:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 84676:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 84677:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 84678:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 84679:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 84680:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 84681:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 84682:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 84683:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 84684:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 84685:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 84686:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 84687:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 84688:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 84689:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 84690:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 84691:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 84692:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 84693:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 84694:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 84695:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 84696:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 84697:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 84698:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 84699:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 84700:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 84701:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 84702:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 84703:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 84704:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 84705:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 84706:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 84707:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 84708:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 84709:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 84710:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 84711:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 84712:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 84713:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 84714:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 84715:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 84716:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 84717:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 84718:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 84719:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 84720:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 84721:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 84722:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 84723:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 84724:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 84725:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 84726:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 84727:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 84728:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 84729:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 84730:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 84731:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 84732:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 84733:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 84734:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 84735:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 84736:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 84737:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 84738:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 84739:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 84740:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 84741:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 84742:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 84743:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 84744:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 84745:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 84746:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 84747:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 84748:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 84749:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 84750:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 84751:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 84752:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 84753:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 84754:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 84755:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 84756:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 84757:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 84758:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 84759:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 84760:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 84761:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 84762:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 84763:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 84764:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 84765:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 84766:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 84767:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 84768:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 84769:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 84770:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 84771:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 84772:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 84773:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 84774:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 84775:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 84776:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 84777:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 84778:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 84779:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 84780:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 84781:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 84782:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 84783:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 84784:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 84785:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 84786:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 84787:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 84788:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 84789:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 84790:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 84791:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 84792:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 84793:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 84794:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 84795:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 84796:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 84797:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 84798:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 84799:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 84800:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 84801:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 84802:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 84803:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 84804:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 84805:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 84806:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 84807:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 84808:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 84809:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 84810:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 84811:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 84812:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 84813:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 84814:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 84815:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 84816:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 84817:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 84818:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 84819:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 84820:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 84821:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 84822:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 84823:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 84824:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 84825:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 84826:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 84827:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 84828:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 84829:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 84830:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 84831:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 84832:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 84833:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 84834:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 84835:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 84836:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 84837:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 84838:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 84839:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 84840:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 84841:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 84842:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 84843:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 84844:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 84845:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 84846:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 84847:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 84848:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 84849:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 84850:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 84851:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 84852:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 84853:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 84854:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 84855:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 84856:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 84857:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 84858:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 84859:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 84860:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 84861:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 84862:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 84863:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 84864:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 84865:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 84866:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 84867:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 84868:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 84869:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 84870:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 84871:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 84872:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 84873:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 84874:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 84875:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 84876:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 84877:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 84878:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 84879:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 84880:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 84881:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 84882:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 84883:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 84884:20]
  assign io_z = ~x60; // @[Snxn100k.scala 84885:16]
endmodule
module SnxnLv3Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst36_io_a; // @[Snxn100k.scala 21988:34]
  wire  inst_SnxnLv4Inst36_io_b; // @[Snxn100k.scala 21988:34]
  wire  inst_SnxnLv4Inst36_io_z; // @[Snxn100k.scala 21988:34]
  wire  inst_SnxnLv4Inst37_io_a; // @[Snxn100k.scala 21992:34]
  wire  inst_SnxnLv4Inst37_io_b; // @[Snxn100k.scala 21992:34]
  wire  inst_SnxnLv4Inst37_io_z; // @[Snxn100k.scala 21992:34]
  wire  inst_SnxnLv4Inst38_io_a; // @[Snxn100k.scala 21996:34]
  wire  inst_SnxnLv4Inst38_io_b; // @[Snxn100k.scala 21996:34]
  wire  inst_SnxnLv4Inst38_io_z; // @[Snxn100k.scala 21996:34]
  wire  inst_SnxnLv4Inst39_io_a; // @[Snxn100k.scala 22000:34]
  wire  inst_SnxnLv4Inst39_io_b; // @[Snxn100k.scala 22000:34]
  wire  inst_SnxnLv4Inst39_io_z; // @[Snxn100k.scala 22000:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst36_io_z + inst_SnxnLv4Inst37_io_z; // @[Snxn100k.scala 22004:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst38_io_z; // @[Snxn100k.scala 22004:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst39_io_z; // @[Snxn100k.scala 22004:89]
  SnxnLv4Inst36 inst_SnxnLv4Inst36 ( // @[Snxn100k.scala 21988:34]
    .io_a(inst_SnxnLv4Inst36_io_a),
    .io_b(inst_SnxnLv4Inst36_io_b),
    .io_z(inst_SnxnLv4Inst36_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst37 ( // @[Snxn100k.scala 21992:34]
    .io_a(inst_SnxnLv4Inst37_io_a),
    .io_b(inst_SnxnLv4Inst37_io_b),
    .io_z(inst_SnxnLv4Inst37_io_z)
  );
  SnxnLv4Inst38 inst_SnxnLv4Inst38 ( // @[Snxn100k.scala 21996:34]
    .io_a(inst_SnxnLv4Inst38_io_a),
    .io_b(inst_SnxnLv4Inst38_io_b),
    .io_z(inst_SnxnLv4Inst38_io_z)
  );
  SnxnLv4Inst39 inst_SnxnLv4Inst39 ( // @[Snxn100k.scala 22000:34]
    .io_a(inst_SnxnLv4Inst39_io_a),
    .io_b(inst_SnxnLv4Inst39_io_b),
    .io_z(inst_SnxnLv4Inst39_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22005:15]
  assign inst_SnxnLv4Inst36_io_a = io_a; // @[Snxn100k.scala 21989:27]
  assign inst_SnxnLv4Inst36_io_b = io_b; // @[Snxn100k.scala 21990:27]
  assign inst_SnxnLv4Inst37_io_a = io_a; // @[Snxn100k.scala 21993:27]
  assign inst_SnxnLv4Inst37_io_b = io_b; // @[Snxn100k.scala 21994:27]
  assign inst_SnxnLv4Inst38_io_a = io_a; // @[Snxn100k.scala 21997:27]
  assign inst_SnxnLv4Inst38_io_b = io_b; // @[Snxn100k.scala 21998:27]
  assign inst_SnxnLv4Inst39_io_a = io_a; // @[Snxn100k.scala 22001:27]
  assign inst_SnxnLv4Inst39_io_b = io_b; // @[Snxn100k.scala 22002:27]
endmodule
module SnxnLv4Inst40(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 86962:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 86963:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 86964:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 86965:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 86966:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 86967:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 86968:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 86969:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 86970:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 86971:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 86972:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 86973:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 86974:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 86975:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 86976:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 86977:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 86978:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 86979:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 86980:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 86981:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 86982:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 86983:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 86984:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 86985:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 86986:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 86987:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 86988:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 86989:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 86990:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 86991:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 86992:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 86993:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 86994:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 86995:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 86996:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 86997:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 86998:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 86999:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 87000:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 87001:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 87002:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 87003:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 87004:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 87005:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 87006:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 87007:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 87008:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 87009:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 87010:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 87011:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 87012:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 87013:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 87014:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 87015:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 87016:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 87017:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 87018:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 87019:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 87020:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 87021:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 87022:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 87023:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 87024:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 87025:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 87026:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 87027:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 87028:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 87029:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 87030:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 87031:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 87032:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 87033:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 87034:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 87035:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 87036:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 87037:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 87038:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 87039:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 87040:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 87041:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 87042:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 87043:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 87044:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 87045:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 87046:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 87047:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 87048:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 87049:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 87050:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 87051:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 87052:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 87053:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 87054:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 87055:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 87056:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 87057:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 87058:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 87059:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 87060:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 87061:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 87062:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 87063:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 87064:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 87065:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 87066:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 87067:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 87068:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 87069:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 87070:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 87071:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 87072:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 87073:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 87074:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 87075:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 87076:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 87077:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 87078:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 87079:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 87080:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 87081:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 87082:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 87083:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 87084:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 87085:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 87086:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 87087:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 87088:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 87089:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 87090:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 87091:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 87092:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 87093:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 87094:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 87095:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 87096:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 87097:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 87098:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 87099:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 87100:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 87101:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 87102:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 87103:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 87104:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 87105:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 87106:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 87107:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 87108:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 87109:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 87110:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 87111:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 87112:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 87113:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 87114:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 87115:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 87116:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 87117:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 87118:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 87119:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 87120:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 87121:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 87122:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 87123:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 87124:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 87125:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 87126:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 87127:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 87128:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 87129:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 87130:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 87131:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 87132:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 87133:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 87134:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 87135:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 87136:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 87137:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 87138:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 87139:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 87140:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 87141:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 87142:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 87143:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 87144:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 87145:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 87146:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 87147:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 87148:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 87149:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 87150:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 87151:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 87152:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 87153:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 87154:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 87155:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 87156:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 87157:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 87158:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 87159:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 87160:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 87161:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 87162:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 87163:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 87164:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 87165:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 87166:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 87167:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 87168:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 87169:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 87170:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 87171:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 87172:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 87173:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 87174:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 87175:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 87176:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 87177:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 87178:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 87179:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 87180:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 87181:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 87182:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 87183:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 87184:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 87185:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 87186:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 87187:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 87188:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 87189:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 87190:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 87191:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 87192:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 87193:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 87194:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 87195:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 87196:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 87197:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 87198:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 87199:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 87200:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 87201:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 87202:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 87203:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 87204:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 87205:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 87206:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 87207:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 87208:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 87209:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 87210:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 87211:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 87212:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 87213:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 87214:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 87215:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 87216:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 87217:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 87218:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 87219:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 87220:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 87221:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 87222:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 87223:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 87224:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 87225:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 87226:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 87227:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 87228:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 87229:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 87230:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 87231:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 87232:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 87233:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 87234:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 87235:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 87236:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 87237:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 87238:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 87239:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 87240:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 87241:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 87242:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 87243:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 87244:20]
  assign io_z = ~x70; // @[Snxn100k.scala 87245:16]
endmodule
module SnxnLv4Inst43(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 87566:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 87567:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 87568:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 87569:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 87570:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 87571:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 87572:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 87573:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 87574:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 87575:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 87576:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 87577:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 87578:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 87579:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 87580:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 87581:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 87582:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 87583:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 87584:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 87585:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 87586:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 87587:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 87588:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 87589:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 87590:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 87591:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 87592:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 87593:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 87594:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 87595:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 87596:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 87597:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 87598:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 87599:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 87600:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 87601:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 87602:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 87603:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 87604:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 87605:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 87606:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 87607:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 87608:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 87609:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 87610:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 87611:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 87612:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 87613:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 87614:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 87615:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 87616:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 87617:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 87618:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 87619:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 87620:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 87621:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 87622:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 87623:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 87624:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 87625:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 87626:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 87627:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 87628:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 87629:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 87630:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 87631:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 87632:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 87633:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 87634:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 87635:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 87636:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 87637:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 87638:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 87639:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 87640:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 87641:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 87642:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 87643:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 87644:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 87645:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 87646:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 87647:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 87648:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 87649:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 87650:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 87651:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 87652:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 87653:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 87654:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 87655:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 87656:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 87657:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 87658:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 87659:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 87660:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 87661:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 87662:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 87663:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 87664:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 87665:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 87666:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 87667:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 87668:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 87669:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 87670:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 87671:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 87672:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 87673:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 87674:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 87675:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 87676:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 87677:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 87678:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 87679:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 87680:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 87681:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 87682:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 87683:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 87684:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 87685:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 87686:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 87687:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 87688:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 87689:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 87690:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 87691:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 87692:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 87693:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 87694:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 87695:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 87696:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 87697:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 87698:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 87699:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 87700:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 87701:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 87702:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 87703:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 87704:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 87705:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 87706:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 87707:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 87708:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 87709:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 87710:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 87711:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 87712:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 87713:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 87714:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 87715:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 87716:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 87717:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 87718:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 87719:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 87720:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 87721:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 87722:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 87723:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 87724:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 87725:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 87726:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 87727:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 87728:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 87729:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 87730:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 87731:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 87732:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 87733:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 87734:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 87735:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 87736:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 87737:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 87738:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 87739:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 87740:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 87741:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 87742:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 87743:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 87744:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 87745:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 87746:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 87747:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 87748:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 87749:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 87750:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 87751:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 87752:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 87753:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 87754:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 87755:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 87756:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 87757:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 87758:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 87759:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 87760:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 87761:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 87762:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 87763:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 87764:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 87765:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 87766:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 87767:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 87768:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 87769:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 87770:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 87771:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 87772:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 87773:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 87774:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 87775:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 87776:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 87777:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 87778:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 87779:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 87780:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 87781:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 87782:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 87783:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 87784:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 87785:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 87786:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 87787:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 87788:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 87789:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 87790:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 87791:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 87792:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 87793:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 87794:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 87795:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 87796:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 87797:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 87798:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 87799:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 87800:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 87801:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 87802:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 87803:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 87804:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 87805:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 87806:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 87807:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 87808:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 87809:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 87810:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 87811:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 87812:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 87813:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 87814:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 87815:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 87816:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 87817:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 87818:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 87819:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 87820:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 87821:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 87822:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 87823:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 87824:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 87825:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 87826:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 87827:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 87828:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 87829:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 87830:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 87831:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 87832:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 87833:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 87834:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 87835:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 87836:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 87837:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 87838:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 87839:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 87840:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 87841:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 87842:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 87843:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 87844:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 87845:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 87846:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 87847:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 87848:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 87849:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 87850:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 87851:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 87852:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 87853:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 87854:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 87855:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 87856:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 87857:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 87858:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 87859:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 87860:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 87861:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 87862:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 87863:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 87864:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 87865:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 87866:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 87867:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 87868:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 87869:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 87870:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 87871:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 87872:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 87873:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 87874:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 87875:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 87876:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 87877:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 87878:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 87879:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 87880:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 87881:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 87882:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 87883:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 87884:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 87885:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 87886:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 87887:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 87888:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 87889:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 87890:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 87891:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 87892:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 87893:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 87894:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 87895:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 87896:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 87897:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 87898:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 87899:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 87900:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 87901:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 87902:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 87903:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 87904:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 87905:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 87906:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 87907:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 87908:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 87909:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 87910:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 87911:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 87912:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 87913:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 87914:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 87915:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 87916:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 87917:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 87918:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 87919:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 87920:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 87921:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 87922:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 87923:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 87924:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 87925:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 87926:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 87927:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 87928:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 87929:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 87930:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 87931:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 87932:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 87933:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 87934:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 87935:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 87936:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 87937:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 87938:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 87939:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 87940:20]
  assign io_z = ~x93; // @[Snxn100k.scala 87941:16]
endmodule
module SnxnLv3Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst40_io_a; // @[Snxn100k.scala 22534:34]
  wire  inst_SnxnLv4Inst40_io_b; // @[Snxn100k.scala 22534:34]
  wire  inst_SnxnLv4Inst40_io_z; // @[Snxn100k.scala 22534:34]
  wire  inst_SnxnLv4Inst41_io_a; // @[Snxn100k.scala 22538:34]
  wire  inst_SnxnLv4Inst41_io_b; // @[Snxn100k.scala 22538:34]
  wire  inst_SnxnLv4Inst41_io_z; // @[Snxn100k.scala 22538:34]
  wire  inst_SnxnLv4Inst42_io_a; // @[Snxn100k.scala 22542:34]
  wire  inst_SnxnLv4Inst42_io_b; // @[Snxn100k.scala 22542:34]
  wire  inst_SnxnLv4Inst42_io_z; // @[Snxn100k.scala 22542:34]
  wire  inst_SnxnLv4Inst43_io_a; // @[Snxn100k.scala 22546:34]
  wire  inst_SnxnLv4Inst43_io_b; // @[Snxn100k.scala 22546:34]
  wire  inst_SnxnLv4Inst43_io_z; // @[Snxn100k.scala 22546:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst40_io_z + inst_SnxnLv4Inst41_io_z; // @[Snxn100k.scala 22550:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst42_io_z; // @[Snxn100k.scala 22550:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst43_io_z; // @[Snxn100k.scala 22550:89]
  SnxnLv4Inst40 inst_SnxnLv4Inst40 ( // @[Snxn100k.scala 22534:34]
    .io_a(inst_SnxnLv4Inst40_io_a),
    .io_b(inst_SnxnLv4Inst40_io_b),
    .io_z(inst_SnxnLv4Inst40_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst41 ( // @[Snxn100k.scala 22538:34]
    .io_a(inst_SnxnLv4Inst41_io_a),
    .io_b(inst_SnxnLv4Inst41_io_b),
    .io_z(inst_SnxnLv4Inst41_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst42 ( // @[Snxn100k.scala 22542:34]
    .io_a(inst_SnxnLv4Inst42_io_a),
    .io_b(inst_SnxnLv4Inst42_io_b),
    .io_z(inst_SnxnLv4Inst42_io_z)
  );
  SnxnLv4Inst43 inst_SnxnLv4Inst43 ( // @[Snxn100k.scala 22546:34]
    .io_a(inst_SnxnLv4Inst43_io_a),
    .io_b(inst_SnxnLv4Inst43_io_b),
    .io_z(inst_SnxnLv4Inst43_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22551:15]
  assign inst_SnxnLv4Inst40_io_a = io_a; // @[Snxn100k.scala 22535:27]
  assign inst_SnxnLv4Inst40_io_b = io_b; // @[Snxn100k.scala 22536:27]
  assign inst_SnxnLv4Inst41_io_a = io_a; // @[Snxn100k.scala 22539:27]
  assign inst_SnxnLv4Inst41_io_b = io_b; // @[Snxn100k.scala 22540:27]
  assign inst_SnxnLv4Inst42_io_a = io_a; // @[Snxn100k.scala 22543:27]
  assign inst_SnxnLv4Inst42_io_b = io_b; // @[Snxn100k.scala 22544:27]
  assign inst_SnxnLv4Inst43_io_a = io_a; // @[Snxn100k.scala 22547:27]
  assign inst_SnxnLv4Inst43_io_b = io_b; // @[Snxn100k.scala 22548:27]
endmodule
module SnxnLv3Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst44_io_a; // @[Snxn100k.scala 22259:34]
  wire  inst_SnxnLv4Inst44_io_b; // @[Snxn100k.scala 22259:34]
  wire  inst_SnxnLv4Inst44_io_z; // @[Snxn100k.scala 22259:34]
  wire  inst_SnxnLv4Inst45_io_a; // @[Snxn100k.scala 22263:34]
  wire  inst_SnxnLv4Inst45_io_b; // @[Snxn100k.scala 22263:34]
  wire  inst_SnxnLv4Inst45_io_z; // @[Snxn100k.scala 22263:34]
  wire  inst_SnxnLv4Inst46_io_a; // @[Snxn100k.scala 22267:34]
  wire  inst_SnxnLv4Inst46_io_b; // @[Snxn100k.scala 22267:34]
  wire  inst_SnxnLv4Inst46_io_z; // @[Snxn100k.scala 22267:34]
  wire  inst_SnxnLv4Inst47_io_a; // @[Snxn100k.scala 22271:34]
  wire  inst_SnxnLv4Inst47_io_b; // @[Snxn100k.scala 22271:34]
  wire  inst_SnxnLv4Inst47_io_z; // @[Snxn100k.scala 22271:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst44_io_z + inst_SnxnLv4Inst45_io_z; // @[Snxn100k.scala 22275:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst46_io_z; // @[Snxn100k.scala 22275:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst47_io_z; // @[Snxn100k.scala 22275:89]
  SnxnLv4Inst33 inst_SnxnLv4Inst44 ( // @[Snxn100k.scala 22259:34]
    .io_a(inst_SnxnLv4Inst44_io_a),
    .io_b(inst_SnxnLv4Inst44_io_b),
    .io_z(inst_SnxnLv4Inst44_io_z)
  );
  SnxnLv4Inst4 inst_SnxnLv4Inst45 ( // @[Snxn100k.scala 22263:34]
    .io_a(inst_SnxnLv4Inst45_io_a),
    .io_b(inst_SnxnLv4Inst45_io_b),
    .io_z(inst_SnxnLv4Inst45_io_z)
  );
  SnxnLv4Inst20 inst_SnxnLv4Inst46 ( // @[Snxn100k.scala 22267:34]
    .io_a(inst_SnxnLv4Inst46_io_a),
    .io_b(inst_SnxnLv4Inst46_io_b),
    .io_z(inst_SnxnLv4Inst46_io_z)
  );
  SnxnLv4Inst20 inst_SnxnLv4Inst47 ( // @[Snxn100k.scala 22271:34]
    .io_a(inst_SnxnLv4Inst47_io_a),
    .io_b(inst_SnxnLv4Inst47_io_b),
    .io_z(inst_SnxnLv4Inst47_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22276:15]
  assign inst_SnxnLv4Inst44_io_a = io_a; // @[Snxn100k.scala 22260:27]
  assign inst_SnxnLv4Inst44_io_b = io_b; // @[Snxn100k.scala 22261:27]
  assign inst_SnxnLv4Inst45_io_a = io_a; // @[Snxn100k.scala 22264:27]
  assign inst_SnxnLv4Inst45_io_b = io_b; // @[Snxn100k.scala 22265:27]
  assign inst_SnxnLv4Inst46_io_a = io_a; // @[Snxn100k.scala 22268:27]
  assign inst_SnxnLv4Inst46_io_b = io_b; // @[Snxn100k.scala 22269:27]
  assign inst_SnxnLv4Inst47_io_a = io_a; // @[Snxn100k.scala 22272:27]
  assign inst_SnxnLv4Inst47_io_b = io_b; // @[Snxn100k.scala 22273:27]
endmodule
module SnxnLv2Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst8_io_a; // @[Snxn100k.scala 5381:33]
  wire  inst_SnxnLv3Inst8_io_b; // @[Snxn100k.scala 5381:33]
  wire  inst_SnxnLv3Inst8_io_z; // @[Snxn100k.scala 5381:33]
  wire  inst_SnxnLv3Inst9_io_a; // @[Snxn100k.scala 5385:33]
  wire  inst_SnxnLv3Inst9_io_b; // @[Snxn100k.scala 5385:33]
  wire  inst_SnxnLv3Inst9_io_z; // @[Snxn100k.scala 5385:33]
  wire  inst_SnxnLv3Inst10_io_a; // @[Snxn100k.scala 5389:34]
  wire  inst_SnxnLv3Inst10_io_b; // @[Snxn100k.scala 5389:34]
  wire  inst_SnxnLv3Inst10_io_z; // @[Snxn100k.scala 5389:34]
  wire  inst_SnxnLv3Inst11_io_a; // @[Snxn100k.scala 5393:34]
  wire  inst_SnxnLv3Inst11_io_b; // @[Snxn100k.scala 5393:34]
  wire  inst_SnxnLv3Inst11_io_z; // @[Snxn100k.scala 5393:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst8_io_z + inst_SnxnLv3Inst9_io_z; // @[Snxn100k.scala 5397:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst10_io_z; // @[Snxn100k.scala 5397:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst11_io_z; // @[Snxn100k.scala 5397:87]
  SnxnLv3Inst8 inst_SnxnLv3Inst8 ( // @[Snxn100k.scala 5381:33]
    .io_a(inst_SnxnLv3Inst8_io_a),
    .io_b(inst_SnxnLv3Inst8_io_b),
    .io_z(inst_SnxnLv3Inst8_io_z)
  );
  SnxnLv3Inst9 inst_SnxnLv3Inst9 ( // @[Snxn100k.scala 5385:33]
    .io_a(inst_SnxnLv3Inst9_io_a),
    .io_b(inst_SnxnLv3Inst9_io_b),
    .io_z(inst_SnxnLv3Inst9_io_z)
  );
  SnxnLv3Inst10 inst_SnxnLv3Inst10 ( // @[Snxn100k.scala 5389:34]
    .io_a(inst_SnxnLv3Inst10_io_a),
    .io_b(inst_SnxnLv3Inst10_io_b),
    .io_z(inst_SnxnLv3Inst10_io_z)
  );
  SnxnLv3Inst11 inst_SnxnLv3Inst11 ( // @[Snxn100k.scala 5393:34]
    .io_a(inst_SnxnLv3Inst11_io_a),
    .io_b(inst_SnxnLv3Inst11_io_b),
    .io_z(inst_SnxnLv3Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 5398:15]
  assign inst_SnxnLv3Inst8_io_a = io_a; // @[Snxn100k.scala 5382:26]
  assign inst_SnxnLv3Inst8_io_b = io_b; // @[Snxn100k.scala 5383:26]
  assign inst_SnxnLv3Inst9_io_a = io_a; // @[Snxn100k.scala 5386:26]
  assign inst_SnxnLv3Inst9_io_b = io_b; // @[Snxn100k.scala 5387:26]
  assign inst_SnxnLv3Inst10_io_a = io_a; // @[Snxn100k.scala 5390:27]
  assign inst_SnxnLv3Inst10_io_b = io_b; // @[Snxn100k.scala 5391:27]
  assign inst_SnxnLv3Inst11_io_a = io_a; // @[Snxn100k.scala 5394:27]
  assign inst_SnxnLv3Inst11_io_b = io_b; // @[Snxn100k.scala 5395:27]
endmodule
module SnxnLv4Inst48(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 73942:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 73943:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 73944:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 73945:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 73946:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 73947:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 73948:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 73949:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 73950:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 73951:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 73952:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 73953:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 73954:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 73955:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 73956:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 73957:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 73958:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 73959:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 73960:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 73961:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 73962:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 73963:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 73964:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 73965:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 73966:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 73967:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 73968:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 73969:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 73970:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 73971:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 73972:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 73973:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 73974:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 73975:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 73976:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 73977:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 73978:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 73979:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 73980:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 73981:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 73982:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 73983:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 73984:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 73985:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 73986:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 73987:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 73988:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 73989:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 73990:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 73991:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 73992:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 73993:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 73994:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 73995:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 73996:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 73997:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 73998:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 73999:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 74000:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 74001:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 74002:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 74003:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 74004:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 74005:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 74006:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 74007:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 74008:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 74009:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 74010:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 74011:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 74012:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 74013:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 74014:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 74015:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 74016:20]
  assign io_z = ~x18; // @[Snxn100k.scala 74017:16]
endmodule
module SnxnLv4Inst50(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72972:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72973:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72974:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72975:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72976:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72977:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72978:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 72979:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 72980:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 72981:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 72982:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 72983:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 72984:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 72985:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 72986:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 72987:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 72988:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 72989:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 72990:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 72991:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 72992:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 72993:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 72994:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 72995:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 72996:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72997:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72998:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72999:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 73000:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 73001:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 73002:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 73003:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 73004:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 73005:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 73006:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 73007:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 73008:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 73009:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 73010:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 73011:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 73012:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 73013:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 73014:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 73015:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 73016:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 73017:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 73018:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 73019:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 73020:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 73021:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 73022:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 73023:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 73024:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 73025:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 73026:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 73027:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 73028:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 73029:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 73030:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 73031:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 73032:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 73033:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 73034:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 73035:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 73036:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 73037:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 73038:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 73039:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 73040:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 73041:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 73042:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 73043:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 73044:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 73045:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 73046:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 73047:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 73048:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 73049:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 73050:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 73051:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 73052:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 73053:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 73054:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 73055:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 73056:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 73057:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 73058:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 73059:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 73060:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 73061:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 73062:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 73063:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 73064:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 73065:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 73066:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 73067:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 73068:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 73069:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 73070:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 73071:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 73072:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 73073:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 73074:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 73075:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 73076:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 73077:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 73078:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 73079:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 73080:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 73081:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 73082:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 73083:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 73084:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 73085:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 73086:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 73087:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 73088:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 73089:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 73090:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 73091:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 73092:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 73093:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 73094:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 73095:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 73096:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 73097:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 73098:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 73099:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 73100:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 73101:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 73102:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 73103:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 73104:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 73105:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 73106:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 73107:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 73108:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 73109:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 73110:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 73111:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 73112:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 73113:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 73114:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 73115:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 73116:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 73117:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 73118:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 73119:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 73120:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 73121:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 73122:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 73123:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 73124:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 73125:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 73126:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 73127:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 73128:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 73129:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 73130:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 73131:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 73132:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 73133:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 73134:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 73135:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 73136:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 73137:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 73138:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 73139:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 73140:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 73141:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 73142:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 73143:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 73144:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 73145:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 73146:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 73147:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 73148:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 73149:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 73150:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 73151:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 73152:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 73153:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 73154:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 73155:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 73156:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 73157:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 73158:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 73159:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 73160:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 73161:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 73162:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 73163:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 73164:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 73165:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 73166:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 73167:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 73168:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 73169:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 73170:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 73171:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 73172:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 73173:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 73174:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 73175:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 73176:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 73177:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 73178:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 73179:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 73180:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 73181:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 73182:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 73183:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 73184:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 73185:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 73186:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 73187:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 73188:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 73189:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 73190:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 73191:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 73192:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 73193:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 73194:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 73195:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 73196:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 73197:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 73198:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 73199:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 73200:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 73201:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 73202:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 73203:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 73204:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 73205:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 73206:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 73207:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 73208:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 73209:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 73210:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 73211:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 73212:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 73213:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 73214:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 73215:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 73216:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 73217:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 73218:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 73219:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 73220:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 73221:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 73222:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 73223:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 73224:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 73225:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 73226:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 73227:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 73228:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 73229:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 73230:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 73231:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 73232:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 73233:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 73234:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 73235:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 73236:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 73237:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 73238:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 73239:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 73240:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 73241:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 73242:20]
  assign io_z = ~x67; // @[Snxn100k.scala 73243:16]
endmodule
module SnxnLv3Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst48_io_a; // @[Snxn100k.scala 19652:34]
  wire  inst_SnxnLv4Inst48_io_b; // @[Snxn100k.scala 19652:34]
  wire  inst_SnxnLv4Inst48_io_z; // @[Snxn100k.scala 19652:34]
  wire  inst_SnxnLv4Inst49_io_a; // @[Snxn100k.scala 19656:34]
  wire  inst_SnxnLv4Inst49_io_b; // @[Snxn100k.scala 19656:34]
  wire  inst_SnxnLv4Inst49_io_z; // @[Snxn100k.scala 19656:34]
  wire  inst_SnxnLv4Inst50_io_a; // @[Snxn100k.scala 19660:34]
  wire  inst_SnxnLv4Inst50_io_b; // @[Snxn100k.scala 19660:34]
  wire  inst_SnxnLv4Inst50_io_z; // @[Snxn100k.scala 19660:34]
  wire  inst_SnxnLv4Inst51_io_a; // @[Snxn100k.scala 19664:34]
  wire  inst_SnxnLv4Inst51_io_b; // @[Snxn100k.scala 19664:34]
  wire  inst_SnxnLv4Inst51_io_z; // @[Snxn100k.scala 19664:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst48_io_z + inst_SnxnLv4Inst49_io_z; // @[Snxn100k.scala 19668:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst50_io_z; // @[Snxn100k.scala 19668:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst51_io_z; // @[Snxn100k.scala 19668:89]
  SnxnLv4Inst48 inst_SnxnLv4Inst48 ( // @[Snxn100k.scala 19652:34]
    .io_a(inst_SnxnLv4Inst48_io_a),
    .io_b(inst_SnxnLv4Inst48_io_b),
    .io_z(inst_SnxnLv4Inst48_io_z)
  );
  SnxnLv4Inst15 inst_SnxnLv4Inst49 ( // @[Snxn100k.scala 19656:34]
    .io_a(inst_SnxnLv4Inst49_io_a),
    .io_b(inst_SnxnLv4Inst49_io_b),
    .io_z(inst_SnxnLv4Inst49_io_z)
  );
  SnxnLv4Inst50 inst_SnxnLv4Inst50 ( // @[Snxn100k.scala 19660:34]
    .io_a(inst_SnxnLv4Inst50_io_a),
    .io_b(inst_SnxnLv4Inst50_io_b),
    .io_z(inst_SnxnLv4Inst50_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst51 ( // @[Snxn100k.scala 19664:34]
    .io_a(inst_SnxnLv4Inst51_io_a),
    .io_b(inst_SnxnLv4Inst51_io_b),
    .io_z(inst_SnxnLv4Inst51_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 19669:15]
  assign inst_SnxnLv4Inst48_io_a = io_a; // @[Snxn100k.scala 19653:27]
  assign inst_SnxnLv4Inst48_io_b = io_b; // @[Snxn100k.scala 19654:27]
  assign inst_SnxnLv4Inst49_io_a = io_a; // @[Snxn100k.scala 19657:27]
  assign inst_SnxnLv4Inst49_io_b = io_b; // @[Snxn100k.scala 19658:27]
  assign inst_SnxnLv4Inst50_io_a = io_a; // @[Snxn100k.scala 19661:27]
  assign inst_SnxnLv4Inst50_io_b = io_b; // @[Snxn100k.scala 19662:27]
  assign inst_SnxnLv4Inst51_io_a = io_a; // @[Snxn100k.scala 19665:27]
  assign inst_SnxnLv4Inst51_io_b = io_b; // @[Snxn100k.scala 19666:27]
endmodule
module SnxnLv4Inst52(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 74306:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 74307:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 74308:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 74309:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 74310:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 74311:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 74312:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 74313:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 74314:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 74315:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 74316:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 74317:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 74318:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 74319:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 74320:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 74321:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 74322:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 74323:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 74324:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 74325:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 74326:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 74327:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 74328:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 74329:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 74330:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 74331:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 74332:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 74333:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 74334:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 74335:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 74336:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 74337:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 74338:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 74339:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 74340:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 74341:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 74342:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 74343:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 74344:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 74345:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 74346:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 74347:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 74348:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 74349:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 74350:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 74351:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 74352:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 74353:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 74354:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 74355:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 74356:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 74357:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 74358:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 74359:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 74360:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 74361:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 74362:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 74363:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 74364:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 74365:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 74366:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 74367:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 74368:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 74369:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 74370:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 74371:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 74372:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 74373:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 74374:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 74375:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 74376:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 74377:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 74378:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 74379:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 74380:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 74381:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 74382:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 74383:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 74384:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 74385:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 74386:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 74387:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 74388:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 74389:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 74390:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 74391:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 74392:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 74393:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 74394:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 74395:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 74396:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 74397:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 74398:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 74399:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 74400:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 74401:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 74402:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 74403:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 74404:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 74405:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 74406:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 74407:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 74408:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 74409:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 74410:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 74411:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 74412:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 74413:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 74414:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 74415:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 74416:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 74417:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 74418:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 74419:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 74420:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 74421:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 74422:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 74423:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 74424:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 74425:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 74426:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 74427:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 74428:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 74429:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 74430:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 74431:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 74432:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 74433:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 74434:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 74435:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 74436:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 74437:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 74438:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 74439:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 74440:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 74441:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 74442:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 74443:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 74444:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 74445:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 74446:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 74447:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 74448:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 74449:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 74450:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 74451:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 74452:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 74453:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 74454:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 74455:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 74456:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 74457:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 74458:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 74459:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 74460:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 74461:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 74462:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 74463:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 74464:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 74465:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 74466:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 74467:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 74468:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 74469:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 74470:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 74471:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 74472:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 74473:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 74474:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 74475:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 74476:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 74477:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 74478:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 74479:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 74480:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 74481:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 74482:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 74483:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 74484:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 74485:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 74486:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 74487:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 74488:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 74489:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 74490:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 74491:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 74492:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 74493:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 74494:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 74495:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 74496:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 74497:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 74498:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 74499:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 74500:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 74501:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 74502:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 74503:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 74504:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 74505:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 74506:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 74507:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 74508:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 74509:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 74510:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 74511:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 74512:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 74513:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 74514:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 74515:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 74516:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 74517:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 74518:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 74519:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 74520:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 74521:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 74522:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 74523:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 74524:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 74525:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 74526:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 74527:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 74528:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 74529:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 74530:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 74531:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 74532:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 74533:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 74534:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 74535:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 74536:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 74537:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 74538:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 74539:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 74540:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 74541:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 74542:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 74543:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 74544:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 74545:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 74546:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 74547:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 74548:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 74549:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 74550:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 74551:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 74552:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 74553:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 74554:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 74555:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 74556:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 74557:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 74558:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 74559:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 74560:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 74561:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 74562:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 74563:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 74564:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 74565:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 74566:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 74567:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 74568:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 74569:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 74570:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 74571:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 74572:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 74573:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 74574:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 74575:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 74576:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 74577:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 74578:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 74579:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 74580:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 74581:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 74582:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 74583:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 74584:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 74585:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 74586:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 74587:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 74588:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 74589:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 74590:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 74591:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 74592:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 74593:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 74594:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 74595:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 74596:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 74597:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 74598:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 74599:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 74600:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 74601:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 74602:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 74603:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 74604:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 74605:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 74606:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 74607:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 74608:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 74609:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 74610:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 74611:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 74612:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 74613:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 74614:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 74615:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 74616:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 74617:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 74618:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 74619:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 74620:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 74621:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 74622:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 74623:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 74624:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 74625:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 74626:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 74627:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 74628:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 74629:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 74630:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 74631:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 74632:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 74633:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 74634:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 74635:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 74636:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 74637:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 74638:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 74639:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 74640:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 74641:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 74642:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 74643:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 74644:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 74645:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 74646:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 74647:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 74648:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 74649:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 74650:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 74651:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 74652:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 74653:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 74654:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 74655:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 74656:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 74657:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 74658:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 74659:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 74660:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 74661:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 74662:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 74663:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 74664:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 74665:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 74666:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 74667:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 74668:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 74669:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 74670:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 74671:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 74672:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 74673:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 74674:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 74675:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 74676:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 74677:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 74678:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 74679:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 74680:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 74681:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 74682:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 74683:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 74684:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 74685:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 74686:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 74687:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 74688:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 74689:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 74690:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 74691:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 74692:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 74693:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 74694:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 74695:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 74696:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 74697:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 74698:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 74699:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 74700:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 74701:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 74702:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 74703:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 74704:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 74705:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 74706:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 74707:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 74708:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 74709:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 74710:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 74711:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 74712:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 74713:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 74714:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 74715:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 74716:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 74717:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 74718:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 74719:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 74720:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 74721:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 74722:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 74723:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 74724:22]
  assign io_z = ~x104; // @[Snxn100k.scala 74725:17]
endmodule
module SnxnLv4Inst54(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75166:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75167:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75168:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75169:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75170:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75171:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75172:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75173:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75174:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75175:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75176:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75177:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75178:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75179:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75180:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75181:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75182:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75183:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75184:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75185:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75186:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75187:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75188:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75189:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75190:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75191:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75192:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75193:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75194:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75195:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75196:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75197:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75198:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 75199:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 75200:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 75201:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 75202:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 75203:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 75204:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 75205:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 75206:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 75207:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 75208:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 75209:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 75210:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 75211:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 75212:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 75213:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 75214:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 75215:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 75216:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 75217:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 75218:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 75219:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 75220:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 75221:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 75222:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 75223:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 75224:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 75225:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 75226:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 75227:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 75228:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 75229:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 75230:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 75231:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 75232:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 75233:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 75234:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 75235:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 75236:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 75237:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 75238:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 75239:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 75240:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 75241:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 75242:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 75243:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 75244:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 75245:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 75246:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 75247:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 75248:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 75249:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 75250:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 75251:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 75252:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 75253:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 75254:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 75255:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 75256:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 75257:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 75258:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 75259:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 75260:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 75261:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 75262:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 75263:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 75264:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 75265:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 75266:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 75267:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 75268:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 75269:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 75270:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 75271:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 75272:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 75273:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 75274:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 75275:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 75276:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 75277:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 75278:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 75279:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 75280:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 75281:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 75282:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 75283:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 75284:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 75285:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 75286:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 75287:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 75288:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 75289:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 75290:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 75291:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 75292:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 75293:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 75294:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 75295:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 75296:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 75297:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 75298:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 75299:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 75300:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 75301:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 75302:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 75303:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 75304:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 75305:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 75306:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 75307:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 75308:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 75309:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 75310:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 75311:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 75312:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 75313:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 75314:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 75315:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 75316:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 75317:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 75318:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 75319:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 75320:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 75321:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 75322:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 75323:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 75324:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 75325:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 75326:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 75327:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 75328:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 75329:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 75330:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 75331:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 75332:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 75333:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 75334:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 75335:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 75336:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 75337:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 75338:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 75339:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 75340:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 75341:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 75342:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 75343:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 75344:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 75345:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 75346:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 75347:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 75348:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 75349:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 75350:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 75351:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 75352:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 75353:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 75354:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 75355:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 75356:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 75357:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 75358:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 75359:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 75360:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 75361:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 75362:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 75363:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 75364:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 75365:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 75366:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 75367:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 75368:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 75369:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 75370:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 75371:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 75372:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 75373:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 75374:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 75375:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 75376:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 75377:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 75378:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 75379:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 75380:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 75381:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 75382:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 75383:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 75384:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 75385:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 75386:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 75387:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 75388:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 75389:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 75390:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 75391:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 75392:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 75393:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 75394:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 75395:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 75396:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 75397:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 75398:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 75399:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 75400:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 75401:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 75402:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 75403:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 75404:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 75405:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 75406:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 75407:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 75408:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 75409:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 75410:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 75411:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 75412:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 75413:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 75414:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 75415:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 75416:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 75417:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 75418:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 75419:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 75420:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 75421:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 75422:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 75423:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 75424:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 75425:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 75426:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 75427:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 75428:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 75429:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 75430:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 75431:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 75432:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 75433:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 75434:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 75435:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 75436:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 75437:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 75438:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 75439:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 75440:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 75441:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 75442:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 75443:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 75444:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 75445:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 75446:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 75447:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 75448:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 75449:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 75450:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 75451:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 75452:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 75453:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 75454:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 75455:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 75456:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 75457:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 75458:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 75459:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 75460:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 75461:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 75462:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 75463:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 75464:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 75465:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 75466:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 75467:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 75468:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 75469:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 75470:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 75471:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 75472:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 75473:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 75474:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 75475:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 75476:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 75477:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 75478:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 75479:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 75480:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 75481:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 75482:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 75483:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 75484:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 75485:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 75486:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 75487:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 75488:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 75489:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 75490:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 75491:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 75492:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 75493:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 75494:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 75495:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 75496:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 75497:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 75498:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 75499:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 75500:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 75501:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 75502:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 75503:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 75504:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 75505:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 75506:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 75507:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 75508:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 75509:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 75510:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 75511:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 75512:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 75513:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 75514:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 75515:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 75516:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 75517:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 75518:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 75519:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 75520:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 75521:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 75522:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 75523:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 75524:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 75525:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 75526:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 75527:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 75528:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 75529:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 75530:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 75531:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 75532:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 75533:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 75534:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 75535:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 75536:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 75537:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 75538:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 75539:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 75540:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 75541:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 75542:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 75543:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 75544:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 75545:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 75546:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 75547:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 75548:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 75549:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 75550:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 75551:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 75552:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 75553:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 75554:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 75555:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 75556:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 75557:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 75558:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 75559:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 75560:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 75561:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 75562:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 75563:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 75564:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 75565:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 75566:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 75567:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 75568:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 75569:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 75570:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 75571:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 75572:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 75573:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 75574:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 75575:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 75576:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 75577:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 75578:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 75579:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 75580:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 75581:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 75582:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 75583:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 75584:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 75585:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 75586:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 75587:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 75588:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 75589:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 75590:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 75591:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 75592:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 75593:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 75594:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 75595:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 75596:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 75597:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 75598:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 75599:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 75600:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 75601:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 75602:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 75603:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 75604:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 75605:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 75606:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 75607:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 75608:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 75609:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 75610:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 75611:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 75612:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 75613:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 75614:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 75615:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 75616:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 75617:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 75618:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 75619:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 75620:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 75621:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 75622:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 75623:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 75624:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 75625:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 75626:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 75627:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 75628:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 75629:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 75630:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 75631:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 75632:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 75633:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 75634:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 75635:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 75636:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 75637:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 75638:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 75639:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 75640:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 75641:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 75642:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 75643:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 75644:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 75645:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 75646:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 75647:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 75648:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 75649:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 75650:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 75651:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 75652:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 75653:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 75654:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 75655:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 75656:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 75657:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 75658:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 75659:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 75660:22]
  assign io_z = ~x123; // @[Snxn100k.scala 75661:17]
endmodule
module SnxnLv3Inst13(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst52_io_a; // @[Snxn100k.scala 19991:34]
  wire  inst_SnxnLv4Inst52_io_b; // @[Snxn100k.scala 19991:34]
  wire  inst_SnxnLv4Inst52_io_z; // @[Snxn100k.scala 19991:34]
  wire  inst_SnxnLv4Inst53_io_a; // @[Snxn100k.scala 19995:34]
  wire  inst_SnxnLv4Inst53_io_b; // @[Snxn100k.scala 19995:34]
  wire  inst_SnxnLv4Inst53_io_z; // @[Snxn100k.scala 19995:34]
  wire  inst_SnxnLv4Inst54_io_a; // @[Snxn100k.scala 19999:34]
  wire  inst_SnxnLv4Inst54_io_b; // @[Snxn100k.scala 19999:34]
  wire  inst_SnxnLv4Inst54_io_z; // @[Snxn100k.scala 19999:34]
  wire  inst_SnxnLv4Inst55_io_a; // @[Snxn100k.scala 20003:34]
  wire  inst_SnxnLv4Inst55_io_b; // @[Snxn100k.scala 20003:34]
  wire  inst_SnxnLv4Inst55_io_z; // @[Snxn100k.scala 20003:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst52_io_z + inst_SnxnLv4Inst53_io_z; // @[Snxn100k.scala 20007:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst54_io_z; // @[Snxn100k.scala 20007:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst55_io_z; // @[Snxn100k.scala 20007:89]
  SnxnLv4Inst52 inst_SnxnLv4Inst52 ( // @[Snxn100k.scala 19991:34]
    .io_a(inst_SnxnLv4Inst52_io_a),
    .io_b(inst_SnxnLv4Inst52_io_b),
    .io_z(inst_SnxnLv4Inst52_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst53 ( // @[Snxn100k.scala 19995:34]
    .io_a(inst_SnxnLv4Inst53_io_a),
    .io_b(inst_SnxnLv4Inst53_io_b),
    .io_z(inst_SnxnLv4Inst53_io_z)
  );
  SnxnLv4Inst54 inst_SnxnLv4Inst54 ( // @[Snxn100k.scala 19999:34]
    .io_a(inst_SnxnLv4Inst54_io_a),
    .io_b(inst_SnxnLv4Inst54_io_b),
    .io_z(inst_SnxnLv4Inst54_io_z)
  );
  SnxnLv4Inst52 inst_SnxnLv4Inst55 ( // @[Snxn100k.scala 20003:34]
    .io_a(inst_SnxnLv4Inst55_io_a),
    .io_b(inst_SnxnLv4Inst55_io_b),
    .io_z(inst_SnxnLv4Inst55_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 20008:15]
  assign inst_SnxnLv4Inst52_io_a = io_a; // @[Snxn100k.scala 19992:27]
  assign inst_SnxnLv4Inst52_io_b = io_b; // @[Snxn100k.scala 19993:27]
  assign inst_SnxnLv4Inst53_io_a = io_a; // @[Snxn100k.scala 19996:27]
  assign inst_SnxnLv4Inst53_io_b = io_b; // @[Snxn100k.scala 19997:27]
  assign inst_SnxnLv4Inst54_io_a = io_a; // @[Snxn100k.scala 20000:27]
  assign inst_SnxnLv4Inst54_io_b = io_b; // @[Snxn100k.scala 20001:27]
  assign inst_SnxnLv4Inst55_io_a = io_a; // @[Snxn100k.scala 20004:27]
  assign inst_SnxnLv4Inst55_io_b = io_b; // @[Snxn100k.scala 20005:27]
endmodule
module SnxnLv4Inst56(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 77796:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 77797:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 77798:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 77799:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 77800:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 77801:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 77802:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 77803:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 77804:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 77805:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 77806:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 77807:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 77808:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 77809:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 77810:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 77811:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 77812:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 77813:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 77814:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 77815:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 77816:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 77817:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 77818:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 77819:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 77820:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 77821:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 77822:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 77823:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 77824:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 77825:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 77826:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 77827:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 77828:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 77829:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 77830:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 77831:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 77832:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 77833:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 77834:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 77835:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 77836:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 77837:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 77838:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 77839:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 77840:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 77841:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 77842:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 77843:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 77844:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 77845:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 77846:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 77847:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 77848:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 77849:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 77850:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 77851:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 77852:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 77853:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 77854:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 77855:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 77856:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 77857:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 77858:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 77859:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 77860:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 77861:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 77862:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 77863:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 77864:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 77865:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 77866:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 77867:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 77868:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 77869:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 77870:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 77871:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 77872:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 77873:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 77874:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 77875:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 77876:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 77877:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 77878:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 77879:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 77880:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 77881:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 77882:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 77883:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 77884:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 77885:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 77886:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 77887:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 77888:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 77889:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 77890:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 77891:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 77892:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 77893:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 77894:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 77895:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 77896:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 77897:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 77898:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 77899:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 77900:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 77901:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 77902:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 77903:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 77904:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 77905:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 77906:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 77907:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 77908:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 77909:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 77910:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 77911:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 77912:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 77913:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 77914:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 77915:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 77916:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 77917:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 77918:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 77919:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 77920:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 77921:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 77922:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 77923:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 77924:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 77925:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 77926:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 77927:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 77928:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 77929:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 77930:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 77931:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 77932:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 77933:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 77934:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 77935:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 77936:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 77937:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 77938:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 77939:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 77940:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 77941:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 77942:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 77943:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 77944:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 77945:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 77946:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 77947:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 77948:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 77949:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 77950:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 77951:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 77952:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 77953:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 77954:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 77955:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 77956:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 77957:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 77958:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 77959:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 77960:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 77961:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 77962:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 77963:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 77964:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 77965:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 77966:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 77967:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 77968:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 77969:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 77970:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 77971:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 77972:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 77973:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 77974:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 77975:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 77976:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 77977:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 77978:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 77979:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 77980:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 77981:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 77982:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 77983:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 77984:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 77985:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 77986:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 77987:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 77988:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 77989:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 77990:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 77991:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 77992:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 77993:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 77994:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 77995:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 77996:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 77997:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 77998:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 77999:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 78000:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 78001:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 78002:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 78003:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 78004:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 78005:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 78006:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 78007:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 78008:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 78009:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 78010:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 78011:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 78012:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 78013:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 78014:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 78015:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 78016:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 78017:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 78018:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 78019:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 78020:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 78021:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 78022:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 78023:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 78024:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 78025:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 78026:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 78027:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 78028:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 78029:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 78030:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 78031:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 78032:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 78033:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 78034:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 78035:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 78036:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 78037:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 78038:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 78039:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 78040:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 78041:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 78042:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 78043:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 78044:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 78045:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 78046:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 78047:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 78048:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 78049:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 78050:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 78051:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 78052:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 78053:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 78054:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 78055:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 78056:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 78057:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 78058:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 78059:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 78060:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 78061:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 78062:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 78063:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 78064:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 78065:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 78066:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 78067:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 78068:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 78069:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 78070:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 78071:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 78072:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 78073:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 78074:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 78075:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 78076:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 78077:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 78078:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 78079:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 78080:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 78081:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 78082:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 78083:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 78084:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 78085:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 78086:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 78087:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 78088:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 78089:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 78090:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 78091:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 78092:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 78093:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 78094:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 78095:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 78096:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 78097:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 78098:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 78099:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 78100:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 78101:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 78102:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 78103:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 78104:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 78105:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 78106:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 78107:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 78108:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 78109:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 78110:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 78111:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 78112:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 78113:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 78114:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 78115:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 78116:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 78117:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 78118:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 78119:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 78120:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 78121:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 78122:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 78123:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 78124:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 78125:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 78126:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 78127:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 78128:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 78129:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 78130:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 78131:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 78132:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 78133:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 78134:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 78135:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 78136:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 78137:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 78138:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 78139:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 78140:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 78141:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 78142:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 78143:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 78144:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 78145:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 78146:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 78147:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 78148:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 78149:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 78150:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 78151:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 78152:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 78153:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 78154:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 78155:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 78156:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 78157:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 78158:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 78159:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 78160:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 78161:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 78162:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 78163:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 78164:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 78165:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 78166:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 78167:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 78168:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 78169:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 78170:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 78171:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 78172:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 78173:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 78174:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 78175:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 78176:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 78177:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 78178:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 78179:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 78180:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 78181:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 78182:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 78183:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 78184:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 78185:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 78186:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 78187:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 78188:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 78189:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 78190:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 78191:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 78192:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 78193:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 78194:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 78195:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 78196:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 78197:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 78198:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 78199:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 78200:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 78201:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 78202:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 78203:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 78204:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 78205:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 78206:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 78207:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 78208:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 78209:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 78210:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 78211:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 78212:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 78213:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 78214:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 78215:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 78216:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 78217:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 78218:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 78219:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 78220:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 78221:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 78222:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 78223:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 78224:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 78225:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 78226:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 78227:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 78228:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 78229:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 78230:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 78231:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 78232:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 78233:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 78234:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 78235:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 78236:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 78237:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 78238:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 78239:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 78240:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 78241:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 78242:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 78243:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 78244:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 78245:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 78246:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 78247:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 78248:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 78249:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 78250:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 78251:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 78252:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 78253:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 78254:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 78255:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 78256:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 78257:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 78258:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 78259:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 78260:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 78261:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 78262:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 78263:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 78264:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 78265:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 78266:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 78267:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 78268:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 78269:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 78270:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 78271:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 78272:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 78273:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 78274:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 78275:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 78276:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 78277:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 78278:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 78279:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 78280:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 78281:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 78282:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 78283:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 78284:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 78285:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 78286:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 78287:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 78288:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 78289:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 78290:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 78291:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 78292:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 78293:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 78294:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 78295:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 78296:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 78297:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 78298:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 78299:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 78300:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 78301:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 78302:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 78303:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 78304:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 78305:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 78306:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 78307:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 78308:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 78309:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 78310:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 78311:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 78312:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 78313:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 78314:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 78315:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 78316:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 78317:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 78318:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 78319:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 78320:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 78321:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 78322:22]
  assign io_z = ~x131; // @[Snxn100k.scala 78323:17]
endmodule
module SnxnLv4Inst58(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78334:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78335:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78336:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78337:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78338:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78339:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78340:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78341:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78342:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78343:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78344:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78345:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78346:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78347:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78348:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78349:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78350:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78351:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78352:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78353:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78354:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78355:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78356:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78357:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78358:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78359:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78360:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78361:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78362:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78363:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78364:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78365:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78366:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78367:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78368:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78369:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78370:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78371:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78372:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78373:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78374:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78375:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78376:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78377:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78378:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78379:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78380:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78381:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78382:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78383:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78384:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78385:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78386:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78387:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78388:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78389:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78390:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78391:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78392:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78393:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78394:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78395:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78396:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78397:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78398:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78399:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78400:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78401:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78402:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78403:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78404:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 78405:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 78406:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 78407:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 78408:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 78409:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 78410:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 78411:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 78412:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 78413:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 78414:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 78415:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 78416:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 78417:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 78418:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 78419:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 78420:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 78421:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 78422:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 78423:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 78424:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 78425:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 78426:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 78427:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 78428:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 78429:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 78430:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 78431:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 78432:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 78433:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 78434:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 78435:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 78436:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 78437:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 78438:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 78439:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 78440:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 78441:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 78442:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 78443:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 78444:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 78445:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 78446:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 78447:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 78448:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 78449:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 78450:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 78451:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 78452:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 78453:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 78454:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 78455:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 78456:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 78457:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 78458:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 78459:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 78460:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 78461:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 78462:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 78463:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 78464:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 78465:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 78466:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 78467:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 78468:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 78469:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 78470:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 78471:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 78472:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 78473:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 78474:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 78475:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 78476:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 78477:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 78478:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 78479:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 78480:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 78481:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 78482:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 78483:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 78484:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 78485:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 78486:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 78487:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 78488:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 78489:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 78490:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 78491:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 78492:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 78493:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 78494:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 78495:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 78496:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 78497:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 78498:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 78499:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 78500:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 78501:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 78502:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 78503:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 78504:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 78505:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 78506:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 78507:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 78508:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 78509:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 78510:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 78511:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 78512:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 78513:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 78514:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 78515:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 78516:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 78517:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 78518:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 78519:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 78520:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 78521:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 78522:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 78523:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 78524:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 78525:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 78526:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 78527:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 78528:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 78529:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 78530:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 78531:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 78532:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 78533:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 78534:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 78535:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 78536:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 78537:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 78538:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 78539:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 78540:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 78541:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 78542:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 78543:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 78544:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 78545:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 78546:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 78547:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 78548:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 78549:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 78550:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 78551:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 78552:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 78553:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 78554:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 78555:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 78556:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 78557:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 78558:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 78559:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 78560:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 78561:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 78562:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 78563:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 78564:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 78565:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 78566:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 78567:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 78568:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 78569:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 78570:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 78571:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 78572:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 78573:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 78574:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 78575:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 78576:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 78577:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 78578:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 78579:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 78580:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 78581:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 78582:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 78583:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 78584:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 78585:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 78586:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 78587:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 78588:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 78589:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 78590:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 78591:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 78592:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 78593:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 78594:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 78595:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 78596:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 78597:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 78598:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 78599:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 78600:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 78601:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 78602:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 78603:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 78604:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 78605:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 78606:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 78607:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 78608:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 78609:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 78610:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 78611:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 78612:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 78613:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 78614:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 78615:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 78616:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 78617:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 78618:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 78619:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 78620:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 78621:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 78622:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 78623:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 78624:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 78625:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 78626:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 78627:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 78628:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 78629:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 78630:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 78631:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 78632:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 78633:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 78634:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 78635:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 78636:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 78637:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 78638:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 78639:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 78640:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 78641:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 78642:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 78643:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 78644:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 78645:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 78646:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 78647:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 78648:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 78649:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 78650:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 78651:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 78652:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 78653:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 78654:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 78655:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 78656:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 78657:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 78658:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 78659:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 78660:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 78661:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 78662:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 78663:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 78664:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 78665:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 78666:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 78667:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 78668:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 78669:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 78670:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 78671:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 78672:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 78673:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 78674:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 78675:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 78676:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 78677:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 78678:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 78679:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 78680:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 78681:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 78682:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 78683:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 78684:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 78685:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 78686:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 78687:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 78688:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 78689:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 78690:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 78691:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 78692:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 78693:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 78694:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 78695:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 78696:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 78697:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 78698:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 78699:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 78700:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 78701:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 78702:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 78703:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 78704:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 78705:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 78706:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 78707:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 78708:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 78709:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 78710:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 78711:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 78712:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 78713:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 78714:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 78715:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 78716:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 78717:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 78718:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 78719:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 78720:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 78721:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 78722:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 78723:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 78724:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 78725:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 78726:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 78727:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 78728:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 78729:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 78730:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 78731:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 78732:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 78733:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 78734:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 78735:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 78736:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 78737:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 78738:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 78739:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 78740:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 78741:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 78742:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 78743:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 78744:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 78745:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 78746:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 78747:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 78748:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 78749:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 78750:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 78751:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 78752:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 78753:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 78754:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 78755:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 78756:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 78757:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 78758:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 78759:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 78760:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 78761:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 78762:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 78763:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 78764:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 78765:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 78766:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 78767:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 78768:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 78769:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 78770:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 78771:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 78772:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 78773:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 78774:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 78775:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 78776:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 78777:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 78778:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 78779:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 78780:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 78781:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 78782:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 78783:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 78784:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 78785:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 78786:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 78787:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 78788:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 78789:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 78790:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 78791:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 78792:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 78793:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 78794:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 78795:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 78796:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 78797:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 78798:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 78799:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 78800:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 78801:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 78802:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 78803:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 78804:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 78805:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 78806:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 78807:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 78808:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 78809:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 78810:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 78811:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 78812:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 78813:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 78814:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 78815:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 78816:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 78817:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 78818:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 78819:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 78820:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 78821:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 78822:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 78823:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 78824:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 78825:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 78826:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 78827:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 78828:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 78829:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 78830:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 78831:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 78832:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 78833:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 78834:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 78835:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 78836:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 78837:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 78838:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 78839:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 78840:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 78841:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 78842:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 78843:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 78844:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 78845:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 78846:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 78847:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 78848:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 78849:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 78850:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 78851:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 78852:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 78853:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 78854:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 78855:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 78856:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 78857:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 78858:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 78859:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 78860:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 78861:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 78862:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 78863:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 78864:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 78865:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 78866:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 78867:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 78868:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 78869:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 78870:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 78871:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 78872:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 78873:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 78874:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 78875:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 78876:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 78877:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 78878:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 78879:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 78880:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 78881:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 78882:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 78883:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 78884:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 78885:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 78886:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 78887:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 78888:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 78889:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 78890:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 78891:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 78892:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 78893:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 78894:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 78895:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 78896:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 78897:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 78898:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 78899:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 78900:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 78901:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 78902:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 78903:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 78904:22]
  wire  invx142 = ~x142; // @[Snxn100k.scala 78905:17]
  wire  t143 = x142 + invx142; // @[Snxn100k.scala 78906:22]
  wire  inv143 = ~t143; // @[Snxn100k.scala 78907:17]
  wire  x143 = t143 ^ inv143; // @[Snxn100k.scala 78908:22]
  wire  invx143 = ~x143; // @[Snxn100k.scala 78909:17]
  wire  t144 = x143 + invx143; // @[Snxn100k.scala 78910:22]
  wire  inv144 = ~t144; // @[Snxn100k.scala 78911:17]
  wire  x144 = t144 ^ inv144; // @[Snxn100k.scala 78912:22]
  wire  invx144 = ~x144; // @[Snxn100k.scala 78913:17]
  wire  t145 = x144 + invx144; // @[Snxn100k.scala 78914:22]
  wire  inv145 = ~t145; // @[Snxn100k.scala 78915:17]
  wire  x145 = t145 ^ inv145; // @[Snxn100k.scala 78916:22]
  wire  invx145 = ~x145; // @[Snxn100k.scala 78917:17]
  wire  t146 = x145 + invx145; // @[Snxn100k.scala 78918:22]
  wire  inv146 = ~t146; // @[Snxn100k.scala 78919:17]
  wire  x146 = t146 ^ inv146; // @[Snxn100k.scala 78920:22]
  wire  invx146 = ~x146; // @[Snxn100k.scala 78921:17]
  wire  t147 = x146 + invx146; // @[Snxn100k.scala 78922:22]
  wire  inv147 = ~t147; // @[Snxn100k.scala 78923:17]
  wire  x147 = t147 ^ inv147; // @[Snxn100k.scala 78924:22]
  assign io_z = ~x147; // @[Snxn100k.scala 78925:17]
endmodule
module SnxnLv3Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst56_io_a; // @[Snxn100k.scala 20709:34]
  wire  inst_SnxnLv4Inst56_io_b; // @[Snxn100k.scala 20709:34]
  wire  inst_SnxnLv4Inst56_io_z; // @[Snxn100k.scala 20709:34]
  wire  inst_SnxnLv4Inst57_io_a; // @[Snxn100k.scala 20713:34]
  wire  inst_SnxnLv4Inst57_io_b; // @[Snxn100k.scala 20713:34]
  wire  inst_SnxnLv4Inst57_io_z; // @[Snxn100k.scala 20713:34]
  wire  inst_SnxnLv4Inst58_io_a; // @[Snxn100k.scala 20717:34]
  wire  inst_SnxnLv4Inst58_io_b; // @[Snxn100k.scala 20717:34]
  wire  inst_SnxnLv4Inst58_io_z; // @[Snxn100k.scala 20717:34]
  wire  inst_SnxnLv4Inst59_io_a; // @[Snxn100k.scala 20721:34]
  wire  inst_SnxnLv4Inst59_io_b; // @[Snxn100k.scala 20721:34]
  wire  inst_SnxnLv4Inst59_io_z; // @[Snxn100k.scala 20721:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst56_io_z + inst_SnxnLv4Inst57_io_z; // @[Snxn100k.scala 20725:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst58_io_z; // @[Snxn100k.scala 20725:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst59_io_z; // @[Snxn100k.scala 20725:89]
  SnxnLv4Inst56 inst_SnxnLv4Inst56 ( // @[Snxn100k.scala 20709:34]
    .io_a(inst_SnxnLv4Inst56_io_a),
    .io_b(inst_SnxnLv4Inst56_io_b),
    .io_z(inst_SnxnLv4Inst56_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst57 ( // @[Snxn100k.scala 20713:34]
    .io_a(inst_SnxnLv4Inst57_io_a),
    .io_b(inst_SnxnLv4Inst57_io_b),
    .io_z(inst_SnxnLv4Inst57_io_z)
  );
  SnxnLv4Inst58 inst_SnxnLv4Inst58 ( // @[Snxn100k.scala 20717:34]
    .io_a(inst_SnxnLv4Inst58_io_a),
    .io_b(inst_SnxnLv4Inst58_io_b),
    .io_z(inst_SnxnLv4Inst58_io_z)
  );
  SnxnLv4Inst35 inst_SnxnLv4Inst59 ( // @[Snxn100k.scala 20721:34]
    .io_a(inst_SnxnLv4Inst59_io_a),
    .io_b(inst_SnxnLv4Inst59_io_b),
    .io_z(inst_SnxnLv4Inst59_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 20726:15]
  assign inst_SnxnLv4Inst56_io_a = io_a; // @[Snxn100k.scala 20710:27]
  assign inst_SnxnLv4Inst56_io_b = io_b; // @[Snxn100k.scala 20711:27]
  assign inst_SnxnLv4Inst57_io_a = io_a; // @[Snxn100k.scala 20714:27]
  assign inst_SnxnLv4Inst57_io_b = io_b; // @[Snxn100k.scala 20715:27]
  assign inst_SnxnLv4Inst58_io_a = io_a; // @[Snxn100k.scala 20718:27]
  assign inst_SnxnLv4Inst58_io_b = io_b; // @[Snxn100k.scala 20719:27]
  assign inst_SnxnLv4Inst59_io_a = io_a; // @[Snxn100k.scala 20722:27]
  assign inst_SnxnLv4Inst59_io_b = io_b; // @[Snxn100k.scala 20723:27]
endmodule
module SnxnLv3Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst60_io_a; // @[Snxn100k.scala 20334:34]
  wire  inst_SnxnLv4Inst60_io_b; // @[Snxn100k.scala 20334:34]
  wire  inst_SnxnLv4Inst60_io_z; // @[Snxn100k.scala 20334:34]
  wire  inst_SnxnLv4Inst61_io_a; // @[Snxn100k.scala 20338:34]
  wire  inst_SnxnLv4Inst61_io_b; // @[Snxn100k.scala 20338:34]
  wire  inst_SnxnLv4Inst61_io_z; // @[Snxn100k.scala 20338:34]
  wire  inst_SnxnLv4Inst62_io_a; // @[Snxn100k.scala 20342:34]
  wire  inst_SnxnLv4Inst62_io_b; // @[Snxn100k.scala 20342:34]
  wire  inst_SnxnLv4Inst62_io_z; // @[Snxn100k.scala 20342:34]
  wire  inst_SnxnLv4Inst63_io_a; // @[Snxn100k.scala 20346:34]
  wire  inst_SnxnLv4Inst63_io_b; // @[Snxn100k.scala 20346:34]
  wire  inst_SnxnLv4Inst63_io_z; // @[Snxn100k.scala 20346:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst60_io_z + inst_SnxnLv4Inst61_io_z; // @[Snxn100k.scala 20350:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst62_io_z; // @[Snxn100k.scala 20350:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst63_io_z; // @[Snxn100k.scala 20350:89]
  SnxnLv4Inst7 inst_SnxnLv4Inst60 ( // @[Snxn100k.scala 20334:34]
    .io_a(inst_SnxnLv4Inst60_io_a),
    .io_b(inst_SnxnLv4Inst60_io_b),
    .io_z(inst_SnxnLv4Inst60_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst61 ( // @[Snxn100k.scala 20338:34]
    .io_a(inst_SnxnLv4Inst61_io_a),
    .io_b(inst_SnxnLv4Inst61_io_b),
    .io_z(inst_SnxnLv4Inst61_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst62 ( // @[Snxn100k.scala 20342:34]
    .io_a(inst_SnxnLv4Inst62_io_a),
    .io_b(inst_SnxnLv4Inst62_io_b),
    .io_z(inst_SnxnLv4Inst62_io_z)
  );
  SnxnLv4Inst15 inst_SnxnLv4Inst63 ( // @[Snxn100k.scala 20346:34]
    .io_a(inst_SnxnLv4Inst63_io_a),
    .io_b(inst_SnxnLv4Inst63_io_b),
    .io_z(inst_SnxnLv4Inst63_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 20351:15]
  assign inst_SnxnLv4Inst60_io_a = io_a; // @[Snxn100k.scala 20335:27]
  assign inst_SnxnLv4Inst60_io_b = io_b; // @[Snxn100k.scala 20336:27]
  assign inst_SnxnLv4Inst61_io_a = io_a; // @[Snxn100k.scala 20339:27]
  assign inst_SnxnLv4Inst61_io_b = io_b; // @[Snxn100k.scala 20340:27]
  assign inst_SnxnLv4Inst62_io_a = io_a; // @[Snxn100k.scala 20343:27]
  assign inst_SnxnLv4Inst62_io_b = io_b; // @[Snxn100k.scala 20344:27]
  assign inst_SnxnLv4Inst63_io_a = io_a; // @[Snxn100k.scala 20347:27]
  assign inst_SnxnLv4Inst63_io_b = io_b; // @[Snxn100k.scala 20348:27]
endmodule
module SnxnLv2Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst12_io_a; // @[Snxn100k.scala 4483:34]
  wire  inst_SnxnLv3Inst12_io_b; // @[Snxn100k.scala 4483:34]
  wire  inst_SnxnLv3Inst12_io_z; // @[Snxn100k.scala 4483:34]
  wire  inst_SnxnLv3Inst13_io_a; // @[Snxn100k.scala 4487:34]
  wire  inst_SnxnLv3Inst13_io_b; // @[Snxn100k.scala 4487:34]
  wire  inst_SnxnLv3Inst13_io_z; // @[Snxn100k.scala 4487:34]
  wire  inst_SnxnLv3Inst14_io_a; // @[Snxn100k.scala 4491:34]
  wire  inst_SnxnLv3Inst14_io_b; // @[Snxn100k.scala 4491:34]
  wire  inst_SnxnLv3Inst14_io_z; // @[Snxn100k.scala 4491:34]
  wire  inst_SnxnLv3Inst15_io_a; // @[Snxn100k.scala 4495:34]
  wire  inst_SnxnLv3Inst15_io_b; // @[Snxn100k.scala 4495:34]
  wire  inst_SnxnLv3Inst15_io_z; // @[Snxn100k.scala 4495:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst12_io_z + inst_SnxnLv3Inst13_io_z; // @[Snxn100k.scala 4499:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst14_io_z; // @[Snxn100k.scala 4499:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst15_io_z; // @[Snxn100k.scala 4499:89]
  SnxnLv3Inst12 inst_SnxnLv3Inst12 ( // @[Snxn100k.scala 4483:34]
    .io_a(inst_SnxnLv3Inst12_io_a),
    .io_b(inst_SnxnLv3Inst12_io_b),
    .io_z(inst_SnxnLv3Inst12_io_z)
  );
  SnxnLv3Inst13 inst_SnxnLv3Inst13 ( // @[Snxn100k.scala 4487:34]
    .io_a(inst_SnxnLv3Inst13_io_a),
    .io_b(inst_SnxnLv3Inst13_io_b),
    .io_z(inst_SnxnLv3Inst13_io_z)
  );
  SnxnLv3Inst14 inst_SnxnLv3Inst14 ( // @[Snxn100k.scala 4491:34]
    .io_a(inst_SnxnLv3Inst14_io_a),
    .io_b(inst_SnxnLv3Inst14_io_b),
    .io_z(inst_SnxnLv3Inst14_io_z)
  );
  SnxnLv3Inst15 inst_SnxnLv3Inst15 ( // @[Snxn100k.scala 4495:34]
    .io_a(inst_SnxnLv3Inst15_io_a),
    .io_b(inst_SnxnLv3Inst15_io_b),
    .io_z(inst_SnxnLv3Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 4500:15]
  assign inst_SnxnLv3Inst12_io_a = io_a; // @[Snxn100k.scala 4484:27]
  assign inst_SnxnLv3Inst12_io_b = io_b; // @[Snxn100k.scala 4485:27]
  assign inst_SnxnLv3Inst13_io_a = io_a; // @[Snxn100k.scala 4488:27]
  assign inst_SnxnLv3Inst13_io_b = io_b; // @[Snxn100k.scala 4489:27]
  assign inst_SnxnLv3Inst14_io_a = io_a; // @[Snxn100k.scala 4492:27]
  assign inst_SnxnLv3Inst14_io_b = io_b; // @[Snxn100k.scala 4493:27]
  assign inst_SnxnLv3Inst15_io_a = io_a; // @[Snxn100k.scala 4496:27]
  assign inst_SnxnLv3Inst15_io_b = io_b; // @[Snxn100k.scala 4497:27]
endmodule
module SnxnLv1Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst0_io_a; // @[Snxn100k.scala 1218:33]
  wire  inst_SnxnLv2Inst0_io_b; // @[Snxn100k.scala 1218:33]
  wire  inst_SnxnLv2Inst0_io_z; // @[Snxn100k.scala 1218:33]
  wire  inst_SnxnLv2Inst1_io_a; // @[Snxn100k.scala 1222:33]
  wire  inst_SnxnLv2Inst1_io_b; // @[Snxn100k.scala 1222:33]
  wire  inst_SnxnLv2Inst1_io_z; // @[Snxn100k.scala 1222:33]
  wire  inst_SnxnLv2Inst2_io_a; // @[Snxn100k.scala 1226:33]
  wire  inst_SnxnLv2Inst2_io_b; // @[Snxn100k.scala 1226:33]
  wire  inst_SnxnLv2Inst2_io_z; // @[Snxn100k.scala 1226:33]
  wire  inst_SnxnLv2Inst3_io_a; // @[Snxn100k.scala 1230:33]
  wire  inst_SnxnLv2Inst3_io_b; // @[Snxn100k.scala 1230:33]
  wire  inst_SnxnLv2Inst3_io_z; // @[Snxn100k.scala 1230:33]
  wire  _sum_T_1 = inst_SnxnLv2Inst0_io_z + inst_SnxnLv2Inst1_io_z; // @[Snxn100k.scala 1234:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst2_io_z; // @[Snxn100k.scala 1234:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst3_io_z; // @[Snxn100k.scala 1234:86]
  SnxnLv2Inst0 inst_SnxnLv2Inst0 ( // @[Snxn100k.scala 1218:33]
    .io_a(inst_SnxnLv2Inst0_io_a),
    .io_b(inst_SnxnLv2Inst0_io_b),
    .io_z(inst_SnxnLv2Inst0_io_z)
  );
  SnxnLv2Inst1 inst_SnxnLv2Inst1 ( // @[Snxn100k.scala 1222:33]
    .io_a(inst_SnxnLv2Inst1_io_a),
    .io_b(inst_SnxnLv2Inst1_io_b),
    .io_z(inst_SnxnLv2Inst1_io_z)
  );
  SnxnLv2Inst2 inst_SnxnLv2Inst2 ( // @[Snxn100k.scala 1226:33]
    .io_a(inst_SnxnLv2Inst2_io_a),
    .io_b(inst_SnxnLv2Inst2_io_b),
    .io_z(inst_SnxnLv2Inst2_io_z)
  );
  SnxnLv2Inst3 inst_SnxnLv2Inst3 ( // @[Snxn100k.scala 1230:33]
    .io_a(inst_SnxnLv2Inst3_io_a),
    .io_b(inst_SnxnLv2Inst3_io_b),
    .io_z(inst_SnxnLv2Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1235:15]
  assign inst_SnxnLv2Inst0_io_a = io_a; // @[Snxn100k.scala 1219:26]
  assign inst_SnxnLv2Inst0_io_b = io_b; // @[Snxn100k.scala 1220:26]
  assign inst_SnxnLv2Inst1_io_a = io_a; // @[Snxn100k.scala 1223:26]
  assign inst_SnxnLv2Inst1_io_b = io_b; // @[Snxn100k.scala 1224:26]
  assign inst_SnxnLv2Inst2_io_a = io_a; // @[Snxn100k.scala 1227:26]
  assign inst_SnxnLv2Inst2_io_b = io_b; // @[Snxn100k.scala 1228:26]
  assign inst_SnxnLv2Inst3_io_a = io_a; // @[Snxn100k.scala 1231:26]
  assign inst_SnxnLv2Inst3_io_b = io_b; // @[Snxn100k.scala 1232:26]
endmodule
module SnxnLv4Inst64(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 34616:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 34617:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 34618:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 34619:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 34620:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 34621:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 34622:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 34623:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 34624:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 34625:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 34626:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 34627:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 34628:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 34629:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 34630:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 34631:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 34632:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 34633:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 34634:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 34635:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 34636:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 34637:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 34638:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 34639:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 34640:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 34641:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 34642:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 34643:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 34644:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 34645:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 34646:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 34647:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 34648:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 34649:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 34650:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 34651:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 34652:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 34653:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 34654:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 34655:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 34656:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 34657:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 34658:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 34659:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 34660:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 34661:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 34662:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 34663:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 34664:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 34665:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 34666:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 34667:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 34668:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 34669:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 34670:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 34671:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 34672:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 34673:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 34674:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 34675:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 34676:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 34677:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 34678:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 34679:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 34680:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 34681:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 34682:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 34683:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 34684:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 34685:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 34686:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 34687:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 34688:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 34689:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 34690:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 34691:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 34692:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 34693:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 34694:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 34695:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 34696:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 34697:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 34698:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 34699:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 34700:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 34701:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 34702:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 34703:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 34704:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 34705:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 34706:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 34707:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 34708:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 34709:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 34710:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 34711:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 34712:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 34713:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 34714:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 34715:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 34716:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 34717:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 34718:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 34719:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 34720:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 34721:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 34722:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 34723:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 34724:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 34725:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 34726:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 34727:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 34728:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 34729:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 34730:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 34731:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 34732:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 34733:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 34734:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 34735:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 34736:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 34737:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 34738:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 34739:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 34740:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 34741:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 34742:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 34743:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 34744:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 34745:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 34746:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 34747:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 34748:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 34749:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 34750:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 34751:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 34752:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 34753:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 34754:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 34755:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 34756:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 34757:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 34758:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 34759:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 34760:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 34761:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 34762:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 34763:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 34764:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 34765:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 34766:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 34767:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 34768:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 34769:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 34770:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 34771:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 34772:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 34773:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 34774:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 34775:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 34776:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 34777:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 34778:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 34779:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 34780:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 34781:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 34782:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 34783:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 34784:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 34785:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 34786:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 34787:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 34788:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 34789:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 34790:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 34791:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 34792:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 34793:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 34794:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 34795:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 34796:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 34797:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 34798:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 34799:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 34800:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 34801:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 34802:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 34803:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 34804:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 34805:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 34806:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 34807:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 34808:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 34809:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 34810:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 34811:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 34812:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 34813:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 34814:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 34815:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 34816:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 34817:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 34818:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 34819:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 34820:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 34821:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 34822:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 34823:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 34824:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 34825:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 34826:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 34827:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 34828:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 34829:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 34830:20]
  assign io_z = ~x53; // @[Snxn100k.scala 34831:16]
endmodule
module SnxnLv3Inst16(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst64_io_a; // @[Snxn100k.scala 9690:34]
  wire  inst_SnxnLv4Inst64_io_b; // @[Snxn100k.scala 9690:34]
  wire  inst_SnxnLv4Inst64_io_z; // @[Snxn100k.scala 9690:34]
  wire  inst_SnxnLv4Inst65_io_a; // @[Snxn100k.scala 9694:34]
  wire  inst_SnxnLv4Inst65_io_b; // @[Snxn100k.scala 9694:34]
  wire  inst_SnxnLv4Inst65_io_z; // @[Snxn100k.scala 9694:34]
  wire  inst_SnxnLv4Inst66_io_a; // @[Snxn100k.scala 9698:34]
  wire  inst_SnxnLv4Inst66_io_b; // @[Snxn100k.scala 9698:34]
  wire  inst_SnxnLv4Inst66_io_z; // @[Snxn100k.scala 9698:34]
  wire  inst_SnxnLv4Inst67_io_a; // @[Snxn100k.scala 9702:34]
  wire  inst_SnxnLv4Inst67_io_b; // @[Snxn100k.scala 9702:34]
  wire  inst_SnxnLv4Inst67_io_z; // @[Snxn100k.scala 9702:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst64_io_z + inst_SnxnLv4Inst65_io_z; // @[Snxn100k.scala 9706:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst66_io_z; // @[Snxn100k.scala 9706:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst67_io_z; // @[Snxn100k.scala 9706:89]
  SnxnLv4Inst64 inst_SnxnLv4Inst64 ( // @[Snxn100k.scala 9690:34]
    .io_a(inst_SnxnLv4Inst64_io_a),
    .io_b(inst_SnxnLv4Inst64_io_b),
    .io_z(inst_SnxnLv4Inst64_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst65 ( // @[Snxn100k.scala 9694:34]
    .io_a(inst_SnxnLv4Inst65_io_a),
    .io_b(inst_SnxnLv4Inst65_io_b),
    .io_z(inst_SnxnLv4Inst65_io_z)
  );
  SnxnLv4Inst19 inst_SnxnLv4Inst66 ( // @[Snxn100k.scala 9698:34]
    .io_a(inst_SnxnLv4Inst66_io_a),
    .io_b(inst_SnxnLv4Inst66_io_b),
    .io_z(inst_SnxnLv4Inst66_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst67 ( // @[Snxn100k.scala 9702:34]
    .io_a(inst_SnxnLv4Inst67_io_a),
    .io_b(inst_SnxnLv4Inst67_io_b),
    .io_z(inst_SnxnLv4Inst67_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 9707:15]
  assign inst_SnxnLv4Inst64_io_a = io_a; // @[Snxn100k.scala 9691:27]
  assign inst_SnxnLv4Inst64_io_b = io_b; // @[Snxn100k.scala 9692:27]
  assign inst_SnxnLv4Inst65_io_a = io_a; // @[Snxn100k.scala 9695:27]
  assign inst_SnxnLv4Inst65_io_b = io_b; // @[Snxn100k.scala 9696:27]
  assign inst_SnxnLv4Inst66_io_a = io_a; // @[Snxn100k.scala 9699:27]
  assign inst_SnxnLv4Inst66_io_b = io_b; // @[Snxn100k.scala 9700:27]
  assign inst_SnxnLv4Inst67_io_a = io_a; // @[Snxn100k.scala 9703:27]
  assign inst_SnxnLv4Inst67_io_b = io_b; // @[Snxn100k.scala 9704:27]
endmodule
module SnxnLv4Inst68(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 32938:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 32939:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 32940:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 32941:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 32942:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 32943:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 32944:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 32945:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 32946:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 32947:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 32948:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 32949:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 32950:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 32951:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 32952:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 32953:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 32954:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 32955:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 32956:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 32957:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 32958:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 32959:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 32960:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 32961:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 32962:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 32963:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 32964:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 32965:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 32966:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 32967:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 32968:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 32969:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 32970:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 32971:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 32972:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 32973:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 32974:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 32975:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 32976:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 32977:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 32978:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 32979:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 32980:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 32981:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 32982:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 32983:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 32984:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 32985:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 32986:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 32987:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 32988:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 32989:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 32990:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 32991:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 32992:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 32993:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 32994:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 32995:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 32996:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 32997:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 32998:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 32999:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 33000:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 33001:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 33002:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 33003:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 33004:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 33005:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 33006:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 33007:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 33008:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 33009:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 33010:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 33011:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 33012:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 33013:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 33014:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 33015:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 33016:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 33017:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 33018:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 33019:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 33020:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 33021:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 33022:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 33023:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 33024:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 33025:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 33026:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 33027:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 33028:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 33029:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 33030:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 33031:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 33032:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 33033:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 33034:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 33035:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 33036:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 33037:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 33038:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 33039:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 33040:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 33041:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 33042:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 33043:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 33044:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 33045:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 33046:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 33047:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 33048:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 33049:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 33050:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 33051:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 33052:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 33053:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 33054:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 33055:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 33056:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 33057:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 33058:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 33059:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 33060:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 33061:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 33062:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 33063:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 33064:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 33065:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 33066:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 33067:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 33068:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 33069:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 33070:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 33071:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 33072:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 33073:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 33074:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 33075:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 33076:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 33077:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 33078:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 33079:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 33080:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 33081:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 33082:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 33083:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 33084:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 33085:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 33086:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 33087:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 33088:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 33089:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 33090:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 33091:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 33092:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 33093:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 33094:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 33095:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 33096:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 33097:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 33098:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 33099:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 33100:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 33101:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 33102:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 33103:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 33104:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 33105:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 33106:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 33107:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 33108:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 33109:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 33110:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 33111:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 33112:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 33113:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 33114:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 33115:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 33116:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 33117:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 33118:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 33119:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 33120:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 33121:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 33122:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 33123:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 33124:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 33125:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 33126:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 33127:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 33128:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 33129:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 33130:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 33131:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 33132:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 33133:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 33134:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 33135:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 33136:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 33137:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 33138:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 33139:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 33140:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 33141:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 33142:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 33143:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 33144:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 33145:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 33146:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 33147:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 33148:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 33149:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 33150:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 33151:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 33152:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 33153:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 33154:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 33155:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 33156:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 33157:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 33158:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 33159:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 33160:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 33161:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 33162:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 33163:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 33164:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 33165:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 33166:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 33167:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 33168:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 33169:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 33170:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 33171:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 33172:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 33173:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 33174:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 33175:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 33176:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 33177:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 33178:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 33179:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 33180:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 33181:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 33182:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 33183:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 33184:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 33185:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 33186:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 33187:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 33188:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 33189:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 33190:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 33191:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 33192:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 33193:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 33194:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 33195:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 33196:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 33197:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 33198:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 33199:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 33200:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 33201:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 33202:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 33203:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 33204:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 33205:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 33206:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 33207:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 33208:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 33209:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 33210:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 33211:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 33212:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 33213:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 33214:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 33215:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 33216:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 33217:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 33218:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 33219:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 33220:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 33221:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 33222:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 33223:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 33224:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 33225:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 33226:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 33227:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 33228:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 33229:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 33230:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 33231:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 33232:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 33233:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 33234:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 33235:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 33236:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 33237:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 33238:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 33239:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 33240:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 33241:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 33242:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 33243:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 33244:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 33245:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 33246:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 33247:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 33248:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 33249:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 33250:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 33251:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 33252:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 33253:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 33254:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 33255:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 33256:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 33257:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 33258:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 33259:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 33260:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 33261:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 33262:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 33263:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 33264:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 33265:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 33266:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 33267:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 33268:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 33269:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 33270:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 33271:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 33272:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 33273:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 33274:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 33275:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 33276:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 33277:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 33278:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 33279:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 33280:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 33281:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 33282:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 33283:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 33284:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 33285:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 33286:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 33287:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 33288:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 33289:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 33290:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 33291:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 33292:20]
  assign io_z = ~x88; // @[Snxn100k.scala 33293:16]
endmodule
module SnxnLv4Inst69(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 32112:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 32113:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 32114:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 32115:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 32116:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 32117:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 32118:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 32119:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 32120:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 32121:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 32122:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 32123:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 32124:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 32125:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 32126:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 32127:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 32128:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 32129:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 32130:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 32131:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 32132:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 32133:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 32134:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 32135:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 32136:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 32137:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 32138:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 32139:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 32140:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 32141:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 32142:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 32143:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 32144:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 32145:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 32146:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 32147:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 32148:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 32149:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 32150:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 32151:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 32152:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 32153:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 32154:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 32155:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 32156:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 32157:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 32158:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 32159:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 32160:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 32161:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 32162:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 32163:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 32164:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 32165:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 32166:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 32167:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 32168:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 32169:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 32170:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 32171:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 32172:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 32173:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 32174:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 32175:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 32176:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 32177:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 32178:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 32179:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 32180:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 32181:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 32182:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 32183:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 32184:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 32185:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 32186:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 32187:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 32188:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 32189:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 32190:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 32191:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 32192:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 32193:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 32194:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 32195:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 32196:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 32197:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 32198:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 32199:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 32200:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 32201:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 32202:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 32203:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 32204:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 32205:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 32206:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 32207:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 32208:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 32209:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 32210:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 32211:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 32212:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 32213:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 32214:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 32215:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 32216:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 32217:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 32218:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 32219:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 32220:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 32221:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 32222:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 32223:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 32224:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 32225:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 32226:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 32227:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 32228:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 32229:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 32230:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 32231:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 32232:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 32233:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 32234:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 32235:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 32236:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 32237:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 32238:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 32239:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 32240:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 32241:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 32242:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 32243:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 32244:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 32245:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 32246:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 32247:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 32248:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 32249:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 32250:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 32251:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 32252:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 32253:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 32254:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 32255:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 32256:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 32257:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 32258:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 32259:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 32260:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 32261:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 32262:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 32263:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 32264:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 32265:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 32266:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 32267:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 32268:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 32269:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 32270:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 32271:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 32272:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 32273:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 32274:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 32275:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 32276:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 32277:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 32278:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 32279:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 32280:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 32281:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 32282:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 32283:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 32284:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 32285:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 32286:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 32287:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 32288:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 32289:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 32290:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 32291:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 32292:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 32293:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 32294:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 32295:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 32296:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 32297:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 32298:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 32299:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 32300:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 32301:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 32302:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 32303:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 32304:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 32305:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 32306:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 32307:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 32308:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 32309:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 32310:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 32311:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 32312:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 32313:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 32314:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 32315:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 32316:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 32317:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 32318:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 32319:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 32320:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 32321:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 32322:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 32323:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 32324:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 32325:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 32326:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 32327:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 32328:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 32329:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 32330:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 32331:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 32332:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 32333:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 32334:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 32335:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 32336:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 32337:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 32338:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 32339:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 32340:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 32341:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 32342:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 32343:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 32344:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 32345:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 32346:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 32347:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 32348:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 32349:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 32350:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 32351:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 32352:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 32353:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 32354:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 32355:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 32356:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 32357:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 32358:20]
  assign io_z = ~x61; // @[Snxn100k.scala 32359:16]
endmodule
module SnxnLv3Inst17(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst68_io_a; // @[Snxn100k.scala 8884:34]
  wire  inst_SnxnLv4Inst68_io_b; // @[Snxn100k.scala 8884:34]
  wire  inst_SnxnLv4Inst68_io_z; // @[Snxn100k.scala 8884:34]
  wire  inst_SnxnLv4Inst69_io_a; // @[Snxn100k.scala 8888:34]
  wire  inst_SnxnLv4Inst69_io_b; // @[Snxn100k.scala 8888:34]
  wire  inst_SnxnLv4Inst69_io_z; // @[Snxn100k.scala 8888:34]
  wire  inst_SnxnLv4Inst70_io_a; // @[Snxn100k.scala 8892:34]
  wire  inst_SnxnLv4Inst70_io_b; // @[Snxn100k.scala 8892:34]
  wire  inst_SnxnLv4Inst70_io_z; // @[Snxn100k.scala 8892:34]
  wire  inst_SnxnLv4Inst71_io_a; // @[Snxn100k.scala 8896:34]
  wire  inst_SnxnLv4Inst71_io_b; // @[Snxn100k.scala 8896:34]
  wire  inst_SnxnLv4Inst71_io_z; // @[Snxn100k.scala 8896:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst68_io_z + inst_SnxnLv4Inst69_io_z; // @[Snxn100k.scala 8900:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst70_io_z; // @[Snxn100k.scala 8900:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst71_io_z; // @[Snxn100k.scala 8900:89]
  SnxnLv4Inst68 inst_SnxnLv4Inst68 ( // @[Snxn100k.scala 8884:34]
    .io_a(inst_SnxnLv4Inst68_io_a),
    .io_b(inst_SnxnLv4Inst68_io_b),
    .io_z(inst_SnxnLv4Inst68_io_z)
  );
  SnxnLv4Inst69 inst_SnxnLv4Inst69 ( // @[Snxn100k.scala 8888:34]
    .io_a(inst_SnxnLv4Inst69_io_a),
    .io_b(inst_SnxnLv4Inst69_io_b),
    .io_z(inst_SnxnLv4Inst69_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst70 ( // @[Snxn100k.scala 8892:34]
    .io_a(inst_SnxnLv4Inst70_io_a),
    .io_b(inst_SnxnLv4Inst70_io_b),
    .io_z(inst_SnxnLv4Inst70_io_z)
  );
  SnxnLv4Inst16 inst_SnxnLv4Inst71 ( // @[Snxn100k.scala 8896:34]
    .io_a(inst_SnxnLv4Inst71_io_a),
    .io_b(inst_SnxnLv4Inst71_io_b),
    .io_z(inst_SnxnLv4Inst71_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 8901:15]
  assign inst_SnxnLv4Inst68_io_a = io_a; // @[Snxn100k.scala 8885:27]
  assign inst_SnxnLv4Inst68_io_b = io_b; // @[Snxn100k.scala 8886:27]
  assign inst_SnxnLv4Inst69_io_a = io_a; // @[Snxn100k.scala 8889:27]
  assign inst_SnxnLv4Inst69_io_b = io_b; // @[Snxn100k.scala 8890:27]
  assign inst_SnxnLv4Inst70_io_a = io_a; // @[Snxn100k.scala 8893:27]
  assign inst_SnxnLv4Inst70_io_b = io_b; // @[Snxn100k.scala 8894:27]
  assign inst_SnxnLv4Inst71_io_a = io_a; // @[Snxn100k.scala 8897:27]
  assign inst_SnxnLv4Inst71_io_b = io_b; // @[Snxn100k.scala 8898:27]
endmodule
module SnxnLv4Inst73(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 34142:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 34143:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 34144:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 34145:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 34146:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 34147:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 34148:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 34149:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 34150:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 34151:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 34152:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 34153:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 34154:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 34155:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 34156:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 34157:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 34158:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 34159:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 34160:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 34161:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 34162:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 34163:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 34164:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 34165:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 34166:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 34167:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 34168:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 34169:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 34170:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 34171:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 34172:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 34173:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 34174:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 34175:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 34176:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 34177:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 34178:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 34179:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 34180:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 34181:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 34182:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 34183:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 34184:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 34185:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 34186:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 34187:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 34188:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 34189:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 34190:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 34191:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 34192:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 34193:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 34194:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 34195:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 34196:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 34197:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 34198:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 34199:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 34200:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 34201:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 34202:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 34203:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 34204:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 34205:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 34206:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 34207:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 34208:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 34209:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 34210:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 34211:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 34212:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 34213:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 34214:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 34215:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 34216:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 34217:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 34218:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 34219:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 34220:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 34221:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 34222:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 34223:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 34224:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 34225:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 34226:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 34227:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 34228:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 34229:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 34230:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 34231:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 34232:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 34233:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 34234:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 34235:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 34236:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 34237:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 34238:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 34239:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 34240:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 34241:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 34242:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 34243:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 34244:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 34245:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 34246:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 34247:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 34248:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 34249:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 34250:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 34251:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 34252:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 34253:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 34254:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 34255:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 34256:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 34257:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 34258:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 34259:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 34260:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 34261:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 34262:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 34263:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 34264:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 34265:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 34266:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 34267:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 34268:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 34269:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 34270:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 34271:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 34272:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 34273:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 34274:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 34275:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 34276:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 34277:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 34278:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 34279:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 34280:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 34281:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 34282:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 34283:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 34284:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 34285:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 34286:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 34287:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 34288:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 34289:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 34290:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 34291:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 34292:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 34293:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 34294:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 34295:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 34296:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 34297:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 34298:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 34299:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 34300:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 34301:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 34302:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 34303:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 34304:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 34305:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 34306:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 34307:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 34308:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 34309:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 34310:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 34311:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 34312:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 34313:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 34314:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 34315:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 34316:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 34317:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 34318:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 34319:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 34320:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 34321:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 34322:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 34323:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 34324:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 34325:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 34326:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 34327:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 34328:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 34329:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 34330:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 34331:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 34332:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 34333:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 34334:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 34335:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 34336:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 34337:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 34338:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 34339:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 34340:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 34341:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 34342:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 34343:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 34344:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 34345:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 34346:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 34347:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 34348:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 34349:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 34350:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 34351:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 34352:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 34353:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 34354:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 34355:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 34356:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 34357:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 34358:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 34359:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 34360:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 34361:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 34362:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 34363:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 34364:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 34365:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 34366:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 34367:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 34368:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 34369:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 34370:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 34371:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 34372:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 34373:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 34374:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 34375:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 34376:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 34377:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 34378:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 34379:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 34380:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 34381:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 34382:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 34383:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 34384:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 34385:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 34386:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 34387:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 34388:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 34389:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 34390:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 34391:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 34392:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 34393:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 34394:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 34395:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 34396:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 34397:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 34398:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 34399:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 34400:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 34401:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 34402:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 34403:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 34404:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 34405:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 34406:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 34407:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 34408:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 34409:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 34410:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 34411:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 34412:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 34413:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 34414:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 34415:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 34416:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 34417:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 34418:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 34419:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 34420:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 34421:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 34422:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 34423:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 34424:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 34425:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 34426:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 34427:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 34428:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 34429:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 34430:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 34431:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 34432:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 34433:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 34434:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 34435:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 34436:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 34437:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 34438:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 34439:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 34440:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 34441:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 34442:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 34443:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 34444:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 34445:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 34446:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 34447:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 34448:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 34449:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 34450:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 34451:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 34452:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 34453:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 34454:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 34455:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 34456:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 34457:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 34458:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 34459:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 34460:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 34461:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 34462:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 34463:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 34464:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 34465:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 34466:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 34467:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 34468:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 34469:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 34470:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 34471:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 34472:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 34473:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 34474:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 34475:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 34476:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 34477:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 34478:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 34479:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 34480:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 34481:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 34482:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 34483:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 34484:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 34485:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 34486:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 34487:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 34488:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 34489:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 34490:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 34491:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 34492:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 34493:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 34494:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 34495:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 34496:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 34497:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 34498:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 34499:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 34500:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 34501:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 34502:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 34503:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 34504:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 34505:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 34506:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 34507:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 34508:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 34509:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 34510:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 34511:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 34512:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 34513:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 34514:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 34515:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 34516:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 34517:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 34518:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 34519:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 34520:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 34521:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 34522:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 34523:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 34524:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 34525:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 34526:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 34527:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 34528:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 34529:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 34530:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 34531:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 34532:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 34533:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 34534:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 34535:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 34536:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 34537:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 34538:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 34539:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 34540:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 34541:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 34542:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 34543:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 34544:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 34545:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 34546:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 34547:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 34548:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 34549:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 34550:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 34551:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 34552:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 34553:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 34554:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 34555:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 34556:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 34557:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 34558:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 34559:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 34560:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 34561:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 34562:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 34563:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 34564:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 34565:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 34566:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 34567:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 34568:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 34569:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 34570:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 34571:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 34572:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 34573:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 34574:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 34575:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 34576:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 34577:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 34578:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 34579:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 34580:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 34581:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 34582:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 34583:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 34584:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 34585:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 34586:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 34587:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 34588:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 34589:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 34590:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 34591:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 34592:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 34593:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 34594:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 34595:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 34596:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 34597:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 34598:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 34599:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 34600:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 34601:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 34602:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 34603:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 34604:22]
  assign io_z = ~x115; // @[Snxn100k.scala 34605:17]
endmodule
module SnxnLv4Inst74(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 33304:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 33305:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 33306:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 33307:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 33308:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 33309:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 33310:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 33311:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 33312:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 33313:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 33314:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 33315:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 33316:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 33317:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 33318:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 33319:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 33320:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 33321:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 33322:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 33323:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 33324:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 33325:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 33326:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 33327:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 33328:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 33329:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 33330:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 33331:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 33332:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 33333:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 33334:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 33335:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 33336:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 33337:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 33338:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 33339:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 33340:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 33341:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 33342:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 33343:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 33344:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 33345:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 33346:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 33347:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 33348:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 33349:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 33350:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 33351:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 33352:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 33353:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 33354:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 33355:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 33356:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 33357:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 33358:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 33359:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 33360:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 33361:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 33362:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 33363:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 33364:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 33365:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 33366:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 33367:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 33368:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 33369:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 33370:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 33371:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 33372:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 33373:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 33374:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 33375:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 33376:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 33377:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 33378:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 33379:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 33380:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 33381:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 33382:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 33383:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 33384:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 33385:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 33386:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 33387:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 33388:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 33389:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 33390:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 33391:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 33392:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 33393:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 33394:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 33395:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 33396:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 33397:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 33398:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 33399:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 33400:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 33401:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 33402:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 33403:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 33404:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 33405:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 33406:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 33407:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 33408:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 33409:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 33410:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 33411:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 33412:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 33413:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 33414:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 33415:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 33416:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 33417:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 33418:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 33419:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 33420:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 33421:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 33422:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 33423:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 33424:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 33425:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 33426:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 33427:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 33428:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 33429:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 33430:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 33431:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 33432:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 33433:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 33434:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 33435:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 33436:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 33437:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 33438:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 33439:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 33440:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 33441:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 33442:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 33443:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 33444:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 33445:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 33446:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 33447:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 33448:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 33449:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 33450:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 33451:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 33452:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 33453:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 33454:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 33455:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 33456:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 33457:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 33458:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 33459:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 33460:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 33461:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 33462:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 33463:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 33464:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 33465:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 33466:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 33467:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 33468:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 33469:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 33470:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 33471:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 33472:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 33473:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 33474:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 33475:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 33476:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 33477:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 33478:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 33479:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 33480:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 33481:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 33482:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 33483:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 33484:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 33485:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 33486:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 33487:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 33488:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 33489:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 33490:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 33491:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 33492:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 33493:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 33494:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 33495:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 33496:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 33497:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 33498:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 33499:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 33500:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 33501:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 33502:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 33503:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 33504:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 33505:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 33506:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 33507:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 33508:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 33509:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 33510:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 33511:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 33512:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 33513:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 33514:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 33515:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 33516:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 33517:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 33518:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 33519:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 33520:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 33521:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 33522:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 33523:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 33524:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 33525:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 33526:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 33527:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 33528:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 33529:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 33530:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 33531:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 33532:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 33533:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 33534:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 33535:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 33536:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 33537:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 33538:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 33539:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 33540:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 33541:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 33542:20]
  assign io_z = ~x59; // @[Snxn100k.scala 33543:16]
endmodule
module SnxnLv4Inst75(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 33554:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 33555:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 33556:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 33557:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 33558:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 33559:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 33560:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 33561:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 33562:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 33563:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 33564:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 33565:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 33566:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 33567:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 33568:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 33569:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 33570:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 33571:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 33572:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 33573:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 33574:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 33575:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 33576:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 33577:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 33578:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 33579:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 33580:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 33581:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 33582:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 33583:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 33584:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 33585:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 33586:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 33587:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 33588:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 33589:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 33590:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 33591:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 33592:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 33593:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 33594:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 33595:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 33596:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 33597:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 33598:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 33599:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 33600:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 33601:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 33602:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 33603:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 33604:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 33605:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 33606:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 33607:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 33608:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 33609:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 33610:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 33611:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 33612:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 33613:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 33614:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 33615:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 33616:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 33617:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 33618:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 33619:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 33620:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 33621:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 33622:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 33623:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 33624:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 33625:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 33626:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 33627:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 33628:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 33629:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 33630:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 33631:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 33632:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 33633:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 33634:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 33635:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 33636:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 33637:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 33638:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 33639:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 33640:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 33641:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 33642:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 33643:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 33644:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 33645:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 33646:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 33647:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 33648:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 33649:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 33650:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 33651:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 33652:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 33653:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 33654:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 33655:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 33656:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 33657:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 33658:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 33659:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 33660:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 33661:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 33662:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 33663:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 33664:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 33665:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 33666:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 33667:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 33668:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 33669:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 33670:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 33671:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 33672:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 33673:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 33674:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 33675:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 33676:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 33677:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 33678:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 33679:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 33680:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 33681:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 33682:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 33683:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 33684:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 33685:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 33686:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 33687:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 33688:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 33689:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 33690:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 33691:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 33692:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 33693:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 33694:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 33695:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 33696:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 33697:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 33698:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 33699:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 33700:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 33701:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 33702:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 33703:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 33704:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 33705:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 33706:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 33707:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 33708:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 33709:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 33710:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 33711:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 33712:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 33713:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 33714:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 33715:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 33716:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 33717:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 33718:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 33719:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 33720:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 33721:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 33722:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 33723:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 33724:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 33725:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 33726:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 33727:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 33728:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 33729:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 33730:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 33731:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 33732:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 33733:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 33734:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 33735:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 33736:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 33737:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 33738:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 33739:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 33740:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 33741:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 33742:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 33743:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 33744:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 33745:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 33746:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 33747:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 33748:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 33749:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 33750:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 33751:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 33752:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 33753:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 33754:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 33755:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 33756:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 33757:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 33758:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 33759:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 33760:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 33761:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 33762:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 33763:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 33764:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 33765:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 33766:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 33767:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 33768:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 33769:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 33770:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 33771:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 33772:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 33773:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 33774:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 33775:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 33776:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 33777:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 33778:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 33779:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 33780:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 33781:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 33782:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 33783:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 33784:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 33785:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 33786:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 33787:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 33788:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 33789:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 33790:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 33791:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 33792:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 33793:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 33794:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 33795:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 33796:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 33797:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 33798:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 33799:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 33800:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 33801:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 33802:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 33803:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 33804:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 33805:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 33806:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 33807:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 33808:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 33809:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 33810:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 33811:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 33812:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 33813:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 33814:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 33815:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 33816:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 33817:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 33818:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 33819:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 33820:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 33821:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 33822:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 33823:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 33824:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 33825:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 33826:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 33827:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 33828:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 33829:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 33830:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 33831:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 33832:20]
  assign io_z = ~x69; // @[Snxn100k.scala 33833:16]
endmodule
module SnxnLv3Inst18(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst72_io_a; // @[Snxn100k.scala 9279:34]
  wire  inst_SnxnLv4Inst72_io_b; // @[Snxn100k.scala 9279:34]
  wire  inst_SnxnLv4Inst72_io_z; // @[Snxn100k.scala 9279:34]
  wire  inst_SnxnLv4Inst73_io_a; // @[Snxn100k.scala 9283:34]
  wire  inst_SnxnLv4Inst73_io_b; // @[Snxn100k.scala 9283:34]
  wire  inst_SnxnLv4Inst73_io_z; // @[Snxn100k.scala 9283:34]
  wire  inst_SnxnLv4Inst74_io_a; // @[Snxn100k.scala 9287:34]
  wire  inst_SnxnLv4Inst74_io_b; // @[Snxn100k.scala 9287:34]
  wire  inst_SnxnLv4Inst74_io_z; // @[Snxn100k.scala 9287:34]
  wire  inst_SnxnLv4Inst75_io_a; // @[Snxn100k.scala 9291:34]
  wire  inst_SnxnLv4Inst75_io_b; // @[Snxn100k.scala 9291:34]
  wire  inst_SnxnLv4Inst75_io_z; // @[Snxn100k.scala 9291:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst72_io_z + inst_SnxnLv4Inst73_io_z; // @[Snxn100k.scala 9295:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst74_io_z; // @[Snxn100k.scala 9295:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst75_io_z; // @[Snxn100k.scala 9295:89]
  SnxnLv4Inst19 inst_SnxnLv4Inst72 ( // @[Snxn100k.scala 9279:34]
    .io_a(inst_SnxnLv4Inst72_io_a),
    .io_b(inst_SnxnLv4Inst72_io_b),
    .io_z(inst_SnxnLv4Inst72_io_z)
  );
  SnxnLv4Inst73 inst_SnxnLv4Inst73 ( // @[Snxn100k.scala 9283:34]
    .io_a(inst_SnxnLv4Inst73_io_a),
    .io_b(inst_SnxnLv4Inst73_io_b),
    .io_z(inst_SnxnLv4Inst73_io_z)
  );
  SnxnLv4Inst74 inst_SnxnLv4Inst74 ( // @[Snxn100k.scala 9287:34]
    .io_a(inst_SnxnLv4Inst74_io_a),
    .io_b(inst_SnxnLv4Inst74_io_b),
    .io_z(inst_SnxnLv4Inst74_io_z)
  );
  SnxnLv4Inst75 inst_SnxnLv4Inst75 ( // @[Snxn100k.scala 9291:34]
    .io_a(inst_SnxnLv4Inst75_io_a),
    .io_b(inst_SnxnLv4Inst75_io_b),
    .io_z(inst_SnxnLv4Inst75_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 9296:15]
  assign inst_SnxnLv4Inst72_io_a = io_a; // @[Snxn100k.scala 9280:27]
  assign inst_SnxnLv4Inst72_io_b = io_b; // @[Snxn100k.scala 9281:27]
  assign inst_SnxnLv4Inst73_io_a = io_a; // @[Snxn100k.scala 9284:27]
  assign inst_SnxnLv4Inst73_io_b = io_b; // @[Snxn100k.scala 9285:27]
  assign inst_SnxnLv4Inst74_io_a = io_a; // @[Snxn100k.scala 9288:27]
  assign inst_SnxnLv4Inst74_io_b = io_b; // @[Snxn100k.scala 9289:27]
  assign inst_SnxnLv4Inst75_io_a = io_a; // @[Snxn100k.scala 9292:27]
  assign inst_SnxnLv4Inst75_io_b = io_b; // @[Snxn100k.scala 9293:27]
endmodule
module SnxnLv4Inst77(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 36102:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 36103:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 36104:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 36105:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 36106:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 36107:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 36108:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 36109:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 36110:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 36111:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 36112:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 36113:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 36114:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 36115:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 36116:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 36117:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 36118:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 36119:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 36120:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 36121:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 36122:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 36123:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 36124:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 36125:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 36126:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 36127:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 36128:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 36129:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 36130:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 36131:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 36132:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 36133:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 36134:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 36135:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 36136:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 36137:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 36138:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 36139:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 36140:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 36141:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 36142:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 36143:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 36144:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 36145:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 36146:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 36147:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 36148:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 36149:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 36150:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 36151:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 36152:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 36153:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 36154:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 36155:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 36156:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 36157:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 36158:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 36159:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 36160:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 36161:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 36162:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 36163:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 36164:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 36165:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 36166:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 36167:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 36168:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 36169:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 36170:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 36171:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 36172:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 36173:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 36174:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 36175:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 36176:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 36177:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 36178:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 36179:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 36180:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 36181:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 36182:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 36183:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 36184:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 36185:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 36186:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 36187:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 36188:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 36189:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 36190:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 36191:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 36192:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 36193:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 36194:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 36195:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 36196:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 36197:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 36198:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 36199:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 36200:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 36201:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 36202:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 36203:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 36204:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 36205:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 36206:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 36207:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 36208:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 36209:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 36210:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 36211:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 36212:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 36213:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 36214:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 36215:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 36216:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 36217:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 36218:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 36219:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 36220:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 36221:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 36222:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 36223:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 36224:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 36225:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 36226:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 36227:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 36228:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 36229:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 36230:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 36231:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 36232:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 36233:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 36234:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 36235:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 36236:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 36237:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 36238:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 36239:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 36240:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 36241:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 36242:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 36243:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 36244:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 36245:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 36246:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 36247:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 36248:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 36249:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 36250:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 36251:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 36252:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 36253:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 36254:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 36255:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 36256:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 36257:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 36258:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 36259:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 36260:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 36261:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 36262:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 36263:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 36264:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 36265:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 36266:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 36267:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 36268:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 36269:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 36270:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 36271:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 36272:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 36273:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 36274:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 36275:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 36276:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 36277:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 36278:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 36279:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 36280:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 36281:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 36282:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 36283:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 36284:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 36285:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 36286:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 36287:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 36288:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 36289:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 36290:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 36291:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 36292:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 36293:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 36294:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 36295:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 36296:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 36297:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 36298:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 36299:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 36300:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 36301:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 36302:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 36303:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 36304:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 36305:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 36306:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 36307:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 36308:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 36309:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 36310:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 36311:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 36312:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 36313:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 36314:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 36315:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 36316:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 36317:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 36318:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 36319:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 36320:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 36321:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 36322:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 36323:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 36324:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 36325:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 36326:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 36327:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 36328:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 36329:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 36330:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 36331:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 36332:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 36333:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 36334:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 36335:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 36336:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 36337:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 36338:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 36339:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 36340:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 36341:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 36342:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 36343:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 36344:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 36345:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 36346:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 36347:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 36348:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 36349:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 36350:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 36351:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 36352:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 36353:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 36354:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 36355:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 36356:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 36357:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 36358:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 36359:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 36360:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 36361:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 36362:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 36363:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 36364:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 36365:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 36366:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 36367:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 36368:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 36369:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 36370:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 36371:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 36372:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 36373:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 36374:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 36375:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 36376:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 36377:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 36378:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 36379:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 36380:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 36381:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 36382:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 36383:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 36384:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 36385:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 36386:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 36387:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 36388:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 36389:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 36390:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 36391:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 36392:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 36393:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 36394:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 36395:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 36396:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 36397:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 36398:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 36399:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 36400:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 36401:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 36402:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 36403:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 36404:20]
  assign io_z = ~x75; // @[Snxn100k.scala 36405:16]
endmodule
module SnxnLv4Inst78(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 36416:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 36417:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 36418:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 36419:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 36420:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 36421:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 36422:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 36423:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 36424:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 36425:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 36426:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 36427:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 36428:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 36429:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 36430:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 36431:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 36432:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 36433:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 36434:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 36435:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 36436:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 36437:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 36438:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 36439:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 36440:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 36441:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 36442:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 36443:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 36444:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 36445:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 36446:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 36447:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 36448:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 36449:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 36450:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 36451:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 36452:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 36453:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 36454:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 36455:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 36456:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 36457:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 36458:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 36459:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 36460:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 36461:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 36462:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 36463:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 36464:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 36465:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 36466:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 36467:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 36468:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 36469:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 36470:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 36471:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 36472:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 36473:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 36474:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 36475:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 36476:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 36477:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 36478:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 36479:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 36480:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 36481:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 36482:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 36483:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 36484:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 36485:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 36486:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 36487:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 36488:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 36489:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 36490:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 36491:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 36492:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 36493:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 36494:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 36495:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 36496:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 36497:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 36498:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 36499:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 36500:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 36501:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 36502:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 36503:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 36504:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 36505:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 36506:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 36507:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 36508:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 36509:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 36510:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 36511:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 36512:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 36513:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 36514:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 36515:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 36516:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 36517:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 36518:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 36519:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 36520:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 36521:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 36522:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 36523:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 36524:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 36525:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 36526:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 36527:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 36528:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 36529:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 36530:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 36531:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 36532:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 36533:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 36534:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 36535:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 36536:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 36537:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 36538:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 36539:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 36540:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 36541:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 36542:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 36543:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 36544:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 36545:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 36546:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 36547:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 36548:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 36549:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 36550:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 36551:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 36552:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 36553:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 36554:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 36555:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 36556:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 36557:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 36558:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 36559:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 36560:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 36561:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 36562:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 36563:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 36564:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 36565:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 36566:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 36567:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 36568:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 36569:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 36570:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 36571:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 36572:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 36573:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 36574:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 36575:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 36576:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 36577:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 36578:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 36579:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 36580:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 36581:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 36582:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 36583:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 36584:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 36585:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 36586:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 36587:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 36588:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 36589:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 36590:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 36591:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 36592:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 36593:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 36594:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 36595:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 36596:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 36597:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 36598:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 36599:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 36600:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 36601:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 36602:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 36603:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 36604:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 36605:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 36606:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 36607:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 36608:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 36609:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 36610:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 36611:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 36612:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 36613:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 36614:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 36615:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 36616:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 36617:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 36618:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 36619:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 36620:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 36621:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 36622:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 36623:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 36624:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 36625:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 36626:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 36627:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 36628:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 36629:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 36630:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 36631:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 36632:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 36633:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 36634:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 36635:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 36636:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 36637:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 36638:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 36639:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 36640:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 36641:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 36642:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 36643:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 36644:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 36645:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 36646:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 36647:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 36648:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 36649:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 36650:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 36651:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 36652:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 36653:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 36654:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 36655:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 36656:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 36657:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 36658:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 36659:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 36660:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 36661:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 36662:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 36663:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 36664:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 36665:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 36666:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 36667:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 36668:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 36669:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 36670:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 36671:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 36672:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 36673:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 36674:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 36675:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 36676:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 36677:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 36678:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 36679:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 36680:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 36681:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 36682:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 36683:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 36684:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 36685:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 36686:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 36687:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 36688:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 36689:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 36690:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 36691:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 36692:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 36693:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 36694:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 36695:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 36696:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 36697:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 36698:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 36699:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 36700:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 36701:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 36702:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 36703:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 36704:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 36705:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 36706:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 36707:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 36708:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 36709:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 36710:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 36711:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 36712:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 36713:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 36714:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 36715:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 36716:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 36717:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 36718:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 36719:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 36720:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 36721:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 36722:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 36723:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 36724:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 36725:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 36726:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 36727:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 36728:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 36729:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 36730:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 36731:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 36732:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 36733:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 36734:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 36735:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 36736:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 36737:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 36738:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 36739:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 36740:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 36741:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 36742:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 36743:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 36744:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 36745:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 36746:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 36747:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 36748:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 36749:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 36750:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 36751:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 36752:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 36753:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 36754:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 36755:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 36756:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 36757:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 36758:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 36759:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 36760:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 36761:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 36762:20]
  assign io_z = ~x86; // @[Snxn100k.scala 36763:16]
endmodule
module SnxnLv3Inst19(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst76_io_a; // @[Snxn100k.scala 10117:34]
  wire  inst_SnxnLv4Inst76_io_b; // @[Snxn100k.scala 10117:34]
  wire  inst_SnxnLv4Inst76_io_z; // @[Snxn100k.scala 10117:34]
  wire  inst_SnxnLv4Inst77_io_a; // @[Snxn100k.scala 10121:34]
  wire  inst_SnxnLv4Inst77_io_b; // @[Snxn100k.scala 10121:34]
  wire  inst_SnxnLv4Inst77_io_z; // @[Snxn100k.scala 10121:34]
  wire  inst_SnxnLv4Inst78_io_a; // @[Snxn100k.scala 10125:34]
  wire  inst_SnxnLv4Inst78_io_b; // @[Snxn100k.scala 10125:34]
  wire  inst_SnxnLv4Inst78_io_z; // @[Snxn100k.scala 10125:34]
  wire  inst_SnxnLv4Inst79_io_a; // @[Snxn100k.scala 10129:34]
  wire  inst_SnxnLv4Inst79_io_b; // @[Snxn100k.scala 10129:34]
  wire  inst_SnxnLv4Inst79_io_z; // @[Snxn100k.scala 10129:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst76_io_z + inst_SnxnLv4Inst77_io_z; // @[Snxn100k.scala 10133:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst78_io_z; // @[Snxn100k.scala 10133:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst79_io_z; // @[Snxn100k.scala 10133:89]
  SnxnLv4Inst9 inst_SnxnLv4Inst76 ( // @[Snxn100k.scala 10117:34]
    .io_a(inst_SnxnLv4Inst76_io_a),
    .io_b(inst_SnxnLv4Inst76_io_b),
    .io_z(inst_SnxnLv4Inst76_io_z)
  );
  SnxnLv4Inst77 inst_SnxnLv4Inst77 ( // @[Snxn100k.scala 10121:34]
    .io_a(inst_SnxnLv4Inst77_io_a),
    .io_b(inst_SnxnLv4Inst77_io_b),
    .io_z(inst_SnxnLv4Inst77_io_z)
  );
  SnxnLv4Inst78 inst_SnxnLv4Inst78 ( // @[Snxn100k.scala 10125:34]
    .io_a(inst_SnxnLv4Inst78_io_a),
    .io_b(inst_SnxnLv4Inst78_io_b),
    .io_z(inst_SnxnLv4Inst78_io_z)
  );
  SnxnLv4Inst43 inst_SnxnLv4Inst79 ( // @[Snxn100k.scala 10129:34]
    .io_a(inst_SnxnLv4Inst79_io_a),
    .io_b(inst_SnxnLv4Inst79_io_b),
    .io_z(inst_SnxnLv4Inst79_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10134:15]
  assign inst_SnxnLv4Inst76_io_a = io_a; // @[Snxn100k.scala 10118:27]
  assign inst_SnxnLv4Inst76_io_b = io_b; // @[Snxn100k.scala 10119:27]
  assign inst_SnxnLv4Inst77_io_a = io_a; // @[Snxn100k.scala 10122:27]
  assign inst_SnxnLv4Inst77_io_b = io_b; // @[Snxn100k.scala 10123:27]
  assign inst_SnxnLv4Inst78_io_a = io_a; // @[Snxn100k.scala 10126:27]
  assign inst_SnxnLv4Inst78_io_b = io_b; // @[Snxn100k.scala 10127:27]
  assign inst_SnxnLv4Inst79_io_a = io_a; // @[Snxn100k.scala 10130:27]
  assign inst_SnxnLv4Inst79_io_b = io_b; // @[Snxn100k.scala 10131:27]
endmodule
module SnxnLv2Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst16_io_a; // @[Snxn100k.scala 1815:34]
  wire  inst_SnxnLv3Inst16_io_b; // @[Snxn100k.scala 1815:34]
  wire  inst_SnxnLv3Inst16_io_z; // @[Snxn100k.scala 1815:34]
  wire  inst_SnxnLv3Inst17_io_a; // @[Snxn100k.scala 1819:34]
  wire  inst_SnxnLv3Inst17_io_b; // @[Snxn100k.scala 1819:34]
  wire  inst_SnxnLv3Inst17_io_z; // @[Snxn100k.scala 1819:34]
  wire  inst_SnxnLv3Inst18_io_a; // @[Snxn100k.scala 1823:34]
  wire  inst_SnxnLv3Inst18_io_b; // @[Snxn100k.scala 1823:34]
  wire  inst_SnxnLv3Inst18_io_z; // @[Snxn100k.scala 1823:34]
  wire  inst_SnxnLv3Inst19_io_a; // @[Snxn100k.scala 1827:34]
  wire  inst_SnxnLv3Inst19_io_b; // @[Snxn100k.scala 1827:34]
  wire  inst_SnxnLv3Inst19_io_z; // @[Snxn100k.scala 1827:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst16_io_z + inst_SnxnLv3Inst17_io_z; // @[Snxn100k.scala 1831:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst18_io_z; // @[Snxn100k.scala 1831:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst19_io_z; // @[Snxn100k.scala 1831:89]
  SnxnLv3Inst16 inst_SnxnLv3Inst16 ( // @[Snxn100k.scala 1815:34]
    .io_a(inst_SnxnLv3Inst16_io_a),
    .io_b(inst_SnxnLv3Inst16_io_b),
    .io_z(inst_SnxnLv3Inst16_io_z)
  );
  SnxnLv3Inst17 inst_SnxnLv3Inst17 ( // @[Snxn100k.scala 1819:34]
    .io_a(inst_SnxnLv3Inst17_io_a),
    .io_b(inst_SnxnLv3Inst17_io_b),
    .io_z(inst_SnxnLv3Inst17_io_z)
  );
  SnxnLv3Inst18 inst_SnxnLv3Inst18 ( // @[Snxn100k.scala 1823:34]
    .io_a(inst_SnxnLv3Inst18_io_a),
    .io_b(inst_SnxnLv3Inst18_io_b),
    .io_z(inst_SnxnLv3Inst18_io_z)
  );
  SnxnLv3Inst19 inst_SnxnLv3Inst19 ( // @[Snxn100k.scala 1827:34]
    .io_a(inst_SnxnLv3Inst19_io_a),
    .io_b(inst_SnxnLv3Inst19_io_b),
    .io_z(inst_SnxnLv3Inst19_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1832:15]
  assign inst_SnxnLv3Inst16_io_a = io_a; // @[Snxn100k.scala 1816:27]
  assign inst_SnxnLv3Inst16_io_b = io_b; // @[Snxn100k.scala 1817:27]
  assign inst_SnxnLv3Inst17_io_a = io_a; // @[Snxn100k.scala 1820:27]
  assign inst_SnxnLv3Inst17_io_b = io_b; // @[Snxn100k.scala 1821:27]
  assign inst_SnxnLv3Inst18_io_a = io_a; // @[Snxn100k.scala 1824:27]
  assign inst_SnxnLv3Inst18_io_b = io_b; // @[Snxn100k.scala 1825:27]
  assign inst_SnxnLv3Inst19_io_a = io_a; // @[Snxn100k.scala 1828:27]
  assign inst_SnxnLv3Inst19_io_b = io_b; // @[Snxn100k.scala 1829:27]
endmodule
module SnxnLv4Inst80(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 40008:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 40009:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 40010:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 40011:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 40012:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 40013:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 40014:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 40015:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 40016:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 40017:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 40018:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 40019:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 40020:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 40021:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 40022:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 40023:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 40024:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 40025:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 40026:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 40027:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 40028:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 40029:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 40030:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 40031:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 40032:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 40033:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 40034:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 40035:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 40036:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 40037:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 40038:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 40039:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 40040:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 40041:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 40042:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 40043:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 40044:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 40045:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 40046:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 40047:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 40048:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 40049:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 40050:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 40051:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 40052:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 40053:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 40054:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 40055:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 40056:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 40057:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 40058:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 40059:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 40060:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 40061:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 40062:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 40063:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 40064:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 40065:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 40066:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 40067:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 40068:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 40069:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 40070:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 40071:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 40072:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 40073:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 40074:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 40075:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 40076:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 40077:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 40078:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 40079:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 40080:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 40081:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 40082:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 40083:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 40084:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 40085:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 40086:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 40087:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 40088:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 40089:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 40090:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 40091:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 40092:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 40093:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 40094:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 40095:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 40096:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 40097:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 40098:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 40099:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 40100:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 40101:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 40102:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 40103:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 40104:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 40105:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 40106:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 40107:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 40108:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 40109:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 40110:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 40111:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 40112:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 40113:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 40114:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 40115:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 40116:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 40117:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 40118:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 40119:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 40120:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 40121:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 40122:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 40123:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 40124:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 40125:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 40126:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 40127:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 40128:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 40129:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 40130:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 40131:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 40132:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 40133:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 40134:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 40135:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 40136:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 40137:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 40138:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 40139:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 40140:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 40141:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 40142:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 40143:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 40144:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 40145:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 40146:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 40147:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 40148:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 40149:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 40150:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 40151:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 40152:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 40153:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 40154:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 40155:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 40156:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 40157:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 40158:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 40159:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 40160:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 40161:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 40162:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 40163:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 40164:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 40165:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 40166:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 40167:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 40168:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 40169:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 40170:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 40171:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 40172:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 40173:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 40174:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 40175:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 40176:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 40177:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 40178:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 40179:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 40180:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 40181:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 40182:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 40183:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 40184:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 40185:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 40186:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 40187:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 40188:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 40189:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 40190:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 40191:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 40192:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 40193:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 40194:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 40195:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 40196:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 40197:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 40198:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 40199:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 40200:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 40201:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 40202:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 40203:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 40204:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 40205:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 40206:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 40207:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 40208:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 40209:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 40210:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 40211:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 40212:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 40213:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 40214:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 40215:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 40216:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 40217:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 40218:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 40219:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 40220:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 40221:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 40222:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 40223:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 40224:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 40225:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 40226:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 40227:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 40228:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 40229:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 40230:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 40231:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 40232:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 40233:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 40234:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 40235:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 40236:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 40237:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 40238:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 40239:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 40240:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 40241:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 40242:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 40243:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 40244:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 40245:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 40246:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 40247:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 40248:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 40249:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 40250:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 40251:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 40252:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 40253:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 40254:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 40255:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 40256:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 40257:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 40258:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 40259:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 40260:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 40261:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 40262:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 40263:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 40264:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 40265:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 40266:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 40267:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 40268:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 40269:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 40270:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 40271:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 40272:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 40273:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 40274:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 40275:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 40276:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 40277:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 40278:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 40279:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 40280:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 40281:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 40282:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 40283:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 40284:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 40285:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 40286:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 40287:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 40288:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 40289:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 40290:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 40291:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 40292:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 40293:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 40294:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 40295:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 40296:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 40297:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 40298:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 40299:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 40300:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 40301:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 40302:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 40303:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 40304:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 40305:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 40306:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 40307:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 40308:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 40309:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 40310:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 40311:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 40312:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 40313:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 40314:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 40315:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 40316:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 40317:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 40318:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 40319:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 40320:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 40321:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 40322:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 40323:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 40324:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 40325:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 40326:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 40327:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 40328:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 40329:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 40330:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 40331:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 40332:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 40333:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 40334:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 40335:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 40336:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 40337:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 40338:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 40339:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 40340:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 40341:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 40342:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 40343:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 40344:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 40345:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 40346:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 40347:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 40348:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 40349:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 40350:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 40351:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 40352:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 40353:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 40354:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 40355:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 40356:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 40357:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 40358:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 40359:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 40360:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 40361:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 40362:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 40363:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 40364:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 40365:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 40366:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 40367:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 40368:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 40369:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 40370:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 40371:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 40372:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 40373:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 40374:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 40375:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 40376:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 40377:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 40378:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 40379:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 40380:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 40381:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 40382:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 40383:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 40384:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 40385:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 40386:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 40387:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 40388:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 40389:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 40390:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 40391:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 40392:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 40393:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 40394:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 40395:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 40396:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 40397:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 40398:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 40399:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 40400:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 40401:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 40402:20]
  assign io_z = ~x98; // @[Snxn100k.scala 40403:16]
endmodule
module SnxnLv4Inst81(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 39476:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 39477:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 39478:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 39479:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 39480:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 39481:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 39482:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 39483:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 39484:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 39485:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 39486:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 39487:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 39488:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 39489:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 39490:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 39491:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 39492:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 39493:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 39494:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 39495:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 39496:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 39497:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 39498:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 39499:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 39500:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 39501:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 39502:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 39503:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 39504:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 39505:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 39506:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 39507:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 39508:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 39509:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 39510:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 39511:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 39512:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 39513:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 39514:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 39515:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 39516:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 39517:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 39518:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 39519:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 39520:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 39521:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 39522:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 39523:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 39524:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 39525:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 39526:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 39527:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 39528:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 39529:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 39530:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 39531:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 39532:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 39533:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 39534:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 39535:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 39536:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 39537:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 39538:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 39539:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 39540:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 39541:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 39542:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 39543:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 39544:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 39545:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 39546:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 39547:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 39548:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 39549:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 39550:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 39551:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 39552:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 39553:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 39554:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 39555:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 39556:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 39557:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 39558:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 39559:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 39560:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 39561:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 39562:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 39563:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 39564:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 39565:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 39566:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 39567:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 39568:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 39569:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 39570:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 39571:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 39572:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 39573:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 39574:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 39575:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 39576:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 39577:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 39578:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 39579:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 39580:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 39581:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 39582:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 39583:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 39584:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 39585:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 39586:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 39587:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 39588:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 39589:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 39590:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 39591:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 39592:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 39593:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 39594:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 39595:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 39596:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 39597:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 39598:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 39599:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 39600:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 39601:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 39602:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 39603:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 39604:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 39605:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 39606:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 39607:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 39608:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 39609:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 39610:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 39611:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 39612:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 39613:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 39614:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 39615:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 39616:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 39617:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 39618:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 39619:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 39620:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 39621:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 39622:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 39623:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 39624:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 39625:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 39626:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 39627:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 39628:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 39629:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 39630:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 39631:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 39632:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 39633:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 39634:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 39635:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 39636:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 39637:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 39638:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 39639:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 39640:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 39641:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 39642:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 39643:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 39644:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 39645:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 39646:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 39647:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 39648:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 39649:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 39650:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 39651:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 39652:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 39653:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 39654:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 39655:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 39656:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 39657:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 39658:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 39659:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 39660:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 39661:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 39662:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 39663:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 39664:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 39665:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 39666:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 39667:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 39668:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 39669:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 39670:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 39671:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 39672:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 39673:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 39674:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 39675:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 39676:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 39677:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 39678:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 39679:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 39680:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 39681:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 39682:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 39683:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 39684:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 39685:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 39686:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 39687:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 39688:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 39689:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 39690:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 39691:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 39692:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 39693:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 39694:20]
  assign io_z = ~x54; // @[Snxn100k.scala 39695:16]
endmodule
module SnxnLv4Inst82(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 40414:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 40415:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 40416:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 40417:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 40418:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 40419:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 40420:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 40421:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 40422:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 40423:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 40424:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 40425:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 40426:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 40427:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 40428:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 40429:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 40430:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 40431:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 40432:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 40433:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 40434:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 40435:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 40436:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 40437:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 40438:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 40439:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 40440:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 40441:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 40442:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 40443:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 40444:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 40445:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 40446:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 40447:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 40448:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 40449:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 40450:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 40451:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 40452:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 40453:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 40454:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 40455:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 40456:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 40457:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 40458:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 40459:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 40460:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 40461:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 40462:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 40463:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 40464:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 40465:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 40466:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 40467:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 40468:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 40469:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 40470:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 40471:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 40472:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 40473:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 40474:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 40475:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 40476:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 40477:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 40478:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 40479:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 40480:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 40481:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 40482:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 40483:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 40484:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 40485:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 40486:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 40487:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 40488:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 40489:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 40490:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 40491:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 40492:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 40493:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 40494:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 40495:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 40496:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 40497:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 40498:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 40499:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 40500:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 40501:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 40502:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 40503:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 40504:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 40505:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 40506:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 40507:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 40508:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 40509:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 40510:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 40511:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 40512:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 40513:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 40514:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 40515:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 40516:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 40517:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 40518:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 40519:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 40520:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 40521:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 40522:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 40523:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 40524:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 40525:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 40526:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 40527:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 40528:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 40529:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 40530:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 40531:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 40532:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 40533:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 40534:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 40535:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 40536:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 40537:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 40538:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 40539:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 40540:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 40541:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 40542:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 40543:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 40544:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 40545:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 40546:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 40547:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 40548:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 40549:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 40550:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 40551:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 40552:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 40553:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 40554:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 40555:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 40556:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 40557:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 40558:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 40559:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 40560:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 40561:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 40562:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 40563:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 40564:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 40565:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 40566:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 40567:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 40568:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 40569:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 40570:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 40571:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 40572:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 40573:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 40574:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 40575:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 40576:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 40577:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 40578:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 40579:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 40580:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 40581:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 40582:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 40583:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 40584:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 40585:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 40586:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 40587:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 40588:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 40589:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 40590:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 40591:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 40592:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 40593:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 40594:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 40595:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 40596:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 40597:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 40598:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 40599:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 40600:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 40601:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 40602:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 40603:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 40604:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 40605:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 40606:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 40607:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 40608:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 40609:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 40610:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 40611:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 40612:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 40613:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 40614:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 40615:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 40616:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 40617:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 40618:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 40619:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 40620:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 40621:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 40622:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 40623:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 40624:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 40625:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 40626:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 40627:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 40628:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 40629:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 40630:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 40631:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 40632:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 40633:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 40634:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 40635:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 40636:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 40637:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 40638:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 40639:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 40640:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 40641:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 40642:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 40643:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 40644:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 40645:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 40646:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 40647:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 40648:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 40649:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 40650:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 40651:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 40652:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 40653:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 40654:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 40655:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 40656:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 40657:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 40658:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 40659:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 40660:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 40661:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 40662:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 40663:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 40664:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 40665:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 40666:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 40667:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 40668:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 40669:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 40670:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 40671:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 40672:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 40673:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 40674:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 40675:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 40676:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 40677:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 40678:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 40679:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 40680:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 40681:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 40682:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 40683:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 40684:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 40685:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 40686:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 40687:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 40688:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 40689:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 40690:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 40691:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 40692:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 40693:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 40694:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 40695:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 40696:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 40697:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 40698:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 40699:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 40700:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 40701:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 40702:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 40703:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 40704:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 40705:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 40706:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 40707:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 40708:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 40709:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 40710:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 40711:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 40712:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 40713:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 40714:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 40715:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 40716:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 40717:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 40718:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 40719:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 40720:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 40721:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 40722:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 40723:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 40724:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 40725:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 40726:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 40727:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 40728:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 40729:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 40730:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 40731:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 40732:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 40733:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 40734:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 40735:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 40736:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 40737:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 40738:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 40739:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 40740:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 40741:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 40742:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 40743:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 40744:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 40745:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 40746:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 40747:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 40748:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 40749:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 40750:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 40751:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 40752:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 40753:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 40754:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 40755:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 40756:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 40757:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 40758:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 40759:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 40760:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 40761:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 40762:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 40763:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 40764:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 40765:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 40766:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 40767:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 40768:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 40769:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 40770:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 40771:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 40772:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 40773:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 40774:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 40775:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 40776:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 40777:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 40778:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 40779:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 40780:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 40781:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 40782:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 40783:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 40784:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 40785:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 40786:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 40787:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 40788:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 40789:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 40790:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 40791:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 40792:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 40793:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 40794:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 40795:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 40796:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 40797:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 40798:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 40799:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 40800:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 40801:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 40802:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 40803:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 40804:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 40805:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 40806:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 40807:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 40808:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 40809:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 40810:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 40811:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 40812:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 40813:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 40814:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 40815:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 40816:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 40817:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 40818:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 40819:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 40820:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 40821:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 40822:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 40823:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 40824:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 40825:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 40826:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 40827:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 40828:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 40829:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 40830:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 40831:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 40832:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 40833:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 40834:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 40835:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 40836:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 40837:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 40838:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 40839:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 40840:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 40841:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 40842:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 40843:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 40844:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 40845:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 40846:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 40847:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 40848:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 40849:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 40850:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 40851:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 40852:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 40853:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 40854:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 40855:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 40856:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 40857:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 40858:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 40859:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 40860:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 40861:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 40862:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 40863:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 40864:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 40865:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 40866:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 40867:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 40868:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 40869:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 40870:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 40871:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 40872:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 40873:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 40874:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 40875:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 40876:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 40877:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 40878:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 40879:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 40880:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 40881:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 40882:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 40883:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 40884:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 40885:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 40886:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 40887:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 40888:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 40889:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 40890:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 40891:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 40892:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 40893:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 40894:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 40895:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 40896:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 40897:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 40898:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 40899:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 40900:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 40901:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 40902:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 40903:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 40904:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 40905:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 40906:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 40907:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 40908:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 40909:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 40910:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 40911:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 40912:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 40913:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 40914:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 40915:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 40916:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 40917:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 40918:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 40919:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 40920:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 40921:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 40922:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 40923:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 40924:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 40925:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 40926:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 40927:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 40928:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 40929:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 40930:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 40931:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 40932:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 40933:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 40934:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 40935:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 40936:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 40937:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 40938:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 40939:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 40940:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 40941:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 40942:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 40943:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 40944:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 40945:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 40946:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 40947:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 40948:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 40949:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 40950:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 40951:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 40952:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 40953:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 40954:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 40955:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 40956:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 40957:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 40958:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 40959:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 40960:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 40961:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 40962:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 40963:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 40964:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 40965:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 40966:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 40967:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 40968:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 40969:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 40970:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 40971:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 40972:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 40973:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 40974:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 40975:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 40976:22]
  assign io_z = ~x140; // @[Snxn100k.scala 40977:17]
endmodule
module SnxnLv4Inst83(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 39706:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 39707:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 39708:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 39709:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 39710:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 39711:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 39712:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 39713:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 39714:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 39715:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 39716:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 39717:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 39718:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 39719:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 39720:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 39721:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 39722:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 39723:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 39724:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 39725:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 39726:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 39727:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 39728:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 39729:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 39730:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 39731:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 39732:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 39733:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 39734:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 39735:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 39736:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 39737:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 39738:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 39739:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 39740:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 39741:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 39742:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 39743:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 39744:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 39745:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 39746:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 39747:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 39748:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 39749:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 39750:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 39751:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 39752:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 39753:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 39754:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 39755:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 39756:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 39757:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 39758:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 39759:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 39760:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 39761:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 39762:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 39763:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 39764:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 39765:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 39766:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 39767:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 39768:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 39769:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 39770:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 39771:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 39772:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 39773:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 39774:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 39775:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 39776:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 39777:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 39778:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 39779:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 39780:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 39781:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 39782:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 39783:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 39784:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 39785:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 39786:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 39787:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 39788:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 39789:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 39790:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 39791:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 39792:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 39793:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 39794:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 39795:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 39796:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 39797:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 39798:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 39799:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 39800:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 39801:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 39802:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 39803:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 39804:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 39805:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 39806:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 39807:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 39808:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 39809:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 39810:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 39811:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 39812:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 39813:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 39814:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 39815:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 39816:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 39817:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 39818:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 39819:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 39820:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 39821:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 39822:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 39823:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 39824:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 39825:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 39826:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 39827:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 39828:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 39829:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 39830:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 39831:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 39832:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 39833:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 39834:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 39835:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 39836:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 39837:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 39838:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 39839:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 39840:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 39841:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 39842:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 39843:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 39844:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 39845:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 39846:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 39847:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 39848:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 39849:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 39850:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 39851:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 39852:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 39853:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 39854:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 39855:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 39856:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 39857:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 39858:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 39859:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 39860:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 39861:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 39862:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 39863:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 39864:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 39865:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 39866:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 39867:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 39868:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 39869:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 39870:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 39871:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 39872:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 39873:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 39874:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 39875:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 39876:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 39877:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 39878:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 39879:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 39880:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 39881:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 39882:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 39883:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 39884:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 39885:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 39886:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 39887:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 39888:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 39889:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 39890:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 39891:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 39892:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 39893:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 39894:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 39895:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 39896:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 39897:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 39898:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 39899:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 39900:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 39901:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 39902:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 39903:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 39904:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 39905:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 39906:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 39907:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 39908:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 39909:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 39910:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 39911:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 39912:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 39913:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 39914:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 39915:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 39916:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 39917:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 39918:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 39919:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 39920:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 39921:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 39922:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 39923:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 39924:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 39925:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 39926:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 39927:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 39928:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 39929:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 39930:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 39931:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 39932:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 39933:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 39934:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 39935:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 39936:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 39937:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 39938:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 39939:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 39940:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 39941:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 39942:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 39943:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 39944:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 39945:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 39946:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 39947:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 39948:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 39949:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 39950:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 39951:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 39952:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 39953:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 39954:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 39955:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 39956:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 39957:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 39958:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 39959:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 39960:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 39961:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 39962:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 39963:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 39964:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 39965:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 39966:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 39967:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 39968:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 39969:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 39970:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 39971:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 39972:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 39973:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 39974:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 39975:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 39976:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 39977:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 39978:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 39979:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 39980:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 39981:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 39982:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 39983:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 39984:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 39985:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 39986:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 39987:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 39988:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 39989:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 39990:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 39991:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 39992:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 39993:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 39994:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 39995:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 39996:20]
  assign io_z = ~x72; // @[Snxn100k.scala 39997:16]
endmodule
module SnxnLv3Inst20(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst80_io_a; // @[Snxn100k.scala 11190:34]
  wire  inst_SnxnLv4Inst80_io_b; // @[Snxn100k.scala 11190:34]
  wire  inst_SnxnLv4Inst80_io_z; // @[Snxn100k.scala 11190:34]
  wire  inst_SnxnLv4Inst81_io_a; // @[Snxn100k.scala 11194:34]
  wire  inst_SnxnLv4Inst81_io_b; // @[Snxn100k.scala 11194:34]
  wire  inst_SnxnLv4Inst81_io_z; // @[Snxn100k.scala 11194:34]
  wire  inst_SnxnLv4Inst82_io_a; // @[Snxn100k.scala 11198:34]
  wire  inst_SnxnLv4Inst82_io_b; // @[Snxn100k.scala 11198:34]
  wire  inst_SnxnLv4Inst82_io_z; // @[Snxn100k.scala 11198:34]
  wire  inst_SnxnLv4Inst83_io_a; // @[Snxn100k.scala 11202:34]
  wire  inst_SnxnLv4Inst83_io_b; // @[Snxn100k.scala 11202:34]
  wire  inst_SnxnLv4Inst83_io_z; // @[Snxn100k.scala 11202:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst80_io_z + inst_SnxnLv4Inst81_io_z; // @[Snxn100k.scala 11206:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst82_io_z; // @[Snxn100k.scala 11206:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst83_io_z; // @[Snxn100k.scala 11206:89]
  SnxnLv4Inst80 inst_SnxnLv4Inst80 ( // @[Snxn100k.scala 11190:34]
    .io_a(inst_SnxnLv4Inst80_io_a),
    .io_b(inst_SnxnLv4Inst80_io_b),
    .io_z(inst_SnxnLv4Inst80_io_z)
  );
  SnxnLv4Inst81 inst_SnxnLv4Inst81 ( // @[Snxn100k.scala 11194:34]
    .io_a(inst_SnxnLv4Inst81_io_a),
    .io_b(inst_SnxnLv4Inst81_io_b),
    .io_z(inst_SnxnLv4Inst81_io_z)
  );
  SnxnLv4Inst82 inst_SnxnLv4Inst82 ( // @[Snxn100k.scala 11198:34]
    .io_a(inst_SnxnLv4Inst82_io_a),
    .io_b(inst_SnxnLv4Inst82_io_b),
    .io_z(inst_SnxnLv4Inst82_io_z)
  );
  SnxnLv4Inst83 inst_SnxnLv4Inst83 ( // @[Snxn100k.scala 11202:34]
    .io_a(inst_SnxnLv4Inst83_io_a),
    .io_b(inst_SnxnLv4Inst83_io_b),
    .io_z(inst_SnxnLv4Inst83_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11207:15]
  assign inst_SnxnLv4Inst80_io_a = io_a; // @[Snxn100k.scala 11191:27]
  assign inst_SnxnLv4Inst80_io_b = io_b; // @[Snxn100k.scala 11192:27]
  assign inst_SnxnLv4Inst81_io_a = io_a; // @[Snxn100k.scala 11195:27]
  assign inst_SnxnLv4Inst81_io_b = io_b; // @[Snxn100k.scala 11196:27]
  assign inst_SnxnLv4Inst82_io_a = io_a; // @[Snxn100k.scala 11199:27]
  assign inst_SnxnLv4Inst82_io_b = io_b; // @[Snxn100k.scala 11200:27]
  assign inst_SnxnLv4Inst83_io_a = io_a; // @[Snxn100k.scala 11203:27]
  assign inst_SnxnLv4Inst83_io_b = io_b; // @[Snxn100k.scala 11204:27]
endmodule
module SnxnLv4Inst84(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 37160:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 37161:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 37162:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 37163:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 37164:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 37165:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 37166:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 37167:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 37168:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 37169:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 37170:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 37171:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 37172:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 37173:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 37174:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 37175:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 37176:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 37177:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 37178:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 37179:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 37180:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 37181:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 37182:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 37183:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 37184:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 37185:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 37186:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 37187:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 37188:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 37189:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 37190:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 37191:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 37192:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 37193:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 37194:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 37195:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 37196:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 37197:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 37198:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 37199:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 37200:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 37201:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 37202:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 37203:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 37204:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 37205:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 37206:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 37207:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 37208:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 37209:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 37210:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 37211:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 37212:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 37213:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 37214:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 37215:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 37216:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 37217:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 37218:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 37219:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 37220:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 37221:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 37222:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 37223:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 37224:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 37225:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 37226:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 37227:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 37228:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 37229:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 37230:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 37231:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 37232:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 37233:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 37234:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 37235:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 37236:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 37237:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 37238:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 37239:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 37240:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 37241:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 37242:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 37243:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 37244:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 37245:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 37246:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 37247:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 37248:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 37249:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 37250:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 37251:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 37252:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 37253:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 37254:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 37255:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 37256:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 37257:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 37258:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 37259:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 37260:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 37261:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 37262:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 37263:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 37264:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 37265:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 37266:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 37267:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 37268:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 37269:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 37270:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 37271:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 37272:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 37273:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 37274:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 37275:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 37276:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 37277:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 37278:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 37279:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 37280:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 37281:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 37282:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 37283:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 37284:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 37285:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 37286:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 37287:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 37288:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 37289:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 37290:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 37291:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 37292:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 37293:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 37294:20]
  assign io_z = ~x33; // @[Snxn100k.scala 37295:16]
endmodule
module SnxnLv4Inst86(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 37898:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 37899:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 37900:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 37901:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 37902:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 37903:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 37904:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 37905:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 37906:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 37907:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 37908:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 37909:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 37910:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 37911:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 37912:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 37913:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 37914:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 37915:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 37916:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 37917:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 37918:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 37919:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 37920:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 37921:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 37922:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 37923:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 37924:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 37925:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 37926:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 37927:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 37928:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 37929:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 37930:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 37931:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 37932:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 37933:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 37934:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 37935:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 37936:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 37937:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 37938:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 37939:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 37940:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 37941:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 37942:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 37943:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 37944:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 37945:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 37946:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 37947:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 37948:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 37949:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 37950:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 37951:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 37952:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 37953:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 37954:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 37955:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 37956:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 37957:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 37958:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 37959:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 37960:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 37961:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 37962:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 37963:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 37964:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 37965:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 37966:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 37967:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 37968:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 37969:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 37970:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 37971:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 37972:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 37973:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 37974:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 37975:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 37976:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 37977:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 37978:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 37979:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 37980:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 37981:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 37982:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 37983:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 37984:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 37985:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 37986:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 37987:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 37988:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 37989:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 37990:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 37991:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 37992:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 37993:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 37994:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 37995:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 37996:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 37997:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 37998:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 37999:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 38000:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 38001:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 38002:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 38003:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 38004:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 38005:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 38006:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 38007:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 38008:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 38009:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 38010:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 38011:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 38012:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 38013:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 38014:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 38015:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 38016:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 38017:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 38018:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 38019:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 38020:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 38021:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 38022:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 38023:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 38024:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 38025:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 38026:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 38027:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 38028:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 38029:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 38030:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 38031:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 38032:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 38033:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 38034:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 38035:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 38036:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 38037:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 38038:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 38039:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 38040:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 38041:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 38042:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 38043:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 38044:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 38045:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 38046:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 38047:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 38048:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 38049:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 38050:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 38051:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 38052:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 38053:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 38054:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 38055:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 38056:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 38057:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 38058:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 38059:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 38060:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 38061:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 38062:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 38063:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 38064:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 38065:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 38066:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 38067:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 38068:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 38069:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 38070:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 38071:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 38072:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 38073:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 38074:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 38075:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 38076:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 38077:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 38078:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 38079:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 38080:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 38081:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 38082:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 38083:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 38084:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 38085:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 38086:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 38087:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 38088:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 38089:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 38090:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 38091:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 38092:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 38093:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 38094:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 38095:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 38096:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 38097:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 38098:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 38099:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 38100:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 38101:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 38102:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 38103:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 38104:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 38105:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 38106:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 38107:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 38108:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 38109:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 38110:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 38111:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 38112:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 38113:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 38114:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 38115:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 38116:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 38117:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 38118:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 38119:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 38120:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 38121:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 38122:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 38123:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 38124:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 38125:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 38126:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 38127:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 38128:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 38129:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 38130:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 38131:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 38132:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 38133:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 38134:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 38135:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 38136:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 38137:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 38138:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 38139:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 38140:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 38141:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 38142:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 38143:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 38144:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 38145:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 38146:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 38147:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 38148:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 38149:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 38150:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 38151:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 38152:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 38153:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 38154:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 38155:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 38156:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 38157:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 38158:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 38159:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 38160:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 38161:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 38162:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 38163:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 38164:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 38165:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 38166:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 38167:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 38168:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 38169:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 38170:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 38171:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 38172:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 38173:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 38174:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 38175:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 38176:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 38177:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 38178:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 38179:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 38180:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 38181:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 38182:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 38183:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 38184:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 38185:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 38186:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 38187:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 38188:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 38189:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 38190:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 38191:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 38192:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 38193:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 38194:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 38195:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 38196:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 38197:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 38198:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 38199:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 38200:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 38201:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 38202:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 38203:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 38204:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 38205:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 38206:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 38207:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 38208:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 38209:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 38210:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 38211:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 38212:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 38213:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 38214:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 38215:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 38216:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 38217:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 38218:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 38219:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 38220:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 38221:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 38222:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 38223:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 38224:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 38225:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 38226:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 38227:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 38228:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 38229:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 38230:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 38231:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 38232:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 38233:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 38234:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 38235:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 38236:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 38237:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 38238:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 38239:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 38240:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 38241:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 38242:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 38243:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 38244:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 38245:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 38246:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 38247:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 38248:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 38249:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 38250:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 38251:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 38252:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 38253:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 38254:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 38255:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 38256:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 38257:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 38258:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 38259:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 38260:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 38261:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 38262:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 38263:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 38264:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 38265:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 38266:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 38267:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 38268:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 38269:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 38270:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 38271:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 38272:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 38273:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 38274:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 38275:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 38276:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 38277:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 38278:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 38279:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 38280:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 38281:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 38282:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 38283:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 38284:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 38285:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 38286:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 38287:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 38288:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 38289:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 38290:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 38291:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 38292:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 38293:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 38294:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 38295:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 38296:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 38297:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 38298:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 38299:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 38300:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 38301:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 38302:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 38303:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 38304:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 38305:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 38306:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 38307:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 38308:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 38309:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 38310:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 38311:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 38312:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 38313:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 38314:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 38315:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 38316:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 38317:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 38318:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 38319:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 38320:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 38321:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 38322:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 38323:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 38324:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 38325:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 38326:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 38327:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 38328:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 38329:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 38330:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 38331:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 38332:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 38333:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 38334:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 38335:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 38336:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 38337:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 38338:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 38339:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 38340:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 38341:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 38342:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 38343:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 38344:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 38345:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 38346:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 38347:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 38348:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 38349:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 38350:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 38351:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 38352:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 38353:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 38354:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 38355:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 38356:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 38357:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 38358:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 38359:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 38360:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 38361:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 38362:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 38363:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 38364:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 38365:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 38366:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 38367:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 38368:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 38369:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 38370:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 38371:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 38372:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 38373:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 38374:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 38375:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 38376:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 38377:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 38378:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 38379:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 38380:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 38381:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 38382:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 38383:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 38384:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 38385:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 38386:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 38387:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 38388:22]
  assign io_z = ~x122; // @[Snxn100k.scala 38389:17]
endmodule
module SnxnLv3Inst21(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst84_io_a; // @[Snxn100k.scala 10392:34]
  wire  inst_SnxnLv4Inst84_io_b; // @[Snxn100k.scala 10392:34]
  wire  inst_SnxnLv4Inst84_io_z; // @[Snxn100k.scala 10392:34]
  wire  inst_SnxnLv4Inst85_io_a; // @[Snxn100k.scala 10396:34]
  wire  inst_SnxnLv4Inst85_io_b; // @[Snxn100k.scala 10396:34]
  wire  inst_SnxnLv4Inst85_io_z; // @[Snxn100k.scala 10396:34]
  wire  inst_SnxnLv4Inst86_io_a; // @[Snxn100k.scala 10400:34]
  wire  inst_SnxnLv4Inst86_io_b; // @[Snxn100k.scala 10400:34]
  wire  inst_SnxnLv4Inst86_io_z; // @[Snxn100k.scala 10400:34]
  wire  inst_SnxnLv4Inst87_io_a; // @[Snxn100k.scala 10404:34]
  wire  inst_SnxnLv4Inst87_io_b; // @[Snxn100k.scala 10404:34]
  wire  inst_SnxnLv4Inst87_io_z; // @[Snxn100k.scala 10404:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst84_io_z + inst_SnxnLv4Inst85_io_z; // @[Snxn100k.scala 10408:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst86_io_z; // @[Snxn100k.scala 10408:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst87_io_z; // @[Snxn100k.scala 10408:89]
  SnxnLv4Inst84 inst_SnxnLv4Inst84 ( // @[Snxn100k.scala 10392:34]
    .io_a(inst_SnxnLv4Inst84_io_a),
    .io_b(inst_SnxnLv4Inst84_io_b),
    .io_z(inst_SnxnLv4Inst84_io_z)
  );
  SnxnLv4Inst83 inst_SnxnLv4Inst85 ( // @[Snxn100k.scala 10396:34]
    .io_a(inst_SnxnLv4Inst85_io_a),
    .io_b(inst_SnxnLv4Inst85_io_b),
    .io_z(inst_SnxnLv4Inst85_io_z)
  );
  SnxnLv4Inst86 inst_SnxnLv4Inst86 ( // @[Snxn100k.scala 10400:34]
    .io_a(inst_SnxnLv4Inst86_io_a),
    .io_b(inst_SnxnLv4Inst86_io_b),
    .io_z(inst_SnxnLv4Inst86_io_z)
  );
  SnxnLv4Inst75 inst_SnxnLv4Inst87 ( // @[Snxn100k.scala 10404:34]
    .io_a(inst_SnxnLv4Inst87_io_a),
    .io_b(inst_SnxnLv4Inst87_io_b),
    .io_z(inst_SnxnLv4Inst87_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10409:15]
  assign inst_SnxnLv4Inst84_io_a = io_a; // @[Snxn100k.scala 10393:27]
  assign inst_SnxnLv4Inst84_io_b = io_b; // @[Snxn100k.scala 10394:27]
  assign inst_SnxnLv4Inst85_io_a = io_a; // @[Snxn100k.scala 10397:27]
  assign inst_SnxnLv4Inst85_io_b = io_b; // @[Snxn100k.scala 10398:27]
  assign inst_SnxnLv4Inst86_io_a = io_a; // @[Snxn100k.scala 10401:27]
  assign inst_SnxnLv4Inst86_io_b = io_b; // @[Snxn100k.scala 10402:27]
  assign inst_SnxnLv4Inst87_io_a = io_a; // @[Snxn100k.scala 10405:27]
  assign inst_SnxnLv4Inst87_io_b = io_b; // @[Snxn100k.scala 10406:27]
endmodule
module SnxnLv3Inst22(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst88_io_a; // @[Snxn100k.scala 11301:34]
  wire  inst_SnxnLv4Inst88_io_b; // @[Snxn100k.scala 11301:34]
  wire  inst_SnxnLv4Inst88_io_z; // @[Snxn100k.scala 11301:34]
  wire  inst_SnxnLv4Inst89_io_a; // @[Snxn100k.scala 11305:34]
  wire  inst_SnxnLv4Inst89_io_b; // @[Snxn100k.scala 11305:34]
  wire  inst_SnxnLv4Inst89_io_z; // @[Snxn100k.scala 11305:34]
  wire  inst_SnxnLv4Inst90_io_a; // @[Snxn100k.scala 11309:34]
  wire  inst_SnxnLv4Inst90_io_b; // @[Snxn100k.scala 11309:34]
  wire  inst_SnxnLv4Inst90_io_z; // @[Snxn100k.scala 11309:34]
  wire  inst_SnxnLv4Inst91_io_a; // @[Snxn100k.scala 11313:34]
  wire  inst_SnxnLv4Inst91_io_b; // @[Snxn100k.scala 11313:34]
  wire  inst_SnxnLv4Inst91_io_z; // @[Snxn100k.scala 11313:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst88_io_z + inst_SnxnLv4Inst89_io_z; // @[Snxn100k.scala 11317:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst90_io_z; // @[Snxn100k.scala 11317:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst91_io_z; // @[Snxn100k.scala 11317:89]
  SnxnLv4Inst23 inst_SnxnLv4Inst88 ( // @[Snxn100k.scala 11301:34]
    .io_a(inst_SnxnLv4Inst88_io_a),
    .io_b(inst_SnxnLv4Inst88_io_b),
    .io_z(inst_SnxnLv4Inst88_io_z)
  );
  SnxnLv4Inst4 inst_SnxnLv4Inst89 ( // @[Snxn100k.scala 11305:34]
    .io_a(inst_SnxnLv4Inst89_io_a),
    .io_b(inst_SnxnLv4Inst89_io_b),
    .io_z(inst_SnxnLv4Inst89_io_z)
  );
  SnxnLv4Inst28 inst_SnxnLv4Inst90 ( // @[Snxn100k.scala 11309:34]
    .io_a(inst_SnxnLv4Inst90_io_a),
    .io_b(inst_SnxnLv4Inst90_io_b),
    .io_z(inst_SnxnLv4Inst90_io_z)
  );
  SnxnLv4Inst78 inst_SnxnLv4Inst91 ( // @[Snxn100k.scala 11313:34]
    .io_a(inst_SnxnLv4Inst91_io_a),
    .io_b(inst_SnxnLv4Inst91_io_b),
    .io_z(inst_SnxnLv4Inst91_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11318:15]
  assign inst_SnxnLv4Inst88_io_a = io_a; // @[Snxn100k.scala 11302:27]
  assign inst_SnxnLv4Inst88_io_b = io_b; // @[Snxn100k.scala 11303:27]
  assign inst_SnxnLv4Inst89_io_a = io_a; // @[Snxn100k.scala 11306:27]
  assign inst_SnxnLv4Inst89_io_b = io_b; // @[Snxn100k.scala 11307:27]
  assign inst_SnxnLv4Inst90_io_a = io_a; // @[Snxn100k.scala 11310:27]
  assign inst_SnxnLv4Inst90_io_b = io_b; // @[Snxn100k.scala 11311:27]
  assign inst_SnxnLv4Inst91_io_a = io_a; // @[Snxn100k.scala 11314:27]
  assign inst_SnxnLv4Inst91_io_b = io_b; // @[Snxn100k.scala 11315:27]
endmodule
module SnxnLv4Inst95(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 38400:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 38401:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 38402:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 38403:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 38404:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 38405:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 38406:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 38407:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 38408:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 38409:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 38410:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 38411:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 38412:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 38413:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 38414:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 38415:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 38416:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 38417:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 38418:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 38419:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 38420:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 38421:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 38422:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 38423:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 38424:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 38425:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 38426:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 38427:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 38428:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 38429:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 38430:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 38431:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 38432:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 38433:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 38434:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 38435:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 38436:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 38437:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 38438:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 38439:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 38440:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 38441:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 38442:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 38443:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 38444:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 38445:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 38446:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 38447:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 38448:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 38449:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 38450:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 38451:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 38452:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 38453:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 38454:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 38455:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 38456:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 38457:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 38458:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 38459:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 38460:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 38461:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 38462:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 38463:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 38464:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 38465:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 38466:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 38467:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 38468:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 38469:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 38470:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 38471:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 38472:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 38473:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 38474:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 38475:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 38476:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 38477:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 38478:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 38479:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 38480:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 38481:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 38482:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 38483:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 38484:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 38485:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 38486:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 38487:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 38488:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 38489:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 38490:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 38491:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 38492:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 38493:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 38494:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 38495:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 38496:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 38497:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 38498:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 38499:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 38500:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 38501:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 38502:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 38503:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 38504:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 38505:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 38506:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 38507:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 38508:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 38509:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 38510:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 38511:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 38512:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 38513:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 38514:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 38515:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 38516:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 38517:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 38518:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 38519:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 38520:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 38521:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 38522:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 38523:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 38524:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 38525:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 38526:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 38527:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 38528:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 38529:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 38530:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 38531:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 38532:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 38533:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 38534:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 38535:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 38536:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 38537:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 38538:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 38539:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 38540:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 38541:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 38542:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 38543:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 38544:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 38545:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 38546:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 38547:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 38548:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 38549:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 38550:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 38551:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 38552:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 38553:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 38554:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 38555:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 38556:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 38557:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 38558:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 38559:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 38560:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 38561:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 38562:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 38563:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 38564:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 38565:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 38566:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 38567:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 38568:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 38569:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 38570:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 38571:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 38572:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 38573:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 38574:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 38575:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 38576:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 38577:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 38578:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 38579:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 38580:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 38581:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 38582:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 38583:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 38584:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 38585:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 38586:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 38587:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 38588:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 38589:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 38590:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 38591:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 38592:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 38593:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 38594:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 38595:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 38596:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 38597:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 38598:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 38599:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 38600:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 38601:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 38602:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 38603:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 38604:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 38605:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 38606:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 38607:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 38608:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 38609:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 38610:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 38611:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 38612:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 38613:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 38614:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 38615:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 38616:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 38617:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 38618:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 38619:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 38620:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 38621:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 38622:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 38623:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 38624:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 38625:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 38626:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 38627:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 38628:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 38629:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 38630:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 38631:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 38632:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 38633:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 38634:20]
  assign io_z = ~x58; // @[Snxn100k.scala 38635:16]
endmodule
module SnxnLv3Inst23(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst92_io_a; // @[Snxn100k.scala 10695:34]
  wire  inst_SnxnLv4Inst92_io_b; // @[Snxn100k.scala 10695:34]
  wire  inst_SnxnLv4Inst92_io_z; // @[Snxn100k.scala 10695:34]
  wire  inst_SnxnLv4Inst93_io_a; // @[Snxn100k.scala 10699:34]
  wire  inst_SnxnLv4Inst93_io_b; // @[Snxn100k.scala 10699:34]
  wire  inst_SnxnLv4Inst93_io_z; // @[Snxn100k.scala 10699:34]
  wire  inst_SnxnLv4Inst94_io_a; // @[Snxn100k.scala 10703:34]
  wire  inst_SnxnLv4Inst94_io_b; // @[Snxn100k.scala 10703:34]
  wire  inst_SnxnLv4Inst94_io_z; // @[Snxn100k.scala 10703:34]
  wire  inst_SnxnLv4Inst95_io_a; // @[Snxn100k.scala 10707:34]
  wire  inst_SnxnLv4Inst95_io_b; // @[Snxn100k.scala 10707:34]
  wire  inst_SnxnLv4Inst95_io_z; // @[Snxn100k.scala 10707:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst92_io_z + inst_SnxnLv4Inst93_io_z; // @[Snxn100k.scala 10711:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst94_io_z; // @[Snxn100k.scala 10711:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst95_io_z; // @[Snxn100k.scala 10711:89]
  SnxnLv4Inst20 inst_SnxnLv4Inst92 ( // @[Snxn100k.scala 10695:34]
    .io_a(inst_SnxnLv4Inst92_io_a),
    .io_b(inst_SnxnLv4Inst92_io_b),
    .io_z(inst_SnxnLv4Inst92_io_z)
  );
  SnxnLv4Inst19 inst_SnxnLv4Inst93 ( // @[Snxn100k.scala 10699:34]
    .io_a(inst_SnxnLv4Inst93_io_a),
    .io_b(inst_SnxnLv4Inst93_io_b),
    .io_z(inst_SnxnLv4Inst93_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst94 ( // @[Snxn100k.scala 10703:34]
    .io_a(inst_SnxnLv4Inst94_io_a),
    .io_b(inst_SnxnLv4Inst94_io_b),
    .io_z(inst_SnxnLv4Inst94_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst95 ( // @[Snxn100k.scala 10707:34]
    .io_a(inst_SnxnLv4Inst95_io_a),
    .io_b(inst_SnxnLv4Inst95_io_b),
    .io_z(inst_SnxnLv4Inst95_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10712:15]
  assign inst_SnxnLv4Inst92_io_a = io_a; // @[Snxn100k.scala 10696:27]
  assign inst_SnxnLv4Inst92_io_b = io_b; // @[Snxn100k.scala 10697:27]
  assign inst_SnxnLv4Inst93_io_a = io_a; // @[Snxn100k.scala 10700:27]
  assign inst_SnxnLv4Inst93_io_b = io_b; // @[Snxn100k.scala 10701:27]
  assign inst_SnxnLv4Inst94_io_a = io_a; // @[Snxn100k.scala 10704:27]
  assign inst_SnxnLv4Inst94_io_b = io_b; // @[Snxn100k.scala 10705:27]
  assign inst_SnxnLv4Inst95_io_a = io_a; // @[Snxn100k.scala 10708:27]
  assign inst_SnxnLv4Inst95_io_b = io_b; // @[Snxn100k.scala 10709:27]
endmodule
module SnxnLv2Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst20_io_a; // @[Snxn100k.scala 2298:34]
  wire  inst_SnxnLv3Inst20_io_b; // @[Snxn100k.scala 2298:34]
  wire  inst_SnxnLv3Inst20_io_z; // @[Snxn100k.scala 2298:34]
  wire  inst_SnxnLv3Inst21_io_a; // @[Snxn100k.scala 2302:34]
  wire  inst_SnxnLv3Inst21_io_b; // @[Snxn100k.scala 2302:34]
  wire  inst_SnxnLv3Inst21_io_z; // @[Snxn100k.scala 2302:34]
  wire  inst_SnxnLv3Inst22_io_a; // @[Snxn100k.scala 2306:34]
  wire  inst_SnxnLv3Inst22_io_b; // @[Snxn100k.scala 2306:34]
  wire  inst_SnxnLv3Inst22_io_z; // @[Snxn100k.scala 2306:34]
  wire  inst_SnxnLv3Inst23_io_a; // @[Snxn100k.scala 2310:34]
  wire  inst_SnxnLv3Inst23_io_b; // @[Snxn100k.scala 2310:34]
  wire  inst_SnxnLv3Inst23_io_z; // @[Snxn100k.scala 2310:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst20_io_z + inst_SnxnLv3Inst21_io_z; // @[Snxn100k.scala 2314:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst22_io_z; // @[Snxn100k.scala 2314:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst23_io_z; // @[Snxn100k.scala 2314:89]
  SnxnLv3Inst20 inst_SnxnLv3Inst20 ( // @[Snxn100k.scala 2298:34]
    .io_a(inst_SnxnLv3Inst20_io_a),
    .io_b(inst_SnxnLv3Inst20_io_b),
    .io_z(inst_SnxnLv3Inst20_io_z)
  );
  SnxnLv3Inst21 inst_SnxnLv3Inst21 ( // @[Snxn100k.scala 2302:34]
    .io_a(inst_SnxnLv3Inst21_io_a),
    .io_b(inst_SnxnLv3Inst21_io_b),
    .io_z(inst_SnxnLv3Inst21_io_z)
  );
  SnxnLv3Inst22 inst_SnxnLv3Inst22 ( // @[Snxn100k.scala 2306:34]
    .io_a(inst_SnxnLv3Inst22_io_a),
    .io_b(inst_SnxnLv3Inst22_io_b),
    .io_z(inst_SnxnLv3Inst22_io_z)
  );
  SnxnLv3Inst23 inst_SnxnLv3Inst23 ( // @[Snxn100k.scala 2310:34]
    .io_a(inst_SnxnLv3Inst23_io_a),
    .io_b(inst_SnxnLv3Inst23_io_b),
    .io_z(inst_SnxnLv3Inst23_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 2315:15]
  assign inst_SnxnLv3Inst20_io_a = io_a; // @[Snxn100k.scala 2299:27]
  assign inst_SnxnLv3Inst20_io_b = io_b; // @[Snxn100k.scala 2300:27]
  assign inst_SnxnLv3Inst21_io_a = io_a; // @[Snxn100k.scala 2303:27]
  assign inst_SnxnLv3Inst21_io_b = io_b; // @[Snxn100k.scala 2304:27]
  assign inst_SnxnLv3Inst22_io_a = io_a; // @[Snxn100k.scala 2307:27]
  assign inst_SnxnLv3Inst22_io_b = io_b; // @[Snxn100k.scala 2308:27]
  assign inst_SnxnLv3Inst23_io_a = io_a; // @[Snxn100k.scala 2311:27]
  assign inst_SnxnLv3Inst23_io_b = io_b; // @[Snxn100k.scala 2312:27]
endmodule
module SnxnLv3Inst24(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst96_io_a; // @[Snxn100k.scala 8509:34]
  wire  inst_SnxnLv4Inst96_io_b; // @[Snxn100k.scala 8509:34]
  wire  inst_SnxnLv4Inst96_io_z; // @[Snxn100k.scala 8509:34]
  wire  inst_SnxnLv4Inst97_io_a; // @[Snxn100k.scala 8513:34]
  wire  inst_SnxnLv4Inst97_io_b; // @[Snxn100k.scala 8513:34]
  wire  inst_SnxnLv4Inst97_io_z; // @[Snxn100k.scala 8513:34]
  wire  inst_SnxnLv4Inst98_io_a; // @[Snxn100k.scala 8517:34]
  wire  inst_SnxnLv4Inst98_io_b; // @[Snxn100k.scala 8517:34]
  wire  inst_SnxnLv4Inst98_io_z; // @[Snxn100k.scala 8517:34]
  wire  inst_SnxnLv4Inst99_io_a; // @[Snxn100k.scala 8521:34]
  wire  inst_SnxnLv4Inst99_io_b; // @[Snxn100k.scala 8521:34]
  wire  inst_SnxnLv4Inst99_io_z; // @[Snxn100k.scala 8521:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst96_io_z + inst_SnxnLv4Inst97_io_z; // @[Snxn100k.scala 8525:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst98_io_z; // @[Snxn100k.scala 8525:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst99_io_z; // @[Snxn100k.scala 8525:89]
  SnxnLv4Inst12 inst_SnxnLv4Inst96 ( // @[Snxn100k.scala 8509:34]
    .io_a(inst_SnxnLv4Inst96_io_a),
    .io_b(inst_SnxnLv4Inst96_io_b),
    .io_z(inst_SnxnLv4Inst96_io_z)
  );
  SnxnLv4Inst38 inst_SnxnLv4Inst97 ( // @[Snxn100k.scala 8513:34]
    .io_a(inst_SnxnLv4Inst97_io_a),
    .io_b(inst_SnxnLv4Inst97_io_b),
    .io_z(inst_SnxnLv4Inst97_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst98 ( // @[Snxn100k.scala 8517:34]
    .io_a(inst_SnxnLv4Inst98_io_a),
    .io_b(inst_SnxnLv4Inst98_io_b),
    .io_z(inst_SnxnLv4Inst98_io_z)
  );
  SnxnLv4Inst10 inst_SnxnLv4Inst99 ( // @[Snxn100k.scala 8521:34]
    .io_a(inst_SnxnLv4Inst99_io_a),
    .io_b(inst_SnxnLv4Inst99_io_b),
    .io_z(inst_SnxnLv4Inst99_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 8526:15]
  assign inst_SnxnLv4Inst96_io_a = io_a; // @[Snxn100k.scala 8510:27]
  assign inst_SnxnLv4Inst96_io_b = io_b; // @[Snxn100k.scala 8511:27]
  assign inst_SnxnLv4Inst97_io_a = io_a; // @[Snxn100k.scala 8514:27]
  assign inst_SnxnLv4Inst97_io_b = io_b; // @[Snxn100k.scala 8515:27]
  assign inst_SnxnLv4Inst98_io_a = io_a; // @[Snxn100k.scala 8518:27]
  assign inst_SnxnLv4Inst98_io_b = io_b; // @[Snxn100k.scala 8519:27]
  assign inst_SnxnLv4Inst99_io_a = io_a; // @[Snxn100k.scala 8522:27]
  assign inst_SnxnLv4Inst99_io_b = io_b; // @[Snxn100k.scala 8523:27]
endmodule
module SnxnLv4Inst101(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 27942:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 27943:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 27944:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 27945:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 27946:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 27947:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 27948:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 27949:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 27950:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 27951:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 27952:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 27953:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 27954:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 27955:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 27956:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 27957:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 27958:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 27959:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 27960:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 27961:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 27962:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 27963:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 27964:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 27965:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 27966:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 27967:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 27968:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 27969:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 27970:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 27971:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 27972:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 27973:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 27974:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 27975:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 27976:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 27977:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 27978:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 27979:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 27980:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 27981:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 27982:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 27983:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 27984:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 27985:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 27986:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 27987:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 27988:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 27989:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 27990:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 27991:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 27992:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 27993:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 27994:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 27995:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 27996:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 27997:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 27998:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 27999:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 28000:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 28001:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 28002:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 28003:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 28004:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 28005:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 28006:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 28007:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 28008:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 28009:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 28010:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 28011:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 28012:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 28013:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 28014:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 28015:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 28016:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 28017:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 28018:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 28019:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 28020:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 28021:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 28022:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 28023:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 28024:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 28025:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 28026:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 28027:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 28028:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 28029:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 28030:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 28031:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 28032:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 28033:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 28034:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 28035:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 28036:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 28037:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 28038:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 28039:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 28040:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 28041:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 28042:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 28043:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 28044:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 28045:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 28046:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 28047:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 28048:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 28049:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 28050:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 28051:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 28052:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 28053:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 28054:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 28055:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 28056:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 28057:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 28058:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 28059:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 28060:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 28061:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 28062:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 28063:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 28064:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 28065:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 28066:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 28067:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 28068:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 28069:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 28070:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 28071:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 28072:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 28073:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 28074:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 28075:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 28076:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 28077:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 28078:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 28079:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 28080:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 28081:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 28082:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 28083:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 28084:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 28085:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 28086:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 28087:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 28088:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 28089:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 28090:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 28091:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 28092:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 28093:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 28094:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 28095:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 28096:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 28097:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 28098:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 28099:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 28100:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 28101:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 28102:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 28103:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 28104:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 28105:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 28106:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 28107:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 28108:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 28109:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 28110:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 28111:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 28112:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 28113:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 28114:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 28115:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 28116:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 28117:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 28118:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 28119:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 28120:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 28121:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 28122:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 28123:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 28124:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 28125:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 28126:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 28127:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 28128:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 28129:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 28130:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 28131:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 28132:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 28133:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 28134:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 28135:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 28136:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 28137:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 28138:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 28139:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 28140:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 28141:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 28142:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 28143:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 28144:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 28145:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 28146:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 28147:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 28148:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 28149:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 28150:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 28151:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 28152:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 28153:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 28154:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 28155:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 28156:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 28157:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 28158:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 28159:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 28160:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 28161:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 28162:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 28163:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 28164:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 28165:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 28166:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 28167:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 28168:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 28169:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 28170:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 28171:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 28172:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 28173:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 28174:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 28175:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 28176:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 28177:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 28178:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 28179:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 28180:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 28181:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 28182:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 28183:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 28184:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 28185:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 28186:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 28187:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 28188:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 28189:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 28190:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 28191:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 28192:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 28193:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 28194:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 28195:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 28196:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 28197:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 28198:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 28199:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 28200:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 28201:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 28202:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 28203:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 28204:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 28205:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 28206:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 28207:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 28208:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 28209:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 28210:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 28211:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 28212:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 28213:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 28214:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 28215:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 28216:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 28217:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 28218:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 28219:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 28220:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 28221:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 28222:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 28223:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 28224:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 28225:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 28226:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 28227:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 28228:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 28229:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 28230:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 28231:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 28232:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 28233:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 28234:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 28235:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 28236:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 28237:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 28238:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 28239:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 28240:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 28241:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 28242:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 28243:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 28244:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 28245:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 28246:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 28247:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 28248:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 28249:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 28250:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 28251:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 28252:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 28253:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 28254:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 28255:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 28256:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 28257:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 28258:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 28259:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 28260:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 28261:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 28262:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 28263:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 28264:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 28265:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 28266:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 28267:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 28268:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 28269:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 28270:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 28271:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 28272:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 28273:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 28274:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 28275:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 28276:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 28277:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 28278:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 28279:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 28280:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 28281:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 28282:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 28283:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 28284:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 28285:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 28286:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 28287:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 28288:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 28289:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 28290:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 28291:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 28292:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 28293:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 28294:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 28295:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 28296:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 28297:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 28298:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 28299:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 28300:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 28301:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 28302:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 28303:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 28304:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 28305:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 28306:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 28307:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 28308:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 28309:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 28310:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 28311:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 28312:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 28313:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 28314:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 28315:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 28316:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 28317:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 28318:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 28319:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 28320:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 28321:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 28322:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 28323:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 28324:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 28325:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 28326:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 28327:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 28328:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 28329:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 28330:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 28331:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 28332:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 28333:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 28334:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 28335:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 28336:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 28337:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 28338:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 28339:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 28340:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 28341:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 28342:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 28343:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 28344:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 28345:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 28346:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 28347:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 28348:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 28349:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 28350:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 28351:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 28352:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 28353:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 28354:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 28355:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 28356:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 28357:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 28358:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 28359:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 28360:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 28361:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 28362:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 28363:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 28364:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 28365:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 28366:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 28367:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 28368:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 28369:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 28370:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 28371:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 28372:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 28373:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 28374:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 28375:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 28376:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 28377:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 28378:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 28379:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 28380:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 28381:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 28382:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 28383:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 28384:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 28385:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 28386:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 28387:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 28388:22]
  assign io_z = ~x111; // @[Snxn100k.scala 28389:17]
endmodule
module SnxnLv4Inst103(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 27676:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 27677:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 27678:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 27679:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 27680:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 27681:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 27682:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 27683:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 27684:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 27685:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 27686:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 27687:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 27688:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 27689:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 27690:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 27691:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 27692:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 27693:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 27694:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 27695:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 27696:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 27697:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 27698:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 27699:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 27700:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 27701:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 27702:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 27703:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 27704:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 27705:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 27706:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 27707:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 27708:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 27709:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 27710:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 27711:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 27712:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 27713:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 27714:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 27715:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 27716:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 27717:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 27718:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 27719:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 27720:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 27721:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 27722:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 27723:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 27724:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 27725:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 27726:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 27727:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 27728:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 27729:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 27730:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 27731:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 27732:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 27733:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 27734:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 27735:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 27736:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 27737:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 27738:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 27739:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 27740:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 27741:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 27742:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 27743:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 27744:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 27745:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 27746:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 27747:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 27748:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 27749:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 27750:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 27751:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 27752:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 27753:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 27754:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 27755:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 27756:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 27757:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 27758:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 27759:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 27760:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 27761:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 27762:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 27763:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 27764:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 27765:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 27766:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 27767:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 27768:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 27769:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 27770:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 27771:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 27772:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 27773:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 27774:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 27775:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 27776:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 27777:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 27778:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 27779:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 27780:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 27781:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 27782:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 27783:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 27784:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 27785:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 27786:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 27787:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 27788:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 27789:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 27790:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 27791:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 27792:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 27793:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 27794:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 27795:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 27796:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 27797:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 27798:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 27799:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 27800:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 27801:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 27802:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 27803:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 27804:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 27805:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 27806:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 27807:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 27808:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 27809:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 27810:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 27811:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 27812:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 27813:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 27814:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 27815:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 27816:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 27817:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 27818:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 27819:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 27820:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 27821:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 27822:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 27823:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 27824:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 27825:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 27826:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 27827:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 27828:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 27829:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 27830:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 27831:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 27832:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 27833:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 27834:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 27835:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 27836:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 27837:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 27838:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 27839:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 27840:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 27841:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 27842:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 27843:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 27844:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 27845:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 27846:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 27847:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 27848:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 27849:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 27850:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 27851:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 27852:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 27853:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 27854:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 27855:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 27856:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 27857:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 27858:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 27859:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 27860:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 27861:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 27862:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 27863:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 27864:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 27865:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 27866:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 27867:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 27868:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 27869:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 27870:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 27871:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 27872:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 27873:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 27874:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 27875:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 27876:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 27877:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 27878:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 27879:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 27880:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 27881:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 27882:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 27883:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 27884:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 27885:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 27886:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 27887:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 27888:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 27889:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 27890:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 27891:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 27892:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 27893:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 27894:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 27895:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 27896:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 27897:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 27898:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 27899:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 27900:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 27901:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 27902:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 27903:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 27904:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 27905:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 27906:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 27907:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 27908:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 27909:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 27910:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 27911:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 27912:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 27913:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 27914:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 27915:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 27916:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 27917:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 27918:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 27919:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 27920:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 27921:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 27922:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 27923:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 27924:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 27925:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 27926:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 27927:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 27928:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 27929:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 27930:20]
  assign io_z = ~x63; // @[Snxn100k.scala 27931:16]
endmodule
module SnxnLv3Inst25(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst100_io_a; // @[Snxn100k.scala 7132:35]
  wire  inst_SnxnLv4Inst100_io_b; // @[Snxn100k.scala 7132:35]
  wire  inst_SnxnLv4Inst100_io_z; // @[Snxn100k.scala 7132:35]
  wire  inst_SnxnLv4Inst101_io_a; // @[Snxn100k.scala 7136:35]
  wire  inst_SnxnLv4Inst101_io_b; // @[Snxn100k.scala 7136:35]
  wire  inst_SnxnLv4Inst101_io_z; // @[Snxn100k.scala 7136:35]
  wire  inst_SnxnLv4Inst102_io_a; // @[Snxn100k.scala 7140:35]
  wire  inst_SnxnLv4Inst102_io_b; // @[Snxn100k.scala 7140:35]
  wire  inst_SnxnLv4Inst102_io_z; // @[Snxn100k.scala 7140:35]
  wire  inst_SnxnLv4Inst103_io_a; // @[Snxn100k.scala 7144:35]
  wire  inst_SnxnLv4Inst103_io_b; // @[Snxn100k.scala 7144:35]
  wire  inst_SnxnLv4Inst103_io_z; // @[Snxn100k.scala 7144:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst100_io_z + inst_SnxnLv4Inst101_io_z; // @[Snxn100k.scala 7148:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst102_io_z; // @[Snxn100k.scala 7148:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst103_io_z; // @[Snxn100k.scala 7148:92]
  SnxnLv4Inst17 inst_SnxnLv4Inst100 ( // @[Snxn100k.scala 7132:35]
    .io_a(inst_SnxnLv4Inst100_io_a),
    .io_b(inst_SnxnLv4Inst100_io_b),
    .io_z(inst_SnxnLv4Inst100_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst101 ( // @[Snxn100k.scala 7136:35]
    .io_a(inst_SnxnLv4Inst101_io_a),
    .io_b(inst_SnxnLv4Inst101_io_b),
    .io_z(inst_SnxnLv4Inst101_io_z)
  );
  SnxnLv4Inst69 inst_SnxnLv4Inst102 ( // @[Snxn100k.scala 7140:35]
    .io_a(inst_SnxnLv4Inst102_io_a),
    .io_b(inst_SnxnLv4Inst102_io_b),
    .io_z(inst_SnxnLv4Inst102_io_z)
  );
  SnxnLv4Inst103 inst_SnxnLv4Inst103 ( // @[Snxn100k.scala 7144:35]
    .io_a(inst_SnxnLv4Inst103_io_a),
    .io_b(inst_SnxnLv4Inst103_io_b),
    .io_z(inst_SnxnLv4Inst103_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7149:15]
  assign inst_SnxnLv4Inst100_io_a = io_a; // @[Snxn100k.scala 7133:28]
  assign inst_SnxnLv4Inst100_io_b = io_b; // @[Snxn100k.scala 7134:28]
  assign inst_SnxnLv4Inst101_io_a = io_a; // @[Snxn100k.scala 7137:28]
  assign inst_SnxnLv4Inst101_io_b = io_b; // @[Snxn100k.scala 7138:28]
  assign inst_SnxnLv4Inst102_io_a = io_a; // @[Snxn100k.scala 7141:28]
  assign inst_SnxnLv4Inst102_io_b = io_b; // @[Snxn100k.scala 7142:28]
  assign inst_SnxnLv4Inst103_io_a = io_a; // @[Snxn100k.scala 7145:28]
  assign inst_SnxnLv4Inst103_io_b = io_b; // @[Snxn100k.scala 7146:28]
endmodule
module SnxnLv4Inst104(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 29032:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 29033:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 29034:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 29035:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 29036:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 29037:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 29038:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 29039:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 29040:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 29041:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 29042:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 29043:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 29044:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 29045:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 29046:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 29047:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 29048:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 29049:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 29050:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 29051:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 29052:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 29053:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 29054:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 29055:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 29056:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 29057:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 29058:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 29059:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 29060:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 29061:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 29062:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 29063:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 29064:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 29065:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 29066:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 29067:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 29068:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 29069:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 29070:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 29071:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 29072:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 29073:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 29074:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 29075:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 29076:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 29077:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 29078:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 29079:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 29080:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 29081:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 29082:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 29083:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 29084:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 29085:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 29086:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 29087:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 29088:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 29089:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 29090:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 29091:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 29092:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 29093:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 29094:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 29095:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 29096:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 29097:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 29098:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 29099:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 29100:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 29101:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 29102:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 29103:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 29104:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 29105:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 29106:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 29107:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 29108:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 29109:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 29110:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 29111:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 29112:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 29113:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 29114:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 29115:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 29116:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 29117:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 29118:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 29119:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 29120:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 29121:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 29122:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 29123:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 29124:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 29125:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 29126:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 29127:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 29128:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 29129:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 29130:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 29131:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 29132:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 29133:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 29134:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 29135:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 29136:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 29137:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 29138:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 29139:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 29140:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 29141:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 29142:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 29143:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 29144:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 29145:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 29146:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 29147:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 29148:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 29149:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 29150:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 29151:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 29152:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 29153:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 29154:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 29155:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 29156:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 29157:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 29158:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 29159:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 29160:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 29161:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 29162:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 29163:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 29164:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 29165:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 29166:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 29167:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 29168:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 29169:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 29170:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 29171:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 29172:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 29173:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 29174:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 29175:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 29176:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 29177:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 29178:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 29179:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 29180:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 29181:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 29182:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 29183:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 29184:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 29185:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 29186:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 29187:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 29188:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 29189:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 29190:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 29191:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 29192:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 29193:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 29194:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 29195:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 29196:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 29197:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 29198:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 29199:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 29200:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 29201:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 29202:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 29203:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 29204:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 29205:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 29206:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 29207:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 29208:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 29209:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 29210:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 29211:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 29212:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 29213:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 29214:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 29215:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 29216:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 29217:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 29218:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 29219:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 29220:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 29221:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 29222:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 29223:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 29224:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 29225:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 29226:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 29227:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 29228:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 29229:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 29230:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 29231:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 29232:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 29233:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 29234:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 29235:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 29236:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 29237:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 29238:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 29239:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 29240:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 29241:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 29242:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 29243:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 29244:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 29245:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 29246:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 29247:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 29248:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 29249:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 29250:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 29251:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 29252:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 29253:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 29254:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 29255:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 29256:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 29257:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 29258:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 29259:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 29260:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 29261:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 29262:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 29263:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 29264:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 29265:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 29266:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 29267:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 29268:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 29269:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 29270:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 29271:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 29272:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 29273:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 29274:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 29275:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 29276:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 29277:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 29278:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 29279:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 29280:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 29281:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 29282:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 29283:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 29284:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 29285:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 29286:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 29287:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 29288:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 29289:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 29290:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 29291:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 29292:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 29293:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 29294:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 29295:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 29296:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 29297:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 29298:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 29299:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 29300:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 29301:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 29302:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 29303:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 29304:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 29305:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 29306:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 29307:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 29308:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 29309:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 29310:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 29311:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 29312:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 29313:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 29314:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 29315:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 29316:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 29317:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 29318:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 29319:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 29320:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 29321:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 29322:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 29323:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 29324:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 29325:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 29326:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 29327:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 29328:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 29329:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 29330:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 29331:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 29332:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 29333:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 29334:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 29335:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 29336:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 29337:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 29338:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 29339:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 29340:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 29341:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 29342:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 29343:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 29344:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 29345:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 29346:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 29347:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 29348:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 29349:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 29350:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 29351:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 29352:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 29353:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 29354:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 29355:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 29356:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 29357:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 29358:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 29359:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 29360:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 29361:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 29362:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 29363:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 29364:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 29365:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 29366:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 29367:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 29368:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 29369:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 29370:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 29371:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 29372:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 29373:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 29374:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 29375:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 29376:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 29377:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 29378:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 29379:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 29380:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 29381:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 29382:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 29383:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 29384:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 29385:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 29386:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 29387:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 29388:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 29389:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 29390:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 29391:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 29392:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 29393:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 29394:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 29395:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 29396:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 29397:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 29398:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 29399:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 29400:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 29401:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 29402:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 29403:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 29404:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 29405:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 29406:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 29407:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 29408:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 29409:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 29410:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 29411:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 29412:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 29413:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 29414:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 29415:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 29416:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 29417:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 29418:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 29419:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 29420:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 29421:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 29422:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 29423:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 29424:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 29425:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 29426:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 29427:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 29428:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 29429:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 29430:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 29431:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 29432:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 29433:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 29434:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 29435:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 29436:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 29437:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 29438:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 29439:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 29440:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 29441:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 29442:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 29443:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 29444:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 29445:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 29446:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 29447:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 29448:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 29449:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 29450:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 29451:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 29452:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 29453:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 29454:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 29455:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 29456:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 29457:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 29458:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 29459:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 29460:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 29461:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 29462:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 29463:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 29464:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 29465:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 29466:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 29467:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 29468:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 29469:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 29470:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 29471:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 29472:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 29473:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 29474:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 29475:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 29476:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 29477:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 29478:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 29479:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 29480:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 29481:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 29482:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 29483:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 29484:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 29485:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 29486:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 29487:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 29488:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 29489:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 29490:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 29491:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 29492:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 29493:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 29494:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 29495:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 29496:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 29497:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 29498:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 29499:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 29500:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 29501:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 29502:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 29503:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 29504:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 29505:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 29506:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 29507:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 29508:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 29509:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 29510:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 29511:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 29512:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 29513:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 29514:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 29515:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 29516:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 29517:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 29518:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 29519:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 29520:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 29521:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 29522:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 29523:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 29524:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 29525:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 29526:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 29527:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 29528:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 29529:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 29530:22]
  assign io_z = ~x124; // @[Snxn100k.scala 29531:17]
endmodule
module SnxnLv4Inst105(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 28566:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 28567:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 28568:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 28569:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 28570:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 28571:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 28572:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 28573:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 28574:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 28575:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 28576:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 28577:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 28578:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 28579:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 28580:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 28581:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 28582:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 28583:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 28584:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 28585:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 28586:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 28587:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 28588:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 28589:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 28590:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 28591:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 28592:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 28593:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 28594:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 28595:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 28596:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 28597:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 28598:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 28599:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 28600:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 28601:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 28602:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 28603:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 28604:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 28605:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 28606:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 28607:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 28608:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 28609:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 28610:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 28611:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 28612:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 28613:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 28614:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 28615:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 28616:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 28617:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 28618:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 28619:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 28620:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 28621:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 28622:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 28623:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 28624:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 28625:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 28626:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 28627:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 28628:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 28629:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 28630:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 28631:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 28632:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 28633:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 28634:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 28635:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 28636:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 28637:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 28638:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 28639:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 28640:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 28641:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 28642:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 28643:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 28644:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 28645:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 28646:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 28647:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 28648:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 28649:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 28650:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 28651:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 28652:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 28653:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 28654:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 28655:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 28656:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 28657:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 28658:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 28659:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 28660:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 28661:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 28662:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 28663:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 28664:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 28665:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 28666:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 28667:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 28668:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 28669:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 28670:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 28671:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 28672:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 28673:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 28674:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 28675:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 28676:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 28677:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 28678:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 28679:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 28680:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 28681:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 28682:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 28683:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 28684:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 28685:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 28686:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 28687:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 28688:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 28689:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 28690:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 28691:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 28692:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 28693:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 28694:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 28695:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 28696:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 28697:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 28698:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 28699:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 28700:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 28701:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 28702:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 28703:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 28704:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 28705:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 28706:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 28707:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 28708:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 28709:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 28710:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 28711:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 28712:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 28713:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 28714:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 28715:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 28716:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 28717:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 28718:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 28719:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 28720:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 28721:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 28722:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 28723:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 28724:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 28725:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 28726:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 28727:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 28728:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 28729:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 28730:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 28731:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 28732:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 28733:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 28734:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 28735:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 28736:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 28737:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 28738:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 28739:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 28740:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 28741:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 28742:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 28743:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 28744:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 28745:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 28746:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 28747:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 28748:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 28749:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 28750:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 28751:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 28752:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 28753:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 28754:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 28755:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 28756:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 28757:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 28758:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 28759:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 28760:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 28761:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 28762:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 28763:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 28764:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 28765:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 28766:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 28767:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 28768:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 28769:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 28770:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 28771:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 28772:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 28773:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 28774:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 28775:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 28776:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 28777:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 28778:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 28779:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 28780:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 28781:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 28782:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 28783:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 28784:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 28785:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 28786:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 28787:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 28788:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 28789:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 28790:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 28791:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 28792:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 28793:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 28794:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 28795:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 28796:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 28797:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 28798:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 28799:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 28800:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 28801:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 28802:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 28803:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 28804:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 28805:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 28806:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 28807:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 28808:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 28809:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 28810:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 28811:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 28812:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 28813:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 28814:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 28815:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 28816:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 28817:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 28818:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 28819:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 28820:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 28821:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 28822:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 28823:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 28824:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 28825:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 28826:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 28827:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 28828:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 28829:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 28830:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 28831:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 28832:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 28833:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 28834:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 28835:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 28836:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 28837:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 28838:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 28839:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 28840:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 28841:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 28842:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 28843:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 28844:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 28845:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 28846:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 28847:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 28848:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 28849:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 28850:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 28851:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 28852:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 28853:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 28854:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 28855:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 28856:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 28857:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 28858:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 28859:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 28860:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 28861:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 28862:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 28863:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 28864:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 28865:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 28866:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 28867:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 28868:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 28869:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 28870:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 28871:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 28872:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 28873:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 28874:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 28875:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 28876:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 28877:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 28878:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 28879:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 28880:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 28881:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 28882:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 28883:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 28884:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 28885:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 28886:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 28887:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 28888:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 28889:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 28890:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 28891:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 28892:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 28893:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 28894:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 28895:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 28896:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 28897:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 28898:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 28899:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 28900:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 28901:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 28902:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 28903:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 28904:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 28905:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 28906:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 28907:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 28908:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 28909:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 28910:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 28911:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 28912:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 28913:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 28914:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 28915:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 28916:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 28917:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 28918:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 28919:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 28920:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 28921:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 28922:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 28923:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 28924:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 28925:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 28926:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 28927:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 28928:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 28929:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 28930:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 28931:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 28932:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 28933:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 28934:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 28935:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 28936:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 28937:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 28938:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 28939:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 28940:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 28941:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 28942:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 28943:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 28944:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 28945:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 28946:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 28947:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 28948:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 28949:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 28950:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 28951:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 28952:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 28953:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 28954:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 28955:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 28956:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 28957:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 28958:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 28959:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 28960:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 28961:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 28962:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 28963:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 28964:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 28965:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 28966:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 28967:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 28968:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 28969:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 28970:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 28971:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 28972:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 28973:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 28974:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 28975:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 28976:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 28977:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 28978:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 28979:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 28980:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 28981:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 28982:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 28983:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 28984:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 28985:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 28986:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 28987:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 28988:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 28989:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 28990:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 28991:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 28992:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 28993:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 28994:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 28995:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 28996:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 28997:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 28998:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 28999:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 29000:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 29001:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 29002:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 29003:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 29004:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 29005:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 29006:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 29007:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 29008:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 29009:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 29010:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 29011:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 29012:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 29013:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 29014:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 29015:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 29016:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 29017:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 29018:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 29019:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 29020:22]
  assign io_z = ~x113; // @[Snxn100k.scala 29021:17]
endmodule
module SnxnLv4Inst106(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 29542:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 29543:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 29544:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 29545:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 29546:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 29547:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 29548:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 29549:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 29550:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 29551:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 29552:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 29553:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 29554:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 29555:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 29556:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 29557:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 29558:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 29559:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 29560:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 29561:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 29562:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 29563:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 29564:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 29565:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 29566:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 29567:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 29568:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 29569:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 29570:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 29571:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 29572:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 29573:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 29574:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 29575:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 29576:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 29577:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 29578:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 29579:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 29580:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 29581:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 29582:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 29583:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 29584:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 29585:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 29586:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 29587:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 29588:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 29589:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 29590:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 29591:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 29592:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 29593:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 29594:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 29595:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 29596:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 29597:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 29598:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 29599:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 29600:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 29601:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 29602:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 29603:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 29604:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 29605:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 29606:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 29607:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 29608:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 29609:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 29610:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 29611:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 29612:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 29613:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 29614:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 29615:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 29616:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 29617:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 29618:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 29619:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 29620:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 29621:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 29622:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 29623:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 29624:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 29625:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 29626:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 29627:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 29628:20]
  assign io_z = ~x21; // @[Snxn100k.scala 29629:16]
endmodule
module SnxnLv4Inst107(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 28400:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 28401:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 28402:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 28403:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 28404:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 28405:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 28406:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 28407:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 28408:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 28409:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 28410:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 28411:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 28412:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 28413:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 28414:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 28415:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 28416:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 28417:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 28418:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 28419:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 28420:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 28421:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 28422:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 28423:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 28424:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 28425:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 28426:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 28427:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 28428:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 28429:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 28430:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 28431:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 28432:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 28433:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 28434:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 28435:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 28436:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 28437:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 28438:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 28439:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 28440:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 28441:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 28442:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 28443:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 28444:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 28445:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 28446:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 28447:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 28448:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 28449:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 28450:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 28451:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 28452:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 28453:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 28454:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 28455:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 28456:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 28457:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 28458:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 28459:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 28460:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 28461:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 28462:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 28463:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 28464:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 28465:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 28466:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 28467:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 28468:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 28469:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 28470:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 28471:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 28472:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 28473:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 28474:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 28475:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 28476:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 28477:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 28478:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 28479:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 28480:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 28481:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 28482:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 28483:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 28484:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 28485:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 28486:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 28487:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 28488:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 28489:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 28490:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 28491:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 28492:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 28493:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 28494:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 28495:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 28496:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 28497:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 28498:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 28499:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 28500:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 28501:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 28502:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 28503:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 28504:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 28505:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 28506:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 28507:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 28508:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 28509:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 28510:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 28511:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 28512:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 28513:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 28514:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 28515:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 28516:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 28517:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 28518:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 28519:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 28520:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 28521:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 28522:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 28523:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 28524:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 28525:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 28526:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 28527:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 28528:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 28529:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 28530:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 28531:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 28532:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 28533:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 28534:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 28535:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 28536:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 28537:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 28538:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 28539:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 28540:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 28541:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 28542:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 28543:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 28544:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 28545:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 28546:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 28547:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 28548:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 28549:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 28550:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 28551:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 28552:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 28553:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 28554:20]
  assign io_z = ~x38; // @[Snxn100k.scala 28555:16]
endmodule
module SnxnLv3Inst26(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst104_io_a; // @[Snxn100k.scala 7531:35]
  wire  inst_SnxnLv4Inst104_io_b; // @[Snxn100k.scala 7531:35]
  wire  inst_SnxnLv4Inst104_io_z; // @[Snxn100k.scala 7531:35]
  wire  inst_SnxnLv4Inst105_io_a; // @[Snxn100k.scala 7535:35]
  wire  inst_SnxnLv4Inst105_io_b; // @[Snxn100k.scala 7535:35]
  wire  inst_SnxnLv4Inst105_io_z; // @[Snxn100k.scala 7535:35]
  wire  inst_SnxnLv4Inst106_io_a; // @[Snxn100k.scala 7539:35]
  wire  inst_SnxnLv4Inst106_io_b; // @[Snxn100k.scala 7539:35]
  wire  inst_SnxnLv4Inst106_io_z; // @[Snxn100k.scala 7539:35]
  wire  inst_SnxnLv4Inst107_io_a; // @[Snxn100k.scala 7543:35]
  wire  inst_SnxnLv4Inst107_io_b; // @[Snxn100k.scala 7543:35]
  wire  inst_SnxnLv4Inst107_io_z; // @[Snxn100k.scala 7543:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst104_io_z + inst_SnxnLv4Inst105_io_z; // @[Snxn100k.scala 7547:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst106_io_z; // @[Snxn100k.scala 7547:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst107_io_z; // @[Snxn100k.scala 7547:92]
  SnxnLv4Inst104 inst_SnxnLv4Inst104 ( // @[Snxn100k.scala 7531:35]
    .io_a(inst_SnxnLv4Inst104_io_a),
    .io_b(inst_SnxnLv4Inst104_io_b),
    .io_z(inst_SnxnLv4Inst104_io_z)
  );
  SnxnLv4Inst105 inst_SnxnLv4Inst105 ( // @[Snxn100k.scala 7535:35]
    .io_a(inst_SnxnLv4Inst105_io_a),
    .io_b(inst_SnxnLv4Inst105_io_b),
    .io_z(inst_SnxnLv4Inst105_io_z)
  );
  SnxnLv4Inst106 inst_SnxnLv4Inst106 ( // @[Snxn100k.scala 7539:35]
    .io_a(inst_SnxnLv4Inst106_io_a),
    .io_b(inst_SnxnLv4Inst106_io_b),
    .io_z(inst_SnxnLv4Inst106_io_z)
  );
  SnxnLv4Inst107 inst_SnxnLv4Inst107 ( // @[Snxn100k.scala 7543:35]
    .io_a(inst_SnxnLv4Inst107_io_a),
    .io_b(inst_SnxnLv4Inst107_io_b),
    .io_z(inst_SnxnLv4Inst107_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7548:15]
  assign inst_SnxnLv4Inst104_io_a = io_a; // @[Snxn100k.scala 7532:28]
  assign inst_SnxnLv4Inst104_io_b = io_b; // @[Snxn100k.scala 7533:28]
  assign inst_SnxnLv4Inst105_io_a = io_a; // @[Snxn100k.scala 7536:28]
  assign inst_SnxnLv4Inst105_io_b = io_b; // @[Snxn100k.scala 7537:28]
  assign inst_SnxnLv4Inst106_io_a = io_a; // @[Snxn100k.scala 7540:28]
  assign inst_SnxnLv4Inst106_io_b = io_b; // @[Snxn100k.scala 7541:28]
  assign inst_SnxnLv4Inst107_io_a = io_a; // @[Snxn100k.scala 7544:28]
  assign inst_SnxnLv4Inst107_io_b = io_b; // @[Snxn100k.scala 7545:28]
endmodule
module SnxnLv4Inst110(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 29640:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 29641:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 29642:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 29643:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 29644:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 29645:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 29646:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 29647:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 29648:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 29649:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 29650:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 29651:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 29652:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 29653:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 29654:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 29655:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 29656:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 29657:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 29658:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 29659:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 29660:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 29661:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 29662:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 29663:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 29664:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 29665:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 29666:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 29667:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 29668:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 29669:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 29670:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 29671:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 29672:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 29673:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 29674:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 29675:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 29676:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 29677:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 29678:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 29679:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 29680:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 29681:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 29682:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 29683:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 29684:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 29685:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 29686:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 29687:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 29688:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 29689:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 29690:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 29691:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 29692:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 29693:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 29694:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 29695:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 29696:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 29697:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 29698:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 29699:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 29700:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 29701:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 29702:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 29703:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 29704:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 29705:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 29706:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 29707:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 29708:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 29709:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 29710:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 29711:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 29712:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 29713:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 29714:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 29715:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 29716:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 29717:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 29718:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 29719:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 29720:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 29721:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 29722:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 29723:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 29724:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 29725:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 29726:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 29727:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 29728:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 29729:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 29730:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 29731:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 29732:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 29733:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 29734:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 29735:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 29736:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 29737:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 29738:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 29739:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 29740:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 29741:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 29742:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 29743:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 29744:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 29745:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 29746:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 29747:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 29748:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 29749:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 29750:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 29751:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 29752:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 29753:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 29754:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 29755:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 29756:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 29757:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 29758:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 29759:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 29760:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 29761:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 29762:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 29763:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 29764:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 29765:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 29766:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 29767:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 29768:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 29769:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 29770:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 29771:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 29772:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 29773:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 29774:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 29775:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 29776:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 29777:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 29778:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 29779:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 29780:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 29781:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 29782:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 29783:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 29784:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 29785:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 29786:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 29787:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 29788:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 29789:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 29790:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 29791:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 29792:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 29793:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 29794:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 29795:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 29796:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 29797:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 29798:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 29799:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 29800:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 29801:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 29802:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 29803:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 29804:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 29805:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 29806:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 29807:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 29808:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 29809:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 29810:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 29811:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 29812:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 29813:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 29814:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 29815:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 29816:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 29817:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 29818:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 29819:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 29820:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 29821:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 29822:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 29823:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 29824:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 29825:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 29826:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 29827:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 29828:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 29829:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 29830:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 29831:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 29832:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 29833:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 29834:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 29835:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 29836:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 29837:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 29838:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 29839:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 29840:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 29841:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 29842:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 29843:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 29844:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 29845:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 29846:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 29847:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 29848:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 29849:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 29850:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 29851:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 29852:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 29853:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 29854:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 29855:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 29856:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 29857:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 29858:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 29859:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 29860:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 29861:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 29862:20]
  assign io_z = ~x55; // @[Snxn100k.scala 29863:16]
endmodule
module SnxnLv3Inst27(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst108_io_a; // @[Snxn100k.scala 7994:35]
  wire  inst_SnxnLv4Inst108_io_b; // @[Snxn100k.scala 7994:35]
  wire  inst_SnxnLv4Inst108_io_z; // @[Snxn100k.scala 7994:35]
  wire  inst_SnxnLv4Inst109_io_a; // @[Snxn100k.scala 7998:35]
  wire  inst_SnxnLv4Inst109_io_b; // @[Snxn100k.scala 7998:35]
  wire  inst_SnxnLv4Inst109_io_z; // @[Snxn100k.scala 7998:35]
  wire  inst_SnxnLv4Inst110_io_a; // @[Snxn100k.scala 8002:35]
  wire  inst_SnxnLv4Inst110_io_b; // @[Snxn100k.scala 8002:35]
  wire  inst_SnxnLv4Inst110_io_z; // @[Snxn100k.scala 8002:35]
  wire  inst_SnxnLv4Inst111_io_a; // @[Snxn100k.scala 8006:35]
  wire  inst_SnxnLv4Inst111_io_b; // @[Snxn100k.scala 8006:35]
  wire  inst_SnxnLv4Inst111_io_z; // @[Snxn100k.scala 8006:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst108_io_z + inst_SnxnLv4Inst109_io_z; // @[Snxn100k.scala 8010:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst110_io_z; // @[Snxn100k.scala 8010:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst111_io_z; // @[Snxn100k.scala 8010:92]
  SnxnLv4Inst0 inst_SnxnLv4Inst108 ( // @[Snxn100k.scala 7994:35]
    .io_a(inst_SnxnLv4Inst108_io_a),
    .io_b(inst_SnxnLv4Inst108_io_b),
    .io_z(inst_SnxnLv4Inst108_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst109 ( // @[Snxn100k.scala 7998:35]
    .io_a(inst_SnxnLv4Inst109_io_a),
    .io_b(inst_SnxnLv4Inst109_io_b),
    .io_z(inst_SnxnLv4Inst109_io_z)
  );
  SnxnLv4Inst110 inst_SnxnLv4Inst110 ( // @[Snxn100k.scala 8002:35]
    .io_a(inst_SnxnLv4Inst110_io_a),
    .io_b(inst_SnxnLv4Inst110_io_b),
    .io_z(inst_SnxnLv4Inst110_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst111 ( // @[Snxn100k.scala 8006:35]
    .io_a(inst_SnxnLv4Inst111_io_a),
    .io_b(inst_SnxnLv4Inst111_io_b),
    .io_z(inst_SnxnLv4Inst111_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 8011:15]
  assign inst_SnxnLv4Inst108_io_a = io_a; // @[Snxn100k.scala 7995:28]
  assign inst_SnxnLv4Inst108_io_b = io_b; // @[Snxn100k.scala 7996:28]
  assign inst_SnxnLv4Inst109_io_a = io_a; // @[Snxn100k.scala 7999:28]
  assign inst_SnxnLv4Inst109_io_b = io_b; // @[Snxn100k.scala 8000:28]
  assign inst_SnxnLv4Inst110_io_a = io_a; // @[Snxn100k.scala 8003:28]
  assign inst_SnxnLv4Inst110_io_b = io_b; // @[Snxn100k.scala 8004:28]
  assign inst_SnxnLv4Inst111_io_a = io_a; // @[Snxn100k.scala 8007:28]
  assign inst_SnxnLv4Inst111_io_b = io_b; // @[Snxn100k.scala 8008:28]
endmodule
module SnxnLv2Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst24_io_a; // @[Snxn100k.scala 1488:34]
  wire  inst_SnxnLv3Inst24_io_b; // @[Snxn100k.scala 1488:34]
  wire  inst_SnxnLv3Inst24_io_z; // @[Snxn100k.scala 1488:34]
  wire  inst_SnxnLv3Inst25_io_a; // @[Snxn100k.scala 1492:34]
  wire  inst_SnxnLv3Inst25_io_b; // @[Snxn100k.scala 1492:34]
  wire  inst_SnxnLv3Inst25_io_z; // @[Snxn100k.scala 1492:34]
  wire  inst_SnxnLv3Inst26_io_a; // @[Snxn100k.scala 1496:34]
  wire  inst_SnxnLv3Inst26_io_b; // @[Snxn100k.scala 1496:34]
  wire  inst_SnxnLv3Inst26_io_z; // @[Snxn100k.scala 1496:34]
  wire  inst_SnxnLv3Inst27_io_a; // @[Snxn100k.scala 1500:34]
  wire  inst_SnxnLv3Inst27_io_b; // @[Snxn100k.scala 1500:34]
  wire  inst_SnxnLv3Inst27_io_z; // @[Snxn100k.scala 1500:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst24_io_z + inst_SnxnLv3Inst25_io_z; // @[Snxn100k.scala 1504:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst26_io_z; // @[Snxn100k.scala 1504:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst27_io_z; // @[Snxn100k.scala 1504:89]
  SnxnLv3Inst24 inst_SnxnLv3Inst24 ( // @[Snxn100k.scala 1488:34]
    .io_a(inst_SnxnLv3Inst24_io_a),
    .io_b(inst_SnxnLv3Inst24_io_b),
    .io_z(inst_SnxnLv3Inst24_io_z)
  );
  SnxnLv3Inst25 inst_SnxnLv3Inst25 ( // @[Snxn100k.scala 1492:34]
    .io_a(inst_SnxnLv3Inst25_io_a),
    .io_b(inst_SnxnLv3Inst25_io_b),
    .io_z(inst_SnxnLv3Inst25_io_z)
  );
  SnxnLv3Inst26 inst_SnxnLv3Inst26 ( // @[Snxn100k.scala 1496:34]
    .io_a(inst_SnxnLv3Inst26_io_a),
    .io_b(inst_SnxnLv3Inst26_io_b),
    .io_z(inst_SnxnLv3Inst26_io_z)
  );
  SnxnLv3Inst27 inst_SnxnLv3Inst27 ( // @[Snxn100k.scala 1500:34]
    .io_a(inst_SnxnLv3Inst27_io_a),
    .io_b(inst_SnxnLv3Inst27_io_b),
    .io_z(inst_SnxnLv3Inst27_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1505:15]
  assign inst_SnxnLv3Inst24_io_a = io_a; // @[Snxn100k.scala 1489:27]
  assign inst_SnxnLv3Inst24_io_b = io_b; // @[Snxn100k.scala 1490:27]
  assign inst_SnxnLv3Inst25_io_a = io_a; // @[Snxn100k.scala 1493:27]
  assign inst_SnxnLv3Inst25_io_b = io_b; // @[Snxn100k.scala 1494:27]
  assign inst_SnxnLv3Inst26_io_a = io_a; // @[Snxn100k.scala 1497:27]
  assign inst_SnxnLv3Inst26_io_b = io_b; // @[Snxn100k.scala 1498:27]
  assign inst_SnxnLv3Inst27_io_a = io_a; // @[Snxn100k.scala 1501:27]
  assign inst_SnxnLv3Inst27_io_b = io_b; // @[Snxn100k.scala 1502:27]
endmodule
module SnxnLv4Inst113(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 43182:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 43183:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 43184:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 43185:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 43186:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 43187:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 43188:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 43189:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 43190:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 43191:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 43192:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 43193:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 43194:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 43195:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 43196:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 43197:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 43198:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 43199:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 43200:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 43201:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 43202:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 43203:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 43204:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 43205:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 43206:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 43207:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 43208:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 43209:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 43210:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 43211:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 43212:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 43213:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 43214:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 43215:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 43216:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 43217:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 43218:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 43219:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 43220:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 43221:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 43222:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 43223:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 43224:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 43225:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 43226:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 43227:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 43228:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 43229:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 43230:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 43231:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 43232:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 43233:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 43234:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 43235:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 43236:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 43237:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 43238:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 43239:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 43240:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 43241:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 43242:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 43243:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 43244:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 43245:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 43246:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 43247:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 43248:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 43249:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 43250:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 43251:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 43252:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 43253:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 43254:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 43255:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 43256:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 43257:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 43258:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 43259:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 43260:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 43261:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 43262:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 43263:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 43264:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 43265:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 43266:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 43267:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 43268:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 43269:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 43270:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 43271:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 43272:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 43273:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 43274:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 43275:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 43276:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 43277:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 43278:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 43279:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 43280:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 43281:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 43282:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 43283:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 43284:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 43285:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 43286:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 43287:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 43288:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 43289:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 43290:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 43291:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 43292:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 43293:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 43294:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 43295:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 43296:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 43297:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 43298:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 43299:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 43300:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 43301:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 43302:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 43303:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 43304:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 43305:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 43306:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 43307:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 43308:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 43309:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 43310:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 43311:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 43312:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 43313:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 43314:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 43315:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 43316:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 43317:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 43318:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 43319:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 43320:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 43321:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 43322:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 43323:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 43324:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 43325:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 43326:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 43327:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 43328:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 43329:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 43330:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 43331:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 43332:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 43333:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 43334:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 43335:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 43336:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 43337:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 43338:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 43339:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 43340:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 43341:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 43342:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 43343:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 43344:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 43345:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 43346:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 43347:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 43348:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 43349:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 43350:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 43351:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 43352:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 43353:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 43354:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 43355:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 43356:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 43357:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 43358:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 43359:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 43360:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 43361:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 43362:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 43363:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 43364:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 43365:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 43366:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 43367:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 43368:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 43369:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 43370:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 43371:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 43372:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 43373:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 43374:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 43375:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 43376:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 43377:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 43378:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 43379:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 43380:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 43381:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 43382:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 43383:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 43384:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 43385:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 43386:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 43387:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 43388:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 43389:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 43390:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 43391:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 43392:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 43393:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 43394:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 43395:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 43396:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 43397:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 43398:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 43399:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 43400:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 43401:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 43402:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 43403:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 43404:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 43405:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 43406:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 43407:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 43408:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 43409:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 43410:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 43411:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 43412:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 43413:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 43414:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 43415:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 43416:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 43417:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 43418:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 43419:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 43420:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 43421:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 43422:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 43423:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 43424:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 43425:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 43426:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 43427:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 43428:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 43429:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 43430:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 43431:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 43432:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 43433:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 43434:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 43435:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 43436:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 43437:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 43438:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 43439:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 43440:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 43441:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 43442:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 43443:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 43444:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 43445:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 43446:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 43447:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 43448:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 43449:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 43450:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 43451:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 43452:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 43453:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 43454:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 43455:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 43456:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 43457:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 43458:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 43459:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 43460:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 43461:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 43462:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 43463:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 43464:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 43465:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 43466:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 43467:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 43468:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 43469:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 43470:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 43471:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 43472:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 43473:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 43474:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 43475:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 43476:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 43477:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 43478:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 43479:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 43480:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 43481:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 43482:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 43483:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 43484:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 43485:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 43486:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 43487:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 43488:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 43489:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 43490:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 43491:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 43492:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 43493:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 43494:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 43495:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 43496:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 43497:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 43498:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 43499:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 43500:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 43501:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 43502:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 43503:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 43504:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 43505:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 43506:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 43507:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 43508:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 43509:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 43510:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 43511:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 43512:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 43513:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 43514:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 43515:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 43516:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 43517:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 43518:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 43519:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 43520:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 43521:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 43522:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 43523:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 43524:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 43525:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 43526:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 43527:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 43528:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 43529:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 43530:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 43531:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 43532:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 43533:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 43534:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 43535:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 43536:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 43537:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 43538:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 43539:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 43540:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 43541:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 43542:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 43543:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 43544:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 43545:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 43546:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 43547:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 43548:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 43549:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 43550:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 43551:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 43552:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 43553:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 43554:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 43555:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 43556:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 43557:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 43558:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 43559:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 43560:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 43561:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 43562:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 43563:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 43564:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 43565:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 43566:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 43567:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 43568:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 43569:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 43570:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 43571:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 43572:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 43573:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 43574:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 43575:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 43576:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 43577:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 43578:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 43579:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 43580:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 43581:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 43582:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 43583:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 43584:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 43585:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 43586:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 43587:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 43588:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 43589:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 43590:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 43591:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 43592:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 43593:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 43594:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 43595:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 43596:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 43597:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 43598:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 43599:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 43600:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 43601:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 43602:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 43603:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 43604:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 43605:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 43606:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 43607:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 43608:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 43609:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 43610:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 43611:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 43612:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 43613:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 43614:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 43615:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 43616:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 43617:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 43618:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 43619:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 43620:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 43621:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 43622:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 43623:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 43624:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 43625:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 43626:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 43627:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 43628:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 43629:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 43630:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 43631:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 43632:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 43633:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 43634:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 43635:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 43636:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 43637:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 43638:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 43639:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 43640:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 43641:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 43642:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 43643:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 43644:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 43645:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 43646:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 43647:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 43648:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 43649:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 43650:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 43651:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 43652:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 43653:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 43654:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 43655:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 43656:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 43657:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 43658:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 43659:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 43660:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 43661:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 43662:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 43663:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 43664:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 43665:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 43666:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 43667:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 43668:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 43669:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 43670:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 43671:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 43672:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 43673:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 43674:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 43675:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 43676:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 43677:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 43678:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 43679:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 43680:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 43681:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 43682:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 43683:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 43684:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 43685:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 43686:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 43687:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 43688:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 43689:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 43690:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 43691:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 43692:22]
  assign io_z = ~x127; // @[Snxn100k.scala 43693:17]
endmodule
module SnxnLv4Inst115(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 42804:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 42805:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 42806:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 42807:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 42808:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 42809:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 42810:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 42811:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 42812:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 42813:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 42814:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 42815:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 42816:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 42817:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 42818:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 42819:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 42820:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 42821:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 42822:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 42823:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 42824:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 42825:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 42826:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 42827:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 42828:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 42829:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 42830:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 42831:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 42832:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 42833:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 42834:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 42835:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 42836:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 42837:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 42838:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 42839:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 42840:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 42841:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 42842:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 42843:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 42844:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 42845:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 42846:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 42847:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 42848:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 42849:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 42850:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 42851:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 42852:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 42853:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 42854:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 42855:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 42856:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 42857:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 42858:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 42859:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 42860:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 42861:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 42862:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 42863:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 42864:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 42865:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 42866:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 42867:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 42868:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 42869:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 42870:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 42871:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 42872:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 42873:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 42874:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 42875:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 42876:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 42877:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 42878:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 42879:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 42880:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 42881:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 42882:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 42883:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 42884:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 42885:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 42886:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 42887:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 42888:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 42889:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 42890:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 42891:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 42892:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 42893:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 42894:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 42895:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 42896:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 42897:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 42898:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 42899:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 42900:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 42901:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 42902:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 42903:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 42904:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 42905:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 42906:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 42907:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 42908:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 42909:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 42910:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 42911:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 42912:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 42913:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 42914:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 42915:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 42916:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 42917:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 42918:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 42919:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 42920:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 42921:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 42922:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 42923:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 42924:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 42925:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 42926:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 42927:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 42928:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 42929:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 42930:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 42931:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 42932:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 42933:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 42934:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 42935:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 42936:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 42937:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 42938:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 42939:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 42940:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 42941:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 42942:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 42943:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 42944:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 42945:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 42946:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 42947:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 42948:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 42949:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 42950:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 42951:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 42952:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 42953:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 42954:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 42955:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 42956:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 42957:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 42958:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 42959:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 42960:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 42961:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 42962:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 42963:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 42964:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 42965:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 42966:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 42967:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 42968:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 42969:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 42970:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 42971:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 42972:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 42973:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 42974:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 42975:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 42976:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 42977:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 42978:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 42979:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 42980:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 42981:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 42982:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 42983:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 42984:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 42985:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 42986:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 42987:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 42988:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 42989:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 42990:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 42991:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 42992:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 42993:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 42994:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 42995:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 42996:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 42997:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 42998:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 42999:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 43000:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 43001:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 43002:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 43003:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 43004:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 43005:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 43006:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 43007:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 43008:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 43009:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 43010:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 43011:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 43012:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 43013:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 43014:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 43015:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 43016:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 43017:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 43018:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 43019:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 43020:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 43021:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 43022:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 43023:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 43024:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 43025:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 43026:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 43027:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 43028:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 43029:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 43030:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 43031:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 43032:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 43033:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 43034:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 43035:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 43036:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 43037:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 43038:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 43039:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 43040:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 43041:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 43042:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 43043:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 43044:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 43045:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 43046:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 43047:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 43048:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 43049:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 43050:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 43051:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 43052:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 43053:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 43054:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 43055:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 43056:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 43057:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 43058:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 43059:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 43060:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 43061:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 43062:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 43063:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 43064:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 43065:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 43066:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 43067:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 43068:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 43069:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 43070:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 43071:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 43072:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 43073:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 43074:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 43075:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 43076:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 43077:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 43078:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 43079:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 43080:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 43081:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 43082:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 43083:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 43084:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 43085:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 43086:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 43087:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 43088:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 43089:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 43090:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 43091:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 43092:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 43093:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 43094:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 43095:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 43096:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 43097:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 43098:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 43099:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 43100:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 43101:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 43102:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 43103:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 43104:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 43105:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 43106:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 43107:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 43108:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 43109:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 43110:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 43111:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 43112:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 43113:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 43114:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 43115:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 43116:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 43117:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 43118:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 43119:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 43120:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 43121:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 43122:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 43123:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 43124:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 43125:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 43126:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 43127:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 43128:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 43129:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 43130:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 43131:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 43132:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 43133:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 43134:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 43135:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 43136:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 43137:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 43138:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 43139:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 43140:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 43141:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 43142:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 43143:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 43144:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 43145:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 43146:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 43147:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 43148:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 43149:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 43150:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 43151:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 43152:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 43153:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 43154:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 43155:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 43156:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 43157:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 43158:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 43159:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 43160:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 43161:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 43162:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 43163:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 43164:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 43165:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 43166:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 43167:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 43168:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 43169:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 43170:20]
  assign io_z = ~x91; // @[Snxn100k.scala 43171:16]
endmodule
module SnxnLv3Inst28(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst112_io_a; // @[Snxn100k.scala 11584:35]
  wire  inst_SnxnLv4Inst112_io_b; // @[Snxn100k.scala 11584:35]
  wire  inst_SnxnLv4Inst112_io_z; // @[Snxn100k.scala 11584:35]
  wire  inst_SnxnLv4Inst113_io_a; // @[Snxn100k.scala 11588:35]
  wire  inst_SnxnLv4Inst113_io_b; // @[Snxn100k.scala 11588:35]
  wire  inst_SnxnLv4Inst113_io_z; // @[Snxn100k.scala 11588:35]
  wire  inst_SnxnLv4Inst114_io_a; // @[Snxn100k.scala 11592:35]
  wire  inst_SnxnLv4Inst114_io_b; // @[Snxn100k.scala 11592:35]
  wire  inst_SnxnLv4Inst114_io_z; // @[Snxn100k.scala 11592:35]
  wire  inst_SnxnLv4Inst115_io_a; // @[Snxn100k.scala 11596:35]
  wire  inst_SnxnLv4Inst115_io_b; // @[Snxn100k.scala 11596:35]
  wire  inst_SnxnLv4Inst115_io_z; // @[Snxn100k.scala 11596:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst112_io_z + inst_SnxnLv4Inst113_io_z; // @[Snxn100k.scala 11600:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst114_io_z; // @[Snxn100k.scala 11600:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst115_io_z; // @[Snxn100k.scala 11600:92]
  SnxnLv4Inst12 inst_SnxnLv4Inst112 ( // @[Snxn100k.scala 11584:35]
    .io_a(inst_SnxnLv4Inst112_io_a),
    .io_b(inst_SnxnLv4Inst112_io_b),
    .io_z(inst_SnxnLv4Inst112_io_z)
  );
  SnxnLv4Inst113 inst_SnxnLv4Inst113 ( // @[Snxn100k.scala 11588:35]
    .io_a(inst_SnxnLv4Inst113_io_a),
    .io_b(inst_SnxnLv4Inst113_io_b),
    .io_z(inst_SnxnLv4Inst113_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst114 ( // @[Snxn100k.scala 11592:35]
    .io_a(inst_SnxnLv4Inst114_io_a),
    .io_b(inst_SnxnLv4Inst114_io_b),
    .io_z(inst_SnxnLv4Inst114_io_z)
  );
  SnxnLv4Inst115 inst_SnxnLv4Inst115 ( // @[Snxn100k.scala 11596:35]
    .io_a(inst_SnxnLv4Inst115_io_a),
    .io_b(inst_SnxnLv4Inst115_io_b),
    .io_z(inst_SnxnLv4Inst115_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11601:15]
  assign inst_SnxnLv4Inst112_io_a = io_a; // @[Snxn100k.scala 11585:28]
  assign inst_SnxnLv4Inst112_io_b = io_b; // @[Snxn100k.scala 11586:28]
  assign inst_SnxnLv4Inst113_io_a = io_a; // @[Snxn100k.scala 11589:28]
  assign inst_SnxnLv4Inst113_io_b = io_b; // @[Snxn100k.scala 11590:28]
  assign inst_SnxnLv4Inst114_io_a = io_a; // @[Snxn100k.scala 11593:28]
  assign inst_SnxnLv4Inst114_io_b = io_b; // @[Snxn100k.scala 11594:28]
  assign inst_SnxnLv4Inst115_io_a = io_a; // @[Snxn100k.scala 11597:28]
  assign inst_SnxnLv4Inst115_io_b = io_b; // @[Snxn100k.scala 11598:28]
endmodule
module SnxnLv4Inst117(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 44792:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 44793:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 44794:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 44795:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 44796:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 44797:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 44798:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 44799:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 44800:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 44801:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 44802:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 44803:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 44804:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 44805:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 44806:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 44807:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 44808:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 44809:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 44810:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 44811:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 44812:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 44813:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 44814:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 44815:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 44816:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 44817:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 44818:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 44819:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 44820:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 44821:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 44822:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 44823:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 44824:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 44825:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 44826:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 44827:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 44828:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 44829:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 44830:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 44831:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 44832:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 44833:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 44834:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 44835:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 44836:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 44837:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 44838:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 44839:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 44840:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 44841:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 44842:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 44843:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 44844:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 44845:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 44846:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 44847:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 44848:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 44849:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 44850:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 44851:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 44852:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 44853:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 44854:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 44855:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 44856:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 44857:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 44858:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 44859:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 44860:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 44861:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 44862:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 44863:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 44864:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 44865:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 44866:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 44867:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 44868:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 44869:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 44870:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 44871:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 44872:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 44873:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 44874:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 44875:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 44876:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 44877:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 44878:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 44879:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 44880:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 44881:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 44882:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 44883:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 44884:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 44885:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 44886:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 44887:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 44888:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 44889:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 44890:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 44891:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 44892:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 44893:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 44894:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 44895:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 44896:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 44897:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 44898:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 44899:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 44900:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 44901:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 44902:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 44903:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 44904:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 44905:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 44906:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 44907:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 44908:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 44909:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 44910:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 44911:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 44912:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 44913:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 44914:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 44915:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 44916:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 44917:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 44918:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 44919:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 44920:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 44921:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 44922:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 44923:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 44924:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 44925:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 44926:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 44927:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 44928:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 44929:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 44930:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 44931:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 44932:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 44933:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 44934:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 44935:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 44936:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 44937:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 44938:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 44939:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 44940:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 44941:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 44942:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 44943:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 44944:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 44945:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 44946:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 44947:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 44948:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 44949:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 44950:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 44951:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 44952:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 44953:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 44954:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 44955:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 44956:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 44957:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 44958:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 44959:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 44960:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 44961:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 44962:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 44963:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 44964:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 44965:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 44966:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 44967:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 44968:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 44969:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 44970:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 44971:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 44972:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 44973:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 44974:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 44975:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 44976:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 44977:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 44978:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 44979:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 44980:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 44981:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 44982:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 44983:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 44984:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 44985:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 44986:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 44987:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 44988:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 44989:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 44990:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 44991:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 44992:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 44993:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 44994:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 44995:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 44996:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 44997:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 44998:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 44999:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 45000:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 45001:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 45002:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 45003:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 45004:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 45005:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 45006:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 45007:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 45008:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 45009:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 45010:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 45011:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 45012:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 45013:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 45014:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 45015:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 45016:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 45017:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 45018:20]
  assign io_z = ~x56; // @[Snxn100k.scala 45019:16]
endmodule
module SnxnLv4Inst118(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 45642:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 45643:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 45644:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 45645:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 45646:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 45647:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 45648:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 45649:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 45650:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 45651:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 45652:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 45653:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 45654:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 45655:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 45656:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 45657:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 45658:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 45659:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 45660:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 45661:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 45662:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 45663:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 45664:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 45665:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 45666:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 45667:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 45668:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 45669:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 45670:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 45671:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 45672:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 45673:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 45674:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 45675:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 45676:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 45677:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 45678:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 45679:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 45680:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 45681:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 45682:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 45683:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 45684:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 45685:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 45686:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 45687:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 45688:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 45689:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 45690:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 45691:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 45692:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 45693:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 45694:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 45695:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 45696:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 45697:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 45698:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 45699:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 45700:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 45701:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 45702:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 45703:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 45704:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 45705:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 45706:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 45707:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 45708:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 45709:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 45710:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 45711:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 45712:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 45713:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 45714:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 45715:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 45716:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 45717:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 45718:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 45719:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 45720:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 45721:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 45722:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 45723:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 45724:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 45725:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 45726:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 45727:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 45728:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 45729:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 45730:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 45731:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 45732:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 45733:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 45734:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 45735:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 45736:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 45737:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 45738:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 45739:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 45740:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 45741:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 45742:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 45743:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 45744:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 45745:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 45746:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 45747:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 45748:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 45749:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 45750:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 45751:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 45752:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 45753:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 45754:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 45755:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 45756:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 45757:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 45758:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 45759:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 45760:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 45761:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 45762:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 45763:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 45764:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 45765:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 45766:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 45767:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 45768:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 45769:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 45770:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 45771:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 45772:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 45773:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 45774:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 45775:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 45776:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 45777:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 45778:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 45779:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 45780:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 45781:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 45782:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 45783:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 45784:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 45785:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 45786:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 45787:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 45788:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 45789:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 45790:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 45791:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 45792:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 45793:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 45794:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 45795:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 45796:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 45797:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 45798:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 45799:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 45800:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 45801:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 45802:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 45803:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 45804:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 45805:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 45806:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 45807:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 45808:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 45809:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 45810:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 45811:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 45812:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 45813:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 45814:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 45815:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 45816:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 45817:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 45818:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 45819:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 45820:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 45821:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 45822:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 45823:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 45824:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 45825:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 45826:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 45827:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 45828:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 45829:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 45830:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 45831:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 45832:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 45833:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 45834:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 45835:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 45836:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 45837:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 45838:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 45839:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 45840:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 45841:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 45842:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 45843:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 45844:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 45845:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 45846:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 45847:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 45848:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 45849:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 45850:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 45851:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 45852:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 45853:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 45854:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 45855:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 45856:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 45857:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 45858:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 45859:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 45860:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 45861:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 45862:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 45863:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 45864:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 45865:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 45866:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 45867:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 45868:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 45869:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 45870:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 45871:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 45872:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 45873:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 45874:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 45875:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 45876:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 45877:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 45878:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 45879:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 45880:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 45881:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 45882:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 45883:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 45884:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 45885:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 45886:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 45887:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 45888:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 45889:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 45890:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 45891:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 45892:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 45893:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 45894:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 45895:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 45896:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 45897:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 45898:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 45899:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 45900:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 45901:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 45902:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 45903:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 45904:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 45905:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 45906:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 45907:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 45908:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 45909:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 45910:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 45911:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 45912:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 45913:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 45914:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 45915:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 45916:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 45917:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 45918:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 45919:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 45920:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 45921:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 45922:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 45923:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 45924:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 45925:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 45926:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 45927:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 45928:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 45929:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 45930:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 45931:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 45932:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 45933:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 45934:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 45935:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 45936:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 45937:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 45938:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 45939:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 45940:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 45941:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 45942:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 45943:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 45944:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 45945:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 45946:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 45947:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 45948:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 45949:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 45950:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 45951:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 45952:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 45953:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 45954:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 45955:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 45956:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 45957:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 45958:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 45959:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 45960:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 45961:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 45962:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 45963:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 45964:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 45965:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 45966:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 45967:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 45968:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 45969:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 45970:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 45971:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 45972:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 45973:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 45974:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 45975:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 45976:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 45977:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 45978:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 45979:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 45980:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 45981:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 45982:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 45983:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 45984:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 45985:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 45986:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 45987:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 45988:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 45989:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 45990:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 45991:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 45992:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 45993:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 45994:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 45995:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 45996:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 45997:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 45998:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 45999:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 46000:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 46001:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 46002:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 46003:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 46004:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 46005:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 46006:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 46007:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 46008:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 46009:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 46010:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 46011:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 46012:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 46013:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 46014:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 46015:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 46016:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 46017:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 46018:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 46019:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 46020:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 46021:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 46022:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 46023:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 46024:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 46025:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 46026:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 46027:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 46028:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 46029:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 46030:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 46031:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 46032:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 46033:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 46034:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 46035:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 46036:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 46037:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 46038:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 46039:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 46040:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 46041:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 46042:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 46043:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 46044:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 46045:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 46046:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 46047:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 46048:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 46049:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 46050:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 46051:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 46052:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 46053:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 46054:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 46055:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 46056:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 46057:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 46058:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 46059:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 46060:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 46061:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 46062:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 46063:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 46064:22]
  assign io_z = ~x105; // @[Snxn100k.scala 46065:17]
endmodule
module SnxnLv3Inst29(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst116_io_a; // @[Snxn100k.scala 12278:35]
  wire  inst_SnxnLv4Inst116_io_b; // @[Snxn100k.scala 12278:35]
  wire  inst_SnxnLv4Inst116_io_z; // @[Snxn100k.scala 12278:35]
  wire  inst_SnxnLv4Inst117_io_a; // @[Snxn100k.scala 12282:35]
  wire  inst_SnxnLv4Inst117_io_b; // @[Snxn100k.scala 12282:35]
  wire  inst_SnxnLv4Inst117_io_z; // @[Snxn100k.scala 12282:35]
  wire  inst_SnxnLv4Inst118_io_a; // @[Snxn100k.scala 12286:35]
  wire  inst_SnxnLv4Inst118_io_b; // @[Snxn100k.scala 12286:35]
  wire  inst_SnxnLv4Inst118_io_z; // @[Snxn100k.scala 12286:35]
  wire  inst_SnxnLv4Inst119_io_a; // @[Snxn100k.scala 12290:35]
  wire  inst_SnxnLv4Inst119_io_b; // @[Snxn100k.scala 12290:35]
  wire  inst_SnxnLv4Inst119_io_z; // @[Snxn100k.scala 12290:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst116_io_z + inst_SnxnLv4Inst117_io_z; // @[Snxn100k.scala 12294:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst118_io_z; // @[Snxn100k.scala 12294:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst119_io_z; // @[Snxn100k.scala 12294:92]
  SnxnLv4Inst50 inst_SnxnLv4Inst116 ( // @[Snxn100k.scala 12278:35]
    .io_a(inst_SnxnLv4Inst116_io_a),
    .io_b(inst_SnxnLv4Inst116_io_b),
    .io_z(inst_SnxnLv4Inst116_io_z)
  );
  SnxnLv4Inst117 inst_SnxnLv4Inst117 ( // @[Snxn100k.scala 12282:35]
    .io_a(inst_SnxnLv4Inst117_io_a),
    .io_b(inst_SnxnLv4Inst117_io_b),
    .io_z(inst_SnxnLv4Inst117_io_z)
  );
  SnxnLv4Inst118 inst_SnxnLv4Inst118 ( // @[Snxn100k.scala 12286:35]
    .io_a(inst_SnxnLv4Inst118_io_a),
    .io_b(inst_SnxnLv4Inst118_io_b),
    .io_z(inst_SnxnLv4Inst118_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst119 ( // @[Snxn100k.scala 12290:35]
    .io_a(inst_SnxnLv4Inst119_io_a),
    .io_b(inst_SnxnLv4Inst119_io_b),
    .io_z(inst_SnxnLv4Inst119_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 12295:15]
  assign inst_SnxnLv4Inst116_io_a = io_a; // @[Snxn100k.scala 12279:28]
  assign inst_SnxnLv4Inst116_io_b = io_b; // @[Snxn100k.scala 12280:28]
  assign inst_SnxnLv4Inst117_io_a = io_a; // @[Snxn100k.scala 12283:28]
  assign inst_SnxnLv4Inst117_io_b = io_b; // @[Snxn100k.scala 12284:28]
  assign inst_SnxnLv4Inst118_io_a = io_a; // @[Snxn100k.scala 12287:28]
  assign inst_SnxnLv4Inst118_io_b = io_b; // @[Snxn100k.scala 12288:28]
  assign inst_SnxnLv4Inst119_io_a = io_a; // @[Snxn100k.scala 12291:28]
  assign inst_SnxnLv4Inst119_io_b = io_b; // @[Snxn100k.scala 12292:28]
endmodule
module SnxnLv4Inst123(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 43704:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 43705:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 43706:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 43707:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 43708:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 43709:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 43710:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 43711:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 43712:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 43713:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 43714:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 43715:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 43716:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 43717:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 43718:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 43719:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 43720:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 43721:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 43722:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 43723:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 43724:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 43725:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 43726:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 43727:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 43728:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 43729:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 43730:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 43731:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 43732:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 43733:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 43734:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 43735:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 43736:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 43737:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 43738:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 43739:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 43740:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 43741:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 43742:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 43743:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 43744:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 43745:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 43746:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 43747:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 43748:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 43749:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 43750:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 43751:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 43752:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 43753:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 43754:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 43755:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 43756:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 43757:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 43758:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 43759:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 43760:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 43761:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 43762:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 43763:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 43764:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 43765:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 43766:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 43767:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 43768:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 43769:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 43770:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 43771:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 43772:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 43773:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 43774:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 43775:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 43776:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 43777:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 43778:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 43779:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 43780:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 43781:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 43782:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 43783:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 43784:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 43785:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 43786:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 43787:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 43788:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 43789:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 43790:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 43791:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 43792:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 43793:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 43794:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 43795:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 43796:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 43797:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 43798:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 43799:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 43800:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 43801:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 43802:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 43803:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 43804:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 43805:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 43806:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 43807:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 43808:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 43809:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 43810:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 43811:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 43812:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 43813:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 43814:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 43815:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 43816:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 43817:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 43818:20]
  assign io_z = ~x28; // @[Snxn100k.scala 43819:16]
endmodule
module SnxnLv3Inst30(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst120_io_a; // @[Snxn100k.scala 11887:35]
  wire  inst_SnxnLv4Inst120_io_b; // @[Snxn100k.scala 11887:35]
  wire  inst_SnxnLv4Inst120_io_z; // @[Snxn100k.scala 11887:35]
  wire  inst_SnxnLv4Inst121_io_a; // @[Snxn100k.scala 11891:35]
  wire  inst_SnxnLv4Inst121_io_b; // @[Snxn100k.scala 11891:35]
  wire  inst_SnxnLv4Inst121_io_z; // @[Snxn100k.scala 11891:35]
  wire  inst_SnxnLv4Inst122_io_a; // @[Snxn100k.scala 11895:35]
  wire  inst_SnxnLv4Inst122_io_b; // @[Snxn100k.scala 11895:35]
  wire  inst_SnxnLv4Inst122_io_z; // @[Snxn100k.scala 11895:35]
  wire  inst_SnxnLv4Inst123_io_a; // @[Snxn100k.scala 11899:35]
  wire  inst_SnxnLv4Inst123_io_b; // @[Snxn100k.scala 11899:35]
  wire  inst_SnxnLv4Inst123_io_z; // @[Snxn100k.scala 11899:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst120_io_z + inst_SnxnLv4Inst121_io_z; // @[Snxn100k.scala 11903:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst122_io_z; // @[Snxn100k.scala 11903:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst123_io_z; // @[Snxn100k.scala 11903:92]
  SnxnLv4Inst52 inst_SnxnLv4Inst120 ( // @[Snxn100k.scala 11887:35]
    .io_a(inst_SnxnLv4Inst120_io_a),
    .io_b(inst_SnxnLv4Inst120_io_b),
    .io_z(inst_SnxnLv4Inst120_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst121 ( // @[Snxn100k.scala 11891:35]
    .io_a(inst_SnxnLv4Inst121_io_a),
    .io_b(inst_SnxnLv4Inst121_io_b),
    .io_z(inst_SnxnLv4Inst121_io_z)
  );
  SnxnLv4Inst12 inst_SnxnLv4Inst122 ( // @[Snxn100k.scala 11895:35]
    .io_a(inst_SnxnLv4Inst122_io_a),
    .io_b(inst_SnxnLv4Inst122_io_b),
    .io_z(inst_SnxnLv4Inst122_io_z)
  );
  SnxnLv4Inst123 inst_SnxnLv4Inst123 ( // @[Snxn100k.scala 11899:35]
    .io_a(inst_SnxnLv4Inst123_io_a),
    .io_b(inst_SnxnLv4Inst123_io_b),
    .io_z(inst_SnxnLv4Inst123_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11904:15]
  assign inst_SnxnLv4Inst120_io_a = io_a; // @[Snxn100k.scala 11888:28]
  assign inst_SnxnLv4Inst120_io_b = io_b; // @[Snxn100k.scala 11889:28]
  assign inst_SnxnLv4Inst121_io_a = io_a; // @[Snxn100k.scala 11892:28]
  assign inst_SnxnLv4Inst121_io_b = io_b; // @[Snxn100k.scala 11893:28]
  assign inst_SnxnLv4Inst122_io_a = io_a; // @[Snxn100k.scala 11896:28]
  assign inst_SnxnLv4Inst122_io_b = io_b; // @[Snxn100k.scala 11897:28]
  assign inst_SnxnLv4Inst123_io_a = io_a; // @[Snxn100k.scala 11900:28]
  assign inst_SnxnLv4Inst123_io_b = io_b; // @[Snxn100k.scala 11901:28]
endmodule
module SnxnLv3Inst31(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst124_io_a; // @[Snxn100k.scala 12765:35]
  wire  inst_SnxnLv4Inst124_io_b; // @[Snxn100k.scala 12765:35]
  wire  inst_SnxnLv4Inst124_io_z; // @[Snxn100k.scala 12765:35]
  wire  inst_SnxnLv4Inst125_io_a; // @[Snxn100k.scala 12769:35]
  wire  inst_SnxnLv4Inst125_io_b; // @[Snxn100k.scala 12769:35]
  wire  inst_SnxnLv4Inst125_io_z; // @[Snxn100k.scala 12769:35]
  wire  inst_SnxnLv4Inst126_io_a; // @[Snxn100k.scala 12773:35]
  wire  inst_SnxnLv4Inst126_io_b; // @[Snxn100k.scala 12773:35]
  wire  inst_SnxnLv4Inst126_io_z; // @[Snxn100k.scala 12773:35]
  wire  inst_SnxnLv4Inst127_io_a; // @[Snxn100k.scala 12777:35]
  wire  inst_SnxnLv4Inst127_io_b; // @[Snxn100k.scala 12777:35]
  wire  inst_SnxnLv4Inst127_io_z; // @[Snxn100k.scala 12777:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst124_io_z + inst_SnxnLv4Inst125_io_z; // @[Snxn100k.scala 12781:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst126_io_z; // @[Snxn100k.scala 12781:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst127_io_z; // @[Snxn100k.scala 12781:92]
  SnxnLv4Inst105 inst_SnxnLv4Inst124 ( // @[Snxn100k.scala 12765:35]
    .io_a(inst_SnxnLv4Inst124_io_a),
    .io_b(inst_SnxnLv4Inst124_io_b),
    .io_z(inst_SnxnLv4Inst124_io_z)
  );
  SnxnLv4Inst107 inst_SnxnLv4Inst125 ( // @[Snxn100k.scala 12769:35]
    .io_a(inst_SnxnLv4Inst125_io_a),
    .io_b(inst_SnxnLv4Inst125_io_b),
    .io_z(inst_SnxnLv4Inst125_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst126 ( // @[Snxn100k.scala 12773:35]
    .io_a(inst_SnxnLv4Inst126_io_a),
    .io_b(inst_SnxnLv4Inst126_io_b),
    .io_z(inst_SnxnLv4Inst126_io_z)
  );
  SnxnLv4Inst74 inst_SnxnLv4Inst127 ( // @[Snxn100k.scala 12777:35]
    .io_a(inst_SnxnLv4Inst127_io_a),
    .io_b(inst_SnxnLv4Inst127_io_b),
    .io_z(inst_SnxnLv4Inst127_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 12782:15]
  assign inst_SnxnLv4Inst124_io_a = io_a; // @[Snxn100k.scala 12766:28]
  assign inst_SnxnLv4Inst124_io_b = io_b; // @[Snxn100k.scala 12767:28]
  assign inst_SnxnLv4Inst125_io_a = io_a; // @[Snxn100k.scala 12770:28]
  assign inst_SnxnLv4Inst125_io_b = io_b; // @[Snxn100k.scala 12771:28]
  assign inst_SnxnLv4Inst126_io_a = io_a; // @[Snxn100k.scala 12774:28]
  assign inst_SnxnLv4Inst126_io_b = io_b; // @[Snxn100k.scala 12775:28]
  assign inst_SnxnLv4Inst127_io_a = io_a; // @[Snxn100k.scala 12778:28]
  assign inst_SnxnLv4Inst127_io_b = io_b; // @[Snxn100k.scala 12779:28]
endmodule
module SnxnLv2Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst28_io_a; // @[Snxn100k.scala 2785:34]
  wire  inst_SnxnLv3Inst28_io_b; // @[Snxn100k.scala 2785:34]
  wire  inst_SnxnLv3Inst28_io_z; // @[Snxn100k.scala 2785:34]
  wire  inst_SnxnLv3Inst29_io_a; // @[Snxn100k.scala 2789:34]
  wire  inst_SnxnLv3Inst29_io_b; // @[Snxn100k.scala 2789:34]
  wire  inst_SnxnLv3Inst29_io_z; // @[Snxn100k.scala 2789:34]
  wire  inst_SnxnLv3Inst30_io_a; // @[Snxn100k.scala 2793:34]
  wire  inst_SnxnLv3Inst30_io_b; // @[Snxn100k.scala 2793:34]
  wire  inst_SnxnLv3Inst30_io_z; // @[Snxn100k.scala 2793:34]
  wire  inst_SnxnLv3Inst31_io_a; // @[Snxn100k.scala 2797:34]
  wire  inst_SnxnLv3Inst31_io_b; // @[Snxn100k.scala 2797:34]
  wire  inst_SnxnLv3Inst31_io_z; // @[Snxn100k.scala 2797:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst28_io_z + inst_SnxnLv3Inst29_io_z; // @[Snxn100k.scala 2801:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst30_io_z; // @[Snxn100k.scala 2801:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst31_io_z; // @[Snxn100k.scala 2801:89]
  SnxnLv3Inst28 inst_SnxnLv3Inst28 ( // @[Snxn100k.scala 2785:34]
    .io_a(inst_SnxnLv3Inst28_io_a),
    .io_b(inst_SnxnLv3Inst28_io_b),
    .io_z(inst_SnxnLv3Inst28_io_z)
  );
  SnxnLv3Inst29 inst_SnxnLv3Inst29 ( // @[Snxn100k.scala 2789:34]
    .io_a(inst_SnxnLv3Inst29_io_a),
    .io_b(inst_SnxnLv3Inst29_io_b),
    .io_z(inst_SnxnLv3Inst29_io_z)
  );
  SnxnLv3Inst30 inst_SnxnLv3Inst30 ( // @[Snxn100k.scala 2793:34]
    .io_a(inst_SnxnLv3Inst30_io_a),
    .io_b(inst_SnxnLv3Inst30_io_b),
    .io_z(inst_SnxnLv3Inst30_io_z)
  );
  SnxnLv3Inst31 inst_SnxnLv3Inst31 ( // @[Snxn100k.scala 2797:34]
    .io_a(inst_SnxnLv3Inst31_io_a),
    .io_b(inst_SnxnLv3Inst31_io_b),
    .io_z(inst_SnxnLv3Inst31_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 2802:15]
  assign inst_SnxnLv3Inst28_io_a = io_a; // @[Snxn100k.scala 2786:27]
  assign inst_SnxnLv3Inst28_io_b = io_b; // @[Snxn100k.scala 2787:27]
  assign inst_SnxnLv3Inst29_io_a = io_a; // @[Snxn100k.scala 2790:27]
  assign inst_SnxnLv3Inst29_io_b = io_b; // @[Snxn100k.scala 2791:27]
  assign inst_SnxnLv3Inst30_io_a = io_a; // @[Snxn100k.scala 2794:27]
  assign inst_SnxnLv3Inst30_io_b = io_b; // @[Snxn100k.scala 2795:27]
  assign inst_SnxnLv3Inst31_io_a = io_a; // @[Snxn100k.scala 2798:27]
  assign inst_SnxnLv3Inst31_io_b = io_b; // @[Snxn100k.scala 2799:27]
endmodule
module SnxnLv1Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst4_io_a; // @[Snxn100k.scala 648:33]
  wire  inst_SnxnLv2Inst4_io_b; // @[Snxn100k.scala 648:33]
  wire  inst_SnxnLv2Inst4_io_z; // @[Snxn100k.scala 648:33]
  wire  inst_SnxnLv2Inst5_io_a; // @[Snxn100k.scala 652:33]
  wire  inst_SnxnLv2Inst5_io_b; // @[Snxn100k.scala 652:33]
  wire  inst_SnxnLv2Inst5_io_z; // @[Snxn100k.scala 652:33]
  wire  inst_SnxnLv2Inst6_io_a; // @[Snxn100k.scala 656:33]
  wire  inst_SnxnLv2Inst6_io_b; // @[Snxn100k.scala 656:33]
  wire  inst_SnxnLv2Inst6_io_z; // @[Snxn100k.scala 656:33]
  wire  inst_SnxnLv2Inst7_io_a; // @[Snxn100k.scala 660:33]
  wire  inst_SnxnLv2Inst7_io_b; // @[Snxn100k.scala 660:33]
  wire  inst_SnxnLv2Inst7_io_z; // @[Snxn100k.scala 660:33]
  wire  _sum_T_1 = inst_SnxnLv2Inst4_io_z + inst_SnxnLv2Inst5_io_z; // @[Snxn100k.scala 664:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst6_io_z; // @[Snxn100k.scala 664:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst7_io_z; // @[Snxn100k.scala 664:86]
  SnxnLv2Inst4 inst_SnxnLv2Inst4 ( // @[Snxn100k.scala 648:33]
    .io_a(inst_SnxnLv2Inst4_io_a),
    .io_b(inst_SnxnLv2Inst4_io_b),
    .io_z(inst_SnxnLv2Inst4_io_z)
  );
  SnxnLv2Inst5 inst_SnxnLv2Inst5 ( // @[Snxn100k.scala 652:33]
    .io_a(inst_SnxnLv2Inst5_io_a),
    .io_b(inst_SnxnLv2Inst5_io_b),
    .io_z(inst_SnxnLv2Inst5_io_z)
  );
  SnxnLv2Inst6 inst_SnxnLv2Inst6 ( // @[Snxn100k.scala 656:33]
    .io_a(inst_SnxnLv2Inst6_io_a),
    .io_b(inst_SnxnLv2Inst6_io_b),
    .io_z(inst_SnxnLv2Inst6_io_z)
  );
  SnxnLv2Inst7 inst_SnxnLv2Inst7 ( // @[Snxn100k.scala 660:33]
    .io_a(inst_SnxnLv2Inst7_io_a),
    .io_b(inst_SnxnLv2Inst7_io_b),
    .io_z(inst_SnxnLv2Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 665:15]
  assign inst_SnxnLv2Inst4_io_a = io_a; // @[Snxn100k.scala 649:26]
  assign inst_SnxnLv2Inst4_io_b = io_b; // @[Snxn100k.scala 650:26]
  assign inst_SnxnLv2Inst5_io_a = io_a; // @[Snxn100k.scala 653:26]
  assign inst_SnxnLv2Inst5_io_b = io_b; // @[Snxn100k.scala 654:26]
  assign inst_SnxnLv2Inst6_io_a = io_a; // @[Snxn100k.scala 657:26]
  assign inst_SnxnLv2Inst6_io_b = io_b; // @[Snxn100k.scala 658:26]
  assign inst_SnxnLv2Inst7_io_a = io_a; // @[Snxn100k.scala 661:26]
  assign inst_SnxnLv2Inst7_io_b = io_b; // @[Snxn100k.scala 662:26]
endmodule
module SnxnLv4Inst129(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 48752:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 48753:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 48754:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 48755:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 48756:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 48757:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 48758:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 48759:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 48760:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 48761:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 48762:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 48763:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 48764:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 48765:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 48766:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 48767:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 48768:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 48769:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 48770:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 48771:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 48772:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 48773:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 48774:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 48775:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 48776:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 48777:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 48778:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 48779:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 48780:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 48781:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 48782:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 48783:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 48784:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 48785:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 48786:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 48787:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 48788:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 48789:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 48790:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 48791:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 48792:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 48793:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 48794:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 48795:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 48796:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 48797:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 48798:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 48799:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 48800:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 48801:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 48802:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 48803:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 48804:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 48805:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 48806:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 48807:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 48808:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 48809:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 48810:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 48811:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 48812:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 48813:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 48814:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 48815:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 48816:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 48817:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 48818:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 48819:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 48820:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 48821:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 48822:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 48823:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 48824:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 48825:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 48826:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 48827:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 48828:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 48829:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 48830:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 48831:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 48832:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 48833:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 48834:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 48835:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 48836:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 48837:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 48838:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 48839:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 48840:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 48841:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 48842:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 48843:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 48844:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 48845:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 48846:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 48847:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 48848:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 48849:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 48850:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 48851:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 48852:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 48853:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 48854:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 48855:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 48856:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 48857:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 48858:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 48859:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 48860:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 48861:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 48862:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 48863:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 48864:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 48865:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 48866:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 48867:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 48868:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 48869:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 48870:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 48871:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 48872:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 48873:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 48874:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 48875:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 48876:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 48877:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 48878:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 48879:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 48880:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 48881:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 48882:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 48883:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 48884:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 48885:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 48886:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 48887:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 48888:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 48889:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 48890:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 48891:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 48892:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 48893:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 48894:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 48895:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 48896:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 48897:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 48898:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 48899:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 48900:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 48901:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 48902:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 48903:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 48904:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 48905:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 48906:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 48907:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 48908:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 48909:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 48910:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 48911:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 48912:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 48913:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 48914:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 48915:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 48916:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 48917:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 48918:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 48919:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 48920:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 48921:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 48922:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 48923:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 48924:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 48925:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 48926:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 48927:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 48928:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 48929:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 48930:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 48931:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 48932:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 48933:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 48934:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 48935:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 48936:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 48937:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 48938:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 48939:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 48940:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 48941:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 48942:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 48943:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 48944:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 48945:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 48946:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 48947:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 48948:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 48949:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 48950:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 48951:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 48952:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 48953:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 48954:20]
  assign io_z = ~x50; // @[Snxn100k.scala 48955:16]
endmodule
module SnxnLv3Inst32(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst128_io_a; // @[Snxn100k.scala 13287:35]
  wire  inst_SnxnLv4Inst128_io_b; // @[Snxn100k.scala 13287:35]
  wire  inst_SnxnLv4Inst128_io_z; // @[Snxn100k.scala 13287:35]
  wire  inst_SnxnLv4Inst129_io_a; // @[Snxn100k.scala 13291:35]
  wire  inst_SnxnLv4Inst129_io_b; // @[Snxn100k.scala 13291:35]
  wire  inst_SnxnLv4Inst129_io_z; // @[Snxn100k.scala 13291:35]
  wire  inst_SnxnLv4Inst130_io_a; // @[Snxn100k.scala 13295:35]
  wire  inst_SnxnLv4Inst130_io_b; // @[Snxn100k.scala 13295:35]
  wire  inst_SnxnLv4Inst130_io_z; // @[Snxn100k.scala 13295:35]
  wire  inst_SnxnLv4Inst131_io_a; // @[Snxn100k.scala 13299:35]
  wire  inst_SnxnLv4Inst131_io_b; // @[Snxn100k.scala 13299:35]
  wire  inst_SnxnLv4Inst131_io_z; // @[Snxn100k.scala 13299:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst128_io_z + inst_SnxnLv4Inst129_io_z; // @[Snxn100k.scala 13303:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst130_io_z; // @[Snxn100k.scala 13303:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst131_io_z; // @[Snxn100k.scala 13303:92]
  SnxnLv4Inst73 inst_SnxnLv4Inst128 ( // @[Snxn100k.scala 13287:35]
    .io_a(inst_SnxnLv4Inst128_io_a),
    .io_b(inst_SnxnLv4Inst128_io_b),
    .io_z(inst_SnxnLv4Inst128_io_z)
  );
  SnxnLv4Inst129 inst_SnxnLv4Inst129 ( // @[Snxn100k.scala 13291:35]
    .io_a(inst_SnxnLv4Inst129_io_a),
    .io_b(inst_SnxnLv4Inst129_io_b),
    .io_z(inst_SnxnLv4Inst129_io_z)
  );
  SnxnLv4Inst20 inst_SnxnLv4Inst130 ( // @[Snxn100k.scala 13295:35]
    .io_a(inst_SnxnLv4Inst130_io_a),
    .io_b(inst_SnxnLv4Inst130_io_b),
    .io_z(inst_SnxnLv4Inst130_io_z)
  );
  SnxnLv4Inst56 inst_SnxnLv4Inst131 ( // @[Snxn100k.scala 13299:35]
    .io_a(inst_SnxnLv4Inst131_io_a),
    .io_b(inst_SnxnLv4Inst131_io_b),
    .io_z(inst_SnxnLv4Inst131_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 13304:15]
  assign inst_SnxnLv4Inst128_io_a = io_a; // @[Snxn100k.scala 13288:28]
  assign inst_SnxnLv4Inst128_io_b = io_b; // @[Snxn100k.scala 13289:28]
  assign inst_SnxnLv4Inst129_io_a = io_a; // @[Snxn100k.scala 13292:28]
  assign inst_SnxnLv4Inst129_io_b = io_b; // @[Snxn100k.scala 13293:28]
  assign inst_SnxnLv4Inst130_io_a = io_a; // @[Snxn100k.scala 13296:28]
  assign inst_SnxnLv4Inst130_io_b = io_b; // @[Snxn100k.scala 13297:28]
  assign inst_SnxnLv4Inst131_io_a = io_a; // @[Snxn100k.scala 13300:28]
  assign inst_SnxnLv4Inst131_io_b = io_b; // @[Snxn100k.scala 13301:28]
endmodule
module SnxnLv4Inst135(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 47976:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 47977:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 47978:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 47979:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 47980:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 47981:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 47982:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 47983:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 47984:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 47985:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 47986:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 47987:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 47988:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 47989:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 47990:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 47991:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 47992:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 47993:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 47994:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 47995:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 47996:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 47997:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 47998:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 47999:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 48000:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 48001:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 48002:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 48003:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 48004:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 48005:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 48006:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 48007:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 48008:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 48009:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 48010:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 48011:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 48012:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 48013:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 48014:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 48015:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 48016:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 48017:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 48018:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 48019:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 48020:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 48021:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 48022:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 48023:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 48024:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 48025:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 48026:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 48027:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 48028:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 48029:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 48030:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 48031:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 48032:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 48033:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 48034:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 48035:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 48036:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 48037:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 48038:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 48039:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 48040:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 48041:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 48042:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 48043:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 48044:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 48045:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 48046:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 48047:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 48048:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 48049:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 48050:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 48051:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 48052:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 48053:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 48054:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 48055:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 48056:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 48057:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 48058:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 48059:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 48060:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 48061:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 48062:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 48063:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 48064:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 48065:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 48066:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 48067:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 48068:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 48069:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 48070:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 48071:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 48072:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 48073:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 48074:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 48075:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 48076:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 48077:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 48078:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 48079:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 48080:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 48081:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 48082:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 48083:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 48084:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 48085:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 48086:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 48087:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 48088:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 48089:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 48090:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 48091:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 48092:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 48093:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 48094:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 48095:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 48096:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 48097:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 48098:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 48099:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 48100:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 48101:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 48102:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 48103:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 48104:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 48105:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 48106:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 48107:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 48108:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 48109:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 48110:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 48111:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 48112:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 48113:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 48114:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 48115:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 48116:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 48117:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 48118:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 48119:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 48120:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 48121:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 48122:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 48123:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 48124:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 48125:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 48126:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 48127:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 48128:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 48129:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 48130:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 48131:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 48132:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 48133:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 48134:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 48135:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 48136:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 48137:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 48138:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 48139:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 48140:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 48141:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 48142:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 48143:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 48144:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 48145:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 48146:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 48147:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 48148:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 48149:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 48150:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 48151:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 48152:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 48153:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 48154:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 48155:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 48156:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 48157:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 48158:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 48159:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 48160:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 48161:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 48162:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 48163:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 48164:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 48165:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 48166:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 48167:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 48168:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 48169:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 48170:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 48171:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 48172:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 48173:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 48174:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 48175:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 48176:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 48177:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 48178:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 48179:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 48180:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 48181:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 48182:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 48183:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 48184:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 48185:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 48186:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 48187:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 48188:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 48189:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 48190:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 48191:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 48192:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 48193:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 48194:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 48195:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 48196:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 48197:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 48198:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 48199:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 48200:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 48201:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 48202:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 48203:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 48204:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 48205:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 48206:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 48207:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 48208:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 48209:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 48210:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 48211:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 48212:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 48213:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 48214:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 48215:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 48216:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 48217:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 48218:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 48219:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 48220:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 48221:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 48222:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 48223:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 48224:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 48225:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 48226:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 48227:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 48228:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 48229:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 48230:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 48231:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 48232:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 48233:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 48234:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 48235:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 48236:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 48237:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 48238:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 48239:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 48240:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 48241:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 48242:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 48243:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 48244:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 48245:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 48246:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 48247:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 48248:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 48249:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 48250:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 48251:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 48252:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 48253:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 48254:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 48255:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 48256:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 48257:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 48258:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 48259:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 48260:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 48261:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 48262:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 48263:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 48264:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 48265:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 48266:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 48267:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 48268:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 48269:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 48270:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 48271:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 48272:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 48273:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 48274:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 48275:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 48276:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 48277:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 48278:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 48279:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 48280:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 48281:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 48282:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 48283:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 48284:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 48285:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 48286:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 48287:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 48288:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 48289:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 48290:20]
  assign io_z = ~x78; // @[Snxn100k.scala 48291:16]
endmodule
module SnxnLv3Inst33(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst132_io_a; // @[Snxn100k.scala 12976:35]
  wire  inst_SnxnLv4Inst132_io_b; // @[Snxn100k.scala 12976:35]
  wire  inst_SnxnLv4Inst132_io_z; // @[Snxn100k.scala 12976:35]
  wire  inst_SnxnLv4Inst133_io_a; // @[Snxn100k.scala 12980:35]
  wire  inst_SnxnLv4Inst133_io_b; // @[Snxn100k.scala 12980:35]
  wire  inst_SnxnLv4Inst133_io_z; // @[Snxn100k.scala 12980:35]
  wire  inst_SnxnLv4Inst134_io_a; // @[Snxn100k.scala 12984:35]
  wire  inst_SnxnLv4Inst134_io_b; // @[Snxn100k.scala 12984:35]
  wire  inst_SnxnLv4Inst134_io_z; // @[Snxn100k.scala 12984:35]
  wire  inst_SnxnLv4Inst135_io_a; // @[Snxn100k.scala 12988:35]
  wire  inst_SnxnLv4Inst135_io_b; // @[Snxn100k.scala 12988:35]
  wire  inst_SnxnLv4Inst135_io_z; // @[Snxn100k.scala 12988:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst132_io_z + inst_SnxnLv4Inst133_io_z; // @[Snxn100k.scala 12992:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst134_io_z; // @[Snxn100k.scala 12992:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst135_io_z; // @[Snxn100k.scala 12992:92]
  SnxnLv4Inst35 inst_SnxnLv4Inst132 ( // @[Snxn100k.scala 12976:35]
    .io_a(inst_SnxnLv4Inst132_io_a),
    .io_b(inst_SnxnLv4Inst132_io_b),
    .io_z(inst_SnxnLv4Inst132_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst133 ( // @[Snxn100k.scala 12980:35]
    .io_a(inst_SnxnLv4Inst133_io_a),
    .io_b(inst_SnxnLv4Inst133_io_b),
    .io_z(inst_SnxnLv4Inst133_io_z)
  );
  SnxnLv4Inst83 inst_SnxnLv4Inst134 ( // @[Snxn100k.scala 12984:35]
    .io_a(inst_SnxnLv4Inst134_io_a),
    .io_b(inst_SnxnLv4Inst134_io_b),
    .io_z(inst_SnxnLv4Inst134_io_z)
  );
  SnxnLv4Inst135 inst_SnxnLv4Inst135 ( // @[Snxn100k.scala 12988:35]
    .io_a(inst_SnxnLv4Inst135_io_a),
    .io_b(inst_SnxnLv4Inst135_io_b),
    .io_z(inst_SnxnLv4Inst135_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 12993:15]
  assign inst_SnxnLv4Inst132_io_a = io_a; // @[Snxn100k.scala 12977:28]
  assign inst_SnxnLv4Inst132_io_b = io_b; // @[Snxn100k.scala 12978:28]
  assign inst_SnxnLv4Inst133_io_a = io_a; // @[Snxn100k.scala 12981:28]
  assign inst_SnxnLv4Inst133_io_b = io_b; // @[Snxn100k.scala 12982:28]
  assign inst_SnxnLv4Inst134_io_a = io_a; // @[Snxn100k.scala 12985:28]
  assign inst_SnxnLv4Inst134_io_b = io_b; // @[Snxn100k.scala 12986:28]
  assign inst_SnxnLv4Inst135_io_a = io_a; // @[Snxn100k.scala 12989:28]
  assign inst_SnxnLv4Inst135_io_b = io_b; // @[Snxn100k.scala 12990:28]
endmodule
module SnxnLv3Inst34(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst136_io_a; // @[Snxn100k.scala 13598:35]
  wire  inst_SnxnLv4Inst136_io_b; // @[Snxn100k.scala 13598:35]
  wire  inst_SnxnLv4Inst136_io_z; // @[Snxn100k.scala 13598:35]
  wire  inst_SnxnLv4Inst137_io_a; // @[Snxn100k.scala 13602:35]
  wire  inst_SnxnLv4Inst137_io_b; // @[Snxn100k.scala 13602:35]
  wire  inst_SnxnLv4Inst137_io_z; // @[Snxn100k.scala 13602:35]
  wire  inst_SnxnLv4Inst138_io_a; // @[Snxn100k.scala 13606:35]
  wire  inst_SnxnLv4Inst138_io_b; // @[Snxn100k.scala 13606:35]
  wire  inst_SnxnLv4Inst138_io_z; // @[Snxn100k.scala 13606:35]
  wire  inst_SnxnLv4Inst139_io_a; // @[Snxn100k.scala 13610:35]
  wire  inst_SnxnLv4Inst139_io_b; // @[Snxn100k.scala 13610:35]
  wire  inst_SnxnLv4Inst139_io_z; // @[Snxn100k.scala 13610:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst136_io_z + inst_SnxnLv4Inst137_io_z; // @[Snxn100k.scala 13614:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst138_io_z; // @[Snxn100k.scala 13614:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst139_io_z; // @[Snxn100k.scala 13614:92]
  SnxnLv4Inst43 inst_SnxnLv4Inst136 ( // @[Snxn100k.scala 13598:35]
    .io_a(inst_SnxnLv4Inst136_io_a),
    .io_b(inst_SnxnLv4Inst136_io_b),
    .io_z(inst_SnxnLv4Inst136_io_z)
  );
  SnxnLv4Inst75 inst_SnxnLv4Inst137 ( // @[Snxn100k.scala 13602:35]
    .io_a(inst_SnxnLv4Inst137_io_a),
    .io_b(inst_SnxnLv4Inst137_io_b),
    .io_z(inst_SnxnLv4Inst137_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst138 ( // @[Snxn100k.scala 13606:35]
    .io_a(inst_SnxnLv4Inst138_io_a),
    .io_b(inst_SnxnLv4Inst138_io_b),
    .io_z(inst_SnxnLv4Inst138_io_z)
  );
  SnxnLv4Inst38 inst_SnxnLv4Inst139 ( // @[Snxn100k.scala 13610:35]
    .io_a(inst_SnxnLv4Inst139_io_a),
    .io_b(inst_SnxnLv4Inst139_io_b),
    .io_z(inst_SnxnLv4Inst139_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 13615:15]
  assign inst_SnxnLv4Inst136_io_a = io_a; // @[Snxn100k.scala 13599:28]
  assign inst_SnxnLv4Inst136_io_b = io_b; // @[Snxn100k.scala 13600:28]
  assign inst_SnxnLv4Inst137_io_a = io_a; // @[Snxn100k.scala 13603:28]
  assign inst_SnxnLv4Inst137_io_b = io_b; // @[Snxn100k.scala 13604:28]
  assign inst_SnxnLv4Inst138_io_a = io_a; // @[Snxn100k.scala 13607:28]
  assign inst_SnxnLv4Inst138_io_b = io_b; // @[Snxn100k.scala 13608:28]
  assign inst_SnxnLv4Inst139_io_a = io_a; // @[Snxn100k.scala 13611:28]
  assign inst_SnxnLv4Inst139_io_b = io_b; // @[Snxn100k.scala 13612:28]
endmodule
module SnxnLv3Inst35(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst140_io_a; // @[Snxn100k.scala 13989:35]
  wire  inst_SnxnLv4Inst140_io_b; // @[Snxn100k.scala 13989:35]
  wire  inst_SnxnLv4Inst140_io_z; // @[Snxn100k.scala 13989:35]
  wire  inst_SnxnLv4Inst141_io_a; // @[Snxn100k.scala 13993:35]
  wire  inst_SnxnLv4Inst141_io_b; // @[Snxn100k.scala 13993:35]
  wire  inst_SnxnLv4Inst141_io_z; // @[Snxn100k.scala 13993:35]
  wire  inst_SnxnLv4Inst142_io_a; // @[Snxn100k.scala 13997:35]
  wire  inst_SnxnLv4Inst142_io_b; // @[Snxn100k.scala 13997:35]
  wire  inst_SnxnLv4Inst142_io_z; // @[Snxn100k.scala 13997:35]
  wire  inst_SnxnLv4Inst143_io_a; // @[Snxn100k.scala 14001:35]
  wire  inst_SnxnLv4Inst143_io_b; // @[Snxn100k.scala 14001:35]
  wire  inst_SnxnLv4Inst143_io_z; // @[Snxn100k.scala 14001:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst140_io_z + inst_SnxnLv4Inst141_io_z; // @[Snxn100k.scala 14005:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst142_io_z; // @[Snxn100k.scala 14005:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst143_io_z; // @[Snxn100k.scala 14005:92]
  SnxnLv4Inst110 inst_SnxnLv4Inst140 ( // @[Snxn100k.scala 13989:35]
    .io_a(inst_SnxnLv4Inst140_io_a),
    .io_b(inst_SnxnLv4Inst140_io_b),
    .io_z(inst_SnxnLv4Inst140_io_z)
  );
  SnxnLv4Inst135 inst_SnxnLv4Inst141 ( // @[Snxn100k.scala 13993:35]
    .io_a(inst_SnxnLv4Inst141_io_a),
    .io_b(inst_SnxnLv4Inst141_io_b),
    .io_z(inst_SnxnLv4Inst141_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst142 ( // @[Snxn100k.scala 13997:35]
    .io_a(inst_SnxnLv4Inst142_io_a),
    .io_b(inst_SnxnLv4Inst142_io_b),
    .io_z(inst_SnxnLv4Inst142_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst143 ( // @[Snxn100k.scala 14001:35]
    .io_a(inst_SnxnLv4Inst143_io_a),
    .io_b(inst_SnxnLv4Inst143_io_b),
    .io_z(inst_SnxnLv4Inst143_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14006:15]
  assign inst_SnxnLv4Inst140_io_a = io_a; // @[Snxn100k.scala 13990:28]
  assign inst_SnxnLv4Inst140_io_b = io_b; // @[Snxn100k.scala 13991:28]
  assign inst_SnxnLv4Inst141_io_a = io_a; // @[Snxn100k.scala 13994:28]
  assign inst_SnxnLv4Inst141_io_b = io_b; // @[Snxn100k.scala 13995:28]
  assign inst_SnxnLv4Inst142_io_a = io_a; // @[Snxn100k.scala 13998:28]
  assign inst_SnxnLv4Inst142_io_b = io_b; // @[Snxn100k.scala 13999:28]
  assign inst_SnxnLv4Inst143_io_a = io_a; // @[Snxn100k.scala 14002:28]
  assign inst_SnxnLv4Inst143_io_b = io_b; // @[Snxn100k.scala 14003:28]
endmodule
module SnxnLv2Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst32_io_a; // @[Snxn100k.scala 2964:34]
  wire  inst_SnxnLv3Inst32_io_b; // @[Snxn100k.scala 2964:34]
  wire  inst_SnxnLv3Inst32_io_z; // @[Snxn100k.scala 2964:34]
  wire  inst_SnxnLv3Inst33_io_a; // @[Snxn100k.scala 2968:34]
  wire  inst_SnxnLv3Inst33_io_b; // @[Snxn100k.scala 2968:34]
  wire  inst_SnxnLv3Inst33_io_z; // @[Snxn100k.scala 2968:34]
  wire  inst_SnxnLv3Inst34_io_a; // @[Snxn100k.scala 2972:34]
  wire  inst_SnxnLv3Inst34_io_b; // @[Snxn100k.scala 2972:34]
  wire  inst_SnxnLv3Inst34_io_z; // @[Snxn100k.scala 2972:34]
  wire  inst_SnxnLv3Inst35_io_a; // @[Snxn100k.scala 2976:34]
  wire  inst_SnxnLv3Inst35_io_b; // @[Snxn100k.scala 2976:34]
  wire  inst_SnxnLv3Inst35_io_z; // @[Snxn100k.scala 2976:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst32_io_z + inst_SnxnLv3Inst33_io_z; // @[Snxn100k.scala 2980:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst34_io_z; // @[Snxn100k.scala 2980:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst35_io_z; // @[Snxn100k.scala 2980:89]
  SnxnLv3Inst32 inst_SnxnLv3Inst32 ( // @[Snxn100k.scala 2964:34]
    .io_a(inst_SnxnLv3Inst32_io_a),
    .io_b(inst_SnxnLv3Inst32_io_b),
    .io_z(inst_SnxnLv3Inst32_io_z)
  );
  SnxnLv3Inst33 inst_SnxnLv3Inst33 ( // @[Snxn100k.scala 2968:34]
    .io_a(inst_SnxnLv3Inst33_io_a),
    .io_b(inst_SnxnLv3Inst33_io_b),
    .io_z(inst_SnxnLv3Inst33_io_z)
  );
  SnxnLv3Inst34 inst_SnxnLv3Inst34 ( // @[Snxn100k.scala 2972:34]
    .io_a(inst_SnxnLv3Inst34_io_a),
    .io_b(inst_SnxnLv3Inst34_io_b),
    .io_z(inst_SnxnLv3Inst34_io_z)
  );
  SnxnLv3Inst35 inst_SnxnLv3Inst35 ( // @[Snxn100k.scala 2976:34]
    .io_a(inst_SnxnLv3Inst35_io_a),
    .io_b(inst_SnxnLv3Inst35_io_b),
    .io_z(inst_SnxnLv3Inst35_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 2981:15]
  assign inst_SnxnLv3Inst32_io_a = io_a; // @[Snxn100k.scala 2965:27]
  assign inst_SnxnLv3Inst32_io_b = io_b; // @[Snxn100k.scala 2966:27]
  assign inst_SnxnLv3Inst33_io_a = io_a; // @[Snxn100k.scala 2969:27]
  assign inst_SnxnLv3Inst33_io_b = io_b; // @[Snxn100k.scala 2970:27]
  assign inst_SnxnLv3Inst34_io_a = io_a; // @[Snxn100k.scala 2973:27]
  assign inst_SnxnLv3Inst34_io_b = io_b; // @[Snxn100k.scala 2974:27]
  assign inst_SnxnLv3Inst35_io_a = io_a; // @[Snxn100k.scala 2977:27]
  assign inst_SnxnLv3Inst35_io_b = io_b; // @[Snxn100k.scala 2978:27]
endmodule
module SnxnLv4Inst146(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 54620:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 54621:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 54622:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 54623:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 54624:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 54625:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 54626:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 54627:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 54628:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 54629:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 54630:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 54631:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 54632:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 54633:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 54634:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 54635:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 54636:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 54637:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 54638:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 54639:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 54640:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 54641:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 54642:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 54643:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 54644:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 54645:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 54646:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 54647:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 54648:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 54649:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 54650:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 54651:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 54652:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 54653:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 54654:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 54655:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 54656:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 54657:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 54658:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 54659:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 54660:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 54661:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 54662:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 54663:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 54664:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 54665:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 54666:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 54667:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 54668:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 54669:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 54670:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 54671:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 54672:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 54673:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 54674:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 54675:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 54676:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 54677:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 54678:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 54679:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 54680:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 54681:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 54682:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 54683:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 54684:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 54685:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 54686:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 54687:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 54688:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 54689:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 54690:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 54691:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 54692:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 54693:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 54694:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 54695:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 54696:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 54697:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 54698:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 54699:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 54700:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 54701:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 54702:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 54703:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 54704:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 54705:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 54706:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 54707:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 54708:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 54709:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 54710:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 54711:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 54712:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 54713:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 54714:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 54715:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 54716:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 54717:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 54718:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 54719:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 54720:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 54721:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 54722:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 54723:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 54724:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 54725:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 54726:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 54727:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 54728:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 54729:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 54730:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 54731:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 54732:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 54733:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 54734:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 54735:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 54736:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 54737:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 54738:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 54739:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 54740:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 54741:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 54742:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 54743:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 54744:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 54745:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 54746:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 54747:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 54748:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 54749:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 54750:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 54751:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 54752:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 54753:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 54754:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 54755:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 54756:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 54757:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 54758:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 54759:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 54760:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 54761:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 54762:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 54763:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 54764:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 54765:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 54766:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 54767:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 54768:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 54769:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 54770:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 54771:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 54772:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 54773:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 54774:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 54775:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 54776:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 54777:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 54778:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 54779:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 54780:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 54781:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 54782:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 54783:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 54784:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 54785:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 54786:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 54787:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 54788:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 54789:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 54790:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 54791:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 54792:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 54793:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 54794:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 54795:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 54796:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 54797:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 54798:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 54799:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 54800:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 54801:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 54802:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 54803:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 54804:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 54805:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 54806:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 54807:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 54808:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 54809:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 54810:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 54811:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 54812:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 54813:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 54814:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 54815:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 54816:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 54817:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 54818:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 54819:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 54820:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 54821:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 54822:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 54823:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 54824:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 54825:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 54826:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 54827:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 54828:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 54829:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 54830:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 54831:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 54832:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 54833:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 54834:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 54835:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 54836:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 54837:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 54838:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 54839:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 54840:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 54841:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 54842:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 54843:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 54844:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 54845:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 54846:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 54847:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 54848:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 54849:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 54850:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 54851:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 54852:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 54853:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 54854:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 54855:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 54856:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 54857:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 54858:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 54859:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 54860:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 54861:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 54862:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 54863:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 54864:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 54865:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 54866:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 54867:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 54868:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 54869:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 54870:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 54871:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 54872:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 54873:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 54874:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 54875:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 54876:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 54877:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 54878:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 54879:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 54880:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 54881:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 54882:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 54883:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 54884:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 54885:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 54886:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 54887:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 54888:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 54889:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 54890:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 54891:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 54892:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 54893:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 54894:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 54895:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 54896:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 54897:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 54898:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 54899:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 54900:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 54901:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 54902:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 54903:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 54904:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 54905:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 54906:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 54907:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 54908:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 54909:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 54910:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 54911:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 54912:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 54913:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 54914:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 54915:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 54916:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 54917:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 54918:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 54919:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 54920:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 54921:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 54922:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 54923:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 54924:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 54925:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 54926:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 54927:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 54928:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 54929:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 54930:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 54931:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 54932:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 54933:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 54934:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 54935:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 54936:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 54937:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 54938:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 54939:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 54940:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 54941:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 54942:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 54943:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 54944:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 54945:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 54946:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 54947:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 54948:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 54949:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 54950:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 54951:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 54952:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 54953:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 54954:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 54955:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 54956:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 54957:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 54958:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 54959:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 54960:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 54961:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 54962:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 54963:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 54964:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 54965:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 54966:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 54967:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 54968:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 54969:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 54970:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 54971:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 54972:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 54973:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 54974:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 54975:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 54976:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 54977:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 54978:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 54979:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 54980:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 54981:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 54982:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 54983:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 54984:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 54985:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 54986:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 54987:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 54988:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 54989:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 54990:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 54991:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 54992:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 54993:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 54994:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 54995:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 54996:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 54997:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 54998:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 54999:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 55000:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 55001:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 55002:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 55003:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 55004:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 55005:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 55006:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 55007:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 55008:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 55009:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 55010:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 55011:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 55012:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 55013:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 55014:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 55015:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 55016:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 55017:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 55018:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 55019:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 55020:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 55021:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 55022:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 55023:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 55024:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 55025:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 55026:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 55027:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 55028:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 55029:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 55030:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 55031:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 55032:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 55033:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 55034:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 55035:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 55036:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 55037:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 55038:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 55039:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 55040:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 55041:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 55042:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 55043:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 55044:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 55045:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 55046:22]
  assign io_z = ~x106; // @[Snxn100k.scala 55047:17]
endmodule
module SnxnLv4Inst147(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 55058:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 55059:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 55060:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 55061:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 55062:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 55063:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 55064:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 55065:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 55066:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 55067:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 55068:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 55069:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 55070:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 55071:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 55072:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 55073:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 55074:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 55075:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 55076:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 55077:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 55078:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 55079:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 55080:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 55081:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 55082:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 55083:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 55084:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 55085:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 55086:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 55087:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 55088:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 55089:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 55090:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 55091:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 55092:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 55093:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 55094:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 55095:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 55096:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 55097:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 55098:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 55099:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 55100:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 55101:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 55102:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 55103:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 55104:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 55105:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 55106:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 55107:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 55108:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 55109:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 55110:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 55111:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 55112:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 55113:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 55114:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 55115:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 55116:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 55117:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 55118:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 55119:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 55120:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 55121:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 55122:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 55123:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 55124:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 55125:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 55126:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 55127:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 55128:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 55129:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 55130:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 55131:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 55132:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 55133:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 55134:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 55135:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 55136:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 55137:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 55138:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 55139:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 55140:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 55141:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 55142:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 55143:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 55144:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 55145:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 55146:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 55147:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 55148:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 55149:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 55150:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 55151:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 55152:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 55153:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 55154:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 55155:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 55156:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 55157:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 55158:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 55159:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 55160:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 55161:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 55162:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 55163:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 55164:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 55165:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 55166:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 55167:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 55168:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 55169:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 55170:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 55171:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 55172:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 55173:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 55174:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 55175:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 55176:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 55177:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 55178:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 55179:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 55180:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 55181:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 55182:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 55183:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 55184:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 55185:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 55186:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 55187:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 55188:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 55189:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 55190:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 55191:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 55192:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 55193:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 55194:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 55195:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 55196:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 55197:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 55198:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 55199:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 55200:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 55201:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 55202:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 55203:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 55204:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 55205:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 55206:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 55207:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 55208:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 55209:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 55210:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 55211:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 55212:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 55213:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 55214:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 55215:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 55216:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 55217:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 55218:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 55219:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 55220:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 55221:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 55222:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 55223:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 55224:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 55225:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 55226:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 55227:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 55228:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 55229:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 55230:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 55231:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 55232:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 55233:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 55234:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 55235:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 55236:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 55237:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 55238:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 55239:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 55240:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 55241:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 55242:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 55243:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 55244:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 55245:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 55246:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 55247:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 55248:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 55249:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 55250:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 55251:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 55252:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 55253:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 55254:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 55255:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 55256:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 55257:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 55258:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 55259:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 55260:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 55261:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 55262:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 55263:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 55264:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 55265:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 55266:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 55267:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 55268:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 55269:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 55270:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 55271:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 55272:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 55273:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 55274:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 55275:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 55276:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 55277:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 55278:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 55279:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 55280:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 55281:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 55282:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 55283:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 55284:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 55285:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 55286:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 55287:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 55288:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 55289:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 55290:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 55291:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 55292:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 55293:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 55294:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 55295:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 55296:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 55297:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 55298:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 55299:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 55300:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 55301:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 55302:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 55303:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 55304:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 55305:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 55306:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 55307:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 55308:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 55309:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 55310:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 55311:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 55312:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 55313:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 55314:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 55315:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 55316:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 55317:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 55318:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 55319:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 55320:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 55321:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 55322:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 55323:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 55324:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 55325:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 55326:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 55327:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 55328:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 55329:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 55330:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 55331:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 55332:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 55333:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 55334:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 55335:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 55336:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 55337:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 55338:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 55339:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 55340:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 55341:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 55342:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 55343:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 55344:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 55345:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 55346:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 55347:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 55348:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 55349:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 55350:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 55351:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 55352:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 55353:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 55354:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 55355:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 55356:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 55357:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 55358:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 55359:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 55360:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 55361:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 55362:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 55363:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 55364:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 55365:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 55366:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 55367:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 55368:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 55369:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 55370:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 55371:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 55372:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 55373:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 55374:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 55375:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 55376:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 55377:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 55378:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 55379:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 55380:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 55381:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 55382:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 55383:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 55384:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 55385:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 55386:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 55387:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 55388:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 55389:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 55390:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 55391:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 55392:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 55393:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 55394:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 55395:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 55396:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 55397:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 55398:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 55399:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 55400:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 55401:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 55402:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 55403:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 55404:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 55405:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 55406:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 55407:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 55408:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 55409:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 55410:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 55411:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 55412:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 55413:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 55414:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 55415:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 55416:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 55417:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 55418:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 55419:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 55420:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 55421:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 55422:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 55423:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 55424:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 55425:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 55426:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 55427:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 55428:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 55429:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 55430:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 55431:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 55432:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 55433:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 55434:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 55435:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 55436:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 55437:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 55438:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 55439:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 55440:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 55441:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 55442:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 55443:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 55444:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 55445:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 55446:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 55447:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 55448:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 55449:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 55450:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 55451:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 55452:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 55453:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 55454:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 55455:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 55456:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 55457:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 55458:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 55459:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 55460:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 55461:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 55462:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 55463:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 55464:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 55465:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 55466:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 55467:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 55468:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 55469:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 55470:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 55471:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 55472:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 55473:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 55474:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 55475:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 55476:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 55477:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 55478:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 55479:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 55480:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 55481:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 55482:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 55483:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 55484:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 55485:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 55486:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 55487:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 55488:22]
  assign io_z = ~x107; // @[Snxn100k.scala 55489:17]
endmodule
module SnxnLv3Inst36(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst144_io_a; // @[Snxn100k.scala 14423:35]
  wire  inst_SnxnLv4Inst144_io_b; // @[Snxn100k.scala 14423:35]
  wire  inst_SnxnLv4Inst144_io_z; // @[Snxn100k.scala 14423:35]
  wire  inst_SnxnLv4Inst145_io_a; // @[Snxn100k.scala 14427:35]
  wire  inst_SnxnLv4Inst145_io_b; // @[Snxn100k.scala 14427:35]
  wire  inst_SnxnLv4Inst145_io_z; // @[Snxn100k.scala 14427:35]
  wire  inst_SnxnLv4Inst146_io_a; // @[Snxn100k.scala 14431:35]
  wire  inst_SnxnLv4Inst146_io_b; // @[Snxn100k.scala 14431:35]
  wire  inst_SnxnLv4Inst146_io_z; // @[Snxn100k.scala 14431:35]
  wire  inst_SnxnLv4Inst147_io_a; // @[Snxn100k.scala 14435:35]
  wire  inst_SnxnLv4Inst147_io_b; // @[Snxn100k.scala 14435:35]
  wire  inst_SnxnLv4Inst147_io_z; // @[Snxn100k.scala 14435:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst144_io_z + inst_SnxnLv4Inst145_io_z; // @[Snxn100k.scala 14439:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst146_io_z; // @[Snxn100k.scala 14439:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst147_io_z; // @[Snxn100k.scala 14439:92]
  SnxnLv4Inst16 inst_SnxnLv4Inst144 ( // @[Snxn100k.scala 14423:35]
    .io_a(inst_SnxnLv4Inst144_io_a),
    .io_b(inst_SnxnLv4Inst144_io_b),
    .io_z(inst_SnxnLv4Inst144_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst145 ( // @[Snxn100k.scala 14427:35]
    .io_a(inst_SnxnLv4Inst145_io_a),
    .io_b(inst_SnxnLv4Inst145_io_b),
    .io_z(inst_SnxnLv4Inst145_io_z)
  );
  SnxnLv4Inst146 inst_SnxnLv4Inst146 ( // @[Snxn100k.scala 14431:35]
    .io_a(inst_SnxnLv4Inst146_io_a),
    .io_b(inst_SnxnLv4Inst146_io_b),
    .io_z(inst_SnxnLv4Inst146_io_z)
  );
  SnxnLv4Inst147 inst_SnxnLv4Inst147 ( // @[Snxn100k.scala 14435:35]
    .io_a(inst_SnxnLv4Inst147_io_a),
    .io_b(inst_SnxnLv4Inst147_io_b),
    .io_z(inst_SnxnLv4Inst147_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14440:15]
  assign inst_SnxnLv4Inst144_io_a = io_a; // @[Snxn100k.scala 14424:28]
  assign inst_SnxnLv4Inst144_io_b = io_b; // @[Snxn100k.scala 14425:28]
  assign inst_SnxnLv4Inst145_io_a = io_a; // @[Snxn100k.scala 14428:28]
  assign inst_SnxnLv4Inst145_io_b = io_b; // @[Snxn100k.scala 14429:28]
  assign inst_SnxnLv4Inst146_io_a = io_a; // @[Snxn100k.scala 14432:28]
  assign inst_SnxnLv4Inst146_io_b = io_b; // @[Snxn100k.scala 14433:28]
  assign inst_SnxnLv4Inst147_io_a = io_a; // @[Snxn100k.scala 14436:28]
  assign inst_SnxnLv4Inst147_io_b = io_b; // @[Snxn100k.scala 14437:28]
endmodule
module SnxnLv4Inst148(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 57174:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 57175:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 57176:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 57177:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 57178:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 57179:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 57180:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 57181:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 57182:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 57183:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 57184:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 57185:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 57186:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 57187:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 57188:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 57189:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 57190:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 57191:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 57192:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 57193:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 57194:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 57195:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 57196:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 57197:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 57198:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 57199:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 57200:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 57201:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 57202:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 57203:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 57204:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 57205:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 57206:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 57207:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 57208:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 57209:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 57210:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 57211:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 57212:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 57213:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 57214:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 57215:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 57216:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 57217:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 57218:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 57219:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 57220:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 57221:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 57222:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 57223:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 57224:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 57225:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 57226:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 57227:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 57228:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 57229:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 57230:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 57231:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 57232:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 57233:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 57234:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 57235:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 57236:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 57237:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 57238:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 57239:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 57240:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 57241:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 57242:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 57243:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 57244:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 57245:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 57246:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 57247:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 57248:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 57249:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 57250:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 57251:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 57252:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 57253:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 57254:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 57255:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 57256:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 57257:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 57258:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 57259:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 57260:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 57261:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 57262:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 57263:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 57264:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 57265:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 57266:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 57267:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 57268:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 57269:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 57270:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 57271:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 57272:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 57273:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 57274:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 57275:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 57276:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 57277:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 57278:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 57279:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 57280:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 57281:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 57282:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 57283:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 57284:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 57285:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 57286:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 57287:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 57288:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 57289:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 57290:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 57291:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 57292:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 57293:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 57294:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 57295:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 57296:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 57297:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 57298:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 57299:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 57300:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 57301:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 57302:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 57303:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 57304:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 57305:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 57306:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 57307:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 57308:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 57309:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 57310:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 57311:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 57312:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 57313:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 57314:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 57315:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 57316:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 57317:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 57318:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 57319:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 57320:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 57321:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 57322:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 57323:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 57324:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 57325:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 57326:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 57327:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 57328:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 57329:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 57330:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 57331:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 57332:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 57333:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 57334:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 57335:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 57336:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 57337:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 57338:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 57339:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 57340:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 57341:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 57342:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 57343:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 57344:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 57345:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 57346:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 57347:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 57348:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 57349:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 57350:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 57351:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 57352:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 57353:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 57354:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 57355:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 57356:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 57357:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 57358:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 57359:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 57360:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 57361:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 57362:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 57363:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 57364:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 57365:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 57366:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 57367:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 57368:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 57369:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 57370:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 57371:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 57372:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 57373:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 57374:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 57375:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 57376:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 57377:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 57378:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 57379:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 57380:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 57381:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 57382:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 57383:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 57384:20]
  assign io_z = ~x52; // @[Snxn100k.scala 57385:16]
endmodule
module SnxnLv4Inst150(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 57016:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 57017:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 57018:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 57019:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 57020:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 57021:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 57022:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 57023:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 57024:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 57025:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 57026:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 57027:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 57028:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 57029:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 57030:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 57031:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 57032:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 57033:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 57034:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 57035:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 57036:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 57037:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 57038:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 57039:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 57040:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 57041:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 57042:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 57043:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 57044:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 57045:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 57046:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 57047:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 57048:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 57049:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 57050:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 57051:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 57052:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 57053:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 57054:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 57055:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 57056:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 57057:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 57058:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 57059:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 57060:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 57061:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 57062:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 57063:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 57064:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 57065:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 57066:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 57067:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 57068:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 57069:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 57070:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 57071:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 57072:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 57073:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 57074:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 57075:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 57076:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 57077:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 57078:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 57079:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 57080:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 57081:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 57082:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 57083:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 57084:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 57085:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 57086:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 57087:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 57088:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 57089:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 57090:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 57091:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 57092:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 57093:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 57094:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 57095:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 57096:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 57097:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 57098:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 57099:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 57100:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 57101:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 57102:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 57103:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 57104:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 57105:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 57106:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 57107:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 57108:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 57109:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 57110:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 57111:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 57112:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 57113:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 57114:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 57115:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 57116:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 57117:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 57118:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 57119:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 57120:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 57121:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 57122:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 57123:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 57124:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 57125:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 57126:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 57127:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 57128:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 57129:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 57130:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 57131:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 57132:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 57133:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 57134:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 57135:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 57136:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 57137:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 57138:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 57139:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 57140:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 57141:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 57142:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 57143:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 57144:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 57145:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 57146:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 57147:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 57148:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 57149:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 57150:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 57151:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 57152:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 57153:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 57154:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 57155:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 57156:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 57157:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 57158:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 57159:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 57160:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 57161:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 57162:20]
  assign io_z = ~x36; // @[Snxn100k.scala 57163:16]
endmodule
module SnxnLv4Inst151(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 57618:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 57619:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 57620:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 57621:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 57622:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 57623:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 57624:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 57625:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 57626:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 57627:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 57628:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 57629:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 57630:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 57631:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 57632:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 57633:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 57634:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 57635:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 57636:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 57637:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 57638:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 57639:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 57640:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 57641:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 57642:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 57643:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 57644:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 57645:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 57646:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 57647:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 57648:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 57649:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 57650:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 57651:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 57652:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 57653:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 57654:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 57655:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 57656:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 57657:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 57658:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 57659:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 57660:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 57661:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 57662:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 57663:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 57664:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 57665:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 57666:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 57667:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 57668:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 57669:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 57670:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 57671:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 57672:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 57673:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 57674:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 57675:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 57676:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 57677:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 57678:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 57679:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 57680:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 57681:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 57682:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 57683:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 57684:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 57685:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 57686:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 57687:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 57688:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 57689:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 57690:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 57691:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 57692:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 57693:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 57694:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 57695:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 57696:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 57697:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 57698:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 57699:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 57700:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 57701:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 57702:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 57703:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 57704:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 57705:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 57706:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 57707:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 57708:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 57709:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 57710:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 57711:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 57712:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 57713:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 57714:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 57715:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 57716:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 57717:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 57718:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 57719:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 57720:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 57721:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 57722:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 57723:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 57724:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 57725:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 57726:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 57727:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 57728:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 57729:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 57730:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 57731:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 57732:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 57733:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 57734:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 57735:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 57736:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 57737:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 57738:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 57739:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 57740:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 57741:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 57742:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 57743:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 57744:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 57745:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 57746:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 57747:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 57748:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 57749:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 57750:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 57751:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 57752:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 57753:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 57754:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 57755:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 57756:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 57757:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 57758:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 57759:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 57760:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 57761:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 57762:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 57763:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 57764:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 57765:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 57766:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 57767:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 57768:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 57769:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 57770:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 57771:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 57772:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 57773:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 57774:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 57775:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 57776:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 57777:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 57778:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 57779:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 57780:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 57781:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 57782:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 57783:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 57784:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 57785:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 57786:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 57787:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 57788:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 57789:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 57790:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 57791:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 57792:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 57793:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 57794:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 57795:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 57796:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 57797:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 57798:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 57799:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 57800:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 57801:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 57802:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 57803:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 57804:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 57805:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 57806:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 57807:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 57808:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 57809:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 57810:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 57811:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 57812:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 57813:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 57814:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 57815:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 57816:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 57817:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 57818:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 57819:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 57820:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 57821:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 57822:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 57823:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 57824:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 57825:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 57826:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 57827:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 57828:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 57829:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 57830:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 57831:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 57832:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 57833:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 57834:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 57835:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 57836:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 57837:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 57838:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 57839:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 57840:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 57841:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 57842:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 57843:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 57844:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 57845:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 57846:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 57847:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 57848:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 57849:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 57850:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 57851:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 57852:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 57853:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 57854:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 57855:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 57856:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 57857:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 57858:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 57859:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 57860:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 57861:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 57862:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 57863:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 57864:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 57865:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 57866:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 57867:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 57868:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 57869:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 57870:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 57871:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 57872:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 57873:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 57874:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 57875:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 57876:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 57877:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 57878:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 57879:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 57880:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 57881:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 57882:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 57883:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 57884:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 57885:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 57886:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 57887:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 57888:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 57889:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 57890:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 57891:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 57892:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 57893:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 57894:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 57895:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 57896:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 57897:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 57898:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 57899:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 57900:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 57901:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 57902:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 57903:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 57904:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 57905:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 57906:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 57907:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 57908:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 57909:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 57910:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 57911:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 57912:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 57913:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 57914:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 57915:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 57916:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 57917:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 57918:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 57919:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 57920:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 57921:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 57922:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 57923:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 57924:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 57925:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 57926:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 57927:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 57928:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 57929:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 57930:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 57931:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 57932:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 57933:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 57934:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 57935:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 57936:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 57937:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 57938:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 57939:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 57940:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 57941:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 57942:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 57943:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 57944:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 57945:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 57946:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 57947:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 57948:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 57949:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 57950:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 57951:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 57952:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 57953:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 57954:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 57955:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 57956:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 57957:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 57958:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 57959:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 57960:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 57961:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 57962:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 57963:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 57964:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 57965:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 57966:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 57967:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 57968:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 57969:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 57970:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 57971:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 57972:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 57973:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 57974:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 57975:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 57976:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 57977:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 57978:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 57979:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 57980:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 57981:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 57982:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 57983:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 57984:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 57985:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 57986:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 57987:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 57988:20]
  assign io_z = ~x92; // @[Snxn100k.scala 57989:16]
endmodule
module SnxnLv3Inst37(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst148_io_a; // @[Snxn100k.scala 15173:35]
  wire  inst_SnxnLv4Inst148_io_b; // @[Snxn100k.scala 15173:35]
  wire  inst_SnxnLv4Inst148_io_z; // @[Snxn100k.scala 15173:35]
  wire  inst_SnxnLv4Inst149_io_a; // @[Snxn100k.scala 15177:35]
  wire  inst_SnxnLv4Inst149_io_b; // @[Snxn100k.scala 15177:35]
  wire  inst_SnxnLv4Inst149_io_z; // @[Snxn100k.scala 15177:35]
  wire  inst_SnxnLv4Inst150_io_a; // @[Snxn100k.scala 15181:35]
  wire  inst_SnxnLv4Inst150_io_b; // @[Snxn100k.scala 15181:35]
  wire  inst_SnxnLv4Inst150_io_z; // @[Snxn100k.scala 15181:35]
  wire  inst_SnxnLv4Inst151_io_a; // @[Snxn100k.scala 15185:35]
  wire  inst_SnxnLv4Inst151_io_b; // @[Snxn100k.scala 15185:35]
  wire  inst_SnxnLv4Inst151_io_z; // @[Snxn100k.scala 15185:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst148_io_z + inst_SnxnLv4Inst149_io_z; // @[Snxn100k.scala 15189:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst150_io_z; // @[Snxn100k.scala 15189:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst151_io_z; // @[Snxn100k.scala 15189:92]
  SnxnLv4Inst148 inst_SnxnLv4Inst148 ( // @[Snxn100k.scala 15173:35]
    .io_a(inst_SnxnLv4Inst148_io_a),
    .io_b(inst_SnxnLv4Inst148_io_b),
    .io_z(inst_SnxnLv4Inst148_io_z)
  );
  SnxnLv4Inst148 inst_SnxnLv4Inst149 ( // @[Snxn100k.scala 15177:35]
    .io_a(inst_SnxnLv4Inst149_io_a),
    .io_b(inst_SnxnLv4Inst149_io_b),
    .io_z(inst_SnxnLv4Inst149_io_z)
  );
  SnxnLv4Inst150 inst_SnxnLv4Inst150 ( // @[Snxn100k.scala 15181:35]
    .io_a(inst_SnxnLv4Inst150_io_a),
    .io_b(inst_SnxnLv4Inst150_io_b),
    .io_z(inst_SnxnLv4Inst150_io_z)
  );
  SnxnLv4Inst151 inst_SnxnLv4Inst151 ( // @[Snxn100k.scala 15185:35]
    .io_a(inst_SnxnLv4Inst151_io_a),
    .io_b(inst_SnxnLv4Inst151_io_b),
    .io_z(inst_SnxnLv4Inst151_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 15190:15]
  assign inst_SnxnLv4Inst148_io_a = io_a; // @[Snxn100k.scala 15174:28]
  assign inst_SnxnLv4Inst148_io_b = io_b; // @[Snxn100k.scala 15175:28]
  assign inst_SnxnLv4Inst149_io_a = io_a; // @[Snxn100k.scala 15178:28]
  assign inst_SnxnLv4Inst149_io_b = io_b; // @[Snxn100k.scala 15179:28]
  assign inst_SnxnLv4Inst150_io_a = io_a; // @[Snxn100k.scala 15182:28]
  assign inst_SnxnLv4Inst150_io_b = io_b; // @[Snxn100k.scala 15183:28]
  assign inst_SnxnLv4Inst151_io_a = io_a; // @[Snxn100k.scala 15186:28]
  assign inst_SnxnLv4Inst151_io_b = io_b; // @[Snxn100k.scala 15187:28]
endmodule
module SnxnLv4Inst153(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 56104:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 56105:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 56106:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 56107:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 56108:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 56109:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 56110:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 56111:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 56112:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 56113:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 56114:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 56115:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 56116:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 56117:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 56118:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 56119:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 56120:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 56121:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 56122:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 56123:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 56124:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 56125:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 56126:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 56127:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 56128:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 56129:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 56130:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 56131:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 56132:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 56133:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 56134:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 56135:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 56136:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 56137:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 56138:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 56139:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 56140:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 56141:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 56142:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 56143:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 56144:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 56145:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 56146:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 56147:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 56148:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 56149:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 56150:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 56151:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 56152:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 56153:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 56154:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 56155:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 56156:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 56157:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 56158:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 56159:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 56160:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 56161:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 56162:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 56163:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 56164:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 56165:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 56166:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 56167:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 56168:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 56169:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 56170:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 56171:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 56172:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 56173:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 56174:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 56175:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 56176:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 56177:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 56178:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 56179:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 56180:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 56181:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 56182:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 56183:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 56184:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 56185:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 56186:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 56187:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 56188:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 56189:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 56190:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 56191:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 56192:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 56193:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 56194:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 56195:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 56196:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 56197:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 56198:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 56199:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 56200:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 56201:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 56202:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 56203:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 56204:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 56205:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 56206:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 56207:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 56208:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 56209:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 56210:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 56211:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 56212:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 56213:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 56214:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 56215:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 56216:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 56217:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 56218:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 56219:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 56220:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 56221:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 56222:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 56223:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 56224:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 56225:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 56226:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 56227:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 56228:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 56229:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 56230:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 56231:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 56232:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 56233:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 56234:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 56235:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 56236:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 56237:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 56238:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 56239:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 56240:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 56241:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 56242:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 56243:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 56244:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 56245:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 56246:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 56247:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 56248:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 56249:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 56250:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 56251:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 56252:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 56253:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 56254:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 56255:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 56256:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 56257:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 56258:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 56259:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 56260:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 56261:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 56262:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 56263:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 56264:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 56265:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 56266:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 56267:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 56268:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 56269:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 56270:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 56271:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 56272:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 56273:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 56274:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 56275:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 56276:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 56277:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 56278:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 56279:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 56280:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 56281:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 56282:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 56283:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 56284:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 56285:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 56286:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 56287:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 56288:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 56289:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 56290:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 56291:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 56292:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 56293:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 56294:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 56295:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 56296:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 56297:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 56298:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 56299:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 56300:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 56301:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 56302:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 56303:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 56304:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 56305:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 56306:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 56307:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 56308:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 56309:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 56310:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 56311:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 56312:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 56313:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 56314:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 56315:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 56316:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 56317:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 56318:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 56319:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 56320:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 56321:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 56322:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 56323:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 56324:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 56325:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 56326:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 56327:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 56328:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 56329:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 56330:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 56331:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 56332:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 56333:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 56334:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 56335:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 56336:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 56337:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 56338:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 56339:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 56340:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 56341:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 56342:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 56343:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 56344:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 56345:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 56346:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 56347:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 56348:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 56349:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 56350:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 56351:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 56352:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 56353:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 56354:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 56355:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 56356:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 56357:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 56358:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 56359:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 56360:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 56361:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 56362:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 56363:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 56364:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 56365:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 56366:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 56367:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 56368:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 56369:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 56370:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 56371:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 56372:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 56373:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 56374:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 56375:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 56376:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 56377:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 56378:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 56379:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 56380:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 56381:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 56382:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 56383:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 56384:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 56385:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 56386:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 56387:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 56388:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 56389:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 56390:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 56391:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 56392:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 56393:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 56394:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 56395:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 56396:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 56397:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 56398:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 56399:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 56400:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 56401:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 56402:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 56403:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 56404:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 56405:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 56406:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 56407:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 56408:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 56409:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 56410:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 56411:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 56412:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 56413:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 56414:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 56415:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 56416:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 56417:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 56418:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 56419:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 56420:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 56421:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 56422:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 56423:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 56424:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 56425:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 56426:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 56427:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 56428:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 56429:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 56430:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 56431:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 56432:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 56433:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 56434:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 56435:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 56436:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 56437:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 56438:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 56439:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 56440:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 56441:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 56442:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 56443:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 56444:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 56445:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 56446:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 56447:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 56448:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 56449:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 56450:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 56451:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 56452:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 56453:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 56454:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 56455:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 56456:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 56457:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 56458:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 56459:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 56460:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 56461:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 56462:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 56463:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 56464:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 56465:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 56466:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 56467:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 56468:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 56469:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 56470:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 56471:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 56472:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 56473:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 56474:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 56475:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 56476:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 56477:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 56478:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 56479:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 56480:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 56481:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 56482:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 56483:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 56484:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 56485:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 56486:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 56487:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 56488:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 56489:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 56490:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 56491:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 56492:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 56493:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 56494:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 56495:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 56496:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 56497:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 56498:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 56499:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 56500:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 56501:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 56502:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 56503:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 56504:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 56505:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 56506:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 56507:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 56508:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 56509:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 56510:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 56511:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 56512:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 56513:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 56514:22]
  assign io_z = ~x102; // @[Snxn100k.scala 56515:17]
endmodule
module SnxnLv4Inst155(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 56526:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 56527:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 56528:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 56529:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 56530:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 56531:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 56532:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 56533:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 56534:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 56535:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 56536:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 56537:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 56538:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 56539:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 56540:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 56541:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 56542:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 56543:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 56544:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 56545:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 56546:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 56547:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 56548:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 56549:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 56550:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 56551:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 56552:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 56553:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 56554:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 56555:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 56556:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 56557:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 56558:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 56559:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 56560:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 56561:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 56562:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 56563:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 56564:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 56565:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 56566:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 56567:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 56568:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 56569:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 56570:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 56571:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 56572:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 56573:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 56574:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 56575:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 56576:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 56577:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 56578:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 56579:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 56580:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 56581:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 56582:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 56583:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 56584:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 56585:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 56586:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 56587:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 56588:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 56589:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 56590:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 56591:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 56592:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 56593:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 56594:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 56595:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 56596:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 56597:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 56598:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 56599:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 56600:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 56601:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 56602:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 56603:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 56604:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 56605:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 56606:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 56607:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 56608:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 56609:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 56610:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 56611:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 56612:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 56613:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 56614:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 56615:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 56616:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 56617:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 56618:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 56619:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 56620:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 56621:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 56622:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 56623:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 56624:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 56625:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 56626:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 56627:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 56628:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 56629:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 56630:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 56631:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 56632:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 56633:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 56634:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 56635:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 56636:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 56637:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 56638:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 56639:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 56640:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 56641:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 56642:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 56643:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 56644:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 56645:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 56646:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 56647:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 56648:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 56649:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 56650:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 56651:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 56652:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 56653:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 56654:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 56655:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 56656:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 56657:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 56658:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 56659:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 56660:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 56661:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 56662:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 56663:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 56664:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 56665:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 56666:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 56667:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 56668:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 56669:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 56670:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 56671:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 56672:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 56673:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 56674:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 56675:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 56676:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 56677:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 56678:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 56679:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 56680:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 56681:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 56682:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 56683:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 56684:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 56685:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 56686:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 56687:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 56688:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 56689:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 56690:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 56691:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 56692:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 56693:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 56694:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 56695:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 56696:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 56697:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 56698:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 56699:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 56700:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 56701:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 56702:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 56703:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 56704:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 56705:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 56706:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 56707:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 56708:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 56709:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 56710:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 56711:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 56712:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 56713:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 56714:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 56715:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 56716:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 56717:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 56718:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 56719:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 56720:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 56721:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 56722:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 56723:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 56724:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 56725:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 56726:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 56727:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 56728:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 56729:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 56730:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 56731:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 56732:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 56733:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 56734:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 56735:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 56736:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 56737:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 56738:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 56739:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 56740:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 56741:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 56742:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 56743:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 56744:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 56745:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 56746:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 56747:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 56748:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 56749:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 56750:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 56751:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 56752:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 56753:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 56754:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 56755:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 56756:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 56757:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 56758:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 56759:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 56760:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 56761:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 56762:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 56763:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 56764:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 56765:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 56766:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 56767:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 56768:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 56769:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 56770:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 56771:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 56772:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 56773:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 56774:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 56775:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 56776:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 56777:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 56778:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 56779:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 56780:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 56781:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 56782:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 56783:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 56784:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 56785:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 56786:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 56787:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 56788:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 56789:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 56790:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 56791:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 56792:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 56793:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 56794:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 56795:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 56796:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 56797:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 56798:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 56799:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 56800:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 56801:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 56802:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 56803:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 56804:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 56805:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 56806:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 56807:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 56808:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 56809:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 56810:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 56811:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 56812:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 56813:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 56814:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 56815:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 56816:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 56817:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 56818:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 56819:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 56820:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 56821:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 56822:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 56823:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 56824:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 56825:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 56826:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 56827:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 56828:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 56829:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 56830:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 56831:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 56832:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 56833:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 56834:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 56835:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 56836:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 56837:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 56838:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 56839:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 56840:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 56841:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 56842:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 56843:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 56844:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 56845:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 56846:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 56847:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 56848:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 56849:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 56850:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 56851:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 56852:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 56853:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 56854:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 56855:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 56856:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 56857:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 56858:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 56859:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 56860:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 56861:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 56862:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 56863:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 56864:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 56865:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 56866:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 56867:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 56868:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 56869:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 56870:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 56871:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 56872:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 56873:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 56874:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 56875:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 56876:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 56877:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 56878:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 56879:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 56880:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 56881:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 56882:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 56883:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 56884:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 56885:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 56886:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 56887:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 56888:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 56889:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 56890:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 56891:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 56892:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 56893:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 56894:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 56895:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 56896:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 56897:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 56898:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 56899:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 56900:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 56901:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 56902:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 56903:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 56904:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 56905:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 56906:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 56907:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 56908:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 56909:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 56910:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 56911:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 56912:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 56913:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 56914:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 56915:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 56916:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 56917:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 56918:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 56919:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 56920:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 56921:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 56922:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 56923:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 56924:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 56925:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 56926:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 56927:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 56928:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 56929:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 56930:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 56931:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 56932:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 56933:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 56934:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 56935:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 56936:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 56937:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 56938:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 56939:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 56940:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 56941:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 56942:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 56943:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 56944:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 56945:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 56946:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 56947:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 56948:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 56949:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 56950:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 56951:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 56952:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 56953:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 56954:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 56955:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 56956:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 56957:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 56958:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 56959:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 56960:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 56961:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 56962:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 56963:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 56964:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 56965:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 56966:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 56967:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 56968:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 56969:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 56970:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 56971:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 56972:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 56973:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 56974:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 56975:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 56976:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 56977:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 56978:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 56979:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 56980:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 56981:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 56982:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 56983:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 56984:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 56985:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 56986:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 56987:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 56988:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 56989:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 56990:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 56991:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 56992:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 56993:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 56994:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 56995:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 56996:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 56997:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 56998:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 56999:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 57000:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 57001:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 57002:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 57003:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 57004:22]
  assign io_z = ~x119; // @[Snxn100k.scala 57005:17]
endmodule
module SnxnLv3Inst38(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst152_io_a; // @[Snxn100k.scala 14766:35]
  wire  inst_SnxnLv4Inst152_io_b; // @[Snxn100k.scala 14766:35]
  wire  inst_SnxnLv4Inst152_io_z; // @[Snxn100k.scala 14766:35]
  wire  inst_SnxnLv4Inst153_io_a; // @[Snxn100k.scala 14770:35]
  wire  inst_SnxnLv4Inst153_io_b; // @[Snxn100k.scala 14770:35]
  wire  inst_SnxnLv4Inst153_io_z; // @[Snxn100k.scala 14770:35]
  wire  inst_SnxnLv4Inst154_io_a; // @[Snxn100k.scala 14774:35]
  wire  inst_SnxnLv4Inst154_io_b; // @[Snxn100k.scala 14774:35]
  wire  inst_SnxnLv4Inst154_io_z; // @[Snxn100k.scala 14774:35]
  wire  inst_SnxnLv4Inst155_io_a; // @[Snxn100k.scala 14778:35]
  wire  inst_SnxnLv4Inst155_io_b; // @[Snxn100k.scala 14778:35]
  wire  inst_SnxnLv4Inst155_io_z; // @[Snxn100k.scala 14778:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst152_io_z + inst_SnxnLv4Inst153_io_z; // @[Snxn100k.scala 14782:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst154_io_z; // @[Snxn100k.scala 14782:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst155_io_z; // @[Snxn100k.scala 14782:92]
  SnxnLv4Inst69 inst_SnxnLv4Inst152 ( // @[Snxn100k.scala 14766:35]
    .io_a(inst_SnxnLv4Inst152_io_a),
    .io_b(inst_SnxnLv4Inst152_io_b),
    .io_z(inst_SnxnLv4Inst152_io_z)
  );
  SnxnLv4Inst153 inst_SnxnLv4Inst153 ( // @[Snxn100k.scala 14770:35]
    .io_a(inst_SnxnLv4Inst153_io_a),
    .io_b(inst_SnxnLv4Inst153_io_b),
    .io_z(inst_SnxnLv4Inst153_io_z)
  );
  SnxnLv4Inst7 inst_SnxnLv4Inst154 ( // @[Snxn100k.scala 14774:35]
    .io_a(inst_SnxnLv4Inst154_io_a),
    .io_b(inst_SnxnLv4Inst154_io_b),
    .io_z(inst_SnxnLv4Inst154_io_z)
  );
  SnxnLv4Inst155 inst_SnxnLv4Inst155 ( // @[Snxn100k.scala 14778:35]
    .io_a(inst_SnxnLv4Inst155_io_a),
    .io_b(inst_SnxnLv4Inst155_io_b),
    .io_z(inst_SnxnLv4Inst155_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14783:15]
  assign inst_SnxnLv4Inst152_io_a = io_a; // @[Snxn100k.scala 14767:28]
  assign inst_SnxnLv4Inst152_io_b = io_b; // @[Snxn100k.scala 14768:28]
  assign inst_SnxnLv4Inst153_io_a = io_a; // @[Snxn100k.scala 14771:28]
  assign inst_SnxnLv4Inst153_io_b = io_b; // @[Snxn100k.scala 14772:28]
  assign inst_SnxnLv4Inst154_io_a = io_a; // @[Snxn100k.scala 14775:28]
  assign inst_SnxnLv4Inst154_io_b = io_b; // @[Snxn100k.scala 14776:28]
  assign inst_SnxnLv4Inst155_io_a = io_a; // @[Snxn100k.scala 14779:28]
  assign inst_SnxnLv4Inst155_io_b = io_b; // @[Snxn100k.scala 14780:28]
endmodule
module SnxnLv3Inst39(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst156_io_a; // @[Snxn100k.scala 14136:35]
  wire  inst_SnxnLv4Inst156_io_b; // @[Snxn100k.scala 14136:35]
  wire  inst_SnxnLv4Inst156_io_z; // @[Snxn100k.scala 14136:35]
  wire  inst_SnxnLv4Inst157_io_a; // @[Snxn100k.scala 14140:35]
  wire  inst_SnxnLv4Inst157_io_b; // @[Snxn100k.scala 14140:35]
  wire  inst_SnxnLv4Inst157_io_z; // @[Snxn100k.scala 14140:35]
  wire  inst_SnxnLv4Inst158_io_a; // @[Snxn100k.scala 14144:35]
  wire  inst_SnxnLv4Inst158_io_b; // @[Snxn100k.scala 14144:35]
  wire  inst_SnxnLv4Inst158_io_z; // @[Snxn100k.scala 14144:35]
  wire  inst_SnxnLv4Inst159_io_a; // @[Snxn100k.scala 14148:35]
  wire  inst_SnxnLv4Inst159_io_b; // @[Snxn100k.scala 14148:35]
  wire  inst_SnxnLv4Inst159_io_z; // @[Snxn100k.scala 14148:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst156_io_z + inst_SnxnLv4Inst157_io_z; // @[Snxn100k.scala 14152:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst158_io_z; // @[Snxn100k.scala 14152:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst159_io_z; // @[Snxn100k.scala 14152:92]
  SnxnLv4Inst7 inst_SnxnLv4Inst156 ( // @[Snxn100k.scala 14136:35]
    .io_a(inst_SnxnLv4Inst156_io_a),
    .io_b(inst_SnxnLv4Inst156_io_b),
    .io_z(inst_SnxnLv4Inst156_io_z)
  );
  SnxnLv4Inst103 inst_SnxnLv4Inst157 ( // @[Snxn100k.scala 14140:35]
    .io_a(inst_SnxnLv4Inst157_io_a),
    .io_b(inst_SnxnLv4Inst157_io_b),
    .io_z(inst_SnxnLv4Inst157_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst158 ( // @[Snxn100k.scala 14144:35]
    .io_a(inst_SnxnLv4Inst158_io_a),
    .io_b(inst_SnxnLv4Inst158_io_b),
    .io_z(inst_SnxnLv4Inst158_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst159 ( // @[Snxn100k.scala 14148:35]
    .io_a(inst_SnxnLv4Inst159_io_a),
    .io_b(inst_SnxnLv4Inst159_io_b),
    .io_z(inst_SnxnLv4Inst159_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14153:15]
  assign inst_SnxnLv4Inst156_io_a = io_a; // @[Snxn100k.scala 14137:28]
  assign inst_SnxnLv4Inst156_io_b = io_b; // @[Snxn100k.scala 14138:28]
  assign inst_SnxnLv4Inst157_io_a = io_a; // @[Snxn100k.scala 14141:28]
  assign inst_SnxnLv4Inst157_io_b = io_b; // @[Snxn100k.scala 14142:28]
  assign inst_SnxnLv4Inst158_io_a = io_a; // @[Snxn100k.scala 14145:28]
  assign inst_SnxnLv4Inst158_io_b = io_b; // @[Snxn100k.scala 14146:28]
  assign inst_SnxnLv4Inst159_io_a = io_a; // @[Snxn100k.scala 14149:28]
  assign inst_SnxnLv4Inst159_io_b = io_b; // @[Snxn100k.scala 14150:28]
endmodule
module SnxnLv2Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst36_io_a; // @[Snxn100k.scala 3243:34]
  wire  inst_SnxnLv3Inst36_io_b; // @[Snxn100k.scala 3243:34]
  wire  inst_SnxnLv3Inst36_io_z; // @[Snxn100k.scala 3243:34]
  wire  inst_SnxnLv3Inst37_io_a; // @[Snxn100k.scala 3247:34]
  wire  inst_SnxnLv3Inst37_io_b; // @[Snxn100k.scala 3247:34]
  wire  inst_SnxnLv3Inst37_io_z; // @[Snxn100k.scala 3247:34]
  wire  inst_SnxnLv3Inst38_io_a; // @[Snxn100k.scala 3251:34]
  wire  inst_SnxnLv3Inst38_io_b; // @[Snxn100k.scala 3251:34]
  wire  inst_SnxnLv3Inst38_io_z; // @[Snxn100k.scala 3251:34]
  wire  inst_SnxnLv3Inst39_io_a; // @[Snxn100k.scala 3255:34]
  wire  inst_SnxnLv3Inst39_io_b; // @[Snxn100k.scala 3255:34]
  wire  inst_SnxnLv3Inst39_io_z; // @[Snxn100k.scala 3255:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst36_io_z + inst_SnxnLv3Inst37_io_z; // @[Snxn100k.scala 3259:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst38_io_z; // @[Snxn100k.scala 3259:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst39_io_z; // @[Snxn100k.scala 3259:89]
  SnxnLv3Inst36 inst_SnxnLv3Inst36 ( // @[Snxn100k.scala 3243:34]
    .io_a(inst_SnxnLv3Inst36_io_a),
    .io_b(inst_SnxnLv3Inst36_io_b),
    .io_z(inst_SnxnLv3Inst36_io_z)
  );
  SnxnLv3Inst37 inst_SnxnLv3Inst37 ( // @[Snxn100k.scala 3247:34]
    .io_a(inst_SnxnLv3Inst37_io_a),
    .io_b(inst_SnxnLv3Inst37_io_b),
    .io_z(inst_SnxnLv3Inst37_io_z)
  );
  SnxnLv3Inst38 inst_SnxnLv3Inst38 ( // @[Snxn100k.scala 3251:34]
    .io_a(inst_SnxnLv3Inst38_io_a),
    .io_b(inst_SnxnLv3Inst38_io_b),
    .io_z(inst_SnxnLv3Inst38_io_z)
  );
  SnxnLv3Inst39 inst_SnxnLv3Inst39 ( // @[Snxn100k.scala 3255:34]
    .io_a(inst_SnxnLv3Inst39_io_a),
    .io_b(inst_SnxnLv3Inst39_io_b),
    .io_z(inst_SnxnLv3Inst39_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 3260:15]
  assign inst_SnxnLv3Inst36_io_a = io_a; // @[Snxn100k.scala 3244:27]
  assign inst_SnxnLv3Inst36_io_b = io_b; // @[Snxn100k.scala 3245:27]
  assign inst_SnxnLv3Inst37_io_a = io_a; // @[Snxn100k.scala 3248:27]
  assign inst_SnxnLv3Inst37_io_b = io_b; // @[Snxn100k.scala 3249:27]
  assign inst_SnxnLv3Inst38_io_a = io_a; // @[Snxn100k.scala 3252:27]
  assign inst_SnxnLv3Inst38_io_b = io_b; // @[Snxn100k.scala 3253:27]
  assign inst_SnxnLv3Inst39_io_a = io_a; // @[Snxn100k.scala 3256:27]
  assign inst_SnxnLv3Inst39_io_b = io_b; // @[Snxn100k.scala 3257:27]
endmodule
module SnxnLv4Inst161(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 66538:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 66539:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 66540:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 66541:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 66542:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 66543:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 66544:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 66545:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 66546:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 66547:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 66548:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 66549:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 66550:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 66551:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 66552:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 66553:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 66554:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 66555:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 66556:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 66557:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 66558:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 66559:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 66560:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 66561:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 66562:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 66563:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 66564:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 66565:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 66566:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 66567:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 66568:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 66569:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 66570:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 66571:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 66572:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 66573:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 66574:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 66575:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 66576:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 66577:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 66578:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 66579:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 66580:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 66581:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 66582:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 66583:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 66584:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 66585:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 66586:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 66587:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 66588:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 66589:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 66590:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 66591:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 66592:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 66593:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 66594:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 66595:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 66596:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 66597:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 66598:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 66599:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 66600:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 66601:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 66602:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 66603:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 66604:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 66605:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 66606:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 66607:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 66608:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 66609:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 66610:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 66611:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 66612:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 66613:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 66614:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 66615:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 66616:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 66617:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 66618:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 66619:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 66620:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 66621:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 66622:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 66623:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 66624:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 66625:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 66626:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 66627:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 66628:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 66629:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 66630:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 66631:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 66632:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 66633:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 66634:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 66635:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 66636:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 66637:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 66638:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 66639:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 66640:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 66641:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 66642:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 66643:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 66644:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 66645:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 66646:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 66647:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 66648:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 66649:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 66650:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 66651:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 66652:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 66653:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 66654:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 66655:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 66656:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 66657:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 66658:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 66659:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 66660:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 66661:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 66662:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 66663:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 66664:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 66665:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 66666:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 66667:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 66668:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 66669:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 66670:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 66671:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 66672:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 66673:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 66674:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 66675:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 66676:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 66677:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 66678:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 66679:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 66680:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 66681:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 66682:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 66683:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 66684:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 66685:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 66686:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 66687:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 66688:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 66689:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 66690:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 66691:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 66692:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 66693:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 66694:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 66695:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 66696:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 66697:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 66698:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 66699:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 66700:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 66701:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 66702:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 66703:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 66704:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 66705:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 66706:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 66707:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 66708:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 66709:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 66710:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 66711:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 66712:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 66713:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 66714:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 66715:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 66716:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 66717:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 66718:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 66719:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 66720:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 66721:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 66722:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 66723:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 66724:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 66725:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 66726:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 66727:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 66728:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 66729:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 66730:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 66731:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 66732:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 66733:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 66734:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 66735:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 66736:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 66737:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 66738:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 66739:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 66740:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 66741:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 66742:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 66743:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 66744:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 66745:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 66746:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 66747:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 66748:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 66749:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 66750:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 66751:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 66752:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 66753:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 66754:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 66755:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 66756:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 66757:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 66758:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 66759:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 66760:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 66761:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 66762:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 66763:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 66764:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 66765:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 66766:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 66767:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 66768:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 66769:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 66770:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 66771:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 66772:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 66773:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 66774:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 66775:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 66776:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 66777:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 66778:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 66779:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 66780:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 66781:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 66782:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 66783:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 66784:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 66785:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 66786:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 66787:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 66788:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 66789:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 66790:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 66791:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 66792:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 66793:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 66794:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 66795:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 66796:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 66797:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 66798:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 66799:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 66800:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 66801:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 66802:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 66803:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 66804:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 66805:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 66806:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 66807:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 66808:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 66809:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 66810:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 66811:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 66812:20]
  assign io_z = ~x68; // @[Snxn100k.scala 66813:16]
endmodule
module SnxnLv3Inst40(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst160_io_a; // @[Snxn100k.scala 17942:35]
  wire  inst_SnxnLv4Inst160_io_b; // @[Snxn100k.scala 17942:35]
  wire  inst_SnxnLv4Inst160_io_z; // @[Snxn100k.scala 17942:35]
  wire  inst_SnxnLv4Inst161_io_a; // @[Snxn100k.scala 17946:35]
  wire  inst_SnxnLv4Inst161_io_b; // @[Snxn100k.scala 17946:35]
  wire  inst_SnxnLv4Inst161_io_z; // @[Snxn100k.scala 17946:35]
  wire  inst_SnxnLv4Inst162_io_a; // @[Snxn100k.scala 17950:35]
  wire  inst_SnxnLv4Inst162_io_b; // @[Snxn100k.scala 17950:35]
  wire  inst_SnxnLv4Inst162_io_z; // @[Snxn100k.scala 17950:35]
  wire  inst_SnxnLv4Inst163_io_a; // @[Snxn100k.scala 17954:35]
  wire  inst_SnxnLv4Inst163_io_b; // @[Snxn100k.scala 17954:35]
  wire  inst_SnxnLv4Inst163_io_z; // @[Snxn100k.scala 17954:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst160_io_z + inst_SnxnLv4Inst161_io_z; // @[Snxn100k.scala 17958:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst162_io_z; // @[Snxn100k.scala 17958:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst163_io_z; // @[Snxn100k.scala 17958:92]
  SnxnLv4Inst68 inst_SnxnLv4Inst160 ( // @[Snxn100k.scala 17942:35]
    .io_a(inst_SnxnLv4Inst160_io_a),
    .io_b(inst_SnxnLv4Inst160_io_b),
    .io_z(inst_SnxnLv4Inst160_io_z)
  );
  SnxnLv4Inst161 inst_SnxnLv4Inst161 ( // @[Snxn100k.scala 17946:35]
    .io_a(inst_SnxnLv4Inst161_io_a),
    .io_b(inst_SnxnLv4Inst161_io_b),
    .io_z(inst_SnxnLv4Inst161_io_z)
  );
  SnxnLv4Inst43 inst_SnxnLv4Inst162 ( // @[Snxn100k.scala 17950:35]
    .io_a(inst_SnxnLv4Inst162_io_a),
    .io_b(inst_SnxnLv4Inst162_io_b),
    .io_z(inst_SnxnLv4Inst162_io_z)
  );
  SnxnLv4Inst129 inst_SnxnLv4Inst163 ( // @[Snxn100k.scala 17954:35]
    .io_a(inst_SnxnLv4Inst163_io_a),
    .io_b(inst_SnxnLv4Inst163_io_b),
    .io_z(inst_SnxnLv4Inst163_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17959:15]
  assign inst_SnxnLv4Inst160_io_a = io_a; // @[Snxn100k.scala 17943:28]
  assign inst_SnxnLv4Inst160_io_b = io_b; // @[Snxn100k.scala 17944:28]
  assign inst_SnxnLv4Inst161_io_a = io_a; // @[Snxn100k.scala 17947:28]
  assign inst_SnxnLv4Inst161_io_b = io_b; // @[Snxn100k.scala 17948:28]
  assign inst_SnxnLv4Inst162_io_a = io_a; // @[Snxn100k.scala 17951:28]
  assign inst_SnxnLv4Inst162_io_b = io_b; // @[Snxn100k.scala 17952:28]
  assign inst_SnxnLv4Inst163_io_a = io_a; // @[Snxn100k.scala 17955:28]
  assign inst_SnxnLv4Inst163_io_b = io_b; // @[Snxn100k.scala 17956:28]
endmodule
module SnxnLv3Inst41(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst164_io_a; // @[Snxn100k.scala 18061:35]
  wire  inst_SnxnLv4Inst164_io_b; // @[Snxn100k.scala 18061:35]
  wire  inst_SnxnLv4Inst164_io_z; // @[Snxn100k.scala 18061:35]
  wire  inst_SnxnLv4Inst165_io_a; // @[Snxn100k.scala 18065:35]
  wire  inst_SnxnLv4Inst165_io_b; // @[Snxn100k.scala 18065:35]
  wire  inst_SnxnLv4Inst165_io_z; // @[Snxn100k.scala 18065:35]
  wire  inst_SnxnLv4Inst166_io_a; // @[Snxn100k.scala 18069:35]
  wire  inst_SnxnLv4Inst166_io_b; // @[Snxn100k.scala 18069:35]
  wire  inst_SnxnLv4Inst166_io_z; // @[Snxn100k.scala 18069:35]
  wire  inst_SnxnLv4Inst167_io_a; // @[Snxn100k.scala 18073:35]
  wire  inst_SnxnLv4Inst167_io_b; // @[Snxn100k.scala 18073:35]
  wire  inst_SnxnLv4Inst167_io_z; // @[Snxn100k.scala 18073:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst164_io_z + inst_SnxnLv4Inst165_io_z; // @[Snxn100k.scala 18077:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst166_io_z; // @[Snxn100k.scala 18077:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst167_io_z; // @[Snxn100k.scala 18077:92]
  SnxnLv4Inst3 inst_SnxnLv4Inst164 ( // @[Snxn100k.scala 18061:35]
    .io_a(inst_SnxnLv4Inst164_io_a),
    .io_b(inst_SnxnLv4Inst164_io_b),
    .io_z(inst_SnxnLv4Inst164_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst165 ( // @[Snxn100k.scala 18065:35]
    .io_a(inst_SnxnLv4Inst165_io_a),
    .io_b(inst_SnxnLv4Inst165_io_b),
    .io_z(inst_SnxnLv4Inst165_io_z)
  );
  SnxnLv4Inst118 inst_SnxnLv4Inst166 ( // @[Snxn100k.scala 18069:35]
    .io_a(inst_SnxnLv4Inst166_io_a),
    .io_b(inst_SnxnLv4Inst166_io_b),
    .io_z(inst_SnxnLv4Inst166_io_z)
  );
  SnxnLv4Inst117 inst_SnxnLv4Inst167 ( // @[Snxn100k.scala 18073:35]
    .io_a(inst_SnxnLv4Inst167_io_a),
    .io_b(inst_SnxnLv4Inst167_io_b),
    .io_z(inst_SnxnLv4Inst167_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 18078:15]
  assign inst_SnxnLv4Inst164_io_a = io_a; // @[Snxn100k.scala 18062:28]
  assign inst_SnxnLv4Inst164_io_b = io_b; // @[Snxn100k.scala 18063:28]
  assign inst_SnxnLv4Inst165_io_a = io_a; // @[Snxn100k.scala 18066:28]
  assign inst_SnxnLv4Inst165_io_b = io_b; // @[Snxn100k.scala 18067:28]
  assign inst_SnxnLv4Inst166_io_a = io_a; // @[Snxn100k.scala 18070:28]
  assign inst_SnxnLv4Inst166_io_b = io_b; // @[Snxn100k.scala 18071:28]
  assign inst_SnxnLv4Inst167_io_a = io_a; // @[Snxn100k.scala 18074:28]
  assign inst_SnxnLv4Inst167_io_b = io_b; // @[Snxn100k.scala 18075:28]
endmodule
module SnxnLv4Inst168(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 65488:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 65489:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 65490:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 65491:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 65492:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 65493:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 65494:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 65495:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 65496:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 65497:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 65498:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 65499:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 65500:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 65501:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 65502:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 65503:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 65504:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 65505:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 65506:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 65507:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 65508:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 65509:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 65510:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 65511:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 65512:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 65513:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 65514:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 65515:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 65516:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 65517:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 65518:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 65519:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 65520:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 65521:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 65522:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 65523:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 65524:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 65525:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 65526:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 65527:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 65528:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 65529:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 65530:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 65531:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 65532:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 65533:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 65534:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 65535:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 65536:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 65537:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 65538:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 65539:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 65540:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 65541:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 65542:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 65543:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 65544:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 65545:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 65546:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 65547:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 65548:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 65549:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 65550:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 65551:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 65552:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 65553:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 65554:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 65555:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 65556:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 65557:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 65558:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 65559:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 65560:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 65561:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 65562:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 65563:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 65564:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 65565:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 65566:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 65567:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 65568:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 65569:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 65570:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 65571:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 65572:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 65573:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 65574:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 65575:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 65576:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 65577:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 65578:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 65579:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 65580:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 65581:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 65582:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 65583:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 65584:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 65585:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 65586:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 65587:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 65588:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 65589:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 65590:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 65591:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 65592:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 65593:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 65594:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 65595:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 65596:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 65597:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 65598:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 65599:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 65600:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 65601:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 65602:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 65603:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 65604:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 65605:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 65606:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 65607:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 65608:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 65609:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 65610:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 65611:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 65612:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 65613:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 65614:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 65615:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 65616:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 65617:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 65618:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 65619:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 65620:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 65621:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 65622:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 65623:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 65624:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 65625:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 65626:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 65627:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 65628:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 65629:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 65630:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 65631:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 65632:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 65633:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 65634:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 65635:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 65636:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 65637:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 65638:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 65639:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 65640:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 65641:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 65642:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 65643:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 65644:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 65645:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 65646:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 65647:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 65648:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 65649:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 65650:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 65651:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 65652:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 65653:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 65654:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 65655:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 65656:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 65657:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 65658:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 65659:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 65660:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 65661:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 65662:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 65663:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 65664:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 65665:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 65666:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 65667:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 65668:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 65669:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 65670:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 65671:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 65672:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 65673:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 65674:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 65675:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 65676:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 65677:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 65678:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 65679:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 65680:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 65681:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 65682:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 65683:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 65684:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 65685:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 65686:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 65687:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 65688:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 65689:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 65690:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 65691:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 65692:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 65693:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 65694:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 65695:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 65696:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 65697:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 65698:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 65699:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 65700:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 65701:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 65702:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 65703:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 65704:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 65705:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 65706:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 65707:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 65708:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 65709:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 65710:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 65711:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 65712:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 65713:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 65714:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 65715:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 65716:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 65717:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 65718:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 65719:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 65720:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 65721:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 65722:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 65723:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 65724:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 65725:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 65726:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 65727:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 65728:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 65729:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 65730:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 65731:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 65732:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 65733:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 65734:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 65735:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 65736:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 65737:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 65738:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 65739:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 65740:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 65741:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 65742:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 65743:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 65744:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 65745:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 65746:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 65747:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 65748:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 65749:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 65750:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 65751:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 65752:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 65753:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 65754:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 65755:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 65756:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 65757:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 65758:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 65759:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 65760:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 65761:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 65762:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 65763:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 65764:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 65765:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 65766:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 65767:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 65768:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 65769:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 65770:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 65771:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 65772:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 65773:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 65774:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 65775:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 65776:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 65777:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 65778:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 65779:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 65780:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 65781:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 65782:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 65783:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 65784:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 65785:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 65786:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 65787:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 65788:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 65789:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 65790:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 65791:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 65792:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 65793:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 65794:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 65795:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 65796:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 65797:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 65798:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 65799:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 65800:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 65801:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 65802:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 65803:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 65804:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 65805:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 65806:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 65807:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 65808:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 65809:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 65810:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 65811:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 65812:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 65813:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 65814:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 65815:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 65816:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 65817:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 65818:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 65819:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 65820:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 65821:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 65822:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 65823:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 65824:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 65825:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 65826:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 65827:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 65828:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 65829:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 65830:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 65831:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 65832:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 65833:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 65834:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 65835:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 65836:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 65837:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 65838:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 65839:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 65840:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 65841:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 65842:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 65843:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 65844:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 65845:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 65846:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 65847:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 65848:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 65849:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 65850:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 65851:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 65852:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 65853:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 65854:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 65855:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 65856:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 65857:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 65858:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 65859:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 65860:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 65861:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 65862:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 65863:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 65864:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 65865:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 65866:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 65867:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 65868:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 65869:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 65870:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 65871:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 65872:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 65873:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 65874:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 65875:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 65876:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 65877:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 65878:20]
  assign io_z = ~x97; // @[Snxn100k.scala 65879:16]
endmodule
module SnxnLv3Inst42(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst168_io_a; // @[Snxn100k.scala 17463:35]
  wire  inst_SnxnLv4Inst168_io_b; // @[Snxn100k.scala 17463:35]
  wire  inst_SnxnLv4Inst168_io_z; // @[Snxn100k.scala 17463:35]
  wire  inst_SnxnLv4Inst169_io_a; // @[Snxn100k.scala 17467:35]
  wire  inst_SnxnLv4Inst169_io_b; // @[Snxn100k.scala 17467:35]
  wire  inst_SnxnLv4Inst169_io_z; // @[Snxn100k.scala 17467:35]
  wire  inst_SnxnLv4Inst170_io_a; // @[Snxn100k.scala 17471:35]
  wire  inst_SnxnLv4Inst170_io_b; // @[Snxn100k.scala 17471:35]
  wire  inst_SnxnLv4Inst170_io_z; // @[Snxn100k.scala 17471:35]
  wire  inst_SnxnLv4Inst171_io_a; // @[Snxn100k.scala 17475:35]
  wire  inst_SnxnLv4Inst171_io_b; // @[Snxn100k.scala 17475:35]
  wire  inst_SnxnLv4Inst171_io_z; // @[Snxn100k.scala 17475:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst168_io_z + inst_SnxnLv4Inst169_io_z; // @[Snxn100k.scala 17479:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst170_io_z; // @[Snxn100k.scala 17479:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst171_io_z; // @[Snxn100k.scala 17479:92]
  SnxnLv4Inst168 inst_SnxnLv4Inst168 ( // @[Snxn100k.scala 17463:35]
    .io_a(inst_SnxnLv4Inst168_io_a),
    .io_b(inst_SnxnLv4Inst168_io_b),
    .io_z(inst_SnxnLv4Inst168_io_z)
  );
  SnxnLv4Inst68 inst_SnxnLv4Inst169 ( // @[Snxn100k.scala 17467:35]
    .io_a(inst_SnxnLv4Inst169_io_a),
    .io_b(inst_SnxnLv4Inst169_io_b),
    .io_z(inst_SnxnLv4Inst169_io_z)
  );
  SnxnLv4Inst118 inst_SnxnLv4Inst170 ( // @[Snxn100k.scala 17471:35]
    .io_a(inst_SnxnLv4Inst170_io_a),
    .io_b(inst_SnxnLv4Inst170_io_b),
    .io_z(inst_SnxnLv4Inst170_io_z)
  );
  SnxnLv4Inst103 inst_SnxnLv4Inst171 ( // @[Snxn100k.scala 17475:35]
    .io_a(inst_SnxnLv4Inst171_io_a),
    .io_b(inst_SnxnLv4Inst171_io_b),
    .io_z(inst_SnxnLv4Inst171_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17480:15]
  assign inst_SnxnLv4Inst168_io_a = io_a; // @[Snxn100k.scala 17464:28]
  assign inst_SnxnLv4Inst168_io_b = io_b; // @[Snxn100k.scala 17465:28]
  assign inst_SnxnLv4Inst169_io_a = io_a; // @[Snxn100k.scala 17468:28]
  assign inst_SnxnLv4Inst169_io_b = io_b; // @[Snxn100k.scala 17469:28]
  assign inst_SnxnLv4Inst170_io_a = io_a; // @[Snxn100k.scala 17472:28]
  assign inst_SnxnLv4Inst170_io_b = io_b; // @[Snxn100k.scala 17473:28]
  assign inst_SnxnLv4Inst171_io_a = io_a; // @[Snxn100k.scala 17476:28]
  assign inst_SnxnLv4Inst171_io_b = io_b; // @[Snxn100k.scala 17477:28]
endmodule
module SnxnLv4Inst173(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 63956:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 63957:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 63958:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 63959:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 63960:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 63961:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 63962:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 63963:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 63964:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 63965:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 63966:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 63967:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 63968:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 63969:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 63970:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 63971:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 63972:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 63973:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 63974:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 63975:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 63976:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 63977:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 63978:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 63979:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 63980:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 63981:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 63982:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 63983:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 63984:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 63985:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 63986:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 63987:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 63988:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 63989:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 63990:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 63991:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 63992:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 63993:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 63994:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 63995:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 63996:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 63997:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 63998:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 63999:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 64000:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 64001:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 64002:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 64003:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 64004:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 64005:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 64006:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 64007:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 64008:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 64009:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 64010:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 64011:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 64012:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 64013:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 64014:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 64015:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 64016:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 64017:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 64018:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 64019:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 64020:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 64021:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 64022:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 64023:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 64024:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 64025:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 64026:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 64027:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 64028:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 64029:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 64030:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 64031:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 64032:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 64033:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 64034:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 64035:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 64036:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 64037:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 64038:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 64039:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 64040:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 64041:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 64042:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 64043:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 64044:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 64045:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 64046:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 64047:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 64048:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 64049:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 64050:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 64051:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 64052:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 64053:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 64054:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 64055:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 64056:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 64057:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 64058:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 64059:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 64060:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 64061:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 64062:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 64063:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 64064:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 64065:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 64066:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 64067:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 64068:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 64069:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 64070:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 64071:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 64072:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 64073:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 64074:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 64075:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 64076:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 64077:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 64078:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 64079:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 64080:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 64081:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 64082:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 64083:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 64084:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 64085:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 64086:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 64087:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 64088:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 64089:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 64090:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 64091:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 64092:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 64093:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 64094:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 64095:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 64096:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 64097:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 64098:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 64099:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 64100:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 64101:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 64102:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 64103:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 64104:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 64105:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 64106:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 64107:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 64108:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 64109:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 64110:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 64111:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 64112:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 64113:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 64114:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 64115:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 64116:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 64117:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 64118:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 64119:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 64120:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 64121:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 64122:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 64123:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 64124:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 64125:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 64126:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 64127:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 64128:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 64129:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 64130:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 64131:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 64132:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 64133:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 64134:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 64135:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 64136:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 64137:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 64138:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 64139:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 64140:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 64141:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 64142:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 64143:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 64144:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 64145:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 64146:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 64147:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 64148:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 64149:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 64150:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 64151:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 64152:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 64153:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 64154:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 64155:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 64156:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 64157:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 64158:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 64159:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 64160:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 64161:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 64162:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 64163:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 64164:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 64165:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 64166:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 64167:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 64168:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 64169:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 64170:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 64171:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 64172:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 64173:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 64174:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 64175:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 64176:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 64177:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 64178:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 64179:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 64180:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 64181:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 64182:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 64183:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 64184:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 64185:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 64186:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 64187:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 64188:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 64189:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 64190:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 64191:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 64192:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 64193:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 64194:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 64195:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 64196:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 64197:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 64198:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 64199:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 64200:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 64201:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 64202:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 64203:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 64204:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 64205:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 64206:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 64207:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 64208:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 64209:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 64210:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 64211:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 64212:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 64213:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 64214:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 64215:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 64216:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 64217:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 64218:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 64219:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 64220:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 64221:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 64222:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 64223:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 64224:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 64225:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 64226:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 64227:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 64228:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 64229:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 64230:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 64231:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 64232:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 64233:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 64234:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 64235:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 64236:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 64237:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 64238:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 64239:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 64240:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 64241:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 64242:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 64243:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 64244:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 64245:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 64246:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 64247:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 64248:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 64249:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 64250:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 64251:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 64252:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 64253:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 64254:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 64255:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 64256:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 64257:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 64258:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 64259:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 64260:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 64261:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 64262:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 64263:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 64264:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 64265:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 64266:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 64267:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 64268:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 64269:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 64270:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 64271:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 64272:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 64273:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 64274:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 64275:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 64276:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 64277:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 64278:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 64279:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 64280:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 64281:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 64282:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 64283:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 64284:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 64285:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 64286:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 64287:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 64288:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 64289:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 64290:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 64291:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 64292:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 64293:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 64294:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 64295:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 64296:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 64297:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 64298:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 64299:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 64300:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 64301:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 64302:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 64303:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 64304:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 64305:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 64306:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 64307:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 64308:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 64309:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 64310:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 64311:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 64312:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 64313:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 64314:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 64315:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 64316:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 64317:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 64318:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 64319:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 64320:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 64321:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 64322:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 64323:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 64324:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 64325:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 64326:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 64327:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 64328:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 64329:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 64330:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 64331:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 64332:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 64333:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 64334:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 64335:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 64336:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 64337:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 64338:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 64339:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 64340:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 64341:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 64342:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 64343:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 64344:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 64345:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 64346:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 64347:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 64348:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 64349:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 64350:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 64351:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 64352:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 64353:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 64354:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 64355:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 64356:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 64357:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 64358:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 64359:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 64360:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 64361:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 64362:22]
  assign io_z = ~x101; // @[Snxn100k.scala 64363:17]
endmodule
module SnxnLv3Inst43(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst172_io_a; // @[Snxn100k.scala 16984:35]
  wire  inst_SnxnLv4Inst172_io_b; // @[Snxn100k.scala 16984:35]
  wire  inst_SnxnLv4Inst172_io_z; // @[Snxn100k.scala 16984:35]
  wire  inst_SnxnLv4Inst173_io_a; // @[Snxn100k.scala 16988:35]
  wire  inst_SnxnLv4Inst173_io_b; // @[Snxn100k.scala 16988:35]
  wire  inst_SnxnLv4Inst173_io_z; // @[Snxn100k.scala 16988:35]
  wire  inst_SnxnLv4Inst174_io_a; // @[Snxn100k.scala 16992:35]
  wire  inst_SnxnLv4Inst174_io_b; // @[Snxn100k.scala 16992:35]
  wire  inst_SnxnLv4Inst174_io_z; // @[Snxn100k.scala 16992:35]
  wire  inst_SnxnLv4Inst175_io_a; // @[Snxn100k.scala 16996:35]
  wire  inst_SnxnLv4Inst175_io_b; // @[Snxn100k.scala 16996:35]
  wire  inst_SnxnLv4Inst175_io_z; // @[Snxn100k.scala 16996:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst172_io_z + inst_SnxnLv4Inst173_io_z; // @[Snxn100k.scala 17000:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst174_io_z; // @[Snxn100k.scala 17000:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst175_io_z; // @[Snxn100k.scala 17000:92]
  SnxnLv4Inst34 inst_SnxnLv4Inst172 ( // @[Snxn100k.scala 16984:35]
    .io_a(inst_SnxnLv4Inst172_io_a),
    .io_b(inst_SnxnLv4Inst172_io_b),
    .io_z(inst_SnxnLv4Inst172_io_z)
  );
  SnxnLv4Inst173 inst_SnxnLv4Inst173 ( // @[Snxn100k.scala 16988:35]
    .io_a(inst_SnxnLv4Inst173_io_a),
    .io_b(inst_SnxnLv4Inst173_io_b),
    .io_z(inst_SnxnLv4Inst173_io_z)
  );
  SnxnLv4Inst43 inst_SnxnLv4Inst174 ( // @[Snxn100k.scala 16992:35]
    .io_a(inst_SnxnLv4Inst174_io_a),
    .io_b(inst_SnxnLv4Inst174_io_b),
    .io_z(inst_SnxnLv4Inst174_io_z)
  );
  SnxnLv4Inst148 inst_SnxnLv4Inst175 ( // @[Snxn100k.scala 16996:35]
    .io_a(inst_SnxnLv4Inst175_io_a),
    .io_b(inst_SnxnLv4Inst175_io_b),
    .io_z(inst_SnxnLv4Inst175_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17001:15]
  assign inst_SnxnLv4Inst172_io_a = io_a; // @[Snxn100k.scala 16985:28]
  assign inst_SnxnLv4Inst172_io_b = io_b; // @[Snxn100k.scala 16986:28]
  assign inst_SnxnLv4Inst173_io_a = io_a; // @[Snxn100k.scala 16989:28]
  assign inst_SnxnLv4Inst173_io_b = io_b; // @[Snxn100k.scala 16990:28]
  assign inst_SnxnLv4Inst174_io_a = io_a; // @[Snxn100k.scala 16993:28]
  assign inst_SnxnLv4Inst174_io_b = io_b; // @[Snxn100k.scala 16994:28]
  assign inst_SnxnLv4Inst175_io_a = io_a; // @[Snxn100k.scala 16997:28]
  assign inst_SnxnLv4Inst175_io_b = io_b; // @[Snxn100k.scala 16998:28]
endmodule
module SnxnLv2Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst40_io_a; // @[Snxn100k.scala 3865:34]
  wire  inst_SnxnLv3Inst40_io_b; // @[Snxn100k.scala 3865:34]
  wire  inst_SnxnLv3Inst40_io_z; // @[Snxn100k.scala 3865:34]
  wire  inst_SnxnLv3Inst41_io_a; // @[Snxn100k.scala 3869:34]
  wire  inst_SnxnLv3Inst41_io_b; // @[Snxn100k.scala 3869:34]
  wire  inst_SnxnLv3Inst41_io_z; // @[Snxn100k.scala 3869:34]
  wire  inst_SnxnLv3Inst42_io_a; // @[Snxn100k.scala 3873:34]
  wire  inst_SnxnLv3Inst42_io_b; // @[Snxn100k.scala 3873:34]
  wire  inst_SnxnLv3Inst42_io_z; // @[Snxn100k.scala 3873:34]
  wire  inst_SnxnLv3Inst43_io_a; // @[Snxn100k.scala 3877:34]
  wire  inst_SnxnLv3Inst43_io_b; // @[Snxn100k.scala 3877:34]
  wire  inst_SnxnLv3Inst43_io_z; // @[Snxn100k.scala 3877:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst40_io_z + inst_SnxnLv3Inst41_io_z; // @[Snxn100k.scala 3881:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst42_io_z; // @[Snxn100k.scala 3881:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst43_io_z; // @[Snxn100k.scala 3881:89]
  SnxnLv3Inst40 inst_SnxnLv3Inst40 ( // @[Snxn100k.scala 3865:34]
    .io_a(inst_SnxnLv3Inst40_io_a),
    .io_b(inst_SnxnLv3Inst40_io_b),
    .io_z(inst_SnxnLv3Inst40_io_z)
  );
  SnxnLv3Inst41 inst_SnxnLv3Inst41 ( // @[Snxn100k.scala 3869:34]
    .io_a(inst_SnxnLv3Inst41_io_a),
    .io_b(inst_SnxnLv3Inst41_io_b),
    .io_z(inst_SnxnLv3Inst41_io_z)
  );
  SnxnLv3Inst42 inst_SnxnLv3Inst42 ( // @[Snxn100k.scala 3873:34]
    .io_a(inst_SnxnLv3Inst42_io_a),
    .io_b(inst_SnxnLv3Inst42_io_b),
    .io_z(inst_SnxnLv3Inst42_io_z)
  );
  SnxnLv3Inst43 inst_SnxnLv3Inst43 ( // @[Snxn100k.scala 3877:34]
    .io_a(inst_SnxnLv3Inst43_io_a),
    .io_b(inst_SnxnLv3Inst43_io_b),
    .io_z(inst_SnxnLv3Inst43_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 3882:15]
  assign inst_SnxnLv3Inst40_io_a = io_a; // @[Snxn100k.scala 3866:27]
  assign inst_SnxnLv3Inst40_io_b = io_b; // @[Snxn100k.scala 3867:27]
  assign inst_SnxnLv3Inst41_io_a = io_a; // @[Snxn100k.scala 3870:27]
  assign inst_SnxnLv3Inst41_io_b = io_b; // @[Snxn100k.scala 3871:27]
  assign inst_SnxnLv3Inst42_io_a = io_a; // @[Snxn100k.scala 3874:27]
  assign inst_SnxnLv3Inst42_io_b = io_b; // @[Snxn100k.scala 3875:27]
  assign inst_SnxnLv3Inst43_io_a = io_a; // @[Snxn100k.scala 3878:27]
  assign inst_SnxnLv3Inst43_io_b = io_b; // @[Snxn100k.scala 3879:27]
endmodule
module SnxnLv3Inst44(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst176_io_a; // @[Snxn100k.scala 16633:35]
  wire  inst_SnxnLv4Inst176_io_b; // @[Snxn100k.scala 16633:35]
  wire  inst_SnxnLv4Inst176_io_z; // @[Snxn100k.scala 16633:35]
  wire  inst_SnxnLv4Inst177_io_a; // @[Snxn100k.scala 16637:35]
  wire  inst_SnxnLv4Inst177_io_b; // @[Snxn100k.scala 16637:35]
  wire  inst_SnxnLv4Inst177_io_z; // @[Snxn100k.scala 16637:35]
  wire  inst_SnxnLv4Inst178_io_a; // @[Snxn100k.scala 16641:35]
  wire  inst_SnxnLv4Inst178_io_b; // @[Snxn100k.scala 16641:35]
  wire  inst_SnxnLv4Inst178_io_z; // @[Snxn100k.scala 16641:35]
  wire  inst_SnxnLv4Inst179_io_a; // @[Snxn100k.scala 16645:35]
  wire  inst_SnxnLv4Inst179_io_b; // @[Snxn100k.scala 16645:35]
  wire  inst_SnxnLv4Inst179_io_z; // @[Snxn100k.scala 16645:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst176_io_z + inst_SnxnLv4Inst177_io_z; // @[Snxn100k.scala 16649:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst178_io_z; // @[Snxn100k.scala 16649:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst179_io_z; // @[Snxn100k.scala 16649:92]
  SnxnLv4Inst15 inst_SnxnLv4Inst176 ( // @[Snxn100k.scala 16633:35]
    .io_a(inst_SnxnLv4Inst176_io_a),
    .io_b(inst_SnxnLv4Inst176_io_b),
    .io_z(inst_SnxnLv4Inst176_io_z)
  );
  SnxnLv4Inst105 inst_SnxnLv4Inst177 ( // @[Snxn100k.scala 16637:35]
    .io_a(inst_SnxnLv4Inst177_io_a),
    .io_b(inst_SnxnLv4Inst177_io_b),
    .io_z(inst_SnxnLv4Inst177_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst178 ( // @[Snxn100k.scala 16641:35]
    .io_a(inst_SnxnLv4Inst178_io_a),
    .io_b(inst_SnxnLv4Inst178_io_b),
    .io_z(inst_SnxnLv4Inst178_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst179 ( // @[Snxn100k.scala 16645:35]
    .io_a(inst_SnxnLv4Inst179_io_a),
    .io_b(inst_SnxnLv4Inst179_io_b),
    .io_z(inst_SnxnLv4Inst179_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 16650:15]
  assign inst_SnxnLv4Inst176_io_a = io_a; // @[Snxn100k.scala 16634:28]
  assign inst_SnxnLv4Inst176_io_b = io_b; // @[Snxn100k.scala 16635:28]
  assign inst_SnxnLv4Inst177_io_a = io_a; // @[Snxn100k.scala 16638:28]
  assign inst_SnxnLv4Inst177_io_b = io_b; // @[Snxn100k.scala 16639:28]
  assign inst_SnxnLv4Inst178_io_a = io_a; // @[Snxn100k.scala 16642:28]
  assign inst_SnxnLv4Inst178_io_b = io_b; // @[Snxn100k.scala 16643:28]
  assign inst_SnxnLv4Inst179_io_a = io_a; // @[Snxn100k.scala 16646:28]
  assign inst_SnxnLv4Inst179_io_b = io_b; // @[Snxn100k.scala 16647:28]
endmodule
module SnxnLv4Inst180(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 59058:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 59059:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 59060:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 59061:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 59062:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 59063:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 59064:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 59065:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 59066:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 59067:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 59068:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 59069:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 59070:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 59071:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 59072:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 59073:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 59074:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 59075:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 59076:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 59077:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 59078:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 59079:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 59080:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 59081:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 59082:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 59083:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 59084:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 59085:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 59086:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 59087:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 59088:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 59089:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 59090:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 59091:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 59092:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 59093:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 59094:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 59095:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 59096:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 59097:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 59098:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 59099:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 59100:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 59101:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 59102:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 59103:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 59104:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 59105:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 59106:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 59107:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 59108:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 59109:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 59110:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 59111:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 59112:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 59113:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 59114:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 59115:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 59116:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 59117:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 59118:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 59119:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 59120:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 59121:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 59122:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 59123:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 59124:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 59125:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 59126:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 59127:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 59128:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 59129:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 59130:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 59131:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 59132:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 59133:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 59134:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 59135:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 59136:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 59137:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 59138:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 59139:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 59140:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 59141:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 59142:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 59143:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 59144:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 59145:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 59146:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 59147:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 59148:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 59149:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 59150:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 59151:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 59152:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 59153:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 59154:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 59155:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 59156:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 59157:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 59158:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 59159:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 59160:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 59161:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 59162:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 59163:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 59164:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 59165:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 59166:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 59167:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 59168:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 59169:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 59170:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 59171:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 59172:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 59173:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 59174:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 59175:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 59176:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 59177:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 59178:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 59179:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 59180:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 59181:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 59182:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 59183:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 59184:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 59185:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 59186:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 59187:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 59188:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 59189:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 59190:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 59191:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 59192:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 59193:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 59194:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 59195:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 59196:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 59197:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 59198:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 59199:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 59200:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 59201:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 59202:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 59203:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 59204:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 59205:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 59206:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 59207:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 59208:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 59209:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 59210:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 59211:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 59212:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 59213:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 59214:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 59215:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 59216:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 59217:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 59218:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 59219:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 59220:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 59221:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 59222:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 59223:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 59224:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 59225:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 59226:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 59227:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 59228:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 59229:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 59230:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 59231:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 59232:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 59233:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 59234:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 59235:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 59236:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 59237:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 59238:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 59239:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 59240:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 59241:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 59242:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 59243:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 59244:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 59245:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 59246:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 59247:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 59248:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 59249:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 59250:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 59251:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 59252:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 59253:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 59254:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 59255:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 59256:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 59257:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 59258:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 59259:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 59260:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 59261:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 59262:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 59263:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 59264:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 59265:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 59266:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 59267:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 59268:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 59269:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 59270:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 59271:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 59272:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 59273:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 59274:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 59275:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 59276:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 59277:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 59278:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 59279:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 59280:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 59281:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 59282:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 59283:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 59284:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 59285:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 59286:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 59287:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 59288:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 59289:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 59290:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 59291:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 59292:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 59293:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 59294:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 59295:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 59296:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 59297:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 59298:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 59299:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 59300:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 59301:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 59302:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 59303:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 59304:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 59305:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 59306:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 59307:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 59308:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 59309:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 59310:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 59311:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 59312:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 59313:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 59314:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 59315:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 59316:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 59317:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 59318:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 59319:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 59320:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 59321:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 59322:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 59323:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 59324:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 59325:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 59326:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 59327:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 59328:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 59329:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 59330:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 59331:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 59332:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 59333:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 59334:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 59335:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 59336:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 59337:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 59338:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 59339:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 59340:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 59341:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 59342:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 59343:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 59344:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 59345:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 59346:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 59347:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 59348:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 59349:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 59350:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 59351:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 59352:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 59353:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 59354:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 59355:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 59356:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 59357:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 59358:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 59359:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 59360:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 59361:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 59362:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 59363:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 59364:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 59365:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 59366:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 59367:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 59368:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 59369:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 59370:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 59371:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 59372:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 59373:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 59374:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 59375:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 59376:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 59377:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 59378:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 59379:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 59380:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 59381:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 59382:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 59383:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 59384:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 59385:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 59386:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 59387:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 59388:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 59389:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 59390:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 59391:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 59392:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 59393:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 59394:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 59395:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 59396:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 59397:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 59398:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 59399:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 59400:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 59401:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 59402:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 59403:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 59404:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 59405:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 59406:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 59407:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 59408:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 59409:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 59410:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 59411:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 59412:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 59413:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 59414:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 59415:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 59416:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 59417:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 59418:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 59419:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 59420:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 59421:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 59422:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 59423:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 59424:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 59425:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 59426:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 59427:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 59428:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 59429:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 59430:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 59431:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 59432:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 59433:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 59434:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 59435:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 59436:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 59437:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 59438:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 59439:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 59440:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 59441:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 59442:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 59443:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 59444:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 59445:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 59446:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 59447:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 59448:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 59449:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 59450:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 59451:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 59452:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 59453:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 59454:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 59455:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 59456:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 59457:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 59458:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 59459:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 59460:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 59461:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 59462:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 59463:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 59464:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 59465:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 59466:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 59467:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 59468:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 59469:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 59470:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 59471:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 59472:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 59473:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 59474:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 59475:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 59476:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 59477:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 59478:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 59479:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 59480:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 59481:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 59482:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 59483:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 59484:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 59485:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 59486:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 59487:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 59488:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 59489:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 59490:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 59491:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 59492:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 59493:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 59494:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 59495:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 59496:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 59497:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 59498:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 59499:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 59500:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 59501:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 59502:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 59503:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 59504:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 59505:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 59506:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 59507:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 59508:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 59509:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 59510:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 59511:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 59512:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 59513:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 59514:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 59515:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 59516:22]
  assign io_z = ~x114; // @[Snxn100k.scala 59517:17]
endmodule
module SnxnLv4Inst181(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 58246:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 58247:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 58248:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 58249:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 58250:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 58251:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 58252:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 58253:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 58254:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 58255:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 58256:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 58257:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 58258:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 58259:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 58260:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 58261:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 58262:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 58263:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 58264:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 58265:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 58266:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 58267:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 58268:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 58269:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 58270:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 58271:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 58272:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 58273:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 58274:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 58275:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 58276:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 58277:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 58278:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 58279:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 58280:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 58281:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 58282:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 58283:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 58284:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 58285:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 58286:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 58287:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 58288:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 58289:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 58290:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 58291:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 58292:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 58293:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 58294:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 58295:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 58296:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 58297:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 58298:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 58299:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 58300:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 58301:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 58302:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 58303:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 58304:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 58305:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 58306:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 58307:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 58308:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 58309:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 58310:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 58311:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 58312:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 58313:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 58314:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 58315:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 58316:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 58317:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 58318:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 58319:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 58320:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 58321:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 58322:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 58323:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 58324:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 58325:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 58326:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 58327:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 58328:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 58329:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 58330:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 58331:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 58332:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 58333:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 58334:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 58335:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 58336:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 58337:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 58338:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 58339:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 58340:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 58341:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 58342:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 58343:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 58344:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 58345:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 58346:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 58347:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 58348:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 58349:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 58350:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 58351:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 58352:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 58353:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 58354:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 58355:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 58356:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 58357:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 58358:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 58359:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 58360:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 58361:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 58362:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 58363:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 58364:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 58365:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 58366:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 58367:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 58368:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 58369:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 58370:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 58371:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 58372:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 58373:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 58374:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 58375:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 58376:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 58377:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 58378:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 58379:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 58380:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 58381:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 58382:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 58383:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 58384:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 58385:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 58386:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 58387:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 58388:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 58389:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 58390:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 58391:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 58392:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 58393:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 58394:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 58395:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 58396:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 58397:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 58398:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 58399:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 58400:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 58401:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 58402:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 58403:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 58404:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 58405:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 58406:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 58407:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 58408:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 58409:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 58410:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 58411:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 58412:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 58413:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 58414:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 58415:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 58416:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 58417:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 58418:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 58419:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 58420:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 58421:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 58422:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 58423:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 58424:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 58425:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 58426:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 58427:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 58428:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 58429:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 58430:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 58431:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 58432:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 58433:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 58434:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 58435:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 58436:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 58437:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 58438:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 58439:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 58440:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 58441:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 58442:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 58443:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 58444:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 58445:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 58446:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 58447:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 58448:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 58449:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 58450:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 58451:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 58452:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 58453:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 58454:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 58455:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 58456:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 58457:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 58458:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 58459:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 58460:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 58461:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 58462:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 58463:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 58464:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 58465:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 58466:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 58467:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 58468:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 58469:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 58470:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 58471:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 58472:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 58473:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 58474:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 58475:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 58476:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 58477:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 58478:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 58479:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 58480:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 58481:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 58482:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 58483:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 58484:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 58485:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 58486:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 58487:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 58488:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 58489:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 58490:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 58491:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 58492:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 58493:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 58494:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 58495:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 58496:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 58497:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 58498:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 58499:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 58500:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 58501:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 58502:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 58503:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 58504:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 58505:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 58506:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 58507:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 58508:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 58509:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 58510:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 58511:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 58512:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 58513:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 58514:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 58515:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 58516:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 58517:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 58518:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 58519:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 58520:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 58521:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 58522:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 58523:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 58524:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 58525:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 58526:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 58527:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 58528:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 58529:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 58530:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 58531:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 58532:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 58533:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 58534:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 58535:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 58536:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 58537:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 58538:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 58539:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 58540:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 58541:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 58542:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 58543:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 58544:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 58545:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 58546:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 58547:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 58548:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 58549:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 58550:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 58551:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 58552:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 58553:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 58554:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 58555:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 58556:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 58557:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 58558:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 58559:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 58560:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 58561:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 58562:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 58563:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 58564:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 58565:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 58566:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 58567:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 58568:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 58569:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 58570:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 58571:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 58572:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 58573:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 58574:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 58575:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 58576:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 58577:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 58578:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 58579:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 58580:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 58581:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 58582:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 58583:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 58584:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 58585:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 58586:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 58587:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 58588:20]
  assign io_z = ~x85; // @[Snxn100k.scala 58589:16]
endmodule
module SnxnLv3Inst45(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst180_io_a; // @[Snxn100k.scala 15460:35]
  wire  inst_SnxnLv4Inst180_io_b; // @[Snxn100k.scala 15460:35]
  wire  inst_SnxnLv4Inst180_io_z; // @[Snxn100k.scala 15460:35]
  wire  inst_SnxnLv4Inst181_io_a; // @[Snxn100k.scala 15464:35]
  wire  inst_SnxnLv4Inst181_io_b; // @[Snxn100k.scala 15464:35]
  wire  inst_SnxnLv4Inst181_io_z; // @[Snxn100k.scala 15464:35]
  wire  inst_SnxnLv4Inst182_io_a; // @[Snxn100k.scala 15468:35]
  wire  inst_SnxnLv4Inst182_io_b; // @[Snxn100k.scala 15468:35]
  wire  inst_SnxnLv4Inst182_io_z; // @[Snxn100k.scala 15468:35]
  wire  inst_SnxnLv4Inst183_io_a; // @[Snxn100k.scala 15472:35]
  wire  inst_SnxnLv4Inst183_io_b; // @[Snxn100k.scala 15472:35]
  wire  inst_SnxnLv4Inst183_io_z; // @[Snxn100k.scala 15472:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst180_io_z + inst_SnxnLv4Inst181_io_z; // @[Snxn100k.scala 15476:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst182_io_z; // @[Snxn100k.scala 15476:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst183_io_z; // @[Snxn100k.scala 15476:92]
  SnxnLv4Inst180 inst_SnxnLv4Inst180 ( // @[Snxn100k.scala 15460:35]
    .io_a(inst_SnxnLv4Inst180_io_a),
    .io_b(inst_SnxnLv4Inst180_io_b),
    .io_z(inst_SnxnLv4Inst180_io_z)
  );
  SnxnLv4Inst181 inst_SnxnLv4Inst181 ( // @[Snxn100k.scala 15464:35]
    .io_a(inst_SnxnLv4Inst181_io_a),
    .io_b(inst_SnxnLv4Inst181_io_b),
    .io_z(inst_SnxnLv4Inst181_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst182 ( // @[Snxn100k.scala 15468:35]
    .io_a(inst_SnxnLv4Inst182_io_a),
    .io_b(inst_SnxnLv4Inst182_io_b),
    .io_z(inst_SnxnLv4Inst182_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst183 ( // @[Snxn100k.scala 15472:35]
    .io_a(inst_SnxnLv4Inst183_io_a),
    .io_b(inst_SnxnLv4Inst183_io_b),
    .io_z(inst_SnxnLv4Inst183_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 15477:15]
  assign inst_SnxnLv4Inst180_io_a = io_a; // @[Snxn100k.scala 15461:28]
  assign inst_SnxnLv4Inst180_io_b = io_b; // @[Snxn100k.scala 15462:28]
  assign inst_SnxnLv4Inst181_io_a = io_a; // @[Snxn100k.scala 15465:28]
  assign inst_SnxnLv4Inst181_io_b = io_b; // @[Snxn100k.scala 15466:28]
  assign inst_SnxnLv4Inst182_io_a = io_a; // @[Snxn100k.scala 15469:28]
  assign inst_SnxnLv4Inst182_io_b = io_b; // @[Snxn100k.scala 15470:28]
  assign inst_SnxnLv4Inst183_io_a = io_a; // @[Snxn100k.scala 15473:28]
  assign inst_SnxnLv4Inst183_io_b = io_b; // @[Snxn100k.scala 15474:28]
endmodule
module SnxnLv4Inst186(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 59984:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 59985:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 59986:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 59987:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 59988:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 59989:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 59990:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 59991:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 59992:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 59993:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 59994:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 59995:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 59996:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 59997:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 59998:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 59999:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 60000:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 60001:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 60002:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 60003:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 60004:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 60005:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 60006:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 60007:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 60008:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 60009:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 60010:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 60011:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 60012:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 60013:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 60014:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 60015:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 60016:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 60017:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 60018:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 60019:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 60020:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 60021:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 60022:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 60023:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 60024:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 60025:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 60026:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 60027:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 60028:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 60029:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 60030:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 60031:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 60032:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 60033:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 60034:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 60035:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 60036:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 60037:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 60038:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 60039:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 60040:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 60041:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 60042:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 60043:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 60044:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 60045:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 60046:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 60047:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 60048:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 60049:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 60050:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 60051:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 60052:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 60053:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 60054:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 60055:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 60056:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 60057:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 60058:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 60059:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 60060:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 60061:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 60062:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 60063:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 60064:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 60065:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 60066:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 60067:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 60068:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 60069:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 60070:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 60071:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 60072:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 60073:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 60074:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 60075:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 60076:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 60077:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 60078:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 60079:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 60080:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 60081:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 60082:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 60083:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 60084:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 60085:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 60086:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 60087:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 60088:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 60089:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 60090:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 60091:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 60092:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 60093:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 60094:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 60095:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 60096:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 60097:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 60098:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 60099:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 60100:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 60101:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 60102:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 60103:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 60104:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 60105:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 60106:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 60107:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 60108:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 60109:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 60110:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 60111:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 60112:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 60113:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 60114:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 60115:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 60116:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 60117:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 60118:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 60119:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 60120:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 60121:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 60122:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 60123:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 60124:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 60125:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 60126:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 60127:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 60128:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 60129:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 60130:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 60131:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 60132:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 60133:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 60134:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 60135:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 60136:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 60137:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 60138:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 60139:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 60140:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 60141:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 60142:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 60143:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 60144:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 60145:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 60146:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 60147:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 60148:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 60149:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 60150:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 60151:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 60152:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 60153:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 60154:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 60155:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 60156:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 60157:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 60158:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 60159:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 60160:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 60161:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 60162:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 60163:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 60164:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 60165:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 60166:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 60167:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 60168:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 60169:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 60170:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 60171:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 60172:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 60173:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 60174:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 60175:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 60176:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 60177:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 60178:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 60179:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 60180:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 60181:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 60182:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 60183:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 60184:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 60185:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 60186:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 60187:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 60188:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 60189:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 60190:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 60191:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 60192:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 60193:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 60194:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 60195:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 60196:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 60197:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 60198:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 60199:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 60200:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 60201:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 60202:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 60203:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 60204:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 60205:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 60206:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 60207:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 60208:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 60209:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 60210:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 60211:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 60212:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 60213:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 60214:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 60215:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 60216:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 60217:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 60218:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 60219:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 60220:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 60221:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 60222:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 60223:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 60224:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 60225:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 60226:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 60227:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 60228:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 60229:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 60230:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 60231:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 60232:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 60233:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 60234:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 60235:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 60236:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 60237:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 60238:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 60239:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 60240:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 60241:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 60242:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 60243:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 60244:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 60245:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 60246:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 60247:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 60248:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 60249:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 60250:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 60251:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 60252:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 60253:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 60254:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 60255:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 60256:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 60257:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 60258:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 60259:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 60260:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 60261:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 60262:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 60263:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 60264:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 60265:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 60266:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 60267:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 60268:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 60269:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 60270:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 60271:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 60272:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 60273:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 60274:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 60275:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 60276:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 60277:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 60278:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 60279:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 60280:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 60281:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 60282:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 60283:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 60284:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 60285:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 60286:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 60287:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 60288:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 60289:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 60290:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 60291:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 60292:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 60293:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 60294:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 60295:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 60296:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 60297:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 60298:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 60299:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 60300:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 60301:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 60302:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 60303:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 60304:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 60305:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 60306:20]
  assign io_z = ~x80; // @[Snxn100k.scala 60307:16]
endmodule
module SnxnLv3Inst46(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst184_io_a; // @[Snxn100k.scala 15751:35]
  wire  inst_SnxnLv4Inst184_io_b; // @[Snxn100k.scala 15751:35]
  wire  inst_SnxnLv4Inst184_io_z; // @[Snxn100k.scala 15751:35]
  wire  inst_SnxnLv4Inst185_io_a; // @[Snxn100k.scala 15755:35]
  wire  inst_SnxnLv4Inst185_io_b; // @[Snxn100k.scala 15755:35]
  wire  inst_SnxnLv4Inst185_io_z; // @[Snxn100k.scala 15755:35]
  wire  inst_SnxnLv4Inst186_io_a; // @[Snxn100k.scala 15759:35]
  wire  inst_SnxnLv4Inst186_io_b; // @[Snxn100k.scala 15759:35]
  wire  inst_SnxnLv4Inst186_io_z; // @[Snxn100k.scala 15759:35]
  wire  inst_SnxnLv4Inst187_io_a; // @[Snxn100k.scala 15763:35]
  wire  inst_SnxnLv4Inst187_io_b; // @[Snxn100k.scala 15763:35]
  wire  inst_SnxnLv4Inst187_io_z; // @[Snxn100k.scala 15763:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst184_io_z + inst_SnxnLv4Inst185_io_z; // @[Snxn100k.scala 15767:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst186_io_z; // @[Snxn100k.scala 15767:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst187_io_z; // @[Snxn100k.scala 15767:92]
  SnxnLv4Inst168 inst_SnxnLv4Inst184 ( // @[Snxn100k.scala 15751:35]
    .io_a(inst_SnxnLv4Inst184_io_a),
    .io_b(inst_SnxnLv4Inst184_io_b),
    .io_z(inst_SnxnLv4Inst184_io_z)
  );
  SnxnLv4Inst75 inst_SnxnLv4Inst185 ( // @[Snxn100k.scala 15755:35]
    .io_a(inst_SnxnLv4Inst185_io_a),
    .io_b(inst_SnxnLv4Inst185_io_b),
    .io_z(inst_SnxnLv4Inst185_io_z)
  );
  SnxnLv4Inst186 inst_SnxnLv4Inst186 ( // @[Snxn100k.scala 15759:35]
    .io_a(inst_SnxnLv4Inst186_io_a),
    .io_b(inst_SnxnLv4Inst186_io_b),
    .io_z(inst_SnxnLv4Inst186_io_z)
  );
  SnxnLv4Inst107 inst_SnxnLv4Inst187 ( // @[Snxn100k.scala 15763:35]
    .io_a(inst_SnxnLv4Inst187_io_a),
    .io_b(inst_SnxnLv4Inst187_io_b),
    .io_z(inst_SnxnLv4Inst187_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 15768:15]
  assign inst_SnxnLv4Inst184_io_a = io_a; // @[Snxn100k.scala 15752:28]
  assign inst_SnxnLv4Inst184_io_b = io_b; // @[Snxn100k.scala 15753:28]
  assign inst_SnxnLv4Inst185_io_a = io_a; // @[Snxn100k.scala 15756:28]
  assign inst_SnxnLv4Inst185_io_b = io_b; // @[Snxn100k.scala 15757:28]
  assign inst_SnxnLv4Inst186_io_a = io_a; // @[Snxn100k.scala 15760:28]
  assign inst_SnxnLv4Inst186_io_b = io_b; // @[Snxn100k.scala 15761:28]
  assign inst_SnxnLv4Inst187_io_a = io_a; // @[Snxn100k.scala 15764:28]
  assign inst_SnxnLv4Inst187_io_b = io_b; // @[Snxn100k.scala 15765:28]
endmodule
module SnxnLv3Inst47(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst188_io_a; // @[Snxn100k.scala 16166:35]
  wire  inst_SnxnLv4Inst188_io_b; // @[Snxn100k.scala 16166:35]
  wire  inst_SnxnLv4Inst188_io_z; // @[Snxn100k.scala 16166:35]
  wire  inst_SnxnLv4Inst189_io_a; // @[Snxn100k.scala 16170:35]
  wire  inst_SnxnLv4Inst189_io_b; // @[Snxn100k.scala 16170:35]
  wire  inst_SnxnLv4Inst189_io_z; // @[Snxn100k.scala 16170:35]
  wire  inst_SnxnLv4Inst190_io_a; // @[Snxn100k.scala 16174:35]
  wire  inst_SnxnLv4Inst190_io_b; // @[Snxn100k.scala 16174:35]
  wire  inst_SnxnLv4Inst190_io_z; // @[Snxn100k.scala 16174:35]
  wire  inst_SnxnLv4Inst191_io_a; // @[Snxn100k.scala 16178:35]
  wire  inst_SnxnLv4Inst191_io_b; // @[Snxn100k.scala 16178:35]
  wire  inst_SnxnLv4Inst191_io_z; // @[Snxn100k.scala 16178:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst188_io_z + inst_SnxnLv4Inst189_io_z; // @[Snxn100k.scala 16182:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst190_io_z; // @[Snxn100k.scala 16182:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst191_io_z; // @[Snxn100k.scala 16182:92]
  SnxnLv4Inst20 inst_SnxnLv4Inst188 ( // @[Snxn100k.scala 16166:35]
    .io_a(inst_SnxnLv4Inst188_io_a),
    .io_b(inst_SnxnLv4Inst188_io_b),
    .io_z(inst_SnxnLv4Inst188_io_z)
  );
  SnxnLv4Inst110 inst_SnxnLv4Inst189 ( // @[Snxn100k.scala 16170:35]
    .io_a(inst_SnxnLv4Inst189_io_a),
    .io_b(inst_SnxnLv4Inst189_io_b),
    .io_z(inst_SnxnLv4Inst189_io_z)
  );
  SnxnLv4Inst161 inst_SnxnLv4Inst190 ( // @[Snxn100k.scala 16174:35]
    .io_a(inst_SnxnLv4Inst190_io_a),
    .io_b(inst_SnxnLv4Inst190_io_b),
    .io_z(inst_SnxnLv4Inst190_io_z)
  );
  SnxnLv4Inst186 inst_SnxnLv4Inst191 ( // @[Snxn100k.scala 16178:35]
    .io_a(inst_SnxnLv4Inst191_io_a),
    .io_b(inst_SnxnLv4Inst191_io_b),
    .io_z(inst_SnxnLv4Inst191_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 16183:15]
  assign inst_SnxnLv4Inst188_io_a = io_a; // @[Snxn100k.scala 16167:28]
  assign inst_SnxnLv4Inst188_io_b = io_b; // @[Snxn100k.scala 16168:28]
  assign inst_SnxnLv4Inst189_io_a = io_a; // @[Snxn100k.scala 16171:28]
  assign inst_SnxnLv4Inst189_io_b = io_b; // @[Snxn100k.scala 16172:28]
  assign inst_SnxnLv4Inst190_io_a = io_a; // @[Snxn100k.scala 16175:28]
  assign inst_SnxnLv4Inst190_io_b = io_b; // @[Snxn100k.scala 16176:28]
  assign inst_SnxnLv4Inst191_io_a = io_a; // @[Snxn100k.scala 16179:28]
  assign inst_SnxnLv4Inst191_io_b = io_b; // @[Snxn100k.scala 16180:28]
endmodule
module SnxnLv2Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst44_io_a; // @[Snxn100k.scala 3550:34]
  wire  inst_SnxnLv3Inst44_io_b; // @[Snxn100k.scala 3550:34]
  wire  inst_SnxnLv3Inst44_io_z; // @[Snxn100k.scala 3550:34]
  wire  inst_SnxnLv3Inst45_io_a; // @[Snxn100k.scala 3554:34]
  wire  inst_SnxnLv3Inst45_io_b; // @[Snxn100k.scala 3554:34]
  wire  inst_SnxnLv3Inst45_io_z; // @[Snxn100k.scala 3554:34]
  wire  inst_SnxnLv3Inst46_io_a; // @[Snxn100k.scala 3558:34]
  wire  inst_SnxnLv3Inst46_io_b; // @[Snxn100k.scala 3558:34]
  wire  inst_SnxnLv3Inst46_io_z; // @[Snxn100k.scala 3558:34]
  wire  inst_SnxnLv3Inst47_io_a; // @[Snxn100k.scala 3562:34]
  wire  inst_SnxnLv3Inst47_io_b; // @[Snxn100k.scala 3562:34]
  wire  inst_SnxnLv3Inst47_io_z; // @[Snxn100k.scala 3562:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst44_io_z + inst_SnxnLv3Inst45_io_z; // @[Snxn100k.scala 3566:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst46_io_z; // @[Snxn100k.scala 3566:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst47_io_z; // @[Snxn100k.scala 3566:89]
  SnxnLv3Inst44 inst_SnxnLv3Inst44 ( // @[Snxn100k.scala 3550:34]
    .io_a(inst_SnxnLv3Inst44_io_a),
    .io_b(inst_SnxnLv3Inst44_io_b),
    .io_z(inst_SnxnLv3Inst44_io_z)
  );
  SnxnLv3Inst45 inst_SnxnLv3Inst45 ( // @[Snxn100k.scala 3554:34]
    .io_a(inst_SnxnLv3Inst45_io_a),
    .io_b(inst_SnxnLv3Inst45_io_b),
    .io_z(inst_SnxnLv3Inst45_io_z)
  );
  SnxnLv3Inst46 inst_SnxnLv3Inst46 ( // @[Snxn100k.scala 3558:34]
    .io_a(inst_SnxnLv3Inst46_io_a),
    .io_b(inst_SnxnLv3Inst46_io_b),
    .io_z(inst_SnxnLv3Inst46_io_z)
  );
  SnxnLv3Inst47 inst_SnxnLv3Inst47 ( // @[Snxn100k.scala 3562:34]
    .io_a(inst_SnxnLv3Inst47_io_a),
    .io_b(inst_SnxnLv3Inst47_io_b),
    .io_z(inst_SnxnLv3Inst47_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 3567:15]
  assign inst_SnxnLv3Inst44_io_a = io_a; // @[Snxn100k.scala 3551:27]
  assign inst_SnxnLv3Inst44_io_b = io_b; // @[Snxn100k.scala 3552:27]
  assign inst_SnxnLv3Inst45_io_a = io_a; // @[Snxn100k.scala 3555:27]
  assign inst_SnxnLv3Inst45_io_b = io_b; // @[Snxn100k.scala 3556:27]
  assign inst_SnxnLv3Inst46_io_a = io_a; // @[Snxn100k.scala 3559:27]
  assign inst_SnxnLv3Inst46_io_b = io_b; // @[Snxn100k.scala 3560:27]
  assign inst_SnxnLv3Inst47_io_a = io_a; // @[Snxn100k.scala 3563:27]
  assign inst_SnxnLv3Inst47_io_b = io_b; // @[Snxn100k.scala 3564:27]
endmodule
module SnxnLv1Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst8_io_a; // @[Snxn100k.scala 875:33]
  wire  inst_SnxnLv2Inst8_io_b; // @[Snxn100k.scala 875:33]
  wire  inst_SnxnLv2Inst8_io_z; // @[Snxn100k.scala 875:33]
  wire  inst_SnxnLv2Inst9_io_a; // @[Snxn100k.scala 879:33]
  wire  inst_SnxnLv2Inst9_io_b; // @[Snxn100k.scala 879:33]
  wire  inst_SnxnLv2Inst9_io_z; // @[Snxn100k.scala 879:33]
  wire  inst_SnxnLv2Inst10_io_a; // @[Snxn100k.scala 883:34]
  wire  inst_SnxnLv2Inst10_io_b; // @[Snxn100k.scala 883:34]
  wire  inst_SnxnLv2Inst10_io_z; // @[Snxn100k.scala 883:34]
  wire  inst_SnxnLv2Inst11_io_a; // @[Snxn100k.scala 887:34]
  wire  inst_SnxnLv2Inst11_io_b; // @[Snxn100k.scala 887:34]
  wire  inst_SnxnLv2Inst11_io_z; // @[Snxn100k.scala 887:34]
  wire  _sum_T_1 = inst_SnxnLv2Inst8_io_z + inst_SnxnLv2Inst9_io_z; // @[Snxn100k.scala 891:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst10_io_z; // @[Snxn100k.scala 891:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst11_io_z; // @[Snxn100k.scala 891:87]
  SnxnLv2Inst8 inst_SnxnLv2Inst8 ( // @[Snxn100k.scala 875:33]
    .io_a(inst_SnxnLv2Inst8_io_a),
    .io_b(inst_SnxnLv2Inst8_io_b),
    .io_z(inst_SnxnLv2Inst8_io_z)
  );
  SnxnLv2Inst9 inst_SnxnLv2Inst9 ( // @[Snxn100k.scala 879:33]
    .io_a(inst_SnxnLv2Inst9_io_a),
    .io_b(inst_SnxnLv2Inst9_io_b),
    .io_z(inst_SnxnLv2Inst9_io_z)
  );
  SnxnLv2Inst10 inst_SnxnLv2Inst10 ( // @[Snxn100k.scala 883:34]
    .io_a(inst_SnxnLv2Inst10_io_a),
    .io_b(inst_SnxnLv2Inst10_io_b),
    .io_z(inst_SnxnLv2Inst10_io_z)
  );
  SnxnLv2Inst11 inst_SnxnLv2Inst11 ( // @[Snxn100k.scala 887:34]
    .io_a(inst_SnxnLv2Inst11_io_a),
    .io_b(inst_SnxnLv2Inst11_io_b),
    .io_z(inst_SnxnLv2Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 892:15]
  assign inst_SnxnLv2Inst8_io_a = io_a; // @[Snxn100k.scala 876:26]
  assign inst_SnxnLv2Inst8_io_b = io_b; // @[Snxn100k.scala 877:26]
  assign inst_SnxnLv2Inst9_io_a = io_a; // @[Snxn100k.scala 880:26]
  assign inst_SnxnLv2Inst9_io_b = io_b; // @[Snxn100k.scala 881:26]
  assign inst_SnxnLv2Inst10_io_a = io_a; // @[Snxn100k.scala 884:27]
  assign inst_SnxnLv2Inst10_io_b = io_b; // @[Snxn100k.scala 885:27]
  assign inst_SnxnLv2Inst11_io_a = io_a; // @[Snxn100k.scala 888:27]
  assign inst_SnxnLv2Inst11_io_b = io_b; // @[Snxn100k.scala 889:27]
endmodule
module SnxnLv3Inst48(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst192_io_a; // @[Snxn100k.scala 23267:35]
  wire  inst_SnxnLv4Inst192_io_b; // @[Snxn100k.scala 23267:35]
  wire  inst_SnxnLv4Inst192_io_z; // @[Snxn100k.scala 23267:35]
  wire  inst_SnxnLv4Inst193_io_a; // @[Snxn100k.scala 23271:35]
  wire  inst_SnxnLv4Inst193_io_b; // @[Snxn100k.scala 23271:35]
  wire  inst_SnxnLv4Inst193_io_z; // @[Snxn100k.scala 23271:35]
  wire  inst_SnxnLv4Inst194_io_a; // @[Snxn100k.scala 23275:35]
  wire  inst_SnxnLv4Inst194_io_b; // @[Snxn100k.scala 23275:35]
  wire  inst_SnxnLv4Inst194_io_z; // @[Snxn100k.scala 23275:35]
  wire  inst_SnxnLv4Inst195_io_a; // @[Snxn100k.scala 23279:35]
  wire  inst_SnxnLv4Inst195_io_b; // @[Snxn100k.scala 23279:35]
  wire  inst_SnxnLv4Inst195_io_z; // @[Snxn100k.scala 23279:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst192_io_z + inst_SnxnLv4Inst193_io_z; // @[Snxn100k.scala 23283:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst194_io_z; // @[Snxn100k.scala 23283:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst195_io_z; // @[Snxn100k.scala 23283:92]
  SnxnLv4Inst50 inst_SnxnLv4Inst192 ( // @[Snxn100k.scala 23267:35]
    .io_a(inst_SnxnLv4Inst192_io_a),
    .io_b(inst_SnxnLv4Inst192_io_b),
    .io_z(inst_SnxnLv4Inst192_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst193 ( // @[Snxn100k.scala 23271:35]
    .io_a(inst_SnxnLv4Inst193_io_a),
    .io_b(inst_SnxnLv4Inst193_io_b),
    .io_z(inst_SnxnLv4Inst193_io_z)
  );
  SnxnLv4Inst129 inst_SnxnLv4Inst194 ( // @[Snxn100k.scala 23275:35]
    .io_a(inst_SnxnLv4Inst194_io_a),
    .io_b(inst_SnxnLv4Inst194_io_b),
    .io_z(inst_SnxnLv4Inst194_io_z)
  );
  SnxnLv4Inst135 inst_SnxnLv4Inst195 ( // @[Snxn100k.scala 23279:35]
    .io_a(inst_SnxnLv4Inst195_io_a),
    .io_b(inst_SnxnLv4Inst195_io_b),
    .io_z(inst_SnxnLv4Inst195_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23284:15]
  assign inst_SnxnLv4Inst192_io_a = io_a; // @[Snxn100k.scala 23268:28]
  assign inst_SnxnLv4Inst192_io_b = io_b; // @[Snxn100k.scala 23269:28]
  assign inst_SnxnLv4Inst193_io_a = io_a; // @[Snxn100k.scala 23272:28]
  assign inst_SnxnLv4Inst193_io_b = io_b; // @[Snxn100k.scala 23273:28]
  assign inst_SnxnLv4Inst194_io_a = io_a; // @[Snxn100k.scala 23276:28]
  assign inst_SnxnLv4Inst194_io_b = io_b; // @[Snxn100k.scala 23277:28]
  assign inst_SnxnLv4Inst195_io_a = io_a; // @[Snxn100k.scala 23280:28]
  assign inst_SnxnLv4Inst195_io_b = io_b; // @[Snxn100k.scala 23281:28]
endmodule
module SnxnLv3Inst49(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst196_io_a; // @[Snxn100k.scala 23649:35]
  wire  inst_SnxnLv4Inst196_io_b; // @[Snxn100k.scala 23649:35]
  wire  inst_SnxnLv4Inst196_io_z; // @[Snxn100k.scala 23649:35]
  wire  inst_SnxnLv4Inst197_io_a; // @[Snxn100k.scala 23653:35]
  wire  inst_SnxnLv4Inst197_io_b; // @[Snxn100k.scala 23653:35]
  wire  inst_SnxnLv4Inst197_io_z; // @[Snxn100k.scala 23653:35]
  wire  inst_SnxnLv4Inst198_io_a; // @[Snxn100k.scala 23657:35]
  wire  inst_SnxnLv4Inst198_io_b; // @[Snxn100k.scala 23657:35]
  wire  inst_SnxnLv4Inst198_io_z; // @[Snxn100k.scala 23657:35]
  wire  inst_SnxnLv4Inst199_io_a; // @[Snxn100k.scala 23661:35]
  wire  inst_SnxnLv4Inst199_io_b; // @[Snxn100k.scala 23661:35]
  wire  inst_SnxnLv4Inst199_io_z; // @[Snxn100k.scala 23661:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst196_io_z + inst_SnxnLv4Inst197_io_z; // @[Snxn100k.scala 23665:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst198_io_z; // @[Snxn100k.scala 23665:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst199_io_z; // @[Snxn100k.scala 23665:92]
  SnxnLv4Inst75 inst_SnxnLv4Inst196 ( // @[Snxn100k.scala 23649:35]
    .io_a(inst_SnxnLv4Inst196_io_a),
    .io_b(inst_SnxnLv4Inst196_io_b),
    .io_z(inst_SnxnLv4Inst196_io_z)
  );
  SnxnLv4Inst7 inst_SnxnLv4Inst197 ( // @[Snxn100k.scala 23653:35]
    .io_a(inst_SnxnLv4Inst197_io_a),
    .io_b(inst_SnxnLv4Inst197_io_b),
    .io_z(inst_SnxnLv4Inst197_io_z)
  );
  SnxnLv4Inst68 inst_SnxnLv4Inst198 ( // @[Snxn100k.scala 23657:35]
    .io_a(inst_SnxnLv4Inst198_io_a),
    .io_b(inst_SnxnLv4Inst198_io_b),
    .io_z(inst_SnxnLv4Inst198_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst199 ( // @[Snxn100k.scala 23661:35]
    .io_a(inst_SnxnLv4Inst199_io_a),
    .io_b(inst_SnxnLv4Inst199_io_b),
    .io_z(inst_SnxnLv4Inst199_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23666:15]
  assign inst_SnxnLv4Inst196_io_a = io_a; // @[Snxn100k.scala 23650:28]
  assign inst_SnxnLv4Inst196_io_b = io_b; // @[Snxn100k.scala 23651:28]
  assign inst_SnxnLv4Inst197_io_a = io_a; // @[Snxn100k.scala 23654:28]
  assign inst_SnxnLv4Inst197_io_b = io_b; // @[Snxn100k.scala 23655:28]
  assign inst_SnxnLv4Inst198_io_a = io_a; // @[Snxn100k.scala 23658:28]
  assign inst_SnxnLv4Inst198_io_b = io_b; // @[Snxn100k.scala 23659:28]
  assign inst_SnxnLv4Inst199_io_a = io_a; // @[Snxn100k.scala 23662:28]
  assign inst_SnxnLv4Inst199_io_b = io_b; // @[Snxn100k.scala 23663:28]
endmodule
module SnxnLv3Inst50(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst200_io_a; // @[Snxn100k.scala 23574:35]
  wire  inst_SnxnLv4Inst200_io_b; // @[Snxn100k.scala 23574:35]
  wire  inst_SnxnLv4Inst200_io_z; // @[Snxn100k.scala 23574:35]
  wire  inst_SnxnLv4Inst201_io_a; // @[Snxn100k.scala 23578:35]
  wire  inst_SnxnLv4Inst201_io_b; // @[Snxn100k.scala 23578:35]
  wire  inst_SnxnLv4Inst201_io_z; // @[Snxn100k.scala 23578:35]
  wire  inst_SnxnLv4Inst202_io_a; // @[Snxn100k.scala 23582:35]
  wire  inst_SnxnLv4Inst202_io_b; // @[Snxn100k.scala 23582:35]
  wire  inst_SnxnLv4Inst202_io_z; // @[Snxn100k.scala 23582:35]
  wire  inst_SnxnLv4Inst203_io_a; // @[Snxn100k.scala 23586:35]
  wire  inst_SnxnLv4Inst203_io_b; // @[Snxn100k.scala 23586:35]
  wire  inst_SnxnLv4Inst203_io_z; // @[Snxn100k.scala 23586:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst200_io_z + inst_SnxnLv4Inst201_io_z; // @[Snxn100k.scala 23590:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst202_io_z; // @[Snxn100k.scala 23590:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst203_io_z; // @[Snxn100k.scala 23590:92]
  SnxnLv4Inst40 inst_SnxnLv4Inst200 ( // @[Snxn100k.scala 23574:35]
    .io_a(inst_SnxnLv4Inst200_io_a),
    .io_b(inst_SnxnLv4Inst200_io_b),
    .io_z(inst_SnxnLv4Inst200_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst201 ( // @[Snxn100k.scala 23578:35]
    .io_a(inst_SnxnLv4Inst201_io_a),
    .io_b(inst_SnxnLv4Inst201_io_b),
    .io_z(inst_SnxnLv4Inst201_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst202 ( // @[Snxn100k.scala 23582:35]
    .io_a(inst_SnxnLv4Inst202_io_a),
    .io_b(inst_SnxnLv4Inst202_io_b),
    .io_z(inst_SnxnLv4Inst202_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst203 ( // @[Snxn100k.scala 23586:35]
    .io_a(inst_SnxnLv4Inst203_io_a),
    .io_b(inst_SnxnLv4Inst203_io_b),
    .io_z(inst_SnxnLv4Inst203_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23591:15]
  assign inst_SnxnLv4Inst200_io_a = io_a; // @[Snxn100k.scala 23575:28]
  assign inst_SnxnLv4Inst200_io_b = io_b; // @[Snxn100k.scala 23576:28]
  assign inst_SnxnLv4Inst201_io_a = io_a; // @[Snxn100k.scala 23579:28]
  assign inst_SnxnLv4Inst201_io_b = io_b; // @[Snxn100k.scala 23580:28]
  assign inst_SnxnLv4Inst202_io_a = io_a; // @[Snxn100k.scala 23583:28]
  assign inst_SnxnLv4Inst202_io_b = io_b; // @[Snxn100k.scala 23584:28]
  assign inst_SnxnLv4Inst203_io_a = io_a; // @[Snxn100k.scala 23587:28]
  assign inst_SnxnLv4Inst203_io_b = io_b; // @[Snxn100k.scala 23588:28]
endmodule
module SnxnLv4Inst205(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 90534:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 90535:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 90536:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 90537:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 90538:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 90539:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 90540:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 90541:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 90542:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 90543:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 90544:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 90545:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 90546:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 90547:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 90548:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 90549:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 90550:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 90551:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 90552:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 90553:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 90554:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 90555:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 90556:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 90557:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 90558:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 90559:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 90560:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 90561:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 90562:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 90563:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 90564:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 90565:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 90566:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 90567:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 90568:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 90569:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 90570:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 90571:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 90572:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 90573:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 90574:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 90575:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 90576:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 90577:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 90578:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 90579:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 90580:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 90581:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 90582:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 90583:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 90584:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 90585:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 90586:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 90587:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 90588:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 90589:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 90590:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 90591:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 90592:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 90593:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 90594:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 90595:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 90596:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 90597:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 90598:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 90599:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 90600:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 90601:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 90602:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 90603:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 90604:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 90605:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 90606:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 90607:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 90608:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 90609:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 90610:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 90611:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 90612:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 90613:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 90614:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 90615:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 90616:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 90617:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 90618:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 90619:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 90620:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 90621:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 90622:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 90623:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 90624:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 90625:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 90626:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 90627:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 90628:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 90629:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 90630:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 90631:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 90632:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 90633:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 90634:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 90635:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 90636:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 90637:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 90638:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 90639:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 90640:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 90641:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 90642:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 90643:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 90644:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 90645:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 90646:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 90647:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 90648:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 90649:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 90650:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 90651:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 90652:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 90653:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 90654:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 90655:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 90656:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 90657:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 90658:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 90659:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 90660:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 90661:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 90662:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 90663:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 90664:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 90665:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 90666:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 90667:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 90668:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 90669:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 90670:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 90671:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 90672:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 90673:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 90674:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 90675:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 90676:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 90677:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 90678:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 90679:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 90680:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 90681:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 90682:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 90683:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 90684:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 90685:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 90686:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 90687:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 90688:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 90689:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 90690:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 90691:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 90692:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 90693:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 90694:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 90695:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 90696:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 90697:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 90698:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 90699:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 90700:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 90701:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 90702:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 90703:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 90704:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 90705:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 90706:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 90707:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 90708:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 90709:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 90710:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 90711:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 90712:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 90713:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 90714:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 90715:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 90716:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 90717:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 90718:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 90719:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 90720:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 90721:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 90722:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 90723:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 90724:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 90725:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 90726:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 90727:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 90728:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 90729:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 90730:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 90731:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 90732:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 90733:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 90734:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 90735:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 90736:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 90737:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 90738:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 90739:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 90740:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 90741:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 90742:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 90743:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 90744:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 90745:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 90746:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 90747:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 90748:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 90749:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 90750:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 90751:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 90752:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 90753:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 90754:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 90755:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 90756:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 90757:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 90758:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 90759:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 90760:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 90761:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 90762:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 90763:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 90764:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 90765:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 90766:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 90767:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 90768:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 90769:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 90770:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 90771:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 90772:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 90773:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 90774:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 90775:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 90776:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 90777:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 90778:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 90779:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 90780:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 90781:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 90782:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 90783:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 90784:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 90785:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 90786:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 90787:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 90788:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 90789:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 90790:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 90791:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 90792:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 90793:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 90794:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 90795:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 90796:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 90797:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 90798:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 90799:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 90800:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 90801:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 90802:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 90803:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 90804:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 90805:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 90806:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 90807:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 90808:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 90809:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 90810:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 90811:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 90812:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 90813:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 90814:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 90815:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 90816:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 90817:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 90818:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 90819:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 90820:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 90821:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 90822:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 90823:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 90824:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 90825:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 90826:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 90827:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 90828:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 90829:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 90830:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 90831:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 90832:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 90833:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 90834:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 90835:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 90836:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 90837:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 90838:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 90839:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 90840:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 90841:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 90842:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 90843:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 90844:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 90845:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 90846:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 90847:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 90848:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 90849:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 90850:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 90851:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 90852:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 90853:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 90854:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 90855:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 90856:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 90857:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 90858:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 90859:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 90860:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 90861:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 90862:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 90863:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 90864:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 90865:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 90866:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 90867:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 90868:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 90869:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 90870:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 90871:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 90872:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 90873:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 90874:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 90875:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 90876:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 90877:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 90878:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 90879:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 90880:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 90881:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 90882:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 90883:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 90884:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 90885:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 90886:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 90887:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 90888:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 90889:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 90890:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 90891:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 90892:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 90893:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 90894:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 90895:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 90896:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 90897:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 90898:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 90899:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 90900:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 90901:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 90902:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 90903:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 90904:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 90905:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 90906:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 90907:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 90908:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 90909:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 90910:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 90911:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 90912:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 90913:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 90914:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 90915:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 90916:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 90917:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 90918:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 90919:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 90920:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 90921:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 90922:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 90923:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 90924:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 90925:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 90926:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 90927:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 90928:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 90929:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 90930:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 90931:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 90932:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 90933:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 90934:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 90935:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 90936:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 90937:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 90938:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 90939:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 90940:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 90941:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 90942:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 90943:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 90944:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 90945:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 90946:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 90947:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 90948:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 90949:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 90950:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 90951:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 90952:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 90953:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 90954:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 90955:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 90956:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 90957:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 90958:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 90959:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 90960:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 90961:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 90962:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 90963:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 90964:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 90965:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 90966:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 90967:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 90968:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 90969:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 90970:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 90971:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 90972:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 90973:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 90974:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 90975:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 90976:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 90977:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 90978:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 90979:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 90980:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 90981:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 90982:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 90983:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 90984:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 90985:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 90986:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 90987:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 90988:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 90989:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 90990:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 90991:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 90992:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 90993:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 90994:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 90995:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 90996:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 90997:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 90998:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 90999:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 91000:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 91001:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 91002:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 91003:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 91004:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 91005:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 91006:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 91007:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 91008:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 91009:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 91010:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 91011:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 91012:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 91013:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 91014:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 91015:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 91016:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 91017:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 91018:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 91019:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 91020:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 91021:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 91022:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 91023:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 91024:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 91025:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 91026:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 91027:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 91028:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 91029:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 91030:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 91031:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 91032:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 91033:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 91034:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 91035:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 91036:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 91037:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 91038:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 91039:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 91040:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 91041:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 91042:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 91043:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 91044:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 91045:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 91046:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 91047:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 91048:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 91049:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 91050:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 91051:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 91052:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 91053:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 91054:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 91055:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 91056:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 91057:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 91058:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 91059:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 91060:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 91061:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 91062:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 91063:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 91064:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 91065:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 91066:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 91067:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 91068:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 91069:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 91070:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 91071:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 91072:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 91073:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 91074:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 91075:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 91076:22]
  assign io_z = ~x135; // @[Snxn100k.scala 91077:17]
endmodule
module SnxnLv4Inst206(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 90144:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 90145:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 90146:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 90147:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 90148:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 90149:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 90150:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 90151:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 90152:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 90153:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 90154:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 90155:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 90156:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 90157:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 90158:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 90159:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 90160:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 90161:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 90162:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 90163:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 90164:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 90165:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 90166:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 90167:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 90168:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 90169:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 90170:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 90171:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 90172:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 90173:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 90174:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 90175:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 90176:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 90177:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 90178:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 90179:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 90180:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 90181:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 90182:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 90183:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 90184:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 90185:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 90186:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 90187:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 90188:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 90189:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 90190:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 90191:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 90192:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 90193:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 90194:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 90195:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 90196:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 90197:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 90198:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 90199:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 90200:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 90201:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 90202:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 90203:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 90204:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 90205:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 90206:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 90207:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 90208:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 90209:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 90210:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 90211:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 90212:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 90213:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 90214:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 90215:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 90216:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 90217:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 90218:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 90219:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 90220:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 90221:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 90222:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 90223:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 90224:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 90225:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 90226:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 90227:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 90228:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 90229:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 90230:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 90231:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 90232:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 90233:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 90234:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 90235:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 90236:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 90237:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 90238:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 90239:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 90240:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 90241:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 90242:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 90243:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 90244:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 90245:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 90246:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 90247:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 90248:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 90249:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 90250:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 90251:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 90252:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 90253:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 90254:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 90255:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 90256:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 90257:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 90258:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 90259:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 90260:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 90261:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 90262:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 90263:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 90264:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 90265:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 90266:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 90267:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 90268:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 90269:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 90270:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 90271:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 90272:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 90273:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 90274:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 90275:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 90276:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 90277:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 90278:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 90279:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 90280:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 90281:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 90282:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 90283:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 90284:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 90285:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 90286:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 90287:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 90288:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 90289:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 90290:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 90291:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 90292:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 90293:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 90294:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 90295:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 90296:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 90297:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 90298:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 90299:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 90300:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 90301:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 90302:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 90303:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 90304:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 90305:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 90306:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 90307:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 90308:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 90309:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 90310:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 90311:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 90312:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 90313:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 90314:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 90315:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 90316:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 90317:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 90318:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 90319:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 90320:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 90321:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 90322:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 90323:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 90324:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 90325:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 90326:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 90327:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 90328:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 90329:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 90330:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 90331:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 90332:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 90333:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 90334:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 90335:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 90336:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 90337:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 90338:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 90339:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 90340:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 90341:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 90342:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 90343:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 90344:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 90345:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 90346:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 90347:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 90348:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 90349:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 90350:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 90351:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 90352:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 90353:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 90354:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 90355:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 90356:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 90357:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 90358:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 90359:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 90360:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 90361:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 90362:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 90363:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 90364:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 90365:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 90366:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 90367:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 90368:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 90369:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 90370:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 90371:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 90372:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 90373:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 90374:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 90375:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 90376:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 90377:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 90378:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 90379:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 90380:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 90381:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 90382:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 90383:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 90384:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 90385:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 90386:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 90387:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 90388:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 90389:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 90390:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 90391:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 90392:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 90393:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 90394:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 90395:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 90396:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 90397:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 90398:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 90399:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 90400:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 90401:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 90402:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 90403:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 90404:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 90405:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 90406:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 90407:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 90408:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 90409:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 90410:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 90411:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 90412:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 90413:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 90414:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 90415:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 90416:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 90417:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 90418:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 90419:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 90420:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 90421:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 90422:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 90423:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 90424:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 90425:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 90426:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 90427:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 90428:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 90429:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 90430:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 90431:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 90432:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 90433:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 90434:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 90435:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 90436:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 90437:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 90438:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 90439:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 90440:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 90441:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 90442:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 90443:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 90444:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 90445:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 90446:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 90447:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 90448:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 90449:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 90450:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 90451:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 90452:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 90453:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 90454:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 90455:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 90456:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 90457:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 90458:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 90459:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 90460:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 90461:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 90462:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 90463:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 90464:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 90465:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 90466:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 90467:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 90468:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 90469:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 90470:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 90471:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 90472:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 90473:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 90474:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 90475:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 90476:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 90477:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 90478:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 90479:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 90480:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 90481:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 90482:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 90483:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 90484:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 90485:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 90486:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 90487:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 90488:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 90489:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 90490:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 90491:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 90492:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 90493:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 90494:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 90495:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 90496:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 90497:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 90498:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 90499:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 90500:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 90501:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 90502:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 90503:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 90504:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 90505:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 90506:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 90507:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 90508:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 90509:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 90510:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 90511:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 90512:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 90513:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 90514:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 90515:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 90516:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 90517:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 90518:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 90519:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 90520:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 90521:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 90522:20]
  assign io_z = ~x94; // @[Snxn100k.scala 90523:16]
endmodule
module SnxnLv4Inst207(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 89592:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 89593:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 89594:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 89595:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 89596:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 89597:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 89598:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 89599:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 89600:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 89601:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 89602:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 89603:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 89604:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 89605:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 89606:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 89607:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 89608:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 89609:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 89610:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 89611:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 89612:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 89613:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 89614:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 89615:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 89616:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 89617:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 89618:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 89619:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 89620:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 89621:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 89622:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 89623:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 89624:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 89625:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 89626:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 89627:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 89628:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 89629:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 89630:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 89631:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 89632:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 89633:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 89634:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 89635:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 89636:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 89637:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 89638:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 89639:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 89640:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 89641:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 89642:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 89643:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 89644:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 89645:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 89646:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 89647:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 89648:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 89649:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 89650:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 89651:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 89652:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 89653:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 89654:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 89655:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 89656:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 89657:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 89658:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 89659:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 89660:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 89661:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 89662:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 89663:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 89664:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 89665:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 89666:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 89667:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 89668:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 89669:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 89670:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 89671:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 89672:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 89673:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 89674:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 89675:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 89676:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 89677:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 89678:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 89679:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 89680:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 89681:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 89682:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 89683:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 89684:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 89685:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 89686:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 89687:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 89688:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 89689:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 89690:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 89691:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 89692:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 89693:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 89694:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 89695:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 89696:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 89697:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 89698:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 89699:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 89700:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 89701:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 89702:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 89703:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 89704:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 89705:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 89706:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 89707:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 89708:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 89709:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 89710:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 89711:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 89712:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 89713:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 89714:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 89715:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 89716:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 89717:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 89718:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 89719:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 89720:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 89721:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 89722:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 89723:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 89724:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 89725:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 89726:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 89727:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 89728:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 89729:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 89730:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 89731:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 89732:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 89733:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 89734:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 89735:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 89736:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 89737:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 89738:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 89739:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 89740:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 89741:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 89742:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 89743:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 89744:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 89745:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 89746:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 89747:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 89748:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 89749:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 89750:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 89751:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 89752:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 89753:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 89754:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 89755:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 89756:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 89757:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 89758:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 89759:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 89760:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 89761:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 89762:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 89763:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 89764:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 89765:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 89766:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 89767:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 89768:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 89769:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 89770:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 89771:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 89772:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 89773:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 89774:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 89775:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 89776:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 89777:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 89778:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 89779:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 89780:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 89781:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 89782:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 89783:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 89784:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 89785:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 89786:20]
  assign io_z = ~x48; // @[Snxn100k.scala 89787:16]
endmodule
module SnxnLv3Inst51(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst204_io_a; // @[Snxn100k.scala 23036:35]
  wire  inst_SnxnLv4Inst204_io_b; // @[Snxn100k.scala 23036:35]
  wire  inst_SnxnLv4Inst204_io_z; // @[Snxn100k.scala 23036:35]
  wire  inst_SnxnLv4Inst205_io_a; // @[Snxn100k.scala 23040:35]
  wire  inst_SnxnLv4Inst205_io_b; // @[Snxn100k.scala 23040:35]
  wire  inst_SnxnLv4Inst205_io_z; // @[Snxn100k.scala 23040:35]
  wire  inst_SnxnLv4Inst206_io_a; // @[Snxn100k.scala 23044:35]
  wire  inst_SnxnLv4Inst206_io_b; // @[Snxn100k.scala 23044:35]
  wire  inst_SnxnLv4Inst206_io_z; // @[Snxn100k.scala 23044:35]
  wire  inst_SnxnLv4Inst207_io_a; // @[Snxn100k.scala 23048:35]
  wire  inst_SnxnLv4Inst207_io_b; // @[Snxn100k.scala 23048:35]
  wire  inst_SnxnLv4Inst207_io_z; // @[Snxn100k.scala 23048:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst204_io_z + inst_SnxnLv4Inst205_io_z; // @[Snxn100k.scala 23052:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst206_io_z; // @[Snxn100k.scala 23052:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst207_io_z; // @[Snxn100k.scala 23052:92]
  SnxnLv4Inst7 inst_SnxnLv4Inst204 ( // @[Snxn100k.scala 23036:35]
    .io_a(inst_SnxnLv4Inst204_io_a),
    .io_b(inst_SnxnLv4Inst204_io_b),
    .io_z(inst_SnxnLv4Inst204_io_z)
  );
  SnxnLv4Inst205 inst_SnxnLv4Inst205 ( // @[Snxn100k.scala 23040:35]
    .io_a(inst_SnxnLv4Inst205_io_a),
    .io_b(inst_SnxnLv4Inst205_io_b),
    .io_z(inst_SnxnLv4Inst205_io_z)
  );
  SnxnLv4Inst206 inst_SnxnLv4Inst206 ( // @[Snxn100k.scala 23044:35]
    .io_a(inst_SnxnLv4Inst206_io_a),
    .io_b(inst_SnxnLv4Inst206_io_b),
    .io_z(inst_SnxnLv4Inst206_io_z)
  );
  SnxnLv4Inst207 inst_SnxnLv4Inst207 ( // @[Snxn100k.scala 23048:35]
    .io_a(inst_SnxnLv4Inst207_io_a),
    .io_b(inst_SnxnLv4Inst207_io_b),
    .io_z(inst_SnxnLv4Inst207_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23053:15]
  assign inst_SnxnLv4Inst204_io_a = io_a; // @[Snxn100k.scala 23037:28]
  assign inst_SnxnLv4Inst204_io_b = io_b; // @[Snxn100k.scala 23038:28]
  assign inst_SnxnLv4Inst205_io_a = io_a; // @[Snxn100k.scala 23041:28]
  assign inst_SnxnLv4Inst205_io_b = io_b; // @[Snxn100k.scala 23042:28]
  assign inst_SnxnLv4Inst206_io_a = io_a; // @[Snxn100k.scala 23045:28]
  assign inst_SnxnLv4Inst206_io_b = io_b; // @[Snxn100k.scala 23046:28]
  assign inst_SnxnLv4Inst207_io_a = io_a; // @[Snxn100k.scala 23049:28]
  assign inst_SnxnLv4Inst207_io_b = io_b; // @[Snxn100k.scala 23050:28]
endmodule
module SnxnLv2Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst48_io_a; // @[Snxn100k.scala 5644:34]
  wire  inst_SnxnLv3Inst48_io_b; // @[Snxn100k.scala 5644:34]
  wire  inst_SnxnLv3Inst48_io_z; // @[Snxn100k.scala 5644:34]
  wire  inst_SnxnLv3Inst49_io_a; // @[Snxn100k.scala 5648:34]
  wire  inst_SnxnLv3Inst49_io_b; // @[Snxn100k.scala 5648:34]
  wire  inst_SnxnLv3Inst49_io_z; // @[Snxn100k.scala 5648:34]
  wire  inst_SnxnLv3Inst50_io_a; // @[Snxn100k.scala 5652:34]
  wire  inst_SnxnLv3Inst50_io_b; // @[Snxn100k.scala 5652:34]
  wire  inst_SnxnLv3Inst50_io_z; // @[Snxn100k.scala 5652:34]
  wire  inst_SnxnLv3Inst51_io_a; // @[Snxn100k.scala 5656:34]
  wire  inst_SnxnLv3Inst51_io_b; // @[Snxn100k.scala 5656:34]
  wire  inst_SnxnLv3Inst51_io_z; // @[Snxn100k.scala 5656:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst48_io_z + inst_SnxnLv3Inst49_io_z; // @[Snxn100k.scala 5660:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst50_io_z; // @[Snxn100k.scala 5660:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst51_io_z; // @[Snxn100k.scala 5660:89]
  SnxnLv3Inst48 inst_SnxnLv3Inst48 ( // @[Snxn100k.scala 5644:34]
    .io_a(inst_SnxnLv3Inst48_io_a),
    .io_b(inst_SnxnLv3Inst48_io_b),
    .io_z(inst_SnxnLv3Inst48_io_z)
  );
  SnxnLv3Inst49 inst_SnxnLv3Inst49 ( // @[Snxn100k.scala 5648:34]
    .io_a(inst_SnxnLv3Inst49_io_a),
    .io_b(inst_SnxnLv3Inst49_io_b),
    .io_z(inst_SnxnLv3Inst49_io_z)
  );
  SnxnLv3Inst50 inst_SnxnLv3Inst50 ( // @[Snxn100k.scala 5652:34]
    .io_a(inst_SnxnLv3Inst50_io_a),
    .io_b(inst_SnxnLv3Inst50_io_b),
    .io_z(inst_SnxnLv3Inst50_io_z)
  );
  SnxnLv3Inst51 inst_SnxnLv3Inst51 ( // @[Snxn100k.scala 5656:34]
    .io_a(inst_SnxnLv3Inst51_io_a),
    .io_b(inst_SnxnLv3Inst51_io_b),
    .io_z(inst_SnxnLv3Inst51_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 5661:15]
  assign inst_SnxnLv3Inst48_io_a = io_a; // @[Snxn100k.scala 5645:27]
  assign inst_SnxnLv3Inst48_io_b = io_b; // @[Snxn100k.scala 5646:27]
  assign inst_SnxnLv3Inst49_io_a = io_a; // @[Snxn100k.scala 5649:27]
  assign inst_SnxnLv3Inst49_io_b = io_b; // @[Snxn100k.scala 5650:27]
  assign inst_SnxnLv3Inst50_io_a = io_a; // @[Snxn100k.scala 5653:27]
  assign inst_SnxnLv3Inst50_io_b = io_b; // @[Snxn100k.scala 5654:27]
  assign inst_SnxnLv3Inst51_io_a = io_a; // @[Snxn100k.scala 5657:27]
  assign inst_SnxnLv3Inst51_io_b = io_b; // @[Snxn100k.scala 5658:27]
endmodule
module SnxnLv3Inst52(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst208_io_a; // @[Snxn100k.scala 26524:35]
  wire  inst_SnxnLv4Inst208_io_b; // @[Snxn100k.scala 26524:35]
  wire  inst_SnxnLv4Inst208_io_z; // @[Snxn100k.scala 26524:35]
  wire  inst_SnxnLv4Inst209_io_a; // @[Snxn100k.scala 26528:35]
  wire  inst_SnxnLv4Inst209_io_b; // @[Snxn100k.scala 26528:35]
  wire  inst_SnxnLv4Inst209_io_z; // @[Snxn100k.scala 26528:35]
  wire  inst_SnxnLv4Inst210_io_a; // @[Snxn100k.scala 26532:35]
  wire  inst_SnxnLv4Inst210_io_b; // @[Snxn100k.scala 26532:35]
  wire  inst_SnxnLv4Inst210_io_z; // @[Snxn100k.scala 26532:35]
  wire  inst_SnxnLv4Inst211_io_a; // @[Snxn100k.scala 26536:35]
  wire  inst_SnxnLv4Inst211_io_b; // @[Snxn100k.scala 26536:35]
  wire  inst_SnxnLv4Inst211_io_z; // @[Snxn100k.scala 26536:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst208_io_z + inst_SnxnLv4Inst209_io_z; // @[Snxn100k.scala 26540:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst210_io_z; // @[Snxn100k.scala 26540:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst211_io_z; // @[Snxn100k.scala 26540:92]
  SnxnLv4Inst4 inst_SnxnLv4Inst208 ( // @[Snxn100k.scala 26524:35]
    .io_a(inst_SnxnLv4Inst208_io_a),
    .io_b(inst_SnxnLv4Inst208_io_b),
    .io_z(inst_SnxnLv4Inst208_io_z)
  );
  SnxnLv4Inst117 inst_SnxnLv4Inst209 ( // @[Snxn100k.scala 26528:35]
    .io_a(inst_SnxnLv4Inst209_io_a),
    .io_b(inst_SnxnLv4Inst209_io_b),
    .io_z(inst_SnxnLv4Inst209_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst210 ( // @[Snxn100k.scala 26532:35]
    .io_a(inst_SnxnLv4Inst210_io_a),
    .io_b(inst_SnxnLv4Inst210_io_b),
    .io_z(inst_SnxnLv4Inst210_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst211 ( // @[Snxn100k.scala 26536:35]
    .io_a(inst_SnxnLv4Inst211_io_a),
    .io_b(inst_SnxnLv4Inst211_io_b),
    .io_z(inst_SnxnLv4Inst211_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26541:15]
  assign inst_SnxnLv4Inst208_io_a = io_a; // @[Snxn100k.scala 26525:28]
  assign inst_SnxnLv4Inst208_io_b = io_b; // @[Snxn100k.scala 26526:28]
  assign inst_SnxnLv4Inst209_io_a = io_a; // @[Snxn100k.scala 26529:28]
  assign inst_SnxnLv4Inst209_io_b = io_b; // @[Snxn100k.scala 26530:28]
  assign inst_SnxnLv4Inst210_io_a = io_a; // @[Snxn100k.scala 26533:28]
  assign inst_SnxnLv4Inst210_io_b = io_b; // @[Snxn100k.scala 26534:28]
  assign inst_SnxnLv4Inst211_io_a = io_a; // @[Snxn100k.scala 26537:28]
  assign inst_SnxnLv4Inst211_io_b = io_b; // @[Snxn100k.scala 26538:28]
endmodule
module SnxnLv3Inst53(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst212_io_a; // @[Snxn100k.scala 26839:35]
  wire  inst_SnxnLv4Inst212_io_b; // @[Snxn100k.scala 26839:35]
  wire  inst_SnxnLv4Inst212_io_z; // @[Snxn100k.scala 26839:35]
  wire  inst_SnxnLv4Inst213_io_a; // @[Snxn100k.scala 26843:35]
  wire  inst_SnxnLv4Inst213_io_b; // @[Snxn100k.scala 26843:35]
  wire  inst_SnxnLv4Inst213_io_z; // @[Snxn100k.scala 26843:35]
  wire  inst_SnxnLv4Inst214_io_a; // @[Snxn100k.scala 26847:35]
  wire  inst_SnxnLv4Inst214_io_b; // @[Snxn100k.scala 26847:35]
  wire  inst_SnxnLv4Inst214_io_z; // @[Snxn100k.scala 26847:35]
  wire  inst_SnxnLv4Inst215_io_a; // @[Snxn100k.scala 26851:35]
  wire  inst_SnxnLv4Inst215_io_b; // @[Snxn100k.scala 26851:35]
  wire  inst_SnxnLv4Inst215_io_z; // @[Snxn100k.scala 26851:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst212_io_z + inst_SnxnLv4Inst213_io_z; // @[Snxn100k.scala 26855:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst214_io_z; // @[Snxn100k.scala 26855:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst215_io_z; // @[Snxn100k.scala 26855:92]
  SnxnLv4Inst103 inst_SnxnLv4Inst212 ( // @[Snxn100k.scala 26839:35]
    .io_a(inst_SnxnLv4Inst212_io_a),
    .io_b(inst_SnxnLv4Inst212_io_b),
    .io_z(inst_SnxnLv4Inst212_io_z)
  );
  SnxnLv4Inst0 inst_SnxnLv4Inst213 ( // @[Snxn100k.scala 26843:35]
    .io_a(inst_SnxnLv4Inst213_io_a),
    .io_b(inst_SnxnLv4Inst213_io_b),
    .io_z(inst_SnxnLv4Inst213_io_z)
  );
  SnxnLv4Inst205 inst_SnxnLv4Inst214 ( // @[Snxn100k.scala 26847:35]
    .io_a(inst_SnxnLv4Inst214_io_a),
    .io_b(inst_SnxnLv4Inst214_io_b),
    .io_z(inst_SnxnLv4Inst214_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst215 ( // @[Snxn100k.scala 26851:35]
    .io_a(inst_SnxnLv4Inst215_io_a),
    .io_b(inst_SnxnLv4Inst215_io_b),
    .io_z(inst_SnxnLv4Inst215_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26856:15]
  assign inst_SnxnLv4Inst212_io_a = io_a; // @[Snxn100k.scala 26840:28]
  assign inst_SnxnLv4Inst212_io_b = io_b; // @[Snxn100k.scala 26841:28]
  assign inst_SnxnLv4Inst213_io_a = io_a; // @[Snxn100k.scala 26844:28]
  assign inst_SnxnLv4Inst213_io_b = io_b; // @[Snxn100k.scala 26845:28]
  assign inst_SnxnLv4Inst214_io_a = io_a; // @[Snxn100k.scala 26848:28]
  assign inst_SnxnLv4Inst214_io_b = io_b; // @[Snxn100k.scala 26849:28]
  assign inst_SnxnLv4Inst215_io_a = io_a; // @[Snxn100k.scala 26852:28]
  assign inst_SnxnLv4Inst215_io_b = io_b; // @[Snxn100k.scala 26853:28]
endmodule
module SnxnLv4Inst217(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 100938:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 100939:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 100940:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 100941:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 100942:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 100943:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 100944:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 100945:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 100946:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 100947:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 100948:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 100949:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 100950:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 100951:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 100952:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 100953:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 100954:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 100955:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 100956:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 100957:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 100958:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 100959:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 100960:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 100961:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 100962:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 100963:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 100964:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 100965:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 100966:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 100967:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 100968:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 100969:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 100970:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 100971:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 100972:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 100973:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 100974:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 100975:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 100976:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 100977:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 100978:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 100979:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 100980:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 100981:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 100982:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 100983:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 100984:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 100985:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 100986:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 100987:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 100988:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 100989:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 100990:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 100991:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 100992:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 100993:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 100994:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 100995:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 100996:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 100997:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 100998:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 100999:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 101000:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 101001:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 101002:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 101003:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 101004:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 101005:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 101006:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 101007:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 101008:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 101009:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 101010:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 101011:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 101012:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 101013:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 101014:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 101015:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 101016:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 101017:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 101018:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 101019:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 101020:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 101021:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 101022:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 101023:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 101024:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 101025:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 101026:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 101027:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 101028:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 101029:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 101030:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 101031:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 101032:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 101033:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 101034:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 101035:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 101036:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 101037:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 101038:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 101039:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 101040:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 101041:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 101042:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 101043:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 101044:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 101045:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 101046:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 101047:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 101048:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 101049:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 101050:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 101051:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 101052:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 101053:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 101054:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 101055:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 101056:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 101057:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 101058:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 101059:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 101060:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 101061:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 101062:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 101063:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 101064:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 101065:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 101066:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 101067:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 101068:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 101069:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 101070:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 101071:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 101072:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 101073:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 101074:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 101075:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 101076:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 101077:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 101078:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 101079:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 101080:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 101081:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 101082:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 101083:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 101084:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 101085:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 101086:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 101087:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 101088:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 101089:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 101090:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 101091:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 101092:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 101093:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 101094:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 101095:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 101096:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 101097:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 101098:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 101099:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 101100:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 101101:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 101102:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 101103:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 101104:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 101105:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 101106:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 101107:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 101108:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 101109:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 101110:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 101111:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 101112:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 101113:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 101114:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 101115:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 101116:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 101117:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 101118:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 101119:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 101120:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 101121:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 101122:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 101123:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 101124:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 101125:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 101126:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 101127:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 101128:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 101129:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 101130:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 101131:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 101132:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 101133:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 101134:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 101135:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 101136:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 101137:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 101138:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 101139:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 101140:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 101141:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 101142:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 101143:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 101144:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 101145:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 101146:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 101147:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 101148:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 101149:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 101150:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 101151:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 101152:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 101153:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 101154:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 101155:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 101156:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 101157:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 101158:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 101159:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 101160:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 101161:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 101162:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 101163:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 101164:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 101165:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 101166:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 101167:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 101168:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 101169:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 101170:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 101171:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 101172:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 101173:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 101174:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 101175:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 101176:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 101177:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 101178:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 101179:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 101180:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 101181:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 101182:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 101183:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 101184:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 101185:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 101186:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 101187:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 101188:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 101189:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 101190:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 101191:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 101192:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 101193:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 101194:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 101195:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 101196:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 101197:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 101198:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 101199:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 101200:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 101201:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 101202:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 101203:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 101204:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 101205:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 101206:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 101207:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 101208:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 101209:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 101210:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 101211:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 101212:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 101213:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 101214:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 101215:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 101216:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 101217:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 101218:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 101219:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 101220:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 101221:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 101222:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 101223:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 101224:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 101225:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 101226:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 101227:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 101228:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 101229:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 101230:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 101231:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 101232:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 101233:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 101234:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 101235:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 101236:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 101237:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 101238:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 101239:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 101240:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 101241:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 101242:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 101243:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 101244:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 101245:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 101246:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 101247:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 101248:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 101249:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 101250:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 101251:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 101252:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 101253:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 101254:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 101255:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 101256:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 101257:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 101258:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 101259:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 101260:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 101261:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 101262:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 101263:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 101264:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 101265:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 101266:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 101267:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 101268:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 101269:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 101270:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 101271:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 101272:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 101273:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 101274:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 101275:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 101276:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 101277:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 101278:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 101279:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 101280:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 101281:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 101282:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 101283:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 101284:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 101285:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 101286:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 101287:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 101288:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 101289:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 101290:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 101291:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 101292:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 101293:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 101294:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 101295:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 101296:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 101297:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 101298:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 101299:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 101300:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 101301:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 101302:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 101303:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 101304:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 101305:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 101306:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 101307:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 101308:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 101309:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 101310:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 101311:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 101312:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 101313:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 101314:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 101315:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 101316:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 101317:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 101318:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 101319:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 101320:20]
  assign io_z = ~x95; // @[Snxn100k.scala 101321:16]
endmodule
module SnxnLv3Inst54(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst216_io_a; // @[Snxn100k.scala 26217:35]
  wire  inst_SnxnLv4Inst216_io_b; // @[Snxn100k.scala 26217:35]
  wire  inst_SnxnLv4Inst216_io_z; // @[Snxn100k.scala 26217:35]
  wire  inst_SnxnLv4Inst217_io_a; // @[Snxn100k.scala 26221:35]
  wire  inst_SnxnLv4Inst217_io_b; // @[Snxn100k.scala 26221:35]
  wire  inst_SnxnLv4Inst217_io_z; // @[Snxn100k.scala 26221:35]
  wire  inst_SnxnLv4Inst218_io_a; // @[Snxn100k.scala 26225:35]
  wire  inst_SnxnLv4Inst218_io_b; // @[Snxn100k.scala 26225:35]
  wire  inst_SnxnLv4Inst218_io_z; // @[Snxn100k.scala 26225:35]
  wire  inst_SnxnLv4Inst219_io_a; // @[Snxn100k.scala 26229:35]
  wire  inst_SnxnLv4Inst219_io_b; // @[Snxn100k.scala 26229:35]
  wire  inst_SnxnLv4Inst219_io_z; // @[Snxn100k.scala 26229:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst216_io_z + inst_SnxnLv4Inst217_io_z; // @[Snxn100k.scala 26233:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst218_io_z; // @[Snxn100k.scala 26233:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst219_io_z; // @[Snxn100k.scala 26233:92]
  SnxnLv4Inst68 inst_SnxnLv4Inst216 ( // @[Snxn100k.scala 26217:35]
    .io_a(inst_SnxnLv4Inst216_io_a),
    .io_b(inst_SnxnLv4Inst216_io_b),
    .io_z(inst_SnxnLv4Inst216_io_z)
  );
  SnxnLv4Inst217 inst_SnxnLv4Inst217 ( // @[Snxn100k.scala 26221:35]
    .io_a(inst_SnxnLv4Inst217_io_a),
    .io_b(inst_SnxnLv4Inst217_io_b),
    .io_z(inst_SnxnLv4Inst217_io_z)
  );
  SnxnLv4Inst39 inst_SnxnLv4Inst218 ( // @[Snxn100k.scala 26225:35]
    .io_a(inst_SnxnLv4Inst218_io_a),
    .io_b(inst_SnxnLv4Inst218_io_b),
    .io_z(inst_SnxnLv4Inst218_io_z)
  );
  SnxnLv4Inst117 inst_SnxnLv4Inst219 ( // @[Snxn100k.scala 26229:35]
    .io_a(inst_SnxnLv4Inst219_io_a),
    .io_b(inst_SnxnLv4Inst219_io_b),
    .io_z(inst_SnxnLv4Inst219_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26234:15]
  assign inst_SnxnLv4Inst216_io_a = io_a; // @[Snxn100k.scala 26218:28]
  assign inst_SnxnLv4Inst216_io_b = io_b; // @[Snxn100k.scala 26219:28]
  assign inst_SnxnLv4Inst217_io_a = io_a; // @[Snxn100k.scala 26222:28]
  assign inst_SnxnLv4Inst217_io_b = io_b; // @[Snxn100k.scala 26223:28]
  assign inst_SnxnLv4Inst218_io_a = io_a; // @[Snxn100k.scala 26226:28]
  assign inst_SnxnLv4Inst218_io_b = io_b; // @[Snxn100k.scala 26227:28]
  assign inst_SnxnLv4Inst219_io_a = io_a; // @[Snxn100k.scala 26230:28]
  assign inst_SnxnLv4Inst219_io_b = io_b; // @[Snxn100k.scala 26231:28]
endmodule
module SnxnLv4Inst221(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 104802:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 104803:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 104804:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 104805:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 104806:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 104807:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 104808:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 104809:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 104810:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 104811:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 104812:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 104813:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 104814:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 104815:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 104816:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 104817:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 104818:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 104819:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 104820:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 104821:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 104822:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 104823:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 104824:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 104825:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 104826:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 104827:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 104828:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 104829:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 104830:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 104831:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 104832:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 104833:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 104834:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 104835:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 104836:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 104837:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 104838:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 104839:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 104840:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 104841:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 104842:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 104843:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 104844:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 104845:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 104846:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 104847:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 104848:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 104849:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 104850:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 104851:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 104852:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 104853:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 104854:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 104855:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 104856:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 104857:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 104858:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 104859:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 104860:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 104861:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 104862:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 104863:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 104864:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 104865:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 104866:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 104867:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 104868:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 104869:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 104870:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 104871:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 104872:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 104873:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 104874:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 104875:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 104876:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 104877:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 104878:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 104879:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 104880:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 104881:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 104882:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 104883:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 104884:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 104885:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 104886:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 104887:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 104888:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 104889:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 104890:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 104891:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 104892:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 104893:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 104894:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 104895:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 104896:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 104897:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 104898:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 104899:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 104900:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 104901:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 104902:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 104903:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 104904:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 104905:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 104906:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 104907:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 104908:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 104909:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 104910:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 104911:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 104912:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 104913:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 104914:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 104915:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 104916:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 104917:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 104918:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 104919:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 104920:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 104921:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 104922:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 104923:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 104924:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 104925:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 104926:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 104927:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 104928:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 104929:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 104930:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 104931:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 104932:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 104933:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 104934:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 104935:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 104936:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 104937:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 104938:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 104939:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 104940:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 104941:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 104942:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 104943:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 104944:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 104945:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 104946:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 104947:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 104948:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 104949:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 104950:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 104951:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 104952:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 104953:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 104954:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 104955:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 104956:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 104957:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 104958:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 104959:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 104960:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 104961:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 104962:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 104963:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 104964:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 104965:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 104966:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 104967:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 104968:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 104969:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 104970:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 104971:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 104972:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 104973:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 104974:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 104975:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 104976:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 104977:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 104978:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 104979:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 104980:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 104981:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 104982:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 104983:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 104984:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 104985:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 104986:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 104987:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 104988:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 104989:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 104990:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 104991:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 104992:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 104993:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 104994:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 104995:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 104996:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 104997:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 104998:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 104999:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 105000:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 105001:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 105002:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 105003:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 105004:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 105005:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 105006:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 105007:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 105008:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 105009:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 105010:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 105011:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 105012:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 105013:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 105014:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 105015:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 105016:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 105017:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 105018:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 105019:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 105020:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 105021:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 105022:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 105023:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 105024:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 105025:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 105026:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 105027:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 105028:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 105029:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 105030:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 105031:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 105032:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 105033:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 105034:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 105035:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 105036:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 105037:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 105038:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 105039:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 105040:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 105041:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 105042:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 105043:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 105044:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 105045:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 105046:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 105047:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 105048:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 105049:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 105050:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 105051:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 105052:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 105053:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 105054:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 105055:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 105056:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 105057:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 105058:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 105059:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 105060:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 105061:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 105062:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 105063:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 105064:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 105065:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 105066:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 105067:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 105068:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 105069:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 105070:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 105071:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 105072:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 105073:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 105074:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 105075:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 105076:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 105077:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 105078:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 105079:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 105080:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 105081:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 105082:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 105083:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 105084:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 105085:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 105086:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 105087:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 105088:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 105089:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 105090:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 105091:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 105092:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 105093:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 105094:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 105095:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 105096:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 105097:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 105098:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 105099:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 105100:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 105101:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 105102:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 105103:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 105104:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 105105:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 105106:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 105107:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 105108:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 105109:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 105110:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 105111:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 105112:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 105113:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 105114:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 105115:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 105116:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 105117:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 105118:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 105119:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 105120:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 105121:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 105122:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 105123:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 105124:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 105125:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 105126:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 105127:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 105128:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 105129:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 105130:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 105131:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 105132:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 105133:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 105134:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 105135:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 105136:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 105137:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 105138:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 105139:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 105140:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 105141:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 105142:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 105143:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 105144:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 105145:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 105146:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 105147:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 105148:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 105149:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 105150:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 105151:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 105152:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 105153:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 105154:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 105155:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 105156:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 105157:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 105158:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 105159:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 105160:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 105161:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 105162:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 105163:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 105164:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 105165:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 105166:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 105167:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 105168:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 105169:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 105170:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 105171:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 105172:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 105173:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 105174:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 105175:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 105176:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 105177:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 105178:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 105179:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 105180:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 105181:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 105182:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 105183:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 105184:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 105185:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 105186:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 105187:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 105188:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 105189:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 105190:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 105191:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 105192:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 105193:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 105194:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 105195:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 105196:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 105197:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 105198:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 105199:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 105200:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 105201:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 105202:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 105203:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 105204:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 105205:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 105206:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 105207:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 105208:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 105209:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 105210:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 105211:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 105212:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 105213:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 105214:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 105215:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 105216:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 105217:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 105218:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 105219:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 105220:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 105221:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 105222:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 105223:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 105224:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 105225:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 105226:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 105227:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 105228:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 105229:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 105230:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 105231:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 105232:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 105233:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 105234:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 105235:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 105236:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 105237:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 105238:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 105239:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 105240:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 105241:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 105242:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 105243:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 105244:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 105245:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 105246:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 105247:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 105248:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 105249:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 105250:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 105251:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 105252:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 105253:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 105254:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 105255:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 105256:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 105257:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 105258:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 105259:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 105260:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 105261:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 105262:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 105263:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 105264:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 105265:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 105266:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 105267:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 105268:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 105269:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 105270:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 105271:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 105272:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 105273:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 105274:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 105275:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 105276:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 105277:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 105278:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 105279:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 105280:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 105281:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 105282:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 105283:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 105284:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 105285:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 105286:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 105287:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 105288:22]
  assign io_z = ~x121; // @[Snxn100k.scala 105289:17]
endmodule
module SnxnLv3Inst55(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst220_io_a; // @[Snxn100k.scala 27190:35]
  wire  inst_SnxnLv4Inst220_io_b; // @[Snxn100k.scala 27190:35]
  wire  inst_SnxnLv4Inst220_io_z; // @[Snxn100k.scala 27190:35]
  wire  inst_SnxnLv4Inst221_io_a; // @[Snxn100k.scala 27194:35]
  wire  inst_SnxnLv4Inst221_io_b; // @[Snxn100k.scala 27194:35]
  wire  inst_SnxnLv4Inst221_io_z; // @[Snxn100k.scala 27194:35]
  wire  inst_SnxnLv4Inst222_io_a; // @[Snxn100k.scala 27198:35]
  wire  inst_SnxnLv4Inst222_io_b; // @[Snxn100k.scala 27198:35]
  wire  inst_SnxnLv4Inst222_io_z; // @[Snxn100k.scala 27198:35]
  wire  inst_SnxnLv4Inst223_io_a; // @[Snxn100k.scala 27202:35]
  wire  inst_SnxnLv4Inst223_io_b; // @[Snxn100k.scala 27202:35]
  wire  inst_SnxnLv4Inst223_io_z; // @[Snxn100k.scala 27202:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst220_io_z + inst_SnxnLv4Inst221_io_z; // @[Snxn100k.scala 27206:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst222_io_z; // @[Snxn100k.scala 27206:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst223_io_z; // @[Snxn100k.scala 27206:92]
  SnxnLv4Inst148 inst_SnxnLv4Inst220 ( // @[Snxn100k.scala 27190:35]
    .io_a(inst_SnxnLv4Inst220_io_a),
    .io_b(inst_SnxnLv4Inst220_io_b),
    .io_z(inst_SnxnLv4Inst220_io_z)
  );
  SnxnLv4Inst221 inst_SnxnLv4Inst221 ( // @[Snxn100k.scala 27194:35]
    .io_a(inst_SnxnLv4Inst221_io_a),
    .io_b(inst_SnxnLv4Inst221_io_b),
    .io_z(inst_SnxnLv4Inst221_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst222 ( // @[Snxn100k.scala 27198:35]
    .io_a(inst_SnxnLv4Inst222_io_a),
    .io_b(inst_SnxnLv4Inst222_io_b),
    .io_z(inst_SnxnLv4Inst222_io_z)
  );
  SnxnLv4Inst68 inst_SnxnLv4Inst223 ( // @[Snxn100k.scala 27202:35]
    .io_a(inst_SnxnLv4Inst223_io_a),
    .io_b(inst_SnxnLv4Inst223_io_b),
    .io_z(inst_SnxnLv4Inst223_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27207:15]
  assign inst_SnxnLv4Inst220_io_a = io_a; // @[Snxn100k.scala 27191:28]
  assign inst_SnxnLv4Inst220_io_b = io_b; // @[Snxn100k.scala 27192:28]
  assign inst_SnxnLv4Inst221_io_a = io_a; // @[Snxn100k.scala 27195:28]
  assign inst_SnxnLv4Inst221_io_b = io_b; // @[Snxn100k.scala 27196:28]
  assign inst_SnxnLv4Inst222_io_a = io_a; // @[Snxn100k.scala 27199:28]
  assign inst_SnxnLv4Inst222_io_b = io_b; // @[Snxn100k.scala 27200:28]
  assign inst_SnxnLv4Inst223_io_a = io_a; // @[Snxn100k.scala 27203:28]
  assign inst_SnxnLv4Inst223_io_b = io_b; // @[Snxn100k.scala 27204:28]
endmodule
module SnxnLv2Inst13(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst52_io_a; // @[Snxn100k.scala 6741:34]
  wire  inst_SnxnLv3Inst52_io_b; // @[Snxn100k.scala 6741:34]
  wire  inst_SnxnLv3Inst52_io_z; // @[Snxn100k.scala 6741:34]
  wire  inst_SnxnLv3Inst53_io_a; // @[Snxn100k.scala 6745:34]
  wire  inst_SnxnLv3Inst53_io_b; // @[Snxn100k.scala 6745:34]
  wire  inst_SnxnLv3Inst53_io_z; // @[Snxn100k.scala 6745:34]
  wire  inst_SnxnLv3Inst54_io_a; // @[Snxn100k.scala 6749:34]
  wire  inst_SnxnLv3Inst54_io_b; // @[Snxn100k.scala 6749:34]
  wire  inst_SnxnLv3Inst54_io_z; // @[Snxn100k.scala 6749:34]
  wire  inst_SnxnLv3Inst55_io_a; // @[Snxn100k.scala 6753:34]
  wire  inst_SnxnLv3Inst55_io_b; // @[Snxn100k.scala 6753:34]
  wire  inst_SnxnLv3Inst55_io_z; // @[Snxn100k.scala 6753:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst52_io_z + inst_SnxnLv3Inst53_io_z; // @[Snxn100k.scala 6757:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst54_io_z; // @[Snxn100k.scala 6757:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst55_io_z; // @[Snxn100k.scala 6757:89]
  SnxnLv3Inst52 inst_SnxnLv3Inst52 ( // @[Snxn100k.scala 6741:34]
    .io_a(inst_SnxnLv3Inst52_io_a),
    .io_b(inst_SnxnLv3Inst52_io_b),
    .io_z(inst_SnxnLv3Inst52_io_z)
  );
  SnxnLv3Inst53 inst_SnxnLv3Inst53 ( // @[Snxn100k.scala 6745:34]
    .io_a(inst_SnxnLv3Inst53_io_a),
    .io_b(inst_SnxnLv3Inst53_io_b),
    .io_z(inst_SnxnLv3Inst53_io_z)
  );
  SnxnLv3Inst54 inst_SnxnLv3Inst54 ( // @[Snxn100k.scala 6749:34]
    .io_a(inst_SnxnLv3Inst54_io_a),
    .io_b(inst_SnxnLv3Inst54_io_b),
    .io_z(inst_SnxnLv3Inst54_io_z)
  );
  SnxnLv3Inst55 inst_SnxnLv3Inst55 ( // @[Snxn100k.scala 6753:34]
    .io_a(inst_SnxnLv3Inst55_io_a),
    .io_b(inst_SnxnLv3Inst55_io_b),
    .io_z(inst_SnxnLv3Inst55_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 6758:15]
  assign inst_SnxnLv3Inst52_io_a = io_a; // @[Snxn100k.scala 6742:27]
  assign inst_SnxnLv3Inst52_io_b = io_b; // @[Snxn100k.scala 6743:27]
  assign inst_SnxnLv3Inst53_io_a = io_a; // @[Snxn100k.scala 6746:27]
  assign inst_SnxnLv3Inst53_io_b = io_b; // @[Snxn100k.scala 6747:27]
  assign inst_SnxnLv3Inst54_io_a = io_a; // @[Snxn100k.scala 6750:27]
  assign inst_SnxnLv3Inst54_io_b = io_b; // @[Snxn100k.scala 6751:27]
  assign inst_SnxnLv3Inst55_io_a = io_a; // @[Snxn100k.scala 6754:27]
  assign inst_SnxnLv3Inst55_io_b = io_b; // @[Snxn100k.scala 6755:27]
endmodule
module SnxnLv3Inst56(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst224_io_a; // @[Snxn100k.scala 25986:35]
  wire  inst_SnxnLv4Inst224_io_b; // @[Snxn100k.scala 25986:35]
  wire  inst_SnxnLv4Inst224_io_z; // @[Snxn100k.scala 25986:35]
  wire  inst_SnxnLv4Inst225_io_a; // @[Snxn100k.scala 25990:35]
  wire  inst_SnxnLv4Inst225_io_b; // @[Snxn100k.scala 25990:35]
  wire  inst_SnxnLv4Inst225_io_z; // @[Snxn100k.scala 25990:35]
  wire  inst_SnxnLv4Inst226_io_a; // @[Snxn100k.scala 25994:35]
  wire  inst_SnxnLv4Inst226_io_b; // @[Snxn100k.scala 25994:35]
  wire  inst_SnxnLv4Inst226_io_z; // @[Snxn100k.scala 25994:35]
  wire  inst_SnxnLv4Inst227_io_a; // @[Snxn100k.scala 25998:35]
  wire  inst_SnxnLv4Inst227_io_b; // @[Snxn100k.scala 25998:35]
  wire  inst_SnxnLv4Inst227_io_z; // @[Snxn100k.scala 25998:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst224_io_z + inst_SnxnLv4Inst225_io_z; // @[Snxn100k.scala 26002:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst226_io_z; // @[Snxn100k.scala 26002:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst227_io_z; // @[Snxn100k.scala 26002:92]
  SnxnLv4Inst117 inst_SnxnLv4Inst224 ( // @[Snxn100k.scala 25986:35]
    .io_a(inst_SnxnLv4Inst224_io_a),
    .io_b(inst_SnxnLv4Inst224_io_b),
    .io_z(inst_SnxnLv4Inst224_io_z)
  );
  SnxnLv4Inst161 inst_SnxnLv4Inst225 ( // @[Snxn100k.scala 25990:35]
    .io_a(inst_SnxnLv4Inst225_io_a),
    .io_b(inst_SnxnLv4Inst225_io_b),
    .io_z(inst_SnxnLv4Inst225_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst226 ( // @[Snxn100k.scala 25994:35]
    .io_a(inst_SnxnLv4Inst226_io_a),
    .io_b(inst_SnxnLv4Inst226_io_b),
    .io_z(inst_SnxnLv4Inst226_io_z)
  );
  SnxnLv4Inst83 inst_SnxnLv4Inst227 ( // @[Snxn100k.scala 25998:35]
    .io_a(inst_SnxnLv4Inst227_io_a),
    .io_b(inst_SnxnLv4Inst227_io_b),
    .io_z(inst_SnxnLv4Inst227_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26003:15]
  assign inst_SnxnLv4Inst224_io_a = io_a; // @[Snxn100k.scala 25987:28]
  assign inst_SnxnLv4Inst224_io_b = io_b; // @[Snxn100k.scala 25988:28]
  assign inst_SnxnLv4Inst225_io_a = io_a; // @[Snxn100k.scala 25991:28]
  assign inst_SnxnLv4Inst225_io_b = io_b; // @[Snxn100k.scala 25992:28]
  assign inst_SnxnLv4Inst226_io_a = io_a; // @[Snxn100k.scala 25995:28]
  assign inst_SnxnLv4Inst226_io_b = io_b; // @[Snxn100k.scala 25996:28]
  assign inst_SnxnLv4Inst227_io_a = io_a; // @[Snxn100k.scala 25999:28]
  assign inst_SnxnLv4Inst227_io_b = io_b; // @[Snxn100k.scala 26000:28]
endmodule
module SnxnLv4Inst229(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 95492:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 95493:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 95494:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 95495:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 95496:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 95497:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 95498:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 95499:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 95500:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 95501:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 95502:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 95503:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 95504:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 95505:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 95506:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 95507:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 95508:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 95509:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 95510:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 95511:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 95512:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 95513:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 95514:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 95515:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 95516:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 95517:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 95518:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 95519:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 95520:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 95521:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 95522:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 95523:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 95524:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 95525:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 95526:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 95527:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 95528:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 95529:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 95530:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 95531:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 95532:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 95533:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 95534:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 95535:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 95536:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 95537:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 95538:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 95539:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 95540:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 95541:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 95542:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 95543:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 95544:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 95545:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 95546:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 95547:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 95548:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 95549:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 95550:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 95551:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 95552:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 95553:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 95554:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 95555:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 95556:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 95557:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 95558:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 95559:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 95560:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 95561:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 95562:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 95563:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 95564:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 95565:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 95566:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 95567:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 95568:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 95569:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 95570:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 95571:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 95572:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 95573:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 95574:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 95575:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 95576:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 95577:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 95578:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 95579:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 95580:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 95581:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 95582:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 95583:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 95584:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 95585:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 95586:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 95587:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 95588:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 95589:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 95590:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 95591:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 95592:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 95593:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 95594:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 95595:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 95596:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 95597:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 95598:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 95599:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 95600:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 95601:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 95602:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 95603:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 95604:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 95605:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 95606:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 95607:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 95608:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 95609:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 95610:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 95611:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 95612:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 95613:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 95614:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 95615:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 95616:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 95617:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 95618:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 95619:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 95620:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 95621:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 95622:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 95623:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 95624:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 95625:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 95626:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 95627:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 95628:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 95629:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 95630:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 95631:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 95632:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 95633:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 95634:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 95635:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 95636:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 95637:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 95638:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 95639:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 95640:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 95641:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 95642:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 95643:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 95644:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 95645:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 95646:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 95647:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 95648:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 95649:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 95650:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 95651:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 95652:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 95653:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 95654:20]
  assign io_z = ~x40; // @[Snxn100k.scala 95655:16]
endmodule
module SnxnLv3Inst57(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst228_io_a; // @[Snxn100k.scala 25065:35]
  wire  inst_SnxnLv4Inst228_io_b; // @[Snxn100k.scala 25065:35]
  wire  inst_SnxnLv4Inst228_io_z; // @[Snxn100k.scala 25065:35]
  wire  inst_SnxnLv4Inst229_io_a; // @[Snxn100k.scala 25069:35]
  wire  inst_SnxnLv4Inst229_io_b; // @[Snxn100k.scala 25069:35]
  wire  inst_SnxnLv4Inst229_io_z; // @[Snxn100k.scala 25069:35]
  wire  inst_SnxnLv4Inst230_io_a; // @[Snxn100k.scala 25073:35]
  wire  inst_SnxnLv4Inst230_io_b; // @[Snxn100k.scala 25073:35]
  wire  inst_SnxnLv4Inst230_io_z; // @[Snxn100k.scala 25073:35]
  wire  inst_SnxnLv4Inst231_io_a; // @[Snxn100k.scala 25077:35]
  wire  inst_SnxnLv4Inst231_io_b; // @[Snxn100k.scala 25077:35]
  wire  inst_SnxnLv4Inst231_io_z; // @[Snxn100k.scala 25077:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst228_io_z + inst_SnxnLv4Inst229_io_z; // @[Snxn100k.scala 25081:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst230_io_z; // @[Snxn100k.scala 25081:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst231_io_z; // @[Snxn100k.scala 25081:92]
  SnxnLv4Inst16 inst_SnxnLv4Inst228 ( // @[Snxn100k.scala 25065:35]
    .io_a(inst_SnxnLv4Inst228_io_a),
    .io_b(inst_SnxnLv4Inst228_io_b),
    .io_z(inst_SnxnLv4Inst228_io_z)
  );
  SnxnLv4Inst229 inst_SnxnLv4Inst229 ( // @[Snxn100k.scala 25069:35]
    .io_a(inst_SnxnLv4Inst229_io_a),
    .io_b(inst_SnxnLv4Inst229_io_b),
    .io_z(inst_SnxnLv4Inst229_io_z)
  );
  SnxnLv4Inst206 inst_SnxnLv4Inst230 ( // @[Snxn100k.scala 25073:35]
    .io_a(inst_SnxnLv4Inst230_io_a),
    .io_b(inst_SnxnLv4Inst230_io_b),
    .io_z(inst_SnxnLv4Inst230_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst231 ( // @[Snxn100k.scala 25077:35]
    .io_a(inst_SnxnLv4Inst231_io_a),
    .io_b(inst_SnxnLv4Inst231_io_b),
    .io_z(inst_SnxnLv4Inst231_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25082:15]
  assign inst_SnxnLv4Inst228_io_a = io_a; // @[Snxn100k.scala 25066:28]
  assign inst_SnxnLv4Inst228_io_b = io_b; // @[Snxn100k.scala 25067:28]
  assign inst_SnxnLv4Inst229_io_a = io_a; // @[Snxn100k.scala 25070:28]
  assign inst_SnxnLv4Inst229_io_b = io_b; // @[Snxn100k.scala 25071:28]
  assign inst_SnxnLv4Inst230_io_a = io_a; // @[Snxn100k.scala 25074:28]
  assign inst_SnxnLv4Inst230_io_b = io_b; // @[Snxn100k.scala 25075:28]
  assign inst_SnxnLv4Inst231_io_a = io_a; // @[Snxn100k.scala 25078:28]
  assign inst_SnxnLv4Inst231_io_b = io_b; // @[Snxn100k.scala 25079:28]
endmodule
module SnxnLv3Inst58(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst232_io_a; // @[Snxn100k.scala 25635:35]
  wire  inst_SnxnLv4Inst232_io_b; // @[Snxn100k.scala 25635:35]
  wire  inst_SnxnLv4Inst232_io_z; // @[Snxn100k.scala 25635:35]
  wire  inst_SnxnLv4Inst233_io_a; // @[Snxn100k.scala 25639:35]
  wire  inst_SnxnLv4Inst233_io_b; // @[Snxn100k.scala 25639:35]
  wire  inst_SnxnLv4Inst233_io_z; // @[Snxn100k.scala 25639:35]
  wire  inst_SnxnLv4Inst234_io_a; // @[Snxn100k.scala 25643:35]
  wire  inst_SnxnLv4Inst234_io_b; // @[Snxn100k.scala 25643:35]
  wire  inst_SnxnLv4Inst234_io_z; // @[Snxn100k.scala 25643:35]
  wire  inst_SnxnLv4Inst235_io_a; // @[Snxn100k.scala 25647:35]
  wire  inst_SnxnLv4Inst235_io_b; // @[Snxn100k.scala 25647:35]
  wire  inst_SnxnLv4Inst235_io_z; // @[Snxn100k.scala 25647:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst232_io_z + inst_SnxnLv4Inst233_io_z; // @[Snxn100k.scala 25651:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst234_io_z; // @[Snxn100k.scala 25651:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst235_io_z; // @[Snxn100k.scala 25651:92]
  SnxnLv4Inst20 inst_SnxnLv4Inst232 ( // @[Snxn100k.scala 25635:35]
    .io_a(inst_SnxnLv4Inst232_io_a),
    .io_b(inst_SnxnLv4Inst232_io_b),
    .io_z(inst_SnxnLv4Inst232_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst233 ( // @[Snxn100k.scala 25639:35]
    .io_a(inst_SnxnLv4Inst233_io_a),
    .io_b(inst_SnxnLv4Inst233_io_b),
    .io_z(inst_SnxnLv4Inst233_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst234 ( // @[Snxn100k.scala 25643:35]
    .io_a(inst_SnxnLv4Inst234_io_a),
    .io_b(inst_SnxnLv4Inst234_io_b),
    .io_z(inst_SnxnLv4Inst234_io_z)
  );
  SnxnLv4Inst115 inst_SnxnLv4Inst235 ( // @[Snxn100k.scala 25647:35]
    .io_a(inst_SnxnLv4Inst235_io_a),
    .io_b(inst_SnxnLv4Inst235_io_b),
    .io_z(inst_SnxnLv4Inst235_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25652:15]
  assign inst_SnxnLv4Inst232_io_a = io_a; // @[Snxn100k.scala 25636:28]
  assign inst_SnxnLv4Inst232_io_b = io_b; // @[Snxn100k.scala 25637:28]
  assign inst_SnxnLv4Inst233_io_a = io_a; // @[Snxn100k.scala 25640:28]
  assign inst_SnxnLv4Inst233_io_b = io_b; // @[Snxn100k.scala 25641:28]
  assign inst_SnxnLv4Inst234_io_a = io_a; // @[Snxn100k.scala 25644:28]
  assign inst_SnxnLv4Inst234_io_b = io_b; // @[Snxn100k.scala 25645:28]
  assign inst_SnxnLv4Inst235_io_a = io_a; // @[Snxn100k.scala 25648:28]
  assign inst_SnxnLv4Inst235_io_b = io_b; // @[Snxn100k.scala 25649:28]
endmodule
module SnxnLv3Inst59(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst236_io_a; // @[Snxn100k.scala 25336:35]
  wire  inst_SnxnLv4Inst236_io_b; // @[Snxn100k.scala 25336:35]
  wire  inst_SnxnLv4Inst236_io_z; // @[Snxn100k.scala 25336:35]
  wire  inst_SnxnLv4Inst237_io_a; // @[Snxn100k.scala 25340:35]
  wire  inst_SnxnLv4Inst237_io_b; // @[Snxn100k.scala 25340:35]
  wire  inst_SnxnLv4Inst237_io_z; // @[Snxn100k.scala 25340:35]
  wire  inst_SnxnLv4Inst238_io_a; // @[Snxn100k.scala 25344:35]
  wire  inst_SnxnLv4Inst238_io_b; // @[Snxn100k.scala 25344:35]
  wire  inst_SnxnLv4Inst238_io_z; // @[Snxn100k.scala 25344:35]
  wire  inst_SnxnLv4Inst239_io_a; // @[Snxn100k.scala 25348:35]
  wire  inst_SnxnLv4Inst239_io_b; // @[Snxn100k.scala 25348:35]
  wire  inst_SnxnLv4Inst239_io_z; // @[Snxn100k.scala 25348:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst236_io_z + inst_SnxnLv4Inst237_io_z; // @[Snxn100k.scala 25352:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst238_io_z; // @[Snxn100k.scala 25352:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst239_io_z; // @[Snxn100k.scala 25352:92]
  SnxnLv4Inst161 inst_SnxnLv4Inst236 ( // @[Snxn100k.scala 25336:35]
    .io_a(inst_SnxnLv4Inst236_io_a),
    .io_b(inst_SnxnLv4Inst236_io_b),
    .io_z(inst_SnxnLv4Inst236_io_z)
  );
  SnxnLv4Inst39 inst_SnxnLv4Inst237 ( // @[Snxn100k.scala 25340:35]
    .io_a(inst_SnxnLv4Inst237_io_a),
    .io_b(inst_SnxnLv4Inst237_io_b),
    .io_z(inst_SnxnLv4Inst237_io_z)
  );
  SnxnLv4Inst50 inst_SnxnLv4Inst238 ( // @[Snxn100k.scala 25344:35]
    .io_a(inst_SnxnLv4Inst238_io_a),
    .io_b(inst_SnxnLv4Inst238_io_b),
    .io_z(inst_SnxnLv4Inst238_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst239 ( // @[Snxn100k.scala 25348:35]
    .io_a(inst_SnxnLv4Inst239_io_a),
    .io_b(inst_SnxnLv4Inst239_io_b),
    .io_z(inst_SnxnLv4Inst239_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25353:15]
  assign inst_SnxnLv4Inst236_io_a = io_a; // @[Snxn100k.scala 25337:28]
  assign inst_SnxnLv4Inst236_io_b = io_b; // @[Snxn100k.scala 25338:28]
  assign inst_SnxnLv4Inst237_io_a = io_a; // @[Snxn100k.scala 25341:28]
  assign inst_SnxnLv4Inst237_io_b = io_b; // @[Snxn100k.scala 25342:28]
  assign inst_SnxnLv4Inst238_io_a = io_a; // @[Snxn100k.scala 25345:28]
  assign inst_SnxnLv4Inst238_io_b = io_b; // @[Snxn100k.scala 25346:28]
  assign inst_SnxnLv4Inst239_io_a = io_a; // @[Snxn100k.scala 25349:28]
  assign inst_SnxnLv4Inst239_io_b = io_b; // @[Snxn100k.scala 25350:28]
endmodule
module SnxnLv2Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst56_io_a; // @[Snxn100k.scala 6306:34]
  wire  inst_SnxnLv3Inst56_io_b; // @[Snxn100k.scala 6306:34]
  wire  inst_SnxnLv3Inst56_io_z; // @[Snxn100k.scala 6306:34]
  wire  inst_SnxnLv3Inst57_io_a; // @[Snxn100k.scala 6310:34]
  wire  inst_SnxnLv3Inst57_io_b; // @[Snxn100k.scala 6310:34]
  wire  inst_SnxnLv3Inst57_io_z; // @[Snxn100k.scala 6310:34]
  wire  inst_SnxnLv3Inst58_io_a; // @[Snxn100k.scala 6314:34]
  wire  inst_SnxnLv3Inst58_io_b; // @[Snxn100k.scala 6314:34]
  wire  inst_SnxnLv3Inst58_io_z; // @[Snxn100k.scala 6314:34]
  wire  inst_SnxnLv3Inst59_io_a; // @[Snxn100k.scala 6318:34]
  wire  inst_SnxnLv3Inst59_io_b; // @[Snxn100k.scala 6318:34]
  wire  inst_SnxnLv3Inst59_io_z; // @[Snxn100k.scala 6318:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst56_io_z + inst_SnxnLv3Inst57_io_z; // @[Snxn100k.scala 6322:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst58_io_z; // @[Snxn100k.scala 6322:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst59_io_z; // @[Snxn100k.scala 6322:89]
  SnxnLv3Inst56 inst_SnxnLv3Inst56 ( // @[Snxn100k.scala 6306:34]
    .io_a(inst_SnxnLv3Inst56_io_a),
    .io_b(inst_SnxnLv3Inst56_io_b),
    .io_z(inst_SnxnLv3Inst56_io_z)
  );
  SnxnLv3Inst57 inst_SnxnLv3Inst57 ( // @[Snxn100k.scala 6310:34]
    .io_a(inst_SnxnLv3Inst57_io_a),
    .io_b(inst_SnxnLv3Inst57_io_b),
    .io_z(inst_SnxnLv3Inst57_io_z)
  );
  SnxnLv3Inst58 inst_SnxnLv3Inst58 ( // @[Snxn100k.scala 6314:34]
    .io_a(inst_SnxnLv3Inst58_io_a),
    .io_b(inst_SnxnLv3Inst58_io_b),
    .io_z(inst_SnxnLv3Inst58_io_z)
  );
  SnxnLv3Inst59 inst_SnxnLv3Inst59 ( // @[Snxn100k.scala 6318:34]
    .io_a(inst_SnxnLv3Inst59_io_a),
    .io_b(inst_SnxnLv3Inst59_io_b),
    .io_z(inst_SnxnLv3Inst59_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 6323:15]
  assign inst_SnxnLv3Inst56_io_a = io_a; // @[Snxn100k.scala 6307:27]
  assign inst_SnxnLv3Inst56_io_b = io_b; // @[Snxn100k.scala 6308:27]
  assign inst_SnxnLv3Inst57_io_a = io_a; // @[Snxn100k.scala 6311:27]
  assign inst_SnxnLv3Inst57_io_b = io_b; // @[Snxn100k.scala 6312:27]
  assign inst_SnxnLv3Inst58_io_a = io_a; // @[Snxn100k.scala 6315:27]
  assign inst_SnxnLv3Inst58_io_b = io_b; // @[Snxn100k.scala 6316:27]
  assign inst_SnxnLv3Inst59_io_a = io_a; // @[Snxn100k.scala 6319:27]
  assign inst_SnxnLv3Inst59_io_b = io_b; // @[Snxn100k.scala 6320:27]
endmodule
module SnxnLv3Inst60(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst240_io_a; // @[Snxn100k.scala 24432:35]
  wire  inst_SnxnLv4Inst240_io_b; // @[Snxn100k.scala 24432:35]
  wire  inst_SnxnLv4Inst240_io_z; // @[Snxn100k.scala 24432:35]
  wire  inst_SnxnLv4Inst241_io_a; // @[Snxn100k.scala 24436:35]
  wire  inst_SnxnLv4Inst241_io_b; // @[Snxn100k.scala 24436:35]
  wire  inst_SnxnLv4Inst241_io_z; // @[Snxn100k.scala 24436:35]
  wire  sum = inst_SnxnLv4Inst240_io_z + inst_SnxnLv4Inst241_io_z; // @[Snxn100k.scala 24440:38]
  SnxnLv4Inst23 inst_SnxnLv4Inst240 ( // @[Snxn100k.scala 24432:35]
    .io_a(inst_SnxnLv4Inst240_io_a),
    .io_b(inst_SnxnLv4Inst240_io_b),
    .io_z(inst_SnxnLv4Inst240_io_z)
  );
  SnxnLv4Inst19 inst_SnxnLv4Inst241 ( // @[Snxn100k.scala 24436:35]
    .io_a(inst_SnxnLv4Inst241_io_a),
    .io_b(inst_SnxnLv4Inst241_io_b),
    .io_z(inst_SnxnLv4Inst241_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 24441:15]
  assign inst_SnxnLv4Inst240_io_a = io_a; // @[Snxn100k.scala 24433:28]
  assign inst_SnxnLv4Inst240_io_b = io_b; // @[Snxn100k.scala 24434:28]
  assign inst_SnxnLv4Inst241_io_a = io_a; // @[Snxn100k.scala 24437:28]
  assign inst_SnxnLv4Inst241_io_b = io_b; // @[Snxn100k.scala 24438:28]
endmodule
module SnxnLv3Inst61(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 23675:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 23676:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 23677:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 23678:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 23679:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 23680:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 23681:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 23682:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 23683:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 23684:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 23685:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 23686:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 23687:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 23688:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 23689:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 23690:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 23691:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 23692:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 23693:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 23694:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 23695:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 23696:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 23697:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 23698:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 23699:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 23700:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 23701:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 23702:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 23703:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 23704:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 23705:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 23706:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 23707:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 23708:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 23709:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 23710:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 23711:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 23712:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 23713:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 23714:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 23715:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 23716:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 23717:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 23718:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 23719:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 23720:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 23721:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 23722:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 23723:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 23724:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 23725:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 23726:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 23727:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 23728:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 23729:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 23730:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 23731:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 23732:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 23733:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 23734:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 23735:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 23736:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 23737:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 23738:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 23739:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 23740:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 23741:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 23742:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 23743:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 23744:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 23745:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 23746:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 23747:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 23748:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 23749:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 23750:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 23751:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 23752:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 23753:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 23754:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 23755:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 23756:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 23757:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 23758:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 23759:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 23760:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 23761:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 23762:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 23763:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 23764:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 23765:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 23766:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 23767:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 23768:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 23769:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 23770:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 23771:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 23772:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 23773:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 23774:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 23775:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 23776:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 23777:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 23778:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 23779:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 23780:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 23781:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 23782:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 23783:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 23784:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 23785:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 23786:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 23787:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 23788:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 23789:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 23790:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 23791:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 23792:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 23793:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 23794:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 23795:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 23796:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 23797:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 23798:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 23799:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 23800:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 23801:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 23802:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 23803:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 23804:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 23805:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 23806:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 23807:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 23808:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 23809:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 23810:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 23811:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 23812:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 23813:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 23814:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 23815:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 23816:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 23817:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 23818:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 23819:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 23820:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 23821:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 23822:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 23823:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 23824:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 23825:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 23826:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 23827:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 23828:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 23829:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 23830:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 23831:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 23832:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 23833:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 23834:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 23835:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 23836:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 23837:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 23838:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 23839:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 23840:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 23841:20]
  assign io_z = ~x41; // @[Snxn100k.scala 23842:16]
endmodule
module SnxnLv2Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst60_io_a; // @[Snxn100k.scala 5955:34]
  wire  inst_SnxnLv3Inst60_io_b; // @[Snxn100k.scala 5955:34]
  wire  inst_SnxnLv3Inst60_io_z; // @[Snxn100k.scala 5955:34]
  wire  inst_SnxnLv3Inst61_io_a; // @[Snxn100k.scala 5959:34]
  wire  inst_SnxnLv3Inst61_io_b; // @[Snxn100k.scala 5959:34]
  wire  inst_SnxnLv3Inst61_io_z; // @[Snxn100k.scala 5959:34]
  wire  inst_SnxnLv3Inst62_io_a; // @[Snxn100k.scala 5963:34]
  wire  inst_SnxnLv3Inst62_io_b; // @[Snxn100k.scala 5963:34]
  wire  inst_SnxnLv3Inst62_io_z; // @[Snxn100k.scala 5963:34]
  wire  inst_SnxnLv3Inst63_io_a; // @[Snxn100k.scala 5967:34]
  wire  inst_SnxnLv3Inst63_io_b; // @[Snxn100k.scala 5967:34]
  wire  inst_SnxnLv3Inst63_io_z; // @[Snxn100k.scala 5967:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst60_io_z + inst_SnxnLv3Inst61_io_z; // @[Snxn100k.scala 5971:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst62_io_z; // @[Snxn100k.scala 5971:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst63_io_z; // @[Snxn100k.scala 5971:89]
  SnxnLv3Inst60 inst_SnxnLv3Inst60 ( // @[Snxn100k.scala 5955:34]
    .io_a(inst_SnxnLv3Inst60_io_a),
    .io_b(inst_SnxnLv3Inst60_io_b),
    .io_z(inst_SnxnLv3Inst60_io_z)
  );
  SnxnLv3Inst61 inst_SnxnLv3Inst61 ( // @[Snxn100k.scala 5959:34]
    .io_a(inst_SnxnLv3Inst61_io_a),
    .io_b(inst_SnxnLv3Inst61_io_b),
    .io_z(inst_SnxnLv3Inst61_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv3Inst62 ( // @[Snxn100k.scala 5963:34]
    .io_a(inst_SnxnLv3Inst62_io_a),
    .io_b(inst_SnxnLv3Inst62_io_b),
    .io_z(inst_SnxnLv3Inst62_io_z)
  );
  SnxnLv4Inst151 inst_SnxnLv3Inst63 ( // @[Snxn100k.scala 5967:34]
    .io_a(inst_SnxnLv3Inst63_io_a),
    .io_b(inst_SnxnLv3Inst63_io_b),
    .io_z(inst_SnxnLv3Inst63_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 5972:15]
  assign inst_SnxnLv3Inst60_io_a = io_a; // @[Snxn100k.scala 5956:27]
  assign inst_SnxnLv3Inst60_io_b = io_b; // @[Snxn100k.scala 5957:27]
  assign inst_SnxnLv3Inst61_io_a = io_a; // @[Snxn100k.scala 5960:27]
  assign inst_SnxnLv3Inst61_io_b = io_b; // @[Snxn100k.scala 5961:27]
  assign inst_SnxnLv3Inst62_io_a = io_a; // @[Snxn100k.scala 5964:27]
  assign inst_SnxnLv3Inst62_io_b = io_b; // @[Snxn100k.scala 5965:27]
  assign inst_SnxnLv3Inst63_io_a = io_a; // @[Snxn100k.scala 5968:27]
  assign inst_SnxnLv3Inst63_io_b = io_b; // @[Snxn100k.scala 5969:27]
endmodule
module SnxnLv1Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst12_io_a; // @[Snxn100k.scala 1341:34]
  wire  inst_SnxnLv2Inst12_io_b; // @[Snxn100k.scala 1341:34]
  wire  inst_SnxnLv2Inst12_io_z; // @[Snxn100k.scala 1341:34]
  wire  inst_SnxnLv2Inst13_io_a; // @[Snxn100k.scala 1345:34]
  wire  inst_SnxnLv2Inst13_io_b; // @[Snxn100k.scala 1345:34]
  wire  inst_SnxnLv2Inst13_io_z; // @[Snxn100k.scala 1345:34]
  wire  inst_SnxnLv2Inst14_io_a; // @[Snxn100k.scala 1349:34]
  wire  inst_SnxnLv2Inst14_io_b; // @[Snxn100k.scala 1349:34]
  wire  inst_SnxnLv2Inst14_io_z; // @[Snxn100k.scala 1349:34]
  wire  inst_SnxnLv2Inst15_io_a; // @[Snxn100k.scala 1353:34]
  wire  inst_SnxnLv2Inst15_io_b; // @[Snxn100k.scala 1353:34]
  wire  inst_SnxnLv2Inst15_io_z; // @[Snxn100k.scala 1353:34]
  wire  _sum_T_1 = inst_SnxnLv2Inst12_io_z + inst_SnxnLv2Inst13_io_z; // @[Snxn100k.scala 1357:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst14_io_z; // @[Snxn100k.scala 1357:63]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst15_io_z; // @[Snxn100k.scala 1357:89]
  SnxnLv2Inst12 inst_SnxnLv2Inst12 ( // @[Snxn100k.scala 1341:34]
    .io_a(inst_SnxnLv2Inst12_io_a),
    .io_b(inst_SnxnLv2Inst12_io_b),
    .io_z(inst_SnxnLv2Inst12_io_z)
  );
  SnxnLv2Inst13 inst_SnxnLv2Inst13 ( // @[Snxn100k.scala 1345:34]
    .io_a(inst_SnxnLv2Inst13_io_a),
    .io_b(inst_SnxnLv2Inst13_io_b),
    .io_z(inst_SnxnLv2Inst13_io_z)
  );
  SnxnLv2Inst14 inst_SnxnLv2Inst14 ( // @[Snxn100k.scala 1349:34]
    .io_a(inst_SnxnLv2Inst14_io_a),
    .io_b(inst_SnxnLv2Inst14_io_b),
    .io_z(inst_SnxnLv2Inst14_io_z)
  );
  SnxnLv2Inst15 inst_SnxnLv2Inst15 ( // @[Snxn100k.scala 1353:34]
    .io_a(inst_SnxnLv2Inst15_io_a),
    .io_b(inst_SnxnLv2Inst15_io_b),
    .io_z(inst_SnxnLv2Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1358:15]
  assign inst_SnxnLv2Inst12_io_a = io_a; // @[Snxn100k.scala 1342:27]
  assign inst_SnxnLv2Inst12_io_b = io_b; // @[Snxn100k.scala 1343:27]
  assign inst_SnxnLv2Inst13_io_a = io_a; // @[Snxn100k.scala 1346:27]
  assign inst_SnxnLv2Inst13_io_b = io_b; // @[Snxn100k.scala 1347:27]
  assign inst_SnxnLv2Inst14_io_a = io_a; // @[Snxn100k.scala 1350:27]
  assign inst_SnxnLv2Inst14_io_b = io_b; // @[Snxn100k.scala 1351:27]
  assign inst_SnxnLv2Inst15_io_a = io_a; // @[Snxn100k.scala 1354:27]
  assign inst_SnxnLv2Inst15_io_b = io_b; // @[Snxn100k.scala 1355:27]
endmodule
module Snxn100k(
  input   clock,
  input   reset,
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv1Inst0_io_a; // @[Snxn100k.scala 421:33]
  wire  inst_SnxnLv1Inst0_io_b; // @[Snxn100k.scala 421:33]
  wire  inst_SnxnLv1Inst0_io_z; // @[Snxn100k.scala 421:33]
  wire  inst_SnxnLv1Inst1_io_a; // @[Snxn100k.scala 425:33]
  wire  inst_SnxnLv1Inst1_io_b; // @[Snxn100k.scala 425:33]
  wire  inst_SnxnLv1Inst1_io_z; // @[Snxn100k.scala 425:33]
  wire  inst_SnxnLv1Inst2_io_a; // @[Snxn100k.scala 429:33]
  wire  inst_SnxnLv1Inst2_io_b; // @[Snxn100k.scala 429:33]
  wire  inst_SnxnLv1Inst2_io_z; // @[Snxn100k.scala 429:33]
  wire  inst_SnxnLv1Inst3_io_a; // @[Snxn100k.scala 433:33]
  wire  inst_SnxnLv1Inst3_io_b; // @[Snxn100k.scala 433:33]
  wire  inst_SnxnLv1Inst3_io_z; // @[Snxn100k.scala 433:33]
  wire  _sum_T_1 = inst_SnxnLv1Inst0_io_z + inst_SnxnLv1Inst1_io_z; // @[Snxn100k.scala 437:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv1Inst2_io_z; // @[Snxn100k.scala 437:61]
  wire  sum = _sum_T_3 + inst_SnxnLv1Inst3_io_z; // @[Snxn100k.scala 437:86]
  SnxnLv1Inst0 inst_SnxnLv1Inst0 ( // @[Snxn100k.scala 421:33]
    .io_a(inst_SnxnLv1Inst0_io_a),
    .io_b(inst_SnxnLv1Inst0_io_b),
    .io_z(inst_SnxnLv1Inst0_io_z)
  );
  SnxnLv1Inst1 inst_SnxnLv1Inst1 ( // @[Snxn100k.scala 425:33]
    .io_a(inst_SnxnLv1Inst1_io_a),
    .io_b(inst_SnxnLv1Inst1_io_b),
    .io_z(inst_SnxnLv1Inst1_io_z)
  );
  SnxnLv1Inst2 inst_SnxnLv1Inst2 ( // @[Snxn100k.scala 429:33]
    .io_a(inst_SnxnLv1Inst2_io_a),
    .io_b(inst_SnxnLv1Inst2_io_b),
    .io_z(inst_SnxnLv1Inst2_io_z)
  );
  SnxnLv1Inst3 inst_SnxnLv1Inst3 ( // @[Snxn100k.scala 433:33]
    .io_a(inst_SnxnLv1Inst3_io_a),
    .io_b(inst_SnxnLv1Inst3_io_b),
    .io_z(inst_SnxnLv1Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 438:15]
  assign inst_SnxnLv1Inst0_io_a = io_a; // @[Snxn100k.scala 422:26]
  assign inst_SnxnLv1Inst0_io_b = io_b; // @[Snxn100k.scala 423:26]
  assign inst_SnxnLv1Inst1_io_a = io_a; // @[Snxn100k.scala 426:26]
  assign inst_SnxnLv1Inst1_io_b = io_b; // @[Snxn100k.scala 427:26]
  assign inst_SnxnLv1Inst2_io_a = io_a; // @[Snxn100k.scala 430:26]
  assign inst_SnxnLv1Inst2_io_b = io_b; // @[Snxn100k.scala 431:26]
  assign inst_SnxnLv1Inst3_io_a = io_a; // @[Snxn100k.scala 434:26]
  assign inst_SnxnLv1Inst3_io_b = io_b; // @[Snxn100k.scala 435:26]
endmodule
