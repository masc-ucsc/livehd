module lhs_wire2 (
  output [1:0] out,
  output [2:0] out2
);

assign out  = 2'd2;
assign out2 = 3'd5;

endmodule 
