module sum2 (
  input  [1:0] a,
  input  [1:0] b,
  output [2:0] o
);

assign o = a + b;

endmodule
