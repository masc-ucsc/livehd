module IntXbar(
   input signed [1:0] reset
  ,input signed clock
  ,input signed \auto_int_in_0 
  ,output reg signed \auto_int_out 
);
always_comb begin
  \auto_int_out  = \auto_int_in_0 ;
end
endmodule
