
module trivial3( \a[0] , \a[1] , \c[0] );
  input \a[0] , \a[1] ;
  output \c[0] ;
  assign \c[0]  = \a[0] ^ \a[1] ;
endmodule

