
module null_port(input a, output b, output c);

assign b = ~a;

endmodule

