module capricious_bits2(
  output [4:0] out
);

assign out = 5'd10;

endmodule
