module SnxnLv4Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 70049:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 70050:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 70051:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 70052:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 70053:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 70054:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 70055:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 70056:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 70057:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 70058:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 70059:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 70060:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 70061:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 70062:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 70063:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 70064:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 70065:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 70066:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 70067:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 70068:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 70069:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 70070:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 70071:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 70072:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 70073:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 70074:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 70075:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 70076:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 70077:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 70078:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 70079:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 70080:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 70081:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 70082:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 70083:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 70084:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 70085:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 70086:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 70087:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 70088:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 70089:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 70090:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 70091:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 70092:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 70093:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 70094:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 70095:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 70096:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 70097:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 70098:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 70099:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 70100:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 70101:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 70102:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 70103:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 70104:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 70105:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 70106:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 70107:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 70108:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 70109:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 70110:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 70111:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 70112:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 70113:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 70114:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 70115:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 70116:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 70117:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 70118:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 70119:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 70120:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 70121:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 70122:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 70123:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 70124:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 70125:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 70126:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 70127:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 70128:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 70129:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 70130:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 70131:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 70132:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 70133:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 70134:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 70135:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 70136:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 70137:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 70138:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 70139:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 70140:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 70141:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 70142:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 70143:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 70144:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 70145:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 70146:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 70147:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 70148:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 70149:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 70150:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 70151:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 70152:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 70153:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 70154:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 70155:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 70156:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 70157:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 70158:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 70159:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 70160:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 70161:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 70162:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 70163:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 70164:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 70165:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 70166:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 70167:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 70168:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 70169:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 70170:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 70171:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 70172:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 70173:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 70174:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 70175:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 70176:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 70177:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 70178:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 70179:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 70180:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 70181:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 70182:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 70183:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 70184:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 70185:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 70186:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 70187:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 70188:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 70189:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 70190:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 70191:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 70192:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 70193:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 70194:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 70195:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 70196:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 70197:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 70198:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 70199:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 70200:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 70201:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 70202:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 70203:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 70204:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 70205:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 70206:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 70207:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 70208:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 70209:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 70210:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 70211:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 70212:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 70213:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 70214:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 70215:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 70216:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 70217:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 70218:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 70219:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 70220:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 70221:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 70222:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 70223:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 70224:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 70225:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 70226:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 70227:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 70228:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 70229:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 70230:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 70231:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 70232:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 70233:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 70234:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 70235:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 70236:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 70237:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 70238:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 70239:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 70240:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 70241:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 70242:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 70243:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 70244:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 70245:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 70246:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 70247:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 70248:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 70249:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 70250:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 70251:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 70252:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 70253:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 70254:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 70255:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 70256:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 70257:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 70258:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 70259:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 70260:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 70261:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 70262:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 70263:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 70264:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 70265:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 70266:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 70267:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 70268:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 70269:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 70270:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 70271:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 70272:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 70273:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 70274:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 70275:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 70276:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 70277:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 70278:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 70279:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 70280:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 70281:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 70282:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 70283:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 70284:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 70285:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 70286:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 70287:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 70288:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 70289:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 70290:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 70291:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 70292:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 70293:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 70294:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 70295:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 70296:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 70297:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 70298:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 70299:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 70300:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 70301:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 70302:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 70303:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 70304:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 70305:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 70306:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 70307:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 70308:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 70309:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 70310:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 70311:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 70312:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 70313:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 70314:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 70315:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 70316:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 70317:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 70318:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 70319:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 70320:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 70321:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 70322:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 70323:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 70324:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 70325:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 70326:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 70327:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 70328:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 70329:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 70330:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 70331:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 70332:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 70333:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 70334:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 70335:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 70336:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 70337:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 70338:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 70339:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 70340:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 70341:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 70342:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 70343:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 70344:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 70345:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 70346:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 70347:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 70348:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 70349:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 70350:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 70351:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 70352:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 70353:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 70354:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 70355:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 70356:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 70357:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 70358:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 70359:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 70360:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 70361:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 70362:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 70363:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 70364:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 70365:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 70366:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 70367:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 70368:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 70369:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 70370:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 70371:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 70372:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 70373:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 70374:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 70375:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 70376:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 70377:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 70378:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 70379:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 70380:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 70381:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 70382:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 70383:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 70384:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 70385:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 70386:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 70387:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 70388:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 70389:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 70390:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 70391:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 70392:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 70393:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 70394:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 70395:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 70396:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 70397:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 70398:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 70399:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 70400:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 70401:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 70402:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 70403:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 70404:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 70405:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 70406:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 70407:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 70408:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 70409:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 70410:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 70411:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 70412:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 70413:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 70414:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 70415:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 70416:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 70417:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 70418:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 70419:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 70420:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 70421:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 70422:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 70423:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 70424:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 70425:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 70426:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 70427:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 70428:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 70429:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 70430:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 70431:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 70432:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 70433:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 70434:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 70435:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 70436:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 70437:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 70438:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 70439:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 70440:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 70441:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 70442:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 70443:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 70444:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 70445:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 70446:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 70447:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 70448:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 70449:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 70450:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 70451:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 70452:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 70453:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 70454:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 70455:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 70456:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 70457:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 70458:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 70459:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 70460:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 70461:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 70462:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 70463:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 70464:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 70465:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 70466:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 70467:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 70468:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 70469:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 70470:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 70471:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 70472:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 70473:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 70474:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 70475:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 70476:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 70477:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 70478:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 70479:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 70480:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 70481:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 70482:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 70483:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 70484:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 70485:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 70486:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 70487:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 70488:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 70489:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 70490:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 70491:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 70492:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 70493:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 70494:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 70495:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 70496:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 70497:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 70498:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 70499:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 70500:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 70501:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 70502:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 70503:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 70504:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 70505:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 70506:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 70507:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 70508:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 70509:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 70510:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 70511:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 70512:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 70513:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 70514:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 70515:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 70516:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 70517:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 70518:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 70519:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 70520:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 70521:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 70522:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 70523:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 70524:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 70525:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 70526:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 70527:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 70528:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 70529:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 70530:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 70531:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 70532:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 70533:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 70534:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 70535:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 70536:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 70537:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 70538:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 70539:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 70540:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 70541:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 70542:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 70543:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 70544:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 70545:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 70546:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 70547:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 70548:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 70549:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 70550:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 70551:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 70552:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 70553:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 70554:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 70555:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 70556:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 70557:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 70558:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 70559:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 70560:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 70561:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 70562:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 70563:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 70564:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 70565:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 70566:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 70567:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 70568:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 70569:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 70570:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 70571:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 70572:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 70573:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 70574:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 70575:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 70576:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 70577:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 70578:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 70579:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 70580:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 70581:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 70582:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 70583:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 70584:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 70585:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 70586:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 70587:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 70588:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 70589:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 70590:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 70591:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 70592:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 70593:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 70594:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 70595:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 70596:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 70597:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 70598:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 70599:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 70600:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 70601:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 70602:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 70603:22]
  assign io_z = ~x138; // @[Snxn100k.scala 70604:17]
endmodule
module SnxnLv4Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 69221:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 69222:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 69223:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 69224:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 69225:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 69226:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 69227:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 69228:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 69229:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 69230:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 69231:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 69232:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 69233:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 69234:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 69235:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 69236:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 69237:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 69238:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 69239:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 69240:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 69241:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 69242:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 69243:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 69244:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 69245:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 69246:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 69247:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 69248:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 69249:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 69250:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 69251:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 69252:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 69253:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 69254:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 69255:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 69256:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 69257:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 69258:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 69259:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 69260:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 69261:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 69262:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 69263:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 69264:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 69265:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 69266:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 69267:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 69268:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 69269:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 69270:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 69271:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 69272:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 69273:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 69274:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 69275:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 69276:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 69277:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 69278:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 69279:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 69280:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 69281:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 69282:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 69283:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 69284:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 69285:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 69286:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 69287:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 69288:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 69289:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 69290:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 69291:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 69292:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 69293:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 69294:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 69295:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 69296:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 69297:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 69298:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 69299:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 69300:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 69301:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 69302:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 69303:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 69304:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 69305:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 69306:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 69307:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 69308:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 69309:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 69310:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 69311:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 69312:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 69313:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 69314:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 69315:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 69316:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 69317:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 69318:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 69319:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 69320:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 69321:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 69322:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 69323:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 69324:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 69325:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 69326:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 69327:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 69328:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 69329:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 69330:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 69331:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 69332:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 69333:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 69334:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 69335:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 69336:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 69337:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 69338:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69339:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69340:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69341:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69342:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69343:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69344:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69345:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69346:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69347:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69348:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69349:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69350:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69351:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69352:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69353:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69354:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69355:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69356:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69357:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69358:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69359:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69360:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69361:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69362:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69363:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69364:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69365:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69366:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69367:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69368:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69369:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69370:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69371:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69372:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69373:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69374:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69375:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69376:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69377:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69378:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69379:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69380:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69381:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69382:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69383:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69384:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69385:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69386:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69387:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69388:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69389:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69390:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69391:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69392:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69393:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69394:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69395:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69396:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69397:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69398:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69399:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69400:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69401:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69402:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69403:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69404:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69405:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69406:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69407:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69408:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69409:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69410:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69411:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 69412:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 69413:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 69414:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 69415:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 69416:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 69417:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 69418:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 69419:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 69420:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 69421:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 69422:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 69423:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 69424:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 69425:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 69426:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 69427:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 69428:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 69429:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 69430:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 69431:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 69432:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 69433:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 69434:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 69435:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 69436:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 69437:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 69438:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 69439:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 69440:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 69441:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 69442:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 69443:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 69444:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 69445:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 69446:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 69447:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 69448:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 69449:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 69450:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 69451:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 69452:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 69453:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 69454:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 69455:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 69456:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 69457:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 69458:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 69459:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 69460:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 69461:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 69462:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 69463:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 69464:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 69465:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 69466:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 69467:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 69468:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 69469:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 69470:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 69471:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 69472:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 69473:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 69474:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 69475:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 69476:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 69477:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 69478:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 69479:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 69480:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 69481:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 69482:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 69483:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 69484:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 69485:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 69486:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 69487:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 69488:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 69489:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 69490:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 69491:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 69492:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 69493:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 69494:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 69495:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 69496:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 69497:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 69498:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 69499:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 69500:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 69501:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 69502:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 69503:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 69504:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 69505:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 69506:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 69507:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 69508:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 69509:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 69510:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 69511:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 69512:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 69513:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 69514:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 69515:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 69516:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 69517:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 69518:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 69519:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 69520:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 69521:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 69522:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 69523:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 69524:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 69525:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 69526:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 69527:20]
  assign io_z = ~x76; // @[Snxn100k.scala 69528:16]
endmodule
module SnxnLv4Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 69539:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 69540:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 69541:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 69542:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 69543:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 69544:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 69545:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 69546:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 69547:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 69548:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 69549:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 69550:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 69551:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 69552:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 69553:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 69554:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 69555:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 69556:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 69557:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 69558:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 69559:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 69560:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 69561:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 69562:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 69563:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 69564:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 69565:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 69566:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 69567:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 69568:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 69569:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 69570:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 69571:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 69572:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 69573:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 69574:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 69575:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 69576:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 69577:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 69578:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 69579:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 69580:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 69581:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 69582:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 69583:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 69584:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 69585:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 69586:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 69587:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 69588:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 69589:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 69590:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 69591:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 69592:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 69593:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 69594:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 69595:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 69596:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 69597:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 69598:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 69599:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 69600:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 69601:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 69602:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 69603:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 69604:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 69605:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 69606:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 69607:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 69608:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 69609:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 69610:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 69611:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 69612:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 69613:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 69614:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 69615:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 69616:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 69617:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 69618:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 69619:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 69620:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 69621:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 69622:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 69623:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 69624:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 69625:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 69626:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 69627:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 69628:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 69629:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 69630:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 69631:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 69632:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 69633:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 69634:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 69635:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 69636:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 69637:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 69638:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 69639:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 69640:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 69641:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 69642:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 69643:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 69644:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 69645:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 69646:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 69647:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 69648:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 69649:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 69650:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 69651:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 69652:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 69653:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 69654:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 69655:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 69656:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69657:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69658:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69659:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69660:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69661:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69662:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69663:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69664:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69665:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69666:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69667:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69668:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69669:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69670:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69671:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69672:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69673:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69674:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69675:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69676:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69677:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69678:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69679:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69680:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69681:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69682:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69683:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69684:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69685:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69686:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69687:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69688:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69689:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69690:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69691:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69692:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69693:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69694:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69695:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69696:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69697:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69698:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69699:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69700:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69701:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69702:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69703:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69704:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69705:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69706:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69707:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69708:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69709:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69710:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69711:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69712:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69713:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69714:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69715:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69716:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69717:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69718:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69719:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69720:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69721:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69722:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69723:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69724:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69725:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69726:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69727:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69728:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69729:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 69730:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 69731:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 69732:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 69733:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 69734:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 69735:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 69736:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 69737:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 69738:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 69739:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 69740:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 69741:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 69742:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 69743:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 69744:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 69745:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 69746:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 69747:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 69748:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 69749:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 69750:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 69751:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 69752:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 69753:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 69754:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 69755:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 69756:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 69757:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 69758:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 69759:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 69760:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 69761:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 69762:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 69763:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 69764:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 69765:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 69766:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 69767:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 69768:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 69769:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 69770:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 69771:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 69772:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 69773:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 69774:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 69775:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 69776:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 69777:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 69778:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 69779:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 69780:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 69781:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 69782:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 69783:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 69784:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 69785:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 69786:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 69787:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 69788:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 69789:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 69790:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 69791:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 69792:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 69793:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 69794:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 69795:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 69796:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 69797:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 69798:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 69799:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 69800:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 69801:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 69802:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 69803:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 69804:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 69805:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 69806:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 69807:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 69808:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 69809:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 69810:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 69811:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 69812:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 69813:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 69814:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 69815:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 69816:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 69817:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 69818:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 69819:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 69820:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 69821:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 69822:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 69823:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 69824:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 69825:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 69826:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 69827:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 69828:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 69829:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 69830:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 69831:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 69832:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 69833:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 69834:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 69835:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 69836:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 69837:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 69838:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 69839:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 69840:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 69841:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 69842:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 69843:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 69844:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 69845:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 69846:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 69847:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 69848:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 69849:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 69850:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 69851:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 69852:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 69853:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 69854:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 69855:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 69856:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 69857:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 69858:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 69859:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 69860:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 69861:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 69862:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 69863:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 69864:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 69865:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 69866:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 69867:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 69868:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 69869:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 69870:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 69871:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 69872:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 69873:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 69874:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 69875:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 69876:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 69877:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 69878:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 69879:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 69880:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 69881:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 69882:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 69883:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 69884:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 69885:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 69886:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 69887:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 69888:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 69889:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 69890:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 69891:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 69892:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 69893:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 69894:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 69895:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 69896:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 69897:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 69898:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 69899:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 69900:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 69901:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 69902:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 69903:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 69904:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 69905:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 69906:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 69907:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 69908:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 69909:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 69910:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 69911:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 69912:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 69913:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 69914:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 69915:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 69916:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 69917:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 69918:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 69919:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 69920:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 69921:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 69922:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 69923:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 69924:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 69925:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 69926:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 69927:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 69928:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 69929:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 69930:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 69931:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 69932:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 69933:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 69934:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 69935:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 69936:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 69937:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 69938:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 69939:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 69940:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 69941:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 69942:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 69943:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 69944:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 69945:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 69946:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 69947:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 69948:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 69949:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 69950:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 69951:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 69952:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 69953:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 69954:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 69955:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 69956:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 69957:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 69958:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 69959:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 69960:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 69961:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 69962:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 69963:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 69964:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 69965:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 69966:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 69967:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 69968:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 69969:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 69970:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 69971:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 69972:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 69973:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 69974:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 69975:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 69976:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 69977:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 69978:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 69979:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 69980:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 69981:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 69982:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 69983:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 69984:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 69985:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 69986:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 69987:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 69988:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 69989:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 69990:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 69991:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 69992:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 69993:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 69994:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 69995:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 69996:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 69997:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 69998:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 69999:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 70000:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 70001:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 70002:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 70003:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 70004:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 70005:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 70006:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 70007:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 70008:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 70009:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 70010:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 70011:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 70012:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 70013:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 70014:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 70015:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 70016:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 70017:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 70018:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 70019:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 70020:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 70021:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 70022:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 70023:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 70024:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 70025:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 70026:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 70027:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 70028:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 70029:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 70030:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 70031:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 70032:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 70033:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 70034:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 70035:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 70036:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 70037:22]
  assign io_z = ~x124; // @[Snxn100k.scala 70038:17]
endmodule
module SnxnLv4Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 68979:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 68980:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 68981:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 68982:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 68983:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 68984:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 68985:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 68986:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 68987:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 68988:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 68989:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 68990:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 68991:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 68992:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 68993:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 68994:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 68995:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 68996:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 68997:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 68998:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 68999:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 69000:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 69001:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 69002:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 69003:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 69004:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 69005:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 69006:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 69007:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 69008:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 69009:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 69010:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 69011:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 69012:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 69013:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 69014:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 69015:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 69016:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 69017:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 69018:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 69019:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 69020:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 69021:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 69022:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 69023:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 69024:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 69025:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 69026:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 69027:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 69028:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 69029:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 69030:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 69031:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 69032:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 69033:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 69034:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 69035:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 69036:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 69037:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 69038:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 69039:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 69040:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 69041:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 69042:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 69043:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 69044:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 69045:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 69046:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 69047:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 69048:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 69049:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 69050:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 69051:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 69052:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 69053:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 69054:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 69055:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 69056:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 69057:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 69058:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 69059:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 69060:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 69061:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 69062:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 69063:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 69064:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 69065:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 69066:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 69067:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 69068:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 69069:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 69070:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 69071:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 69072:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 69073:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 69074:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 69075:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 69076:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 69077:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 69078:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 69079:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 69080:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 69081:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 69082:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 69083:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 69084:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 69085:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 69086:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 69087:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 69088:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 69089:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 69090:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 69091:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 69092:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 69093:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 69094:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 69095:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 69096:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 69097:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 69098:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 69099:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 69100:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 69101:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 69102:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 69103:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 69104:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 69105:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 69106:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 69107:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 69108:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 69109:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 69110:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 69111:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 69112:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 69113:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 69114:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 69115:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 69116:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 69117:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 69118:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 69119:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 69120:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 69121:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 69122:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 69123:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 69124:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 69125:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 69126:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 69127:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 69128:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 69129:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 69130:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 69131:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 69132:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 69133:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 69134:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 69135:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 69136:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 69137:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 69138:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 69139:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 69140:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 69141:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 69142:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 69143:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 69144:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 69145:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 69146:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 69147:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 69148:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 69149:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 69150:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 69151:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 69152:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 69153:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 69154:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 69155:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 69156:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 69157:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 69158:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 69159:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 69160:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 69161:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 69162:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 69163:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 69164:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 69165:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 69166:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 69167:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 69168:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 69169:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 69170:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 69171:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 69172:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 69173:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 69174:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 69175:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 69176:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 69177:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 69178:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 69179:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 69180:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 69181:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 69182:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 69183:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 69184:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 69185:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 69186:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 69187:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 69188:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 69189:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 69190:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 69191:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 69192:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 69193:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 69194:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 69195:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 69196:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 69197:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 69198:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 69199:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 69200:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 69201:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 69202:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 69203:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 69204:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 69205:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 69206:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 69207:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 69208:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 69209:20]
  assign io_z = ~x57; // @[Snxn100k.scala 69210:16]
endmodule
module SnxnLv3Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst0_io_a; // @[Snxn100k.scala 21950:33]
  wire  inst_SnxnLv4Inst0_io_b; // @[Snxn100k.scala 21950:33]
  wire  inst_SnxnLv4Inst0_io_z; // @[Snxn100k.scala 21950:33]
  wire  inst_SnxnLv4Inst1_io_a; // @[Snxn100k.scala 21954:33]
  wire  inst_SnxnLv4Inst1_io_b; // @[Snxn100k.scala 21954:33]
  wire  inst_SnxnLv4Inst1_io_z; // @[Snxn100k.scala 21954:33]
  wire  inst_SnxnLv4Inst2_io_a; // @[Snxn100k.scala 21958:33]
  wire  inst_SnxnLv4Inst2_io_b; // @[Snxn100k.scala 21958:33]
  wire  inst_SnxnLv4Inst2_io_z; // @[Snxn100k.scala 21958:33]
  wire  inst_SnxnLv4Inst3_io_a; // @[Snxn100k.scala 21962:33]
  wire  inst_SnxnLv4Inst3_io_b; // @[Snxn100k.scala 21962:33]
  wire  inst_SnxnLv4Inst3_io_z; // @[Snxn100k.scala 21962:33]
  wire  _sum_T_1 = inst_SnxnLv4Inst0_io_z + inst_SnxnLv4Inst1_io_z; // @[Snxn100k.scala 21966:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst2_io_z; // @[Snxn100k.scala 21966:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst3_io_z; // @[Snxn100k.scala 21966:86]
  SnxnLv4Inst0 inst_SnxnLv4Inst0 ( // @[Snxn100k.scala 21950:33]
    .io_a(inst_SnxnLv4Inst0_io_a),
    .io_b(inst_SnxnLv4Inst0_io_b),
    .io_z(inst_SnxnLv4Inst0_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst1 ( // @[Snxn100k.scala 21954:33]
    .io_a(inst_SnxnLv4Inst1_io_a),
    .io_b(inst_SnxnLv4Inst1_io_b),
    .io_z(inst_SnxnLv4Inst1_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst2 ( // @[Snxn100k.scala 21958:33]
    .io_a(inst_SnxnLv4Inst2_io_a),
    .io_b(inst_SnxnLv4Inst2_io_b),
    .io_z(inst_SnxnLv4Inst2_io_z)
  );
  SnxnLv4Inst3 inst_SnxnLv4Inst3 ( // @[Snxn100k.scala 21962:33]
    .io_a(inst_SnxnLv4Inst3_io_a),
    .io_b(inst_SnxnLv4Inst3_io_b),
    .io_z(inst_SnxnLv4Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21967:15]
  assign inst_SnxnLv4Inst0_io_a = io_a; // @[Snxn100k.scala 21951:26]
  assign inst_SnxnLv4Inst0_io_b = io_b; // @[Snxn100k.scala 21952:26]
  assign inst_SnxnLv4Inst1_io_a = io_a; // @[Snxn100k.scala 21955:26]
  assign inst_SnxnLv4Inst1_io_b = io_b; // @[Snxn100k.scala 21956:26]
  assign inst_SnxnLv4Inst2_io_a = io_a; // @[Snxn100k.scala 21959:26]
  assign inst_SnxnLv4Inst2_io_b = io_b; // @[Snxn100k.scala 21960:26]
  assign inst_SnxnLv4Inst3_io_a = io_a; // @[Snxn100k.scala 21963:26]
  assign inst_SnxnLv4Inst3_io_b = io_b; // @[Snxn100k.scala 21964:26]
endmodule
module SnxnLv4Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72281:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72282:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72283:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72284:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72285:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72286:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72287:18]
  assign io_z = ~x1; // @[Snxn100k.scala 72288:15]
endmodule
module SnxnLv4Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71575:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71576:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71577:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71578:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71579:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71580:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71581:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71582:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71583:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71584:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71585:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71586:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71587:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71588:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71589:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71590:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71591:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71592:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71593:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71594:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71595:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71596:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71597:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71598:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71599:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71600:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71601:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71602:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71603:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71604:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71605:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71606:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71607:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71608:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71609:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71610:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71611:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71612:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71613:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71614:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71615:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71616:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71617:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71618:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71619:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71620:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71621:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71622:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71623:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71624:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71625:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71626:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71627:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71628:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71629:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71630:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71631:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71632:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71633:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71634:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71635:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71636:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71637:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71638:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71639:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71640:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71641:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71642:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71643:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71644:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71645:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71646:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71647:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71648:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71649:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71650:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71651:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71652:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71653:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71654:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71655:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71656:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71657:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71658:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71659:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71660:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71661:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71662:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71663:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71664:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71665:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71666:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71667:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71668:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71669:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71670:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71671:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71672:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71673:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71674:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71675:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71676:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71677:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71678:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71679:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71680:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71681:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71682:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71683:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71684:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71685:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71686:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71687:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71688:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71689:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71690:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71691:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71692:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71693:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71694:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71695:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71696:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71697:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71698:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71699:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71700:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71701:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71702:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71703:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71704:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71705:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71706:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71707:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71708:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71709:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71710:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71711:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71712:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71713:20]
  assign io_z = ~x34; // @[Snxn100k.scala 71714:16]
endmodule
module SnxnLv4Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71975:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71976:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71977:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71978:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71979:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71980:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71981:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71982:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71983:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71984:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71985:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71986:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71987:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71988:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71989:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71990:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71991:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71992:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71993:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71994:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71995:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71996:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71997:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71998:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71999:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72000:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72001:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72002:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 72003:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 72004:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 72005:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 72006:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 72007:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 72008:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 72009:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 72010:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 72011:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 72012:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 72013:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 72014:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72015:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72016:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72017:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72018:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72019:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72020:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72021:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72022:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72023:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72024:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72025:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72026:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72027:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72028:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72029:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72030:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72031:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72032:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72033:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72034:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72035:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72036:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72037:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72038:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72039:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72040:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72041:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72042:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72043:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72044:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72045:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72046:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72047:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72048:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72049:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72050:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72051:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72052:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72053:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72054:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72055:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72056:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72057:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72058:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72059:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72060:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72061:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72062:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72063:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72064:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72065:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72066:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72067:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72068:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72069:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72070:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72071:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72072:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72073:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 72074:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 72075:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 72076:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 72077:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 72078:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 72079:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 72080:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 72081:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 72082:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 72083:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 72084:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 72085:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 72086:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 72087:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 72088:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 72089:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 72090:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 72091:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 72092:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 72093:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 72094:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 72095:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 72096:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 72097:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 72098:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 72099:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 72100:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 72101:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 72102:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 72103:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 72104:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 72105:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 72106:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 72107:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 72108:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 72109:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 72110:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 72111:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 72112:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 72113:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 72114:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 72115:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 72116:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 72117:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 72118:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 72119:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 72120:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 72121:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 72122:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 72123:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 72124:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 72125:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 72126:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 72127:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 72128:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 72129:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 72130:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 72131:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 72132:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 72133:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 72134:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 72135:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 72136:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 72137:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 72138:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 72139:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 72140:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 72141:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 72142:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 72143:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 72144:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 72145:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 72146:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 72147:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 72148:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 72149:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 72150:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 72151:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 72152:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 72153:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 72154:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 72155:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 72156:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 72157:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 72158:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 72159:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 72160:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 72161:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 72162:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 72163:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 72164:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 72165:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 72166:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 72167:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 72168:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 72169:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 72170:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 72171:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 72172:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 72173:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 72174:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 72175:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 72176:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 72177:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 72178:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 72179:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 72180:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 72181:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 72182:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 72183:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 72184:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 72185:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 72186:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 72187:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 72188:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 72189:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 72190:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 72191:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 72192:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 72193:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 72194:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 72195:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 72196:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 72197:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 72198:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 72199:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 72200:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 72201:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 72202:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 72203:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 72204:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 72205:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 72206:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 72207:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 72208:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 72209:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 72210:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 72211:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 72212:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 72213:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 72214:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 72215:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 72216:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 72217:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 72218:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 72219:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 72220:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 72221:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 72222:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 72223:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 72224:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 72225:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 72226:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 72227:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 72228:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 72229:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 72230:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 72231:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 72232:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 72233:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 72234:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 72235:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 72236:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 72237:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 72238:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 72239:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 72240:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 72241:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 72242:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 72243:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 72244:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 72245:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 72246:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 72247:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 72248:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 72249:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 72250:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 72251:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 72252:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 72253:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 72254:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 72255:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 72256:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 72257:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 72258:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 72259:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 72260:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 72261:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 72262:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 72263:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 72264:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 72265:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 72266:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 72267:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 72268:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 72269:20]
  assign io_z = ~x73; // @[Snxn100k.scala 72270:16]
endmodule
module SnxnLv4Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71725:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71726:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71727:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71728:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71729:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71730:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71731:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71732:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71733:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71734:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71735:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71736:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71737:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71738:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71739:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71740:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71741:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71742:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71743:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71744:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71745:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71746:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71747:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71748:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71749:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71750:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71751:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71752:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71753:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71754:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71755:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71756:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71757:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71758:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71759:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71760:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71761:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71762:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71763:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71764:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71765:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71766:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71767:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71768:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71769:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71770:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71771:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71772:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71773:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71774:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71775:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71776:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71777:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71778:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71779:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71780:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71781:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71782:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71783:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71784:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71785:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71786:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71787:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71788:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71789:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71790:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71791:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71792:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71793:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71794:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71795:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71796:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71797:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71798:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71799:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71800:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71801:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71802:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71803:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71804:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71805:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71806:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71807:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71808:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71809:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71810:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71811:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71812:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71813:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71814:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71815:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71816:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71817:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71818:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71819:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71820:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71821:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71822:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71823:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71824:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71825:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71826:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71827:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71828:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71829:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71830:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71831:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71832:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71833:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71834:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71835:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71836:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71837:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71838:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71839:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71840:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71841:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71842:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71843:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71844:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71845:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71846:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71847:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71848:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71849:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71850:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71851:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71852:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71853:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71854:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71855:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71856:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71857:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71858:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71859:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71860:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71861:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71862:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71863:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 71864:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 71865:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 71866:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 71867:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 71868:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 71869:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 71870:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 71871:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 71872:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 71873:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 71874:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 71875:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 71876:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 71877:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 71878:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 71879:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 71880:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 71881:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 71882:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 71883:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 71884:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 71885:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 71886:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 71887:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 71888:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 71889:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 71890:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 71891:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 71892:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 71893:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 71894:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 71895:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 71896:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 71897:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 71898:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 71899:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 71900:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 71901:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 71902:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 71903:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 71904:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 71905:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 71906:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 71907:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 71908:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 71909:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 71910:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 71911:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 71912:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 71913:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 71914:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 71915:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 71916:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 71917:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 71918:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 71919:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 71920:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 71921:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 71922:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 71923:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 71924:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 71925:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 71926:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 71927:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 71928:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 71929:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 71930:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 71931:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 71932:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 71933:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 71934:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 71935:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 71936:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 71937:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 71938:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 71939:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 71940:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 71941:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 71942:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 71943:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 71944:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 71945:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 71946:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 71947:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 71948:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 71949:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 71950:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 71951:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 71952:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 71953:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 71954:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 71955:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 71956:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 71957:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 71958:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 71959:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 71960:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 71961:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 71962:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 71963:20]
  assign io_z = ~x59; // @[Snxn100k.scala 71964:16]
endmodule
module SnxnLv3Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst4_io_a; // @[Snxn100k.scala 22416:33]
  wire  inst_SnxnLv4Inst4_io_b; // @[Snxn100k.scala 22416:33]
  wire  inst_SnxnLv4Inst4_io_z; // @[Snxn100k.scala 22416:33]
  wire  inst_SnxnLv4Inst5_io_a; // @[Snxn100k.scala 22420:33]
  wire  inst_SnxnLv4Inst5_io_b; // @[Snxn100k.scala 22420:33]
  wire  inst_SnxnLv4Inst5_io_z; // @[Snxn100k.scala 22420:33]
  wire  inst_SnxnLv4Inst6_io_a; // @[Snxn100k.scala 22424:33]
  wire  inst_SnxnLv4Inst6_io_b; // @[Snxn100k.scala 22424:33]
  wire  inst_SnxnLv4Inst6_io_z; // @[Snxn100k.scala 22424:33]
  wire  inst_SnxnLv4Inst7_io_a; // @[Snxn100k.scala 22428:33]
  wire  inst_SnxnLv4Inst7_io_b; // @[Snxn100k.scala 22428:33]
  wire  inst_SnxnLv4Inst7_io_z; // @[Snxn100k.scala 22428:33]
  wire  _sum_T_1 = inst_SnxnLv4Inst4_io_z + inst_SnxnLv4Inst5_io_z; // @[Snxn100k.scala 22432:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst6_io_z; // @[Snxn100k.scala 22432:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst7_io_z; // @[Snxn100k.scala 22432:86]
  SnxnLv4Inst4 inst_SnxnLv4Inst4 ( // @[Snxn100k.scala 22416:33]
    .io_a(inst_SnxnLv4Inst4_io_a),
    .io_b(inst_SnxnLv4Inst4_io_b),
    .io_z(inst_SnxnLv4Inst4_io_z)
  );
  SnxnLv4Inst5 inst_SnxnLv4Inst5 ( // @[Snxn100k.scala 22420:33]
    .io_a(inst_SnxnLv4Inst5_io_a),
    .io_b(inst_SnxnLv4Inst5_io_b),
    .io_z(inst_SnxnLv4Inst5_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst6 ( // @[Snxn100k.scala 22424:33]
    .io_a(inst_SnxnLv4Inst6_io_a),
    .io_b(inst_SnxnLv4Inst6_io_b),
    .io_z(inst_SnxnLv4Inst6_io_z)
  );
  SnxnLv4Inst7 inst_SnxnLv4Inst7 ( // @[Snxn100k.scala 22428:33]
    .io_a(inst_SnxnLv4Inst7_io_a),
    .io_b(inst_SnxnLv4Inst7_io_b),
    .io_z(inst_SnxnLv4Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22433:15]
  assign inst_SnxnLv4Inst4_io_a = io_a; // @[Snxn100k.scala 22417:26]
  assign inst_SnxnLv4Inst4_io_b = io_b; // @[Snxn100k.scala 22418:26]
  assign inst_SnxnLv4Inst5_io_a = io_a; // @[Snxn100k.scala 22421:26]
  assign inst_SnxnLv4Inst5_io_b = io_b; // @[Snxn100k.scala 22422:26]
  assign inst_SnxnLv4Inst6_io_a = io_a; // @[Snxn100k.scala 22425:26]
  assign inst_SnxnLv4Inst6_io_b = io_b; // @[Snxn100k.scala 22426:26]
  assign inst_SnxnLv4Inst7_io_a = io_a; // @[Snxn100k.scala 22429:26]
  assign inst_SnxnLv4Inst7_io_b = io_b; // @[Snxn100k.scala 22430:26]
endmodule
module SnxnLv4Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71011:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71012:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71013:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71014:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71015:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71016:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71017:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71018:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71019:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71020:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71021:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71022:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71023:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71024:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71025:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71026:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71027:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71028:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71029:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71030:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71031:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71032:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71033:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71034:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71035:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71036:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71037:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71038:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71039:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71040:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71041:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71042:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71043:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71044:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71045:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71046:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71047:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71048:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71049:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71050:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71051:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71052:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71053:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71054:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71055:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71056:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71057:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71058:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71059:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71060:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71061:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71062:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71063:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71064:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71065:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71066:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71067:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71068:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71069:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71070:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71071:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71072:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71073:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71074:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71075:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71076:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71077:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71078:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71079:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71080:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71081:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71082:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71083:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71084:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71085:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71086:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71087:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71088:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71089:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71090:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71091:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71092:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71093:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 71094:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 71095:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 71096:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 71097:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 71098:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 71099:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 71100:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 71101:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 71102:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 71103:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 71104:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 71105:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 71106:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 71107:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 71108:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 71109:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 71110:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 71111:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 71112:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 71113:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 71114:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 71115:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 71116:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 71117:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 71118:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 71119:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 71120:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 71121:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 71122:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 71123:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 71124:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 71125:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 71126:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 71127:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 71128:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 71129:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 71130:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 71131:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 71132:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 71133:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 71134:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 71135:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 71136:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 71137:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 71138:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 71139:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 71140:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 71141:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 71142:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 71143:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 71144:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 71145:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 71146:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 71147:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 71148:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 71149:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 71150:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 71151:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 71152:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 71153:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 71154:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 71155:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 71156:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 71157:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 71158:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 71159:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 71160:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 71161:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 71162:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 71163:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 71164:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 71165:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 71166:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 71167:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 71168:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 71169:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 71170:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 71171:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 71172:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 71173:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 71174:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 71175:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 71176:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 71177:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 71178:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 71179:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 71180:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 71181:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 71182:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 71183:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 71184:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 71185:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 71186:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 71187:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 71188:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 71189:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 71190:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 71191:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 71192:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 71193:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 71194:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 71195:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 71196:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 71197:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 71198:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 71199:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 71200:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 71201:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 71202:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 71203:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 71204:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 71205:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 71206:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 71207:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 71208:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 71209:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 71210:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 71211:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 71212:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 71213:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 71214:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 71215:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 71216:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 71217:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 71218:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 71219:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 71220:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 71221:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 71222:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 71223:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 71224:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 71225:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 71226:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 71227:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 71228:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 71229:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 71230:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 71231:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 71232:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 71233:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 71234:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 71235:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 71236:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 71237:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 71238:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 71239:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 71240:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 71241:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 71242:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 71243:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 71244:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 71245:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 71246:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 71247:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 71248:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 71249:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 71250:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 71251:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 71252:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 71253:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 71254:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 71255:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 71256:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 71257:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 71258:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 71259:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 71260:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 71261:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 71262:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 71263:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 71264:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 71265:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 71266:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 71267:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 71268:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 71269:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 71270:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 71271:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 71272:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 71273:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 71274:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 71275:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 71276:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 71277:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 71278:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 71279:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 71280:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 71281:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 71282:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 71283:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 71284:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 71285:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 71286:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 71287:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 71288:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 71289:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 71290:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 71291:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 71292:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 71293:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 71294:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 71295:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 71296:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 71297:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 71298:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 71299:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 71300:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 71301:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 71302:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 71303:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 71304:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 71305:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 71306:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 71307:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 71308:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 71309:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 71310:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 71311:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 71312:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 71313:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 71314:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 71315:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 71316:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 71317:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 71318:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 71319:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 71320:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 71321:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 71322:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 71323:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 71324:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 71325:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 71326:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 71327:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 71328:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 71329:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 71330:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 71331:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 71332:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 71333:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 71334:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 71335:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 71336:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 71337:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 71338:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 71339:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 71340:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 71341:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 71342:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 71343:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 71344:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 71345:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 71346:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 71347:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 71348:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 71349:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 71350:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 71351:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 71352:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 71353:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 71354:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 71355:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 71356:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 71357:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 71358:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 71359:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 71360:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 71361:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 71362:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 71363:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 71364:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 71365:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 71366:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 71367:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 71368:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 71369:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 71370:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 71371:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 71372:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 71373:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 71374:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 71375:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 71376:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 71377:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 71378:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 71379:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 71380:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 71381:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 71382:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 71383:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 71384:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 71385:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 71386:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 71387:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 71388:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 71389:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 71390:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 71391:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 71392:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 71393:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 71394:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 71395:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 71396:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 71397:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 71398:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 71399:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 71400:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 71401:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 71402:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 71403:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 71404:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 71405:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 71406:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 71407:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 71408:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 71409:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 71410:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 71411:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 71412:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 71413:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 71414:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 71415:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 71416:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 71417:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 71418:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 71419:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 71420:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 71421:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 71422:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 71423:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 71424:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 71425:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 71426:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 71427:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 71428:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 71429:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 71430:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 71431:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 71432:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 71433:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 71434:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 71435:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 71436:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 71437:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 71438:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 71439:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 71440:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 71441:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 71442:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 71443:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 71444:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 71445:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 71446:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 71447:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 71448:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 71449:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 71450:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 71451:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 71452:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 71453:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 71454:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 71455:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 71456:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 71457:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 71458:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 71459:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 71460:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 71461:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 71462:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 71463:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 71464:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 71465:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 71466:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 71467:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 71468:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 71469:22]
  assign io_z = ~x114; // @[Snxn100k.scala 71470:17]
endmodule
module SnxnLv4Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 70615:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 70616:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 70617:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 70618:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 70619:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 70620:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 70621:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 70622:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 70623:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 70624:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 70625:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 70626:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 70627:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 70628:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 70629:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 70630:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 70631:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 70632:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 70633:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 70634:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 70635:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 70636:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 70637:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 70638:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 70639:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 70640:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 70641:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 70642:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 70643:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 70644:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 70645:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 70646:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 70647:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 70648:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 70649:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 70650:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 70651:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 70652:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 70653:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 70654:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 70655:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 70656:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 70657:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 70658:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 70659:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 70660:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 70661:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 70662:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 70663:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 70664:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 70665:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 70666:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 70667:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 70668:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 70669:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 70670:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 70671:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 70672:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 70673:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 70674:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 70675:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 70676:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 70677:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 70678:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 70679:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 70680:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 70681:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 70682:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 70683:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 70684:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 70685:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 70686:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 70687:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 70688:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 70689:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 70690:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 70691:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 70692:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 70693:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 70694:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 70695:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 70696:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 70697:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 70698:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 70699:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 70700:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 70701:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 70702:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 70703:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 70704:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 70705:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 70706:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 70707:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 70708:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 70709:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 70710:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 70711:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 70712:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 70713:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 70714:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 70715:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 70716:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 70717:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 70718:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 70719:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 70720:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 70721:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 70722:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 70723:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 70724:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 70725:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 70726:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 70727:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 70728:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 70729:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 70730:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 70731:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 70732:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 70733:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 70734:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 70735:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 70736:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 70737:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 70738:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 70739:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 70740:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 70741:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 70742:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 70743:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 70744:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 70745:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 70746:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 70747:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 70748:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 70749:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 70750:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 70751:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 70752:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 70753:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 70754:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 70755:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 70756:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 70757:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 70758:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 70759:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 70760:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 70761:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 70762:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 70763:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 70764:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 70765:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 70766:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 70767:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 70768:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 70769:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 70770:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 70771:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 70772:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 70773:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 70774:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 70775:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 70776:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 70777:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 70778:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 70779:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 70780:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 70781:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 70782:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 70783:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 70784:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 70785:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 70786:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 70787:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 70788:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 70789:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 70790:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 70791:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 70792:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 70793:20]
  assign io_z = ~x44; // @[Snxn100k.scala 70794:16]
endmodule
module SnxnLv4Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 71481:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 71482:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 71483:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 71484:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 71485:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 71486:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 71487:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 71488:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 71489:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 71490:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 71491:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 71492:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 71493:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 71494:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 71495:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 71496:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 71497:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 71498:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 71499:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 71500:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 71501:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 71502:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 71503:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 71504:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 71505:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 71506:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 71507:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 71508:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 71509:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 71510:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 71511:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 71512:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 71513:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 71514:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 71515:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 71516:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 71517:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 71518:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 71519:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 71520:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 71521:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 71522:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 71523:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 71524:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 71525:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 71526:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 71527:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 71528:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 71529:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 71530:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 71531:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 71532:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 71533:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 71534:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 71535:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 71536:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 71537:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 71538:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 71539:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 71540:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 71541:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 71542:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 71543:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 71544:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 71545:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 71546:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 71547:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 71548:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 71549:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 71550:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 71551:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 71552:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 71553:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 71554:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 71555:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 71556:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 71557:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 71558:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 71559:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 71560:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 71561:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 71562:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 71563:20]
  assign io_z = ~x20; // @[Snxn100k.scala 71564:16]
endmodule
module SnxnLv4Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 70805:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 70806:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 70807:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 70808:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 70809:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 70810:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 70811:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 70812:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 70813:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 70814:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 70815:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 70816:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 70817:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 70818:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 70819:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 70820:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 70821:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 70822:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 70823:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 70824:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 70825:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 70826:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 70827:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 70828:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 70829:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 70830:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 70831:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 70832:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 70833:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 70834:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 70835:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 70836:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 70837:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 70838:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 70839:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 70840:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 70841:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 70842:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 70843:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 70844:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 70845:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 70846:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 70847:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 70848:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 70849:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 70850:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 70851:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 70852:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 70853:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 70854:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 70855:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 70856:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 70857:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 70858:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 70859:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 70860:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 70861:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 70862:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 70863:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 70864:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 70865:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 70866:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 70867:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 70868:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 70869:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 70870:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 70871:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 70872:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 70873:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 70874:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 70875:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 70876:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 70877:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 70878:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 70879:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 70880:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 70881:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 70882:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 70883:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 70884:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 70885:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 70886:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 70887:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 70888:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 70889:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 70890:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 70891:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 70892:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 70893:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 70894:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 70895:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 70896:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 70897:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 70898:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 70899:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 70900:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 70901:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 70902:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 70903:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 70904:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 70905:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 70906:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 70907:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 70908:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 70909:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 70910:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 70911:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 70912:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 70913:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 70914:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 70915:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 70916:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 70917:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 70918:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 70919:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 70920:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 70921:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 70922:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 70923:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 70924:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 70925:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 70926:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 70927:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 70928:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 70929:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 70930:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 70931:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 70932:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 70933:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 70934:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 70935:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 70936:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 70937:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 70938:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 70939:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 70940:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 70941:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 70942:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 70943:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 70944:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 70945:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 70946:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 70947:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 70948:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 70949:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 70950:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 70951:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 70952:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 70953:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 70954:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 70955:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 70956:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 70957:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 70958:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 70959:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 70960:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 70961:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 70962:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 70963:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 70964:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 70965:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 70966:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 70967:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 70968:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 70969:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 70970:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 70971:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 70972:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 70973:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 70974:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 70975:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 70976:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 70977:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 70978:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 70979:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 70980:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 70981:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 70982:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 70983:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 70984:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 70985:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 70986:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 70987:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 70988:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 70989:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 70990:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 70991:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 70992:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 70993:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 70994:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 70995:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 70996:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 70997:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 70998:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 70999:20]
  assign io_z = ~x48; // @[Snxn100k.scala 71000:16]
endmodule
module SnxnLv3Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst8_io_a; // @[Snxn100k.scala 22349:33]
  wire  inst_SnxnLv4Inst8_io_b; // @[Snxn100k.scala 22349:33]
  wire  inst_SnxnLv4Inst8_io_z; // @[Snxn100k.scala 22349:33]
  wire  inst_SnxnLv4Inst9_io_a; // @[Snxn100k.scala 22353:33]
  wire  inst_SnxnLv4Inst9_io_b; // @[Snxn100k.scala 22353:33]
  wire  inst_SnxnLv4Inst9_io_z; // @[Snxn100k.scala 22353:33]
  wire  inst_SnxnLv4Inst10_io_a; // @[Snxn100k.scala 22357:34]
  wire  inst_SnxnLv4Inst10_io_b; // @[Snxn100k.scala 22357:34]
  wire  inst_SnxnLv4Inst10_io_z; // @[Snxn100k.scala 22357:34]
  wire  inst_SnxnLv4Inst11_io_a; // @[Snxn100k.scala 22361:34]
  wire  inst_SnxnLv4Inst11_io_b; // @[Snxn100k.scala 22361:34]
  wire  inst_SnxnLv4Inst11_io_z; // @[Snxn100k.scala 22361:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst8_io_z + inst_SnxnLv4Inst9_io_z; // @[Snxn100k.scala 22365:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst10_io_z; // @[Snxn100k.scala 22365:61]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst11_io_z; // @[Snxn100k.scala 22365:87]
  SnxnLv4Inst8 inst_SnxnLv4Inst8 ( // @[Snxn100k.scala 22349:33]
    .io_a(inst_SnxnLv4Inst8_io_a),
    .io_b(inst_SnxnLv4Inst8_io_b),
    .io_z(inst_SnxnLv4Inst8_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst9 ( // @[Snxn100k.scala 22353:33]
    .io_a(inst_SnxnLv4Inst9_io_a),
    .io_b(inst_SnxnLv4Inst9_io_b),
    .io_z(inst_SnxnLv4Inst9_io_z)
  );
  SnxnLv4Inst10 inst_SnxnLv4Inst10 ( // @[Snxn100k.scala 22357:34]
    .io_a(inst_SnxnLv4Inst10_io_a),
    .io_b(inst_SnxnLv4Inst10_io_b),
    .io_z(inst_SnxnLv4Inst10_io_z)
  );
  SnxnLv4Inst11 inst_SnxnLv4Inst11 ( // @[Snxn100k.scala 22361:34]
    .io_a(inst_SnxnLv4Inst11_io_a),
    .io_b(inst_SnxnLv4Inst11_io_b),
    .io_z(inst_SnxnLv4Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22366:15]
  assign inst_SnxnLv4Inst8_io_a = io_a; // @[Snxn100k.scala 22350:26]
  assign inst_SnxnLv4Inst8_io_b = io_b; // @[Snxn100k.scala 22351:26]
  assign inst_SnxnLv4Inst9_io_a = io_a; // @[Snxn100k.scala 22354:26]
  assign inst_SnxnLv4Inst9_io_b = io_b; // @[Snxn100k.scala 22355:26]
  assign inst_SnxnLv4Inst10_io_a = io_a; // @[Snxn100k.scala 22358:27]
  assign inst_SnxnLv4Inst10_io_b = io_b; // @[Snxn100k.scala 22359:27]
  assign inst_SnxnLv4Inst11_io_a = io_a; // @[Snxn100k.scala 22362:27]
  assign inst_SnxnLv4Inst11_io_b = io_b; // @[Snxn100k.scala 22363:27]
endmodule
module SnxnLv4Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72645:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72646:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72647:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72648:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72649:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72650:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72651:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 72652:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 72653:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 72654:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 72655:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 72656:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 72657:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 72658:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 72659:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 72660:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 72661:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 72662:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 72663:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 72664:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 72665:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 72666:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 72667:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 72668:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 72669:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72670:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72671:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72672:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 72673:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 72674:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 72675:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 72676:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 72677:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 72678:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 72679:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 72680:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 72681:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 72682:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 72683:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 72684:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72685:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72686:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72687:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72688:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72689:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72690:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72691:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72692:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72693:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72694:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72695:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72696:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72697:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72698:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72699:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72700:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72701:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72702:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72703:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72704:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72705:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72706:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72707:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72708:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72709:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72710:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72711:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72712:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72713:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72714:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72715:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72716:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72717:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72718:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72719:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72720:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72721:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72722:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72723:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72724:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72725:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72726:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72727:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72728:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72729:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72730:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72731:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72732:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72733:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72734:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72735:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72736:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72737:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72738:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72739:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72740:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72741:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72742:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72743:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 72744:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 72745:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 72746:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 72747:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 72748:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 72749:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 72750:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 72751:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 72752:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 72753:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 72754:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 72755:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 72756:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 72757:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 72758:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 72759:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 72760:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 72761:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 72762:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 72763:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 72764:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 72765:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 72766:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 72767:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 72768:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 72769:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 72770:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 72771:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 72772:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 72773:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 72774:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 72775:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 72776:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 72777:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 72778:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 72779:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 72780:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 72781:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 72782:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 72783:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 72784:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 72785:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 72786:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 72787:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 72788:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 72789:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 72790:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 72791:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 72792:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 72793:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 72794:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 72795:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 72796:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 72797:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 72798:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 72799:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 72800:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 72801:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 72802:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 72803:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 72804:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 72805:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 72806:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 72807:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 72808:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 72809:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 72810:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 72811:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 72812:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 72813:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 72814:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 72815:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 72816:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 72817:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 72818:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 72819:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 72820:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 72821:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 72822:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 72823:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 72824:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 72825:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 72826:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 72827:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 72828:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 72829:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 72830:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 72831:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 72832:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 72833:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 72834:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 72835:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 72836:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 72837:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 72838:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 72839:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 72840:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 72841:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 72842:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 72843:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 72844:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 72845:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 72846:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 72847:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 72848:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 72849:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 72850:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 72851:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 72852:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 72853:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 72854:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 72855:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 72856:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 72857:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 72858:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 72859:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 72860:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 72861:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 72862:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 72863:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 72864:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 72865:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 72866:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 72867:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 72868:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 72869:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 72870:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 72871:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 72872:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 72873:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 72874:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 72875:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 72876:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 72877:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 72878:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 72879:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 72880:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 72881:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 72882:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 72883:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 72884:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 72885:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 72886:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 72887:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 72888:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 72889:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 72890:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 72891:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 72892:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 72893:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 72894:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 72895:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 72896:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 72897:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 72898:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 72899:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 72900:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 72901:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 72902:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 72903:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 72904:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 72905:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 72906:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 72907:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 72908:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 72909:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 72910:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 72911:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 72912:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 72913:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 72914:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 72915:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 72916:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 72917:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 72918:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 72919:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 72920:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 72921:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 72922:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 72923:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 72924:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 72925:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 72926:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 72927:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 72928:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 72929:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 72930:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 72931:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 72932:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 72933:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 72934:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 72935:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 72936:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 72937:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 72938:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 72939:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 72940:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 72941:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 72942:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 72943:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 72944:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 72945:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 72946:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 72947:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 72948:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 72949:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 72950:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 72951:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 72952:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 72953:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 72954:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 72955:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 72956:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 72957:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 72958:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 72959:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 72960:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 72961:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 72962:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 72963:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 72964:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 72965:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 72966:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 72967:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 72968:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 72969:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 72970:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 72971:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 72972:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 72973:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 72974:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 72975:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 72976:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 72977:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 72978:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 72979:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 72980:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 72981:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 72982:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 72983:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 72984:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 72985:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 72986:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 72987:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 72988:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 72989:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 72990:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 72991:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 72992:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 72993:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 72994:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 72995:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 72996:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 72997:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 72998:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 72999:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 73000:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 73001:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 73002:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 73003:20]
  assign io_z = ~x89; // @[Snxn100k.scala 73004:16]
endmodule
module SnxnLv4Inst13(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 72299:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 72300:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 72301:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 72302:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 72303:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 72304:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 72305:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 72306:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 72307:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 72308:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 72309:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 72310:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 72311:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 72312:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 72313:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 72314:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 72315:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 72316:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 72317:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 72318:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 72319:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 72320:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 72321:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 72322:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 72323:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 72324:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 72325:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 72326:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 72327:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 72328:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 72329:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 72330:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 72331:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 72332:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 72333:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 72334:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 72335:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 72336:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 72337:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 72338:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 72339:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 72340:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 72341:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 72342:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 72343:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 72344:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 72345:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 72346:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 72347:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 72348:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 72349:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 72350:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 72351:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 72352:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 72353:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 72354:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 72355:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 72356:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 72357:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 72358:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 72359:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 72360:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 72361:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 72362:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 72363:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 72364:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 72365:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 72366:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 72367:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 72368:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 72369:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 72370:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 72371:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 72372:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 72373:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 72374:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 72375:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 72376:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 72377:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 72378:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 72379:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 72380:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 72381:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 72382:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 72383:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 72384:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 72385:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 72386:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 72387:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 72388:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 72389:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 72390:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 72391:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 72392:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 72393:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 72394:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 72395:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 72396:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 72397:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 72398:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 72399:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 72400:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 72401:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 72402:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 72403:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 72404:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 72405:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 72406:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 72407:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 72408:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 72409:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 72410:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 72411:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 72412:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 72413:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 72414:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 72415:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 72416:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 72417:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 72418:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 72419:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 72420:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 72421:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 72422:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 72423:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 72424:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 72425:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 72426:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 72427:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 72428:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 72429:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 72430:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 72431:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 72432:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 72433:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 72434:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 72435:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 72436:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 72437:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 72438:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 72439:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 72440:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 72441:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 72442:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 72443:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 72444:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 72445:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 72446:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 72447:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 72448:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 72449:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 72450:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 72451:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 72452:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 72453:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 72454:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 72455:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 72456:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 72457:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 72458:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 72459:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 72460:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 72461:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 72462:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 72463:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 72464:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 72465:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 72466:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 72467:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 72468:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 72469:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 72470:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 72471:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 72472:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 72473:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 72474:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 72475:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 72476:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 72477:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 72478:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 72479:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 72480:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 72481:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 72482:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 72483:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 72484:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 72485:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 72486:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 72487:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 72488:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 72489:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 72490:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 72491:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 72492:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 72493:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 72494:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 72495:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 72496:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 72497:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 72498:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 72499:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 72500:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 72501:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 72502:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 72503:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 72504:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 72505:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 72506:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 72507:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 72508:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 72509:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 72510:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 72511:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 72512:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 72513:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 72514:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 72515:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 72516:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 72517:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 72518:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 72519:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 72520:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 72521:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 72522:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 72523:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 72524:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 72525:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 72526:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 72527:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 72528:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 72529:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 72530:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 72531:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 72532:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 72533:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 72534:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 72535:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 72536:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 72537:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 72538:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 72539:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 72540:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 72541:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 72542:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 72543:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 72544:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 72545:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 72546:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 72547:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 72548:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 72549:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 72550:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 72551:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 72552:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 72553:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 72554:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 72555:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 72556:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 72557:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 72558:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 72559:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 72560:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 72561:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 72562:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 72563:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 72564:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 72565:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 72566:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 72567:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 72568:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 72569:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 72570:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 72571:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 72572:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 72573:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 72574:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 72575:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 72576:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 72577:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 72578:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 72579:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 72580:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 72581:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 72582:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 72583:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 72584:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 72585:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 72586:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 72587:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 72588:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 72589:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 72590:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 72591:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 72592:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 72593:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 72594:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 72595:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 72596:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 72597:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 72598:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 72599:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 72600:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 72601:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 72602:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 72603:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 72604:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 72605:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 72606:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 72607:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 72608:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 72609:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 72610:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 72611:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 72612:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 72613:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 72614:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 72615:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 72616:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 72617:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 72618:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 72619:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 72620:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 72621:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 72622:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 72623:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 72624:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 72625:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 72626:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 72627:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 72628:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 72629:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 72630:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 72631:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 72632:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 72633:20]
  assign io_z = ~x83; // @[Snxn100k.scala 72634:16]
endmodule
module SnxnLv4Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 73015:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 73016:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 73017:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 73018:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 73019:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 73020:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 73021:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 73022:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 73023:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 73024:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 73025:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 73026:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 73027:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 73028:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 73029:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 73030:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 73031:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 73032:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 73033:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 73034:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 73035:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 73036:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 73037:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 73038:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 73039:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 73040:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 73041:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 73042:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 73043:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 73044:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 73045:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 73046:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 73047:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 73048:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 73049:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 73050:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 73051:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 73052:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 73053:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 73054:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 73055:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 73056:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 73057:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 73058:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 73059:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 73060:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 73061:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 73062:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 73063:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 73064:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 73065:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 73066:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 73067:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 73068:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 73069:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 73070:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 73071:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 73072:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 73073:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 73074:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 73075:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 73076:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 73077:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 73078:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 73079:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 73080:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 73081:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 73082:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 73083:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 73084:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 73085:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 73086:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 73087:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 73088:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 73089:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 73090:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 73091:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 73092:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 73093:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 73094:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 73095:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 73096:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 73097:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 73098:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 73099:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 73100:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 73101:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 73102:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 73103:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 73104:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 73105:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 73106:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 73107:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 73108:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 73109:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 73110:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 73111:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 73112:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 73113:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 73114:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 73115:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 73116:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 73117:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 73118:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 73119:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 73120:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 73121:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 73122:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 73123:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 73124:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 73125:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 73126:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 73127:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 73128:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 73129:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 73130:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 73131:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 73132:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 73133:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 73134:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 73135:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 73136:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 73137:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 73138:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 73139:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 73140:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 73141:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 73142:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 73143:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 73144:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 73145:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 73146:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 73147:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 73148:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 73149:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 73150:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 73151:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 73152:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 73153:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 73154:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 73155:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 73156:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 73157:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 73158:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 73159:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 73160:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 73161:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 73162:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 73163:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 73164:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 73165:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 73166:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 73167:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 73168:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 73169:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 73170:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 73171:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 73172:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 73173:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 73174:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 73175:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 73176:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 73177:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 73178:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 73179:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 73180:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 73181:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 73182:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 73183:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 73184:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 73185:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 73186:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 73187:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 73188:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 73189:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 73190:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 73191:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 73192:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 73193:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 73194:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 73195:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 73196:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 73197:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 73198:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 73199:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 73200:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 73201:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 73202:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 73203:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 73204:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 73205:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 73206:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 73207:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 73208:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 73209:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 73210:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 73211:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 73212:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 73213:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 73214:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 73215:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 73216:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 73217:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 73218:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 73219:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 73220:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 73221:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 73222:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 73223:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 73224:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 73225:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 73226:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 73227:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 73228:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 73229:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 73230:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 73231:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 73232:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 73233:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 73234:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 73235:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 73236:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 73237:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 73238:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 73239:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 73240:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 73241:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 73242:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 73243:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 73244:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 73245:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 73246:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 73247:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 73248:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 73249:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 73250:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 73251:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 73252:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 73253:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 73254:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 73255:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 73256:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 73257:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 73258:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 73259:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 73260:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 73261:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 73262:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 73263:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 73264:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 73265:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 73266:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 73267:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 73268:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 73269:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 73270:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 73271:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 73272:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 73273:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 73274:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 73275:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 73276:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 73277:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 73278:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 73279:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 73280:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 73281:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 73282:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 73283:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 73284:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 73285:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 73286:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 73287:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 73288:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 73289:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 73290:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 73291:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 73292:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 73293:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 73294:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 73295:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 73296:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 73297:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 73298:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 73299:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 73300:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 73301:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 73302:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 73303:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 73304:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 73305:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 73306:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 73307:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 73308:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 73309:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 73310:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 73311:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 73312:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 73313:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 73314:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 73315:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 73316:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 73317:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 73318:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 73319:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 73320:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 73321:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 73322:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 73323:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 73324:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 73325:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 73326:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 73327:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 73328:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 73329:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 73330:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 73331:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 73332:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 73333:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 73334:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 73335:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 73336:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 73337:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 73338:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 73339:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 73340:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 73341:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 73342:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 73343:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 73344:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 73345:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 73346:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 73347:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 73348:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 73349:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 73350:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 73351:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 73352:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 73353:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 73354:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 73355:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 73356:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 73357:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 73358:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 73359:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 73360:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 73361:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 73362:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 73363:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 73364:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 73365:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 73366:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 73367:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 73368:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 73369:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 73370:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 73371:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 73372:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 73373:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 73374:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 73375:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 73376:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 73377:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 73378:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 73379:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 73380:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 73381:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 73382:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 73383:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 73384:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 73385:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 73386:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 73387:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 73388:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 73389:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 73390:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 73391:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 73392:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 73393:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 73394:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 73395:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 73396:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 73397:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 73398:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 73399:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 73400:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 73401:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 73402:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 73403:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 73404:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 73405:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 73406:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 73407:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 73408:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 73409:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 73410:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 73411:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 73412:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 73413:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 73414:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 73415:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 73416:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 73417:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 73418:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 73419:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 73420:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 73421:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 73422:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 73423:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 73424:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 73425:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 73426:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 73427:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 73428:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 73429:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 73430:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 73431:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 73432:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 73433:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 73434:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 73435:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 73436:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 73437:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 73438:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 73439:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 73440:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 73441:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 73442:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 73443:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 73444:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 73445:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 73446:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 73447:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 73448:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 73449:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 73450:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 73451:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 73452:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 73453:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 73454:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 73455:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 73456:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 73457:22]
  assign io_z = ~x110; // @[Snxn100k.scala 73458:17]
endmodule
module SnxnLv4Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 73469:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 73470:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 73471:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 73472:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 73473:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 73474:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 73475:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 73476:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 73477:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 73478:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 73479:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 73480:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 73481:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 73482:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 73483:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 73484:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 73485:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 73486:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 73487:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 73488:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 73489:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 73490:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 73491:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 73492:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 73493:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 73494:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 73495:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 73496:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 73497:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 73498:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 73499:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 73500:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 73501:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 73502:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 73503:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 73504:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 73505:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 73506:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 73507:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 73508:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 73509:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 73510:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 73511:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 73512:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 73513:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 73514:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 73515:20]
  assign io_z = ~x11; // @[Snxn100k.scala 73516:16]
endmodule
module SnxnLv3Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst12_io_a; // @[Snxn100k.scala 22947:34]
  wire  inst_SnxnLv4Inst12_io_b; // @[Snxn100k.scala 22947:34]
  wire  inst_SnxnLv4Inst12_io_z; // @[Snxn100k.scala 22947:34]
  wire  inst_SnxnLv4Inst13_io_a; // @[Snxn100k.scala 22951:34]
  wire  inst_SnxnLv4Inst13_io_b; // @[Snxn100k.scala 22951:34]
  wire  inst_SnxnLv4Inst13_io_z; // @[Snxn100k.scala 22951:34]
  wire  inst_SnxnLv4Inst14_io_a; // @[Snxn100k.scala 22955:34]
  wire  inst_SnxnLv4Inst14_io_b; // @[Snxn100k.scala 22955:34]
  wire  inst_SnxnLv4Inst14_io_z; // @[Snxn100k.scala 22955:34]
  wire  inst_SnxnLv4Inst15_io_a; // @[Snxn100k.scala 22959:34]
  wire  inst_SnxnLv4Inst15_io_b; // @[Snxn100k.scala 22959:34]
  wire  inst_SnxnLv4Inst15_io_z; // @[Snxn100k.scala 22959:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst12_io_z + inst_SnxnLv4Inst13_io_z; // @[Snxn100k.scala 22963:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst14_io_z; // @[Snxn100k.scala 22963:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst15_io_z; // @[Snxn100k.scala 22963:89]
  SnxnLv4Inst12 inst_SnxnLv4Inst12 ( // @[Snxn100k.scala 22947:34]
    .io_a(inst_SnxnLv4Inst12_io_a),
    .io_b(inst_SnxnLv4Inst12_io_b),
    .io_z(inst_SnxnLv4Inst12_io_z)
  );
  SnxnLv4Inst13 inst_SnxnLv4Inst13 ( // @[Snxn100k.scala 22951:34]
    .io_a(inst_SnxnLv4Inst13_io_a),
    .io_b(inst_SnxnLv4Inst13_io_b),
    .io_z(inst_SnxnLv4Inst13_io_z)
  );
  SnxnLv4Inst14 inst_SnxnLv4Inst14 ( // @[Snxn100k.scala 22955:34]
    .io_a(inst_SnxnLv4Inst14_io_a),
    .io_b(inst_SnxnLv4Inst14_io_b),
    .io_z(inst_SnxnLv4Inst14_io_z)
  );
  SnxnLv4Inst15 inst_SnxnLv4Inst15 ( // @[Snxn100k.scala 22959:34]
    .io_a(inst_SnxnLv4Inst15_io_a),
    .io_b(inst_SnxnLv4Inst15_io_b),
    .io_z(inst_SnxnLv4Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 22964:15]
  assign inst_SnxnLv4Inst12_io_a = io_a; // @[Snxn100k.scala 22948:27]
  assign inst_SnxnLv4Inst12_io_b = io_b; // @[Snxn100k.scala 22949:27]
  assign inst_SnxnLv4Inst13_io_a = io_a; // @[Snxn100k.scala 22952:27]
  assign inst_SnxnLv4Inst13_io_b = io_b; // @[Snxn100k.scala 22953:27]
  assign inst_SnxnLv4Inst14_io_a = io_a; // @[Snxn100k.scala 22956:27]
  assign inst_SnxnLv4Inst14_io_b = io_b; // @[Snxn100k.scala 22957:27]
  assign inst_SnxnLv4Inst15_io_a = io_a; // @[Snxn100k.scala 22960:27]
  assign inst_SnxnLv4Inst15_io_b = io_b; // @[Snxn100k.scala 22961:27]
endmodule
module SnxnLv2Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst0_io_a; // @[Snxn100k.scala 6483:33]
  wire  inst_SnxnLv3Inst0_io_b; // @[Snxn100k.scala 6483:33]
  wire  inst_SnxnLv3Inst0_io_z; // @[Snxn100k.scala 6483:33]
  wire  inst_SnxnLv3Inst1_io_a; // @[Snxn100k.scala 6487:33]
  wire  inst_SnxnLv3Inst1_io_b; // @[Snxn100k.scala 6487:33]
  wire  inst_SnxnLv3Inst1_io_z; // @[Snxn100k.scala 6487:33]
  wire  inst_SnxnLv3Inst2_io_a; // @[Snxn100k.scala 6491:33]
  wire  inst_SnxnLv3Inst2_io_b; // @[Snxn100k.scala 6491:33]
  wire  inst_SnxnLv3Inst2_io_z; // @[Snxn100k.scala 6491:33]
  wire  inst_SnxnLv3Inst3_io_a; // @[Snxn100k.scala 6495:33]
  wire  inst_SnxnLv3Inst3_io_b; // @[Snxn100k.scala 6495:33]
  wire  inst_SnxnLv3Inst3_io_z; // @[Snxn100k.scala 6495:33]
  wire  _sum_T_1 = inst_SnxnLv3Inst0_io_z + inst_SnxnLv3Inst1_io_z; // @[Snxn100k.scala 6499:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst2_io_z; // @[Snxn100k.scala 6499:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst3_io_z; // @[Snxn100k.scala 6499:86]
  SnxnLv3Inst0 inst_SnxnLv3Inst0 ( // @[Snxn100k.scala 6483:33]
    .io_a(inst_SnxnLv3Inst0_io_a),
    .io_b(inst_SnxnLv3Inst0_io_b),
    .io_z(inst_SnxnLv3Inst0_io_z)
  );
  SnxnLv3Inst1 inst_SnxnLv3Inst1 ( // @[Snxn100k.scala 6487:33]
    .io_a(inst_SnxnLv3Inst1_io_a),
    .io_b(inst_SnxnLv3Inst1_io_b),
    .io_z(inst_SnxnLv3Inst1_io_z)
  );
  SnxnLv3Inst2 inst_SnxnLv3Inst2 ( // @[Snxn100k.scala 6491:33]
    .io_a(inst_SnxnLv3Inst2_io_a),
    .io_b(inst_SnxnLv3Inst2_io_b),
    .io_z(inst_SnxnLv3Inst2_io_z)
  );
  SnxnLv3Inst3 inst_SnxnLv3Inst3 ( // @[Snxn100k.scala 6495:33]
    .io_a(inst_SnxnLv3Inst3_io_a),
    .io_b(inst_SnxnLv3Inst3_io_b),
    .io_z(inst_SnxnLv3Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 6500:15]
  assign inst_SnxnLv3Inst0_io_a = io_a; // @[Snxn100k.scala 6484:26]
  assign inst_SnxnLv3Inst0_io_b = io_b; // @[Snxn100k.scala 6485:26]
  assign inst_SnxnLv3Inst1_io_a = io_a; // @[Snxn100k.scala 6488:26]
  assign inst_SnxnLv3Inst1_io_b = io_b; // @[Snxn100k.scala 6489:26]
  assign inst_SnxnLv3Inst2_io_a = io_a; // @[Snxn100k.scala 6492:26]
  assign inst_SnxnLv3Inst2_io_b = io_b; // @[Snxn100k.scala 6493:26]
  assign inst_SnxnLv3Inst3_io_a = io_a; // @[Snxn100k.scala 6496:26]
  assign inst_SnxnLv3Inst3_io_b = io_b; // @[Snxn100k.scala 6497:26]
endmodule
module SnxnLv4Inst16(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 79999:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 80000:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 80001:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 80002:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 80003:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 80004:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 80005:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 80006:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 80007:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 80008:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 80009:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 80010:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 80011:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 80012:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 80013:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 80014:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 80015:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 80016:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 80017:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 80018:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 80019:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 80020:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 80021:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 80022:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 80023:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 80024:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 80025:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 80026:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 80027:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 80028:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 80029:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 80030:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 80031:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 80032:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 80033:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 80034:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 80035:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 80036:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 80037:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 80038:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 80039:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 80040:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 80041:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 80042:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 80043:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 80044:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 80045:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 80046:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 80047:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 80048:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 80049:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 80050:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 80051:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 80052:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 80053:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 80054:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 80055:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 80056:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 80057:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 80058:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 80059:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 80060:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 80061:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 80062:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 80063:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 80064:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 80065:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 80066:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 80067:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 80068:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 80069:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 80070:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 80071:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 80072:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 80073:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 80074:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 80075:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 80076:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 80077:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 80078:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 80079:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 80080:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 80081:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 80082:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 80083:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 80084:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 80085:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 80086:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 80087:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 80088:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 80089:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 80090:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 80091:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 80092:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 80093:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 80094:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 80095:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 80096:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 80097:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 80098:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 80099:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 80100:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 80101:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 80102:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 80103:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 80104:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 80105:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 80106:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 80107:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 80108:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 80109:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 80110:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 80111:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 80112:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 80113:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 80114:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 80115:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 80116:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 80117:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 80118:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 80119:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 80120:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 80121:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 80122:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 80123:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 80124:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 80125:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 80126:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 80127:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 80128:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 80129:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 80130:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 80131:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 80132:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 80133:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 80134:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 80135:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 80136:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 80137:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 80138:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 80139:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 80140:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 80141:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 80142:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 80143:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 80144:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 80145:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 80146:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 80147:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 80148:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 80149:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 80150:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 80151:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 80152:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 80153:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 80154:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 80155:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 80156:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 80157:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 80158:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 80159:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 80160:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 80161:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 80162:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 80163:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 80164:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 80165:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 80166:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 80167:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 80168:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 80169:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 80170:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 80171:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 80172:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 80173:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 80174:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 80175:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 80176:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 80177:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 80178:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 80179:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 80180:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 80181:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 80182:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 80183:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 80184:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 80185:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 80186:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 80187:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 80188:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 80189:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 80190:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 80191:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 80192:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 80193:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 80194:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 80195:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 80196:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 80197:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 80198:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 80199:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 80200:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 80201:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 80202:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 80203:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 80204:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 80205:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 80206:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 80207:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 80208:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 80209:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 80210:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 80211:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 80212:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 80213:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 80214:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 80215:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 80216:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 80217:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 80218:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 80219:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 80220:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 80221:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 80222:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 80223:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 80224:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 80225:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 80226:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 80227:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 80228:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 80229:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 80230:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 80231:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 80232:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 80233:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 80234:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 80235:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 80236:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 80237:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 80238:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 80239:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 80240:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 80241:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 80242:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 80243:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 80244:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 80245:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 80246:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 80247:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 80248:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 80249:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 80250:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 80251:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 80252:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 80253:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 80254:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 80255:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 80256:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 80257:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 80258:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 80259:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 80260:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 80261:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 80262:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 80263:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 80264:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 80265:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 80266:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 80267:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 80268:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 80269:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 80270:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 80271:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 80272:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 80273:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 80274:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 80275:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 80276:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 80277:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 80278:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 80279:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 80280:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 80281:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 80282:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 80283:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 80284:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 80285:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 80286:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 80287:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 80288:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 80289:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 80290:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 80291:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 80292:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 80293:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 80294:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 80295:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 80296:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 80297:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 80298:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 80299:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 80300:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 80301:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 80302:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 80303:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 80304:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 80305:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 80306:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 80307:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 80308:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 80309:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 80310:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 80311:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 80312:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 80313:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 80314:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 80315:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 80316:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 80317:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 80318:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 80319:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 80320:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 80321:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 80322:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 80323:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 80324:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 80325:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 80326:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 80327:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 80328:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 80329:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 80330:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 80331:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 80332:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 80333:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 80334:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 80335:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 80336:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 80337:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 80338:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 80339:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 80340:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 80341:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 80342:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 80343:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 80344:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 80345:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 80346:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 80347:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 80348:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 80349:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 80350:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 80351:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 80352:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 80353:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 80354:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 80355:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 80356:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 80357:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 80358:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 80359:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 80360:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 80361:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 80362:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 80363:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 80364:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 80365:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 80366:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 80367:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 80368:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 80369:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 80370:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 80371:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 80372:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 80373:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 80374:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 80375:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 80376:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 80377:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 80378:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 80379:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 80380:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 80381:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 80382:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 80383:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 80384:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 80385:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 80386:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 80387:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 80388:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 80389:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 80390:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 80391:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 80392:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 80393:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 80394:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 80395:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 80396:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 80397:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 80398:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 80399:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 80400:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 80401:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 80402:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 80403:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 80404:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 80405:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 80406:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 80407:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 80408:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 80409:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 80410:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 80411:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 80412:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 80413:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 80414:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 80415:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 80416:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 80417:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 80418:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 80419:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 80420:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 80421:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 80422:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 80423:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 80424:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 80425:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 80426:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 80427:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 80428:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 80429:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 80430:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 80431:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 80432:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 80433:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 80434:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 80435:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 80436:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 80437:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 80438:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 80439:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 80440:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 80441:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 80442:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 80443:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 80444:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 80445:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 80446:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 80447:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 80448:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 80449:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 80450:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 80451:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 80452:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 80453:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 80454:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 80455:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 80456:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 80457:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 80458:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 80459:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 80460:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 80461:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 80462:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 80463:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 80464:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 80465:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 80466:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 80467:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 80468:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 80469:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 80470:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 80471:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 80472:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 80473:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 80474:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 80475:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 80476:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 80477:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 80478:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 80479:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 80480:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 80481:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 80482:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 80483:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 80484:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 80485:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 80486:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 80487:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 80488:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 80489:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 80490:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 80491:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 80492:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 80493:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 80494:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 80495:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 80496:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 80497:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 80498:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 80499:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 80500:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 80501:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 80502:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 80503:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 80504:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 80505:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 80506:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 80507:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 80508:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 80509:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 80510:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 80511:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 80512:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 80513:22]
  assign io_z = ~x128; // @[Snxn100k.scala 80514:17]
endmodule
module SnxnLv4Inst17(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 79481:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 79482:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 79483:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 79484:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 79485:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 79486:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 79487:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 79488:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 79489:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 79490:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 79491:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 79492:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 79493:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 79494:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 79495:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 79496:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 79497:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 79498:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 79499:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 79500:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 79501:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 79502:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 79503:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 79504:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 79505:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 79506:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 79507:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 79508:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 79509:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 79510:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 79511:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 79512:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 79513:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 79514:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 79515:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 79516:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 79517:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 79518:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 79519:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 79520:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 79521:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 79522:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 79523:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 79524:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 79525:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 79526:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 79527:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 79528:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 79529:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 79530:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 79531:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 79532:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 79533:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 79534:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 79535:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 79536:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 79537:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 79538:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 79539:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 79540:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 79541:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 79542:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 79543:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 79544:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 79545:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 79546:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 79547:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 79548:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 79549:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 79550:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 79551:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 79552:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 79553:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 79554:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 79555:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 79556:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 79557:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 79558:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 79559:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 79560:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 79561:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 79562:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 79563:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 79564:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 79565:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 79566:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 79567:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 79568:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 79569:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 79570:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 79571:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 79572:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 79573:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 79574:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 79575:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 79576:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 79577:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 79578:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 79579:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 79580:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 79581:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 79582:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 79583:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 79584:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 79585:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 79586:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 79587:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 79588:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 79589:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 79590:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 79591:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 79592:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 79593:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 79594:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 79595:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 79596:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 79597:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 79598:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 79599:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 79600:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 79601:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 79602:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 79603:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 79604:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 79605:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 79606:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 79607:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79608:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79609:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79610:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79611:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79612:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79613:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79614:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79615:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79616:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79617:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79618:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79619:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79620:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79621:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79622:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79623:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79624:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79625:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79626:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79627:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79628:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79629:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79630:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79631:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79632:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79633:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79634:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79635:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79636:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79637:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79638:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79639:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79640:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79641:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79642:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79643:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79644:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79645:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79646:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79647:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79648:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79649:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79650:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79651:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79652:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79653:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79654:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79655:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79656:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79657:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79658:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79659:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79660:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79661:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79662:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79663:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79664:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79665:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79666:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79667:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79668:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79669:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79670:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79671:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79672:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79673:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79674:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79675:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79676:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79677:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79678:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79679:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 79680:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 79681:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 79682:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 79683:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 79684:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 79685:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 79686:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 79687:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 79688:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 79689:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 79690:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 79691:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 79692:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 79693:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 79694:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 79695:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 79696:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 79697:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 79698:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 79699:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 79700:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 79701:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 79702:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 79703:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 79704:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 79705:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 79706:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 79707:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 79708:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 79709:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 79710:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 79711:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 79712:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 79713:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 79714:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 79715:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 79716:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 79717:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 79718:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 79719:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 79720:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 79721:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 79722:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 79723:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 79724:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 79725:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 79726:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 79727:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 79728:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 79729:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 79730:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 79731:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 79732:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 79733:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 79734:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 79735:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 79736:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 79737:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 79738:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 79739:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 79740:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 79741:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 79742:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 79743:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 79744:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 79745:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 79746:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 79747:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 79748:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 79749:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 79750:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 79751:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 79752:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 79753:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 79754:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 79755:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 79756:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 79757:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 79758:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 79759:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 79760:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 79761:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 79762:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 79763:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 79764:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 79765:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 79766:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 79767:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 79768:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 79769:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 79770:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 79771:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 79772:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 79773:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 79774:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 79775:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 79776:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 79777:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 79778:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 79779:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 79780:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 79781:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 79782:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 79783:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 79784:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 79785:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 79786:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 79787:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 79788:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 79789:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 79790:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 79791:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 79792:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 79793:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 79794:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 79795:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 79796:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 79797:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 79798:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 79799:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 79800:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 79801:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 79802:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 79803:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 79804:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 79805:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 79806:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 79807:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 79808:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 79809:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 79810:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 79811:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 79812:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 79813:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 79814:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 79815:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 79816:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 79817:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 79818:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 79819:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 79820:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 79821:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 79822:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 79823:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 79824:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 79825:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 79826:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 79827:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 79828:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 79829:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 79830:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 79831:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 79832:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 79833:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 79834:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 79835:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 79836:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 79837:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 79838:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 79839:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 79840:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 79841:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 79842:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 79843:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 79844:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 79845:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 79846:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 79847:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 79848:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 79849:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 79850:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 79851:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 79852:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 79853:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 79854:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 79855:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 79856:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 79857:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 79858:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 79859:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 79860:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 79861:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 79862:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 79863:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 79864:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 79865:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 79866:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 79867:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 79868:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 79869:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 79870:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 79871:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 79872:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 79873:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 79874:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 79875:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 79876:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 79877:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 79878:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 79879:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 79880:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 79881:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 79882:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 79883:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 79884:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 79885:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 79886:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 79887:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 79888:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 79889:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 79890:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 79891:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 79892:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 79893:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 79894:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 79895:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 79896:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 79897:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 79898:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 79899:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 79900:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 79901:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 79902:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 79903:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 79904:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 79905:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 79906:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 79907:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 79908:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 79909:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 79910:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 79911:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 79912:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 79913:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 79914:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 79915:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 79916:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 79917:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 79918:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 79919:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 79920:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 79921:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 79922:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 79923:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 79924:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 79925:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 79926:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 79927:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 79928:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 79929:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 79930:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 79931:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 79932:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 79933:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 79934:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 79935:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 79936:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 79937:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 79938:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 79939:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 79940:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 79941:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 79942:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 79943:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 79944:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 79945:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 79946:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 79947:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 79948:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 79949:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 79950:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 79951:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 79952:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 79953:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 79954:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 79955:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 79956:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 79957:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 79958:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 79959:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 79960:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 79961:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 79962:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 79963:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 79964:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 79965:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 79966:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 79967:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 79968:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 79969:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 79970:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 79971:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 79972:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 79973:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 79974:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 79975:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 79976:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 79977:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 79978:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 79979:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 79980:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 79981:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 79982:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 79983:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 79984:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 79985:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 79986:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 79987:22]
  assign io_z = ~x126; // @[Snxn100k.scala 79988:17]
endmodule
module SnxnLv4Inst18(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 80525:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 80526:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 80527:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 80528:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 80529:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 80530:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 80531:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 80532:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 80533:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 80534:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 80535:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 80536:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 80537:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 80538:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 80539:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 80540:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 80541:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 80542:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 80543:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 80544:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 80545:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 80546:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 80547:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 80548:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 80549:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 80550:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 80551:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 80552:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 80553:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 80554:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 80555:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 80556:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 80557:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 80558:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 80559:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 80560:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 80561:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 80562:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 80563:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 80564:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 80565:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 80566:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 80567:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 80568:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 80569:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 80570:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 80571:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 80572:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 80573:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 80574:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 80575:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 80576:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 80577:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 80578:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 80579:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 80580:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 80581:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 80582:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 80583:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 80584:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 80585:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 80586:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 80587:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 80588:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 80589:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 80590:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 80591:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 80592:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 80593:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 80594:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 80595:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 80596:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 80597:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 80598:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 80599:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 80600:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 80601:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 80602:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 80603:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 80604:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 80605:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 80606:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 80607:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 80608:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 80609:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 80610:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 80611:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 80612:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 80613:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 80614:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 80615:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 80616:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 80617:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 80618:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 80619:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 80620:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 80621:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 80622:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 80623:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 80624:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 80625:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 80626:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 80627:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 80628:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 80629:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 80630:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 80631:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 80632:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 80633:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 80634:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 80635:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 80636:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 80637:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 80638:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 80639:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 80640:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 80641:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 80642:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 80643:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 80644:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 80645:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 80646:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 80647:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 80648:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 80649:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 80650:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 80651:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 80652:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 80653:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 80654:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 80655:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 80656:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 80657:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 80658:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 80659:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 80660:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 80661:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 80662:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 80663:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 80664:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 80665:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 80666:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 80667:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 80668:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 80669:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 80670:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 80671:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 80672:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 80673:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 80674:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 80675:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 80676:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 80677:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 80678:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 80679:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 80680:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 80681:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 80682:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 80683:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 80684:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 80685:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 80686:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 80687:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 80688:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 80689:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 80690:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 80691:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 80692:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 80693:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 80694:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 80695:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 80696:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 80697:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 80698:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 80699:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 80700:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 80701:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 80702:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 80703:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 80704:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 80705:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 80706:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 80707:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 80708:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 80709:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 80710:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 80711:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 80712:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 80713:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 80714:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 80715:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 80716:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 80717:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 80718:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 80719:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 80720:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 80721:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 80722:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 80723:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 80724:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 80725:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 80726:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 80727:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 80728:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 80729:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 80730:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 80731:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 80732:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 80733:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 80734:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 80735:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 80736:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 80737:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 80738:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 80739:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 80740:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 80741:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 80742:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 80743:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 80744:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 80745:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 80746:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 80747:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 80748:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 80749:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 80750:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 80751:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 80752:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 80753:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 80754:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 80755:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 80756:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 80757:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 80758:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 80759:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 80760:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 80761:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 80762:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 80763:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 80764:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 80765:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 80766:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 80767:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 80768:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 80769:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 80770:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 80771:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 80772:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 80773:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 80774:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 80775:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 80776:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 80777:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 80778:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 80779:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 80780:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 80781:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 80782:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 80783:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 80784:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 80785:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 80786:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 80787:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 80788:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 80789:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 80790:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 80791:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 80792:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 80793:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 80794:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 80795:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 80796:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 80797:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 80798:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 80799:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 80800:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 80801:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 80802:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 80803:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 80804:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 80805:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 80806:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 80807:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 80808:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 80809:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 80810:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 80811:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 80812:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 80813:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 80814:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 80815:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 80816:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 80817:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 80818:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 80819:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 80820:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 80821:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 80822:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 80823:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 80824:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 80825:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 80826:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 80827:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 80828:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 80829:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 80830:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 80831:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 80832:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 80833:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 80834:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 80835:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 80836:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 80837:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 80838:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 80839:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 80840:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 80841:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 80842:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 80843:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 80844:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 80845:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 80846:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 80847:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 80848:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 80849:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 80850:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 80851:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 80852:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 80853:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 80854:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 80855:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 80856:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 80857:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 80858:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 80859:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 80860:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 80861:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 80862:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 80863:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 80864:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 80865:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 80866:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 80867:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 80868:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 80869:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 80870:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 80871:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 80872:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 80873:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 80874:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 80875:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 80876:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 80877:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 80878:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 80879:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 80880:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 80881:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 80882:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 80883:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 80884:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 80885:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 80886:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 80887:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 80888:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 80889:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 80890:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 80891:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 80892:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 80893:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 80894:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 80895:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 80896:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 80897:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 80898:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 80899:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 80900:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 80901:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 80902:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 80903:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 80904:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 80905:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 80906:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 80907:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 80908:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 80909:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 80910:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 80911:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 80912:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 80913:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 80914:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 80915:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 80916:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 80917:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 80918:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 80919:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 80920:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 80921:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 80922:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 80923:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 80924:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 80925:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 80926:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 80927:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 80928:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 80929:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 80930:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 80931:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 80932:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 80933:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 80934:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 80935:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 80936:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 80937:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 80938:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 80939:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 80940:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 80941:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 80942:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 80943:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 80944:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 80945:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 80946:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 80947:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 80948:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 80949:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 80950:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 80951:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 80952:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 80953:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 80954:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 80955:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 80956:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 80957:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 80958:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 80959:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 80960:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 80961:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 80962:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 80963:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 80964:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 80965:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 80966:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 80967:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 80968:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 80969:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 80970:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 80971:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 80972:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 80973:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 80974:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 80975:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 80976:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 80977:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 80978:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 80979:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 80980:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 80981:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 80982:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 80983:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 80984:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 80985:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 80986:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 80987:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 80988:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 80989:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 80990:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 80991:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 80992:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 80993:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 80994:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 80995:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 80996:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 80997:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 80998:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 80999:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 81000:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 81001:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 81002:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 81003:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 81004:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 81005:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 81006:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 81007:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 81008:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 81009:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 81010:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 81011:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 81012:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 81013:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 81014:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 81015:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 81016:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 81017:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 81018:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 81019:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 81020:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 81021:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 81022:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 81023:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 81024:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 81025:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 81026:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 81027:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 81028:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 81029:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 81030:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 81031:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 81032:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 81033:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 81034:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 81035:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 81036:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 81037:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 81038:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 81039:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 81040:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 81041:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 81042:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 81043:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 81044:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 81045:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 81046:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 81047:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 81048:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 81049:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 81050:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 81051:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 81052:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 81053:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 81054:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 81055:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 81056:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 81057:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 81058:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 81059:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 81060:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 81061:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 81062:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 81063:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 81064:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 81065:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 81066:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 81067:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 81068:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 81069:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 81070:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 81071:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 81072:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 81073:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 81074:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 81075:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 81076:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 81077:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 81078:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 81079:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 81080:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 81081:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 81082:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 81083:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 81084:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 81085:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 81086:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 81087:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 81088:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 81089:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 81090:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 81091:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 81092:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 81093:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 81094:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 81095:22]
  wire  invx142 = ~x142; // @[Snxn100k.scala 81096:17]
  wire  t143 = x142 + invx142; // @[Snxn100k.scala 81097:22]
  wire  inv143 = ~t143; // @[Snxn100k.scala 81098:17]
  wire  x143 = t143 ^ inv143; // @[Snxn100k.scala 81099:22]
  wire  invx143 = ~x143; // @[Snxn100k.scala 81100:17]
  wire  t144 = x143 + invx143; // @[Snxn100k.scala 81101:22]
  wire  inv144 = ~t144; // @[Snxn100k.scala 81102:17]
  wire  x144 = t144 ^ inv144; // @[Snxn100k.scala 81103:22]
  wire  invx144 = ~x144; // @[Snxn100k.scala 81104:17]
  wire  t145 = x144 + invx144; // @[Snxn100k.scala 81105:22]
  wire  inv145 = ~t145; // @[Snxn100k.scala 81106:17]
  wire  x145 = t145 ^ inv145; // @[Snxn100k.scala 81107:22]
  wire  invx145 = ~x145; // @[Snxn100k.scala 81108:17]
  wire  t146 = x145 + invx145; // @[Snxn100k.scala 81109:22]
  wire  inv146 = ~t146; // @[Snxn100k.scala 81110:17]
  wire  x146 = t146 ^ inv146; // @[Snxn100k.scala 81111:22]
  assign io_z = ~x146; // @[Snxn100k.scala 81112:17]
endmodule
module SnxnLv4Inst19(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 79271:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 79272:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 79273:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 79274:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 79275:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 79276:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 79277:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 79278:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 79279:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 79280:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 79281:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 79282:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 79283:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 79284:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 79285:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 79286:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 79287:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 79288:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 79289:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 79290:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 79291:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 79292:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 79293:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 79294:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 79295:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 79296:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 79297:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 79298:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 79299:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 79300:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 79301:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 79302:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 79303:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 79304:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 79305:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 79306:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 79307:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 79308:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 79309:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 79310:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 79311:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 79312:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 79313:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 79314:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 79315:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 79316:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 79317:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 79318:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 79319:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 79320:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 79321:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 79322:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 79323:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 79324:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 79325:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 79326:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 79327:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 79328:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 79329:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 79330:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 79331:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 79332:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 79333:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 79334:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 79335:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 79336:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 79337:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 79338:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 79339:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 79340:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 79341:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 79342:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 79343:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 79344:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 79345:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 79346:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 79347:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 79348:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 79349:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 79350:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 79351:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 79352:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 79353:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 79354:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 79355:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 79356:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 79357:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 79358:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 79359:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 79360:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 79361:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 79362:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 79363:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 79364:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 79365:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 79366:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 79367:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 79368:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 79369:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 79370:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 79371:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 79372:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 79373:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 79374:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 79375:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 79376:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 79377:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 79378:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 79379:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 79380:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 79381:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 79382:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 79383:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 79384:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 79385:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 79386:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 79387:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 79388:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 79389:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 79390:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 79391:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 79392:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 79393:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 79394:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 79395:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 79396:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 79397:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79398:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79399:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79400:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79401:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79402:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79403:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79404:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79405:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79406:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79407:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79408:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79409:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79410:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79411:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79412:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79413:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79414:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79415:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79416:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79417:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79418:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79419:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79420:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79421:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79422:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79423:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79424:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79425:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79426:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79427:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79428:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79429:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79430:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79431:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79432:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79433:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79434:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79435:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79436:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79437:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79438:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79439:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79440:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79441:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79442:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79443:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79444:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79445:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79446:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79447:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79448:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79449:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79450:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79451:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79452:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79453:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79454:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79455:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79456:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79457:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79458:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79459:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79460:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79461:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79462:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79463:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79464:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79465:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79466:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79467:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79468:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79469:20]
  assign io_z = ~x49; // @[Snxn100k.scala 79470:16]
endmodule
module SnxnLv3Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst16_io_a; // @[Snxn100k.scala 24189:34]
  wire  inst_SnxnLv4Inst16_io_b; // @[Snxn100k.scala 24189:34]
  wire  inst_SnxnLv4Inst16_io_z; // @[Snxn100k.scala 24189:34]
  wire  inst_SnxnLv4Inst17_io_a; // @[Snxn100k.scala 24193:34]
  wire  inst_SnxnLv4Inst17_io_b; // @[Snxn100k.scala 24193:34]
  wire  inst_SnxnLv4Inst17_io_z; // @[Snxn100k.scala 24193:34]
  wire  inst_SnxnLv4Inst18_io_a; // @[Snxn100k.scala 24197:34]
  wire  inst_SnxnLv4Inst18_io_b; // @[Snxn100k.scala 24197:34]
  wire  inst_SnxnLv4Inst18_io_z; // @[Snxn100k.scala 24197:34]
  wire  inst_SnxnLv4Inst19_io_a; // @[Snxn100k.scala 24201:34]
  wire  inst_SnxnLv4Inst19_io_b; // @[Snxn100k.scala 24201:34]
  wire  inst_SnxnLv4Inst19_io_z; // @[Snxn100k.scala 24201:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst16_io_z + inst_SnxnLv4Inst17_io_z; // @[Snxn100k.scala 24205:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst18_io_z; // @[Snxn100k.scala 24205:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst19_io_z; // @[Snxn100k.scala 24205:89]
  SnxnLv4Inst16 inst_SnxnLv4Inst16 ( // @[Snxn100k.scala 24189:34]
    .io_a(inst_SnxnLv4Inst16_io_a),
    .io_b(inst_SnxnLv4Inst16_io_b),
    .io_z(inst_SnxnLv4Inst16_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst17 ( // @[Snxn100k.scala 24193:34]
    .io_a(inst_SnxnLv4Inst17_io_a),
    .io_b(inst_SnxnLv4Inst17_io_b),
    .io_z(inst_SnxnLv4Inst17_io_z)
  );
  SnxnLv4Inst18 inst_SnxnLv4Inst18 ( // @[Snxn100k.scala 24197:34]
    .io_a(inst_SnxnLv4Inst18_io_a),
    .io_b(inst_SnxnLv4Inst18_io_b),
    .io_z(inst_SnxnLv4Inst18_io_z)
  );
  SnxnLv4Inst19 inst_SnxnLv4Inst19 ( // @[Snxn100k.scala 24201:34]
    .io_a(inst_SnxnLv4Inst19_io_a),
    .io_b(inst_SnxnLv4Inst19_io_b),
    .io_z(inst_SnxnLv4Inst19_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 24206:15]
  assign inst_SnxnLv4Inst16_io_a = io_a; // @[Snxn100k.scala 24190:27]
  assign inst_SnxnLv4Inst16_io_b = io_b; // @[Snxn100k.scala 24191:27]
  assign inst_SnxnLv4Inst17_io_a = io_a; // @[Snxn100k.scala 24194:27]
  assign inst_SnxnLv4Inst17_io_b = io_b; // @[Snxn100k.scala 24195:27]
  assign inst_SnxnLv4Inst18_io_a = io_a; // @[Snxn100k.scala 24198:27]
  assign inst_SnxnLv4Inst18_io_b = io_b; // @[Snxn100k.scala 24199:27]
  assign inst_SnxnLv4Inst19_io_a = io_a; // @[Snxn100k.scala 24202:27]
  assign inst_SnxnLv4Inst19_io_b = io_b; // @[Snxn100k.scala 24203:27]
endmodule
module SnxnLv4Inst21(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78419:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78420:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78421:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78422:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78423:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78424:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78425:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78426:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78427:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78428:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78429:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78430:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78431:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78432:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78433:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78434:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78435:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78436:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78437:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78438:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78439:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78440:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78441:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78442:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78443:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78444:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78445:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78446:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78447:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78448:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78449:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78450:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78451:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78452:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78453:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78454:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78455:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78456:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78457:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78458:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78459:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78460:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78461:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78462:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78463:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78464:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78465:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78466:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78467:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78468:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78469:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78470:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78471:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78472:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78473:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78474:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78475:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78476:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78477:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78478:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78479:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78480:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78481:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78482:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78483:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78484:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78485:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78486:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78487:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78488:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78489:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 78490:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 78491:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 78492:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 78493:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 78494:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 78495:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 78496:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 78497:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 78498:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 78499:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 78500:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 78501:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 78502:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 78503:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 78504:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 78505:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 78506:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 78507:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 78508:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 78509:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 78510:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 78511:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 78512:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 78513:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 78514:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 78515:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 78516:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 78517:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 78518:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 78519:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 78520:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 78521:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 78522:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 78523:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 78524:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 78525:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 78526:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 78527:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 78528:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 78529:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 78530:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 78531:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 78532:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 78533:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 78534:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 78535:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 78536:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 78537:20]
  assign io_z = ~x29; // @[Snxn100k.scala 78538:16]
endmodule
module SnxnLv4Inst22(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78873:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78874:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78875:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78876:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78877:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78878:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78879:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78880:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78881:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78882:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78883:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78884:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78885:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78886:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78887:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78888:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78889:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78890:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78891:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78892:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78893:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78894:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78895:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78896:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78897:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78898:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78899:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78900:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78901:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78902:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78903:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78904:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78905:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78906:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78907:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78908:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78909:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78910:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78911:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78912:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78913:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78914:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78915:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78916:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78917:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78918:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78919:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78920:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78921:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78922:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78923:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78924:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78925:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78926:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78927:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78928:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78929:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78930:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78931:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78932:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78933:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78934:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78935:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78936:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78937:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78938:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78939:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78940:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78941:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78942:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78943:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 78944:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 78945:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 78946:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 78947:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 78948:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 78949:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 78950:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 78951:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 78952:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 78953:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 78954:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 78955:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 78956:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 78957:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 78958:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 78959:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 78960:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 78961:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 78962:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 78963:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 78964:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 78965:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 78966:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 78967:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 78968:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 78969:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 78970:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 78971:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 78972:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 78973:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 78974:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 78975:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 78976:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 78977:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 78978:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 78979:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 78980:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 78981:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 78982:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 78983:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 78984:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 78985:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 78986:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 78987:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 78988:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 78989:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 78990:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 78991:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 78992:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 78993:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 78994:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 78995:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 78996:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 78997:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 78998:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 78999:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 79000:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 79001:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 79002:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 79003:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 79004:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 79005:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 79006:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 79007:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 79008:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 79009:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 79010:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 79011:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 79012:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 79013:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 79014:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 79015:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 79016:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 79017:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 79018:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 79019:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 79020:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 79021:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 79022:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 79023:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 79024:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 79025:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 79026:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 79027:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 79028:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 79029:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 79030:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 79031:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 79032:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 79033:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 79034:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 79035:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 79036:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 79037:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 79038:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 79039:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 79040:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 79041:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 79042:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 79043:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 79044:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 79045:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 79046:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 79047:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 79048:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 79049:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 79050:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 79051:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 79052:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 79053:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 79054:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 79055:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 79056:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 79057:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 79058:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 79059:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 79060:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 79061:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 79062:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 79063:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 79064:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 79065:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 79066:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 79067:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 79068:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 79069:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 79070:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 79071:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 79072:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 79073:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 79074:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 79075:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 79076:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 79077:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 79078:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 79079:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 79080:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 79081:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 79082:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 79083:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 79084:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 79085:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 79086:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 79087:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 79088:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 79089:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 79090:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 79091:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 79092:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 79093:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 79094:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 79095:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 79096:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 79097:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 79098:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 79099:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 79100:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 79101:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 79102:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 79103:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 79104:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 79105:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 79106:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 79107:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 79108:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 79109:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 79110:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 79111:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 79112:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 79113:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 79114:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 79115:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 79116:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 79117:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 79118:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 79119:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 79120:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 79121:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 79122:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 79123:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 79124:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 79125:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 79126:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 79127:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 79128:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 79129:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 79130:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 79131:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 79132:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 79133:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 79134:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 79135:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 79136:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 79137:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 79138:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 79139:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 79140:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 79141:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 79142:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 79143:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 79144:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 79145:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 79146:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 79147:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 79148:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 79149:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 79150:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 79151:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 79152:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 79153:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 79154:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 79155:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 79156:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 79157:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 79158:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 79159:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 79160:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 79161:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 79162:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 79163:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 79164:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 79165:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 79166:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 79167:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 79168:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 79169:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 79170:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 79171:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 79172:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 79173:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 79174:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 79175:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 79176:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 79177:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 79178:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 79179:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 79180:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 79181:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 79182:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 79183:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 79184:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 79185:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 79186:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 79187:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 79188:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 79189:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 79190:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 79191:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 79192:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 79193:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 79194:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 79195:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 79196:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 79197:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 79198:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 79199:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 79200:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 79201:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 79202:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 79203:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 79204:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 79205:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 79206:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 79207:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 79208:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 79209:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 79210:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 79211:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 79212:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 79213:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 79214:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 79215:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 79216:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 79217:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 79218:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 79219:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 79220:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 79221:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 79222:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 79223:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 79224:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 79225:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 79226:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 79227:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 79228:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 79229:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 79230:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 79231:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 79232:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 79233:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 79234:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 79235:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 79236:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 79237:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 79238:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 79239:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 79240:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 79241:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 79242:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 79243:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 79244:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 79245:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 79246:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 79247:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 79248:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 79249:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 79250:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 79251:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 79252:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 79253:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 79254:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 79255:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 79256:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 79257:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 79258:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 79259:20]
  assign io_z = ~x96; // @[Snxn100k.scala 79260:16]
endmodule
module SnxnLv4Inst23(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78549:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78550:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78551:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78552:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78553:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78554:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78555:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78556:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78557:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78558:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78559:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78560:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78561:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78562:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78563:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78564:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78565:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78566:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78567:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78568:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78569:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78570:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78571:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78572:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78573:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78574:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78575:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78576:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78577:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78578:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78579:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78580:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78581:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78582:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78583:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78584:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78585:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78586:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78587:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78588:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78589:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78590:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78591:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78592:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78593:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78594:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78595:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78596:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78597:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78598:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78599:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78600:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78601:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78602:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78603:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78604:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78605:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78606:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78607:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78608:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78609:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78610:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78611:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78612:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78613:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78614:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78615:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78616:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78617:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78618:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78619:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 78620:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 78621:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 78622:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 78623:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 78624:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 78625:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 78626:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 78627:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 78628:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 78629:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 78630:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 78631:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 78632:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 78633:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 78634:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 78635:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 78636:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 78637:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 78638:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 78639:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 78640:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 78641:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 78642:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 78643:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 78644:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 78645:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 78646:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 78647:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 78648:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 78649:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 78650:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 78651:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 78652:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 78653:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 78654:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 78655:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 78656:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 78657:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 78658:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 78659:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 78660:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 78661:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 78662:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 78663:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 78664:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 78665:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 78666:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 78667:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 78668:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 78669:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 78670:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 78671:20]
  assign io_z = ~x30; // @[Snxn100k.scala 78672:16]
endmodule
module SnxnLv3Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst20_io_a; // @[Snxn100k.scala 24046:34]
  wire  inst_SnxnLv4Inst20_io_b; // @[Snxn100k.scala 24046:34]
  wire  inst_SnxnLv4Inst20_io_z; // @[Snxn100k.scala 24046:34]
  wire  inst_SnxnLv4Inst21_io_a; // @[Snxn100k.scala 24050:34]
  wire  inst_SnxnLv4Inst21_io_b; // @[Snxn100k.scala 24050:34]
  wire  inst_SnxnLv4Inst21_io_z; // @[Snxn100k.scala 24050:34]
  wire  inst_SnxnLv4Inst22_io_a; // @[Snxn100k.scala 24054:34]
  wire  inst_SnxnLv4Inst22_io_b; // @[Snxn100k.scala 24054:34]
  wire  inst_SnxnLv4Inst22_io_z; // @[Snxn100k.scala 24054:34]
  wire  inst_SnxnLv4Inst23_io_a; // @[Snxn100k.scala 24058:34]
  wire  inst_SnxnLv4Inst23_io_b; // @[Snxn100k.scala 24058:34]
  wire  inst_SnxnLv4Inst23_io_z; // @[Snxn100k.scala 24058:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst20_io_z + inst_SnxnLv4Inst21_io_z; // @[Snxn100k.scala 24062:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst22_io_z; // @[Snxn100k.scala 24062:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst23_io_z; // @[Snxn100k.scala 24062:89]
  SnxnLv4Inst9 inst_SnxnLv4Inst20 ( // @[Snxn100k.scala 24046:34]
    .io_a(inst_SnxnLv4Inst20_io_a),
    .io_b(inst_SnxnLv4Inst20_io_b),
    .io_z(inst_SnxnLv4Inst20_io_z)
  );
  SnxnLv4Inst21 inst_SnxnLv4Inst21 ( // @[Snxn100k.scala 24050:34]
    .io_a(inst_SnxnLv4Inst21_io_a),
    .io_b(inst_SnxnLv4Inst21_io_b),
    .io_z(inst_SnxnLv4Inst21_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst22 ( // @[Snxn100k.scala 24054:34]
    .io_a(inst_SnxnLv4Inst22_io_a),
    .io_b(inst_SnxnLv4Inst22_io_b),
    .io_z(inst_SnxnLv4Inst22_io_z)
  );
  SnxnLv4Inst23 inst_SnxnLv4Inst23 ( // @[Snxn100k.scala 24058:34]
    .io_a(inst_SnxnLv4Inst23_io_a),
    .io_b(inst_SnxnLv4Inst23_io_b),
    .io_z(inst_SnxnLv4Inst23_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 24063:15]
  assign inst_SnxnLv4Inst20_io_a = io_a; // @[Snxn100k.scala 24047:27]
  assign inst_SnxnLv4Inst20_io_b = io_b; // @[Snxn100k.scala 24048:27]
  assign inst_SnxnLv4Inst21_io_a = io_a; // @[Snxn100k.scala 24051:27]
  assign inst_SnxnLv4Inst21_io_b = io_b; // @[Snxn100k.scala 24052:27]
  assign inst_SnxnLv4Inst22_io_a = io_a; // @[Snxn100k.scala 24055:27]
  assign inst_SnxnLv4Inst22_io_b = io_b; // @[Snxn100k.scala 24056:27]
  assign inst_SnxnLv4Inst23_io_a = io_a; // @[Snxn100k.scala 24059:27]
  assign inst_SnxnLv4Inst23_io_b = io_b; // @[Snxn100k.scala 24060:27]
endmodule
module SnxnLv4Inst24(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82577:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82578:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82579:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82580:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82581:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82582:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82583:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82584:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82585:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82586:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82587:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82588:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82589:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82590:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82591:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82592:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82593:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82594:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82595:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 82596:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 82597:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 82598:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 82599:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 82600:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 82601:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 82602:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 82603:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 82604:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 82605:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 82606:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 82607:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 82608:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 82609:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 82610:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 82611:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 82612:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 82613:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 82614:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 82615:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 82616:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 82617:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 82618:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 82619:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 82620:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 82621:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 82622:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 82623:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 82624:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 82625:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 82626:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 82627:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 82628:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 82629:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 82630:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 82631:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 82632:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 82633:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 82634:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 82635:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 82636:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 82637:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 82638:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 82639:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 82640:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 82641:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 82642:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 82643:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 82644:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 82645:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 82646:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 82647:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 82648:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 82649:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 82650:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 82651:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 82652:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 82653:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 82654:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 82655:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 82656:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82657:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82658:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82659:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82660:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82661:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82662:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82663:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82664:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82665:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82666:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82667:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82668:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82669:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82670:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82671:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82672:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82673:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82674:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82675:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82676:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82677:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82678:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82679:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82680:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82681:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82682:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82683:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82684:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82685:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82686:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82687:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82688:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82689:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82690:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82691:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82692:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82693:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82694:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82695:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82696:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82697:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82698:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82699:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82700:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82701:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82702:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82703:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82704:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82705:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82706:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82707:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82708:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82709:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82710:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82711:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82712:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82713:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82714:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82715:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82716:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82717:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82718:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82719:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82720:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82721:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82722:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82723:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82724:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82725:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82726:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82727:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82728:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82729:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82730:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82731:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82732:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82733:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82734:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82735:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82736:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82737:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82738:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82739:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82740:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82741:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82742:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82743:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82744:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82745:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82746:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82747:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82748:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82749:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82750:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82751:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 82752:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 82753:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 82754:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 82755:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 82756:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 82757:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 82758:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 82759:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 82760:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 82761:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 82762:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 82763:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 82764:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 82765:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 82766:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 82767:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 82768:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 82769:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 82770:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 82771:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 82772:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 82773:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 82774:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 82775:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 82776:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 82777:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 82778:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 82779:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 82780:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 82781:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 82782:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 82783:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 82784:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 82785:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 82786:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 82787:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 82788:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 82789:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 82790:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 82791:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 82792:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 82793:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 82794:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 82795:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 82796:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 82797:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 82798:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 82799:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 82800:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 82801:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 82802:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 82803:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 82804:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 82805:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 82806:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 82807:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 82808:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 82809:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 82810:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 82811:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 82812:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 82813:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 82814:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 82815:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 82816:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 82817:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 82818:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 82819:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 82820:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 82821:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 82822:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 82823:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 82824:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 82825:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 82826:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 82827:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 82828:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 82829:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 82830:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 82831:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 82832:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 82833:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 82834:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 82835:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 82836:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 82837:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 82838:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 82839:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 82840:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 82841:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 82842:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 82843:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 82844:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 82845:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 82846:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 82847:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 82848:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 82849:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 82850:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 82851:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 82852:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 82853:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 82854:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 82855:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 82856:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 82857:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 82858:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 82859:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 82860:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 82861:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 82862:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 82863:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 82864:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 82865:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 82866:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 82867:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 82868:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 82869:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 82870:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 82871:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 82872:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 82873:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 82874:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 82875:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 82876:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 82877:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 82878:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 82879:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 82880:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 82881:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 82882:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 82883:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 82884:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 82885:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 82886:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 82887:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 82888:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 82889:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 82890:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 82891:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 82892:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 82893:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 82894:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 82895:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 82896:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 82897:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 82898:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 82899:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 82900:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 82901:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 82902:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 82903:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 82904:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 82905:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 82906:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 82907:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 82908:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 82909:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 82910:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 82911:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 82912:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 82913:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 82914:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 82915:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 82916:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 82917:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 82918:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 82919:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 82920:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 82921:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 82922:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 82923:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 82924:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 82925:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 82926:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 82927:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 82928:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 82929:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 82930:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 82931:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 82932:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 82933:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 82934:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 82935:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 82936:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 82937:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 82938:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 82939:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 82940:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 82941:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 82942:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 82943:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 82944:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 82945:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 82946:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 82947:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 82948:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 82949:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 82950:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 82951:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 82952:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 82953:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 82954:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 82955:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 82956:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 82957:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 82958:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 82959:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 82960:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 82961:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 82962:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 82963:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 82964:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 82965:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 82966:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 82967:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 82968:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 82969:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 82970:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 82971:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 82972:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 82973:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 82974:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 82975:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 82976:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 82977:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 82978:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 82979:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 82980:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 82981:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 82982:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 82983:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 82984:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 82985:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 82986:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 82987:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 82988:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 82989:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 82990:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 82991:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 82992:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 82993:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 82994:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 82995:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 82996:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 82997:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 82998:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 82999:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 83000:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 83001:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 83002:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 83003:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 83004:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 83005:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 83006:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 83007:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 83008:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 83009:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 83010:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 83011:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 83012:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 83013:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 83014:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 83015:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 83016:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 83017:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 83018:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 83019:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 83020:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 83021:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 83022:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 83023:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 83024:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 83025:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 83026:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 83027:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 83028:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 83029:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 83030:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 83031:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 83032:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 83033:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 83034:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 83035:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 83036:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 83037:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 83038:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 83039:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 83040:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 83041:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 83042:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 83043:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 83044:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 83045:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 83046:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 83047:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 83048:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 83049:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 83050:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 83051:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 83052:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 83053:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 83054:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 83055:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 83056:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 83057:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 83058:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 83059:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 83060:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 83061:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 83062:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 83063:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 83064:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 83065:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 83066:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 83067:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 83068:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 83069:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 83070:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 83071:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 83072:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 83073:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 83074:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 83075:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 83076:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 83077:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 83078:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 83079:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 83080:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 83081:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 83082:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 83083:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 83084:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 83085:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 83086:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 83087:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 83088:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 83089:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 83090:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 83091:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 83092:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 83093:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 83094:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 83095:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 83096:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 83097:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 83098:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 83099:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 83100:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 83101:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 83102:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 83103:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 83104:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 83105:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 83106:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 83107:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 83108:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 83109:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 83110:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 83111:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 83112:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 83113:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 83114:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 83115:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 83116:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 83117:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 83118:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 83119:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 83120:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 83121:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 83122:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 83123:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 83124:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 83125:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 83126:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 83127:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 83128:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 83129:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 83130:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 83131:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 83132:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 83133:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 83134:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 83135:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 83136:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 83137:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 83138:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 83139:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 83140:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 83141:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 83142:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 83143:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 83144:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 83145:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 83146:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 83147:22]
  assign io_z = ~x142; // @[Snxn100k.scala 83148:17]
endmodule
module SnxnLv4Inst25(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82343:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82344:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82345:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82346:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82347:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82348:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82349:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82350:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82351:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82352:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82353:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82354:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82355:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82356:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82357:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82358:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82359:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82360:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82361:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 82362:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 82363:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 82364:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 82365:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 82366:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 82367:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 82368:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 82369:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 82370:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 82371:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 82372:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 82373:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 82374:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 82375:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 82376:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 82377:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 82378:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 82379:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 82380:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 82381:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 82382:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 82383:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 82384:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 82385:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 82386:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 82387:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 82388:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 82389:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 82390:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 82391:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 82392:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 82393:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 82394:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 82395:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 82396:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 82397:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 82398:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 82399:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 82400:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 82401:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 82402:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 82403:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 82404:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 82405:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 82406:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 82407:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 82408:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 82409:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 82410:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 82411:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 82412:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 82413:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 82414:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 82415:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 82416:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 82417:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 82418:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 82419:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 82420:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 82421:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 82422:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82423:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82424:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82425:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82426:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82427:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82428:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82429:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82430:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82431:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82432:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82433:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82434:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82435:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82436:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82437:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82438:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82439:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82440:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82441:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82442:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82443:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82444:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82445:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82446:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82447:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82448:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82449:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82450:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82451:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82452:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82453:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82454:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82455:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82456:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82457:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82458:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82459:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82460:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82461:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82462:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82463:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82464:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82465:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82466:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82467:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82468:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82469:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82470:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82471:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82472:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82473:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82474:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82475:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82476:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82477:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82478:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82479:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82480:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82481:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82482:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82483:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82484:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82485:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82486:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82487:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82488:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82489:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82490:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82491:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82492:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82493:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82494:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82495:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82496:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82497:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82498:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82499:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82500:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82501:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82502:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82503:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82504:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82505:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82506:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82507:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82508:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82509:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82510:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82511:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82512:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82513:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82514:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82515:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82516:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82517:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 82518:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 82519:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 82520:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 82521:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 82522:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 82523:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 82524:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 82525:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 82526:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 82527:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 82528:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 82529:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 82530:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 82531:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 82532:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 82533:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 82534:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 82535:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 82536:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 82537:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 82538:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 82539:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 82540:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 82541:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 82542:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 82543:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 82544:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 82545:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 82546:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 82547:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 82548:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 82549:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 82550:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 82551:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 82552:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 82553:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 82554:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 82555:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 82556:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 82557:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 82558:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 82559:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 82560:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 82561:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 82562:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 82563:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 82564:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 82565:20]
  assign io_z = ~x55; // @[Snxn100k.scala 82566:16]
endmodule
module SnxnLv4Inst26(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82313:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82314:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82315:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82316:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82317:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82318:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82319:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82320:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82321:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82322:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82323:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82324:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82325:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82326:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82327:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82328:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82329:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82330:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82331:18]
  assign io_z = ~x4; // @[Snxn100k.scala 82332:15]
endmodule
module SnxnLv4Inst27(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 82127:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 82128:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 82129:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 82130:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 82131:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 82132:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 82133:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 82134:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 82135:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 82136:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 82137:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 82138:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 82139:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 82140:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 82141:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 82142:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 82143:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 82144:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 82145:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 82146:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 82147:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 82148:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 82149:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 82150:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 82151:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 82152:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 82153:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 82154:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 82155:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 82156:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 82157:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 82158:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 82159:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 82160:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 82161:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 82162:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 82163:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 82164:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 82165:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 82166:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 82167:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 82168:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 82169:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 82170:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 82171:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 82172:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 82173:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 82174:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 82175:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 82176:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 82177:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 82178:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 82179:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 82180:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 82181:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 82182:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 82183:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 82184:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 82185:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 82186:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 82187:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 82188:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 82189:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 82190:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 82191:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 82192:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 82193:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 82194:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 82195:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 82196:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 82197:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 82198:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 82199:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 82200:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 82201:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 82202:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 82203:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 82204:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 82205:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 82206:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 82207:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 82208:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 82209:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 82210:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 82211:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 82212:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 82213:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 82214:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 82215:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 82216:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 82217:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 82218:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 82219:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 82220:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 82221:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 82222:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 82223:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 82224:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 82225:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 82226:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 82227:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 82228:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 82229:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 82230:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 82231:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 82232:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 82233:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 82234:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 82235:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 82236:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 82237:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 82238:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 82239:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 82240:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 82241:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 82242:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 82243:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 82244:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 82245:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 82246:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 82247:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 82248:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 82249:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 82250:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 82251:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 82252:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 82253:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 82254:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 82255:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 82256:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 82257:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 82258:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 82259:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 82260:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 82261:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 82262:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 82263:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 82264:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 82265:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 82266:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 82267:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 82268:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 82269:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 82270:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 82271:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 82272:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 82273:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 82274:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 82275:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 82276:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 82277:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 82278:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 82279:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 82280:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 82281:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82282:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82283:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82284:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82285:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82286:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82287:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82288:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82289:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82290:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82291:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82292:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82293:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82294:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82295:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82296:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82297:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82298:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82299:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82300:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82301:20]
  assign io_z = ~x43; // @[Snxn100k.scala 82302:16]
endmodule
module SnxnLv3Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst24_io_a; // @[Snxn100k.scala 25015:34]
  wire  inst_SnxnLv4Inst24_io_b; // @[Snxn100k.scala 25015:34]
  wire  inst_SnxnLv4Inst24_io_z; // @[Snxn100k.scala 25015:34]
  wire  inst_SnxnLv4Inst25_io_a; // @[Snxn100k.scala 25019:34]
  wire  inst_SnxnLv4Inst25_io_b; // @[Snxn100k.scala 25019:34]
  wire  inst_SnxnLv4Inst25_io_z; // @[Snxn100k.scala 25019:34]
  wire  inst_SnxnLv4Inst26_io_a; // @[Snxn100k.scala 25023:34]
  wire  inst_SnxnLv4Inst26_io_b; // @[Snxn100k.scala 25023:34]
  wire  inst_SnxnLv4Inst26_io_z; // @[Snxn100k.scala 25023:34]
  wire  inst_SnxnLv4Inst27_io_a; // @[Snxn100k.scala 25027:34]
  wire  inst_SnxnLv4Inst27_io_b; // @[Snxn100k.scala 25027:34]
  wire  inst_SnxnLv4Inst27_io_z; // @[Snxn100k.scala 25027:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst24_io_z + inst_SnxnLv4Inst25_io_z; // @[Snxn100k.scala 25031:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst26_io_z; // @[Snxn100k.scala 25031:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst27_io_z; // @[Snxn100k.scala 25031:89]
  SnxnLv4Inst24 inst_SnxnLv4Inst24 ( // @[Snxn100k.scala 25015:34]
    .io_a(inst_SnxnLv4Inst24_io_a),
    .io_b(inst_SnxnLv4Inst24_io_b),
    .io_z(inst_SnxnLv4Inst24_io_z)
  );
  SnxnLv4Inst25 inst_SnxnLv4Inst25 ( // @[Snxn100k.scala 25019:34]
    .io_a(inst_SnxnLv4Inst25_io_a),
    .io_b(inst_SnxnLv4Inst25_io_b),
    .io_z(inst_SnxnLv4Inst25_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst26 ( // @[Snxn100k.scala 25023:34]
    .io_a(inst_SnxnLv4Inst26_io_a),
    .io_b(inst_SnxnLv4Inst26_io_b),
    .io_z(inst_SnxnLv4Inst26_io_z)
  );
  SnxnLv4Inst27 inst_SnxnLv4Inst27 ( // @[Snxn100k.scala 25027:34]
    .io_a(inst_SnxnLv4Inst27_io_a),
    .io_b(inst_SnxnLv4Inst27_io_b),
    .io_z(inst_SnxnLv4Inst27_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25032:15]
  assign inst_SnxnLv4Inst24_io_a = io_a; // @[Snxn100k.scala 25016:27]
  assign inst_SnxnLv4Inst24_io_b = io_b; // @[Snxn100k.scala 25017:27]
  assign inst_SnxnLv4Inst25_io_a = io_a; // @[Snxn100k.scala 25020:27]
  assign inst_SnxnLv4Inst25_io_b = io_b; // @[Snxn100k.scala 25021:27]
  assign inst_SnxnLv4Inst26_io_a = io_a; // @[Snxn100k.scala 25024:27]
  assign inst_SnxnLv4Inst26_io_b = io_b; // @[Snxn100k.scala 25025:27]
  assign inst_SnxnLv4Inst27_io_a = io_a; // @[Snxn100k.scala 25028:27]
  assign inst_SnxnLv4Inst27_io_b = io_b; // @[Snxn100k.scala 25029:27]
endmodule
module SnxnLv4Inst29(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81349:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81350:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81351:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81352:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81353:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81354:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81355:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81356:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81357:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81358:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81359:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81360:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81361:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81362:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81363:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81364:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81365:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81366:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81367:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81368:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81369:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81370:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81371:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81372:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81373:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81374:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81375:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81376:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81377:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81378:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81379:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81380:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81381:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81382:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81383:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81384:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81385:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81386:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81387:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81388:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81389:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81390:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81391:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81392:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81393:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81394:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81395:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81396:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81397:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81398:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81399:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81400:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81401:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81402:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81403:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81404:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81405:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81406:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81407:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81408:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81409:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81410:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81411:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81412:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81413:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81414:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81415:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81416:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81417:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81418:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81419:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81420:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81421:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81422:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81423:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81424:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81425:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81426:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81427:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81428:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 81429:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 81430:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 81431:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 81432:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 81433:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 81434:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 81435:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 81436:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 81437:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 81438:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 81439:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 81440:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 81441:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 81442:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 81443:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 81444:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 81445:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 81446:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 81447:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 81448:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 81449:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 81450:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 81451:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 81452:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 81453:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 81454:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 81455:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 81456:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 81457:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 81458:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 81459:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 81460:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 81461:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 81462:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 81463:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 81464:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 81465:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 81466:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 81467:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 81468:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 81469:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 81470:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 81471:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 81472:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 81473:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 81474:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 81475:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 81476:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 81477:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 81478:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 81479:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 81480:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 81481:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 81482:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 81483:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 81484:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 81485:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 81486:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 81487:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 81488:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 81489:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 81490:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 81491:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 81492:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 81493:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 81494:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 81495:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 81496:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 81497:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 81498:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 81499:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 81500:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 81501:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 81502:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81503:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 81504:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 81505:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 81506:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 81507:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 81508:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 81509:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 81510:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 81511:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 81512:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 81513:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 81514:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 81515:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 81516:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 81517:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 81518:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 81519:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 81520:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 81521:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 81522:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 81523:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 81524:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 81525:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 81526:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 81527:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 81528:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 81529:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 81530:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 81531:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 81532:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 81533:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 81534:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 81535:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 81536:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 81537:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 81538:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 81539:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 81540:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 81541:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 81542:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 81543:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 81544:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 81545:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 81546:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 81547:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 81548:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 81549:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 81550:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 81551:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 81552:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 81553:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 81554:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 81555:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 81556:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 81557:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 81558:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 81559:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 81560:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 81561:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 81562:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 81563:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 81564:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 81565:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 81566:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 81567:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 81568:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 81569:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 81570:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 81571:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 81572:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 81573:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 81574:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 81575:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 81576:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 81577:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 81578:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 81579:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 81580:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 81581:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 81582:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 81583:20]
  assign io_z = ~x58; // @[Snxn100k.scala 81584:16]
endmodule
module SnxnLv4Inst30(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81845:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81846:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81847:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81848:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81849:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81850:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81851:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81852:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81853:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81854:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81855:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81856:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81857:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81858:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81859:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81860:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81861:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81862:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81863:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81864:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81865:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81866:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81867:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81868:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81869:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81870:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81871:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81872:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81873:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81874:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81875:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81876:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81877:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81878:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81879:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81880:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81881:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81882:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81883:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81884:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81885:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81886:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81887:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81888:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81889:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81890:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81891:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81892:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81893:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81894:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81895:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81896:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81897:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81898:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81899:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81900:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81901:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81902:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81903:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81904:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81905:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81906:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81907:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81908:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81909:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81910:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81911:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81912:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81913:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81914:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81915:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81916:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81917:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81918:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81919:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81920:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81921:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81922:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81923:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81924:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 81925:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 81926:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 81927:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 81928:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 81929:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 81930:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 81931:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 81932:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 81933:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 81934:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 81935:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 81936:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 81937:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 81938:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 81939:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 81940:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 81941:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 81942:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 81943:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 81944:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 81945:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 81946:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 81947:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 81948:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 81949:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 81950:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 81951:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 81952:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 81953:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 81954:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 81955:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 81956:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 81957:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 81958:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 81959:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 81960:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 81961:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 81962:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 81963:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 81964:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 81965:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 81966:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 81967:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 81968:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 81969:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 81970:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 81971:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 81972:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 81973:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 81974:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 81975:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 81976:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 81977:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 81978:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 81979:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 81980:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 81981:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 81982:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 81983:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 81984:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 81985:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 81986:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 81987:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 81988:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 81989:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 81990:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 81991:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 81992:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 81993:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 81994:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 81995:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 81996:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 81997:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 81998:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81999:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 82000:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 82001:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 82002:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 82003:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 82004:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 82005:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 82006:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 82007:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 82008:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 82009:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 82010:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 82011:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 82012:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 82013:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 82014:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 82015:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 82016:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 82017:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 82018:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 82019:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 82020:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 82021:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 82022:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 82023:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 82024:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 82025:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 82026:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 82027:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 82028:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 82029:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 82030:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 82031:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 82032:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 82033:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 82034:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 82035:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 82036:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 82037:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 82038:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 82039:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 82040:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 82041:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 82042:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 82043:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 82044:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 82045:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 82046:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 82047:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 82048:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 82049:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 82050:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 82051:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 82052:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 82053:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 82054:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 82055:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 82056:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 82057:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 82058:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 82059:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 82060:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 82061:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 82062:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 82063:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 82064:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 82065:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 82066:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 82067:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 82068:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 82069:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 82070:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 82071:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 82072:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 82073:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 82074:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 82075:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 82076:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 82077:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 82078:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 82079:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 82080:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 82081:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 82082:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 82083:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 82084:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 82085:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 82086:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 82087:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 82088:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 82089:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 82090:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 82091:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 82092:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 82093:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 82094:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 82095:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 82096:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 82097:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 82098:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 82099:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 82100:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 82101:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 82102:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 82103:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 82104:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 82105:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 82106:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 82107:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 82108:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 82109:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 82110:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 82111:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 82112:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 82113:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 82114:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 82115:20]
  assign io_z = ~x67; // @[Snxn100k.scala 82116:16]
endmodule
module SnxnLv4Inst31(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 81123:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 81124:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 81125:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 81126:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 81127:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 81128:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 81129:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 81130:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 81131:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 81132:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 81133:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 81134:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 81135:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 81136:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 81137:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 81138:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 81139:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 81140:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 81141:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 81142:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 81143:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 81144:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 81145:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 81146:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 81147:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 81148:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 81149:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 81150:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 81151:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 81152:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 81153:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 81154:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 81155:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 81156:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 81157:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 81158:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 81159:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 81160:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 81161:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 81162:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 81163:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 81164:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 81165:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 81166:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 81167:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 81168:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 81169:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 81170:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 81171:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 81172:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 81173:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 81174:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 81175:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 81176:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 81177:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 81178:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 81179:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 81180:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 81181:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 81182:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 81183:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 81184:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 81185:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 81186:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 81187:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 81188:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 81189:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 81190:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 81191:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 81192:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 81193:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 81194:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 81195:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 81196:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 81197:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 81198:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 81199:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 81200:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 81201:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 81202:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 81203:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 81204:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 81205:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 81206:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 81207:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 81208:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 81209:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 81210:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 81211:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 81212:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 81213:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 81214:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 81215:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 81216:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 81217:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 81218:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 81219:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 81220:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 81221:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 81222:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 81223:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 81224:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 81225:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 81226:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 81227:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 81228:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 81229:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 81230:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 81231:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 81232:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 81233:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 81234:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 81235:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 81236:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 81237:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 81238:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 81239:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 81240:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 81241:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 81242:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 81243:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 81244:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 81245:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 81246:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 81247:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 81248:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 81249:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 81250:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 81251:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 81252:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 81253:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 81254:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 81255:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 81256:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 81257:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 81258:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 81259:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 81260:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 81261:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 81262:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 81263:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 81264:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 81265:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 81266:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 81267:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 81268:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 81269:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 81270:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 81271:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 81272:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 81273:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 81274:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 81275:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 81276:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 81277:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 81278:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 81279:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 81280:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 81281:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 81282:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 81283:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 81284:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 81285:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 81286:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 81287:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 81288:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 81289:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 81290:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 81291:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 81292:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 81293:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 81294:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 81295:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 81296:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 81297:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 81298:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 81299:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 81300:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 81301:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 81302:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 81303:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 81304:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 81305:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 81306:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 81307:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 81308:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 81309:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 81310:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 81311:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 81312:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 81313:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 81314:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 81315:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 81316:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 81317:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 81318:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 81319:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 81320:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 81321:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 81322:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 81323:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 81324:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 81325:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 81326:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 81327:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 81328:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 81329:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 81330:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 81331:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 81332:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 81333:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 81334:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 81335:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 81336:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 81337:20]
  assign io_z = ~x53; // @[Snxn100k.scala 81338:16]
endmodule
module SnxnLv3Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst28_io_a; // @[Snxn100k.scala 24436:34]
  wire  inst_SnxnLv4Inst28_io_b; // @[Snxn100k.scala 24436:34]
  wire  inst_SnxnLv4Inst28_io_z; // @[Snxn100k.scala 24436:34]
  wire  inst_SnxnLv4Inst29_io_a; // @[Snxn100k.scala 24440:34]
  wire  inst_SnxnLv4Inst29_io_b; // @[Snxn100k.scala 24440:34]
  wire  inst_SnxnLv4Inst29_io_z; // @[Snxn100k.scala 24440:34]
  wire  inst_SnxnLv4Inst30_io_a; // @[Snxn100k.scala 24444:34]
  wire  inst_SnxnLv4Inst30_io_b; // @[Snxn100k.scala 24444:34]
  wire  inst_SnxnLv4Inst30_io_z; // @[Snxn100k.scala 24444:34]
  wire  inst_SnxnLv4Inst31_io_a; // @[Snxn100k.scala 24448:34]
  wire  inst_SnxnLv4Inst31_io_b; // @[Snxn100k.scala 24448:34]
  wire  inst_SnxnLv4Inst31_io_z; // @[Snxn100k.scala 24448:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst28_io_z + inst_SnxnLv4Inst29_io_z; // @[Snxn100k.scala 24452:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst30_io_z; // @[Snxn100k.scala 24452:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst31_io_z; // @[Snxn100k.scala 24452:89]
  SnxnLv4Inst7 inst_SnxnLv4Inst28 ( // @[Snxn100k.scala 24436:34]
    .io_a(inst_SnxnLv4Inst28_io_a),
    .io_b(inst_SnxnLv4Inst28_io_b),
    .io_z(inst_SnxnLv4Inst28_io_z)
  );
  SnxnLv4Inst29 inst_SnxnLv4Inst29 ( // @[Snxn100k.scala 24440:34]
    .io_a(inst_SnxnLv4Inst29_io_a),
    .io_b(inst_SnxnLv4Inst29_io_b),
    .io_z(inst_SnxnLv4Inst29_io_z)
  );
  SnxnLv4Inst30 inst_SnxnLv4Inst30 ( // @[Snxn100k.scala 24444:34]
    .io_a(inst_SnxnLv4Inst30_io_a),
    .io_b(inst_SnxnLv4Inst30_io_b),
    .io_z(inst_SnxnLv4Inst30_io_z)
  );
  SnxnLv4Inst31 inst_SnxnLv4Inst31 ( // @[Snxn100k.scala 24448:34]
    .io_a(inst_SnxnLv4Inst31_io_a),
    .io_b(inst_SnxnLv4Inst31_io_b),
    .io_z(inst_SnxnLv4Inst31_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 24453:15]
  assign inst_SnxnLv4Inst28_io_a = io_a; // @[Snxn100k.scala 24437:27]
  assign inst_SnxnLv4Inst28_io_b = io_b; // @[Snxn100k.scala 24438:27]
  assign inst_SnxnLv4Inst29_io_a = io_a; // @[Snxn100k.scala 24441:27]
  assign inst_SnxnLv4Inst29_io_b = io_b; // @[Snxn100k.scala 24442:27]
  assign inst_SnxnLv4Inst30_io_a = io_a; // @[Snxn100k.scala 24445:27]
  assign inst_SnxnLv4Inst30_io_b = io_b; // @[Snxn100k.scala 24446:27]
  assign inst_SnxnLv4Inst31_io_a = io_a; // @[Snxn100k.scala 24449:27]
  assign inst_SnxnLv4Inst31_io_b = io_b; // @[Snxn100k.scala 24450:27]
endmodule
module SnxnLv2Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst4_io_a; // @[Snxn100k.scala 7217:33]
  wire  inst_SnxnLv3Inst4_io_b; // @[Snxn100k.scala 7217:33]
  wire  inst_SnxnLv3Inst4_io_z; // @[Snxn100k.scala 7217:33]
  wire  inst_SnxnLv3Inst5_io_a; // @[Snxn100k.scala 7221:33]
  wire  inst_SnxnLv3Inst5_io_b; // @[Snxn100k.scala 7221:33]
  wire  inst_SnxnLv3Inst5_io_z; // @[Snxn100k.scala 7221:33]
  wire  inst_SnxnLv3Inst6_io_a; // @[Snxn100k.scala 7225:33]
  wire  inst_SnxnLv3Inst6_io_b; // @[Snxn100k.scala 7225:33]
  wire  inst_SnxnLv3Inst6_io_z; // @[Snxn100k.scala 7225:33]
  wire  inst_SnxnLv3Inst7_io_a; // @[Snxn100k.scala 7229:33]
  wire  inst_SnxnLv3Inst7_io_b; // @[Snxn100k.scala 7229:33]
  wire  inst_SnxnLv3Inst7_io_z; // @[Snxn100k.scala 7229:33]
  wire  _sum_T_1 = inst_SnxnLv3Inst4_io_z + inst_SnxnLv3Inst5_io_z; // @[Snxn100k.scala 7233:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst6_io_z; // @[Snxn100k.scala 7233:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst7_io_z; // @[Snxn100k.scala 7233:86]
  SnxnLv3Inst4 inst_SnxnLv3Inst4 ( // @[Snxn100k.scala 7217:33]
    .io_a(inst_SnxnLv3Inst4_io_a),
    .io_b(inst_SnxnLv3Inst4_io_b),
    .io_z(inst_SnxnLv3Inst4_io_z)
  );
  SnxnLv3Inst5 inst_SnxnLv3Inst5 ( // @[Snxn100k.scala 7221:33]
    .io_a(inst_SnxnLv3Inst5_io_a),
    .io_b(inst_SnxnLv3Inst5_io_b),
    .io_z(inst_SnxnLv3Inst5_io_z)
  );
  SnxnLv3Inst6 inst_SnxnLv3Inst6 ( // @[Snxn100k.scala 7225:33]
    .io_a(inst_SnxnLv3Inst6_io_a),
    .io_b(inst_SnxnLv3Inst6_io_b),
    .io_z(inst_SnxnLv3Inst6_io_z)
  );
  SnxnLv3Inst7 inst_SnxnLv3Inst7 ( // @[Snxn100k.scala 7229:33]
    .io_a(inst_SnxnLv3Inst7_io_a),
    .io_b(inst_SnxnLv3Inst7_io_b),
    .io_z(inst_SnxnLv3Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7234:15]
  assign inst_SnxnLv3Inst4_io_a = io_a; // @[Snxn100k.scala 7218:26]
  assign inst_SnxnLv3Inst4_io_b = io_b; // @[Snxn100k.scala 7219:26]
  assign inst_SnxnLv3Inst5_io_a = io_a; // @[Snxn100k.scala 7222:26]
  assign inst_SnxnLv3Inst5_io_b = io_b; // @[Snxn100k.scala 7223:26]
  assign inst_SnxnLv3Inst6_io_a = io_a; // @[Snxn100k.scala 7226:26]
  assign inst_SnxnLv3Inst6_io_b = io_b; // @[Snxn100k.scala 7227:26]
  assign inst_SnxnLv3Inst7_io_a = io_a; // @[Snxn100k.scala 7230:26]
  assign inst_SnxnLv3Inst7_io_b = io_b; // @[Snxn100k.scala 7231:26]
endmodule
module SnxnLv4Inst32(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 73527:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 73528:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 73529:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 73530:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 73531:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 73532:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 73533:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 73534:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 73535:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 73536:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 73537:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 73538:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 73539:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 73540:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 73541:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 73542:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 73543:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 73544:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 73545:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 73546:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 73547:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 73548:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 73549:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 73550:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 73551:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 73552:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 73553:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 73554:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 73555:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 73556:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 73557:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 73558:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 73559:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 73560:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 73561:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 73562:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 73563:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 73564:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 73565:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 73566:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 73567:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 73568:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 73569:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 73570:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 73571:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 73572:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 73573:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 73574:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 73575:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 73576:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 73577:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 73578:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 73579:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 73580:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 73581:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 73582:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 73583:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 73584:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 73585:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 73586:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 73587:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 73588:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 73589:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 73590:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 73591:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 73592:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 73593:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 73594:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 73595:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 73596:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 73597:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 73598:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 73599:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 73600:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 73601:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 73602:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 73603:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 73604:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 73605:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 73606:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 73607:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 73608:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 73609:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 73610:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 73611:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 73612:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 73613:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 73614:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 73615:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 73616:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 73617:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 73618:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 73619:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 73620:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 73621:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 73622:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 73623:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 73624:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 73625:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 73626:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 73627:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 73628:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 73629:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 73630:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 73631:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 73632:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 73633:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 73634:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 73635:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 73636:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 73637:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 73638:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 73639:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 73640:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 73641:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 73642:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 73643:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 73644:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 73645:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 73646:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 73647:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 73648:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 73649:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 73650:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 73651:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 73652:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 73653:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 73654:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 73655:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 73656:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 73657:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 73658:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 73659:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 73660:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 73661:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 73662:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 73663:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 73664:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 73665:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 73666:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 73667:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 73668:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 73669:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 73670:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 73671:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 73672:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 73673:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 73674:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 73675:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 73676:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 73677:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 73678:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 73679:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 73680:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 73681:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 73682:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 73683:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 73684:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 73685:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 73686:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 73687:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 73688:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 73689:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 73690:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 73691:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 73692:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 73693:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 73694:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 73695:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 73696:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 73697:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 73698:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 73699:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 73700:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 73701:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 73702:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 73703:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 73704:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 73705:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 73706:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 73707:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 73708:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 73709:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 73710:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 73711:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 73712:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 73713:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 73714:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 73715:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 73716:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 73717:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 73718:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 73719:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 73720:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 73721:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 73722:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 73723:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 73724:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 73725:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 73726:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 73727:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 73728:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 73729:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 73730:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 73731:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 73732:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 73733:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 73734:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 73735:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 73736:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 73737:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 73738:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 73739:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 73740:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 73741:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 73742:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 73743:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 73744:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 73745:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 73746:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 73747:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 73748:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 73749:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 73750:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 73751:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 73752:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 73753:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 73754:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 73755:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 73756:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 73757:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 73758:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 73759:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 73760:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 73761:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 73762:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 73763:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 73764:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 73765:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 73766:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 73767:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 73768:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 73769:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 73770:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 73771:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 73772:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 73773:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 73774:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 73775:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 73776:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 73777:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 73778:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 73779:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 73780:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 73781:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 73782:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 73783:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 73784:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 73785:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 73786:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 73787:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 73788:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 73789:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 73790:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 73791:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 73792:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 73793:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 73794:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 73795:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 73796:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 73797:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 73798:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 73799:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 73800:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 73801:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 73802:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 73803:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 73804:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 73805:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 73806:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 73807:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 73808:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 73809:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 73810:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 73811:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 73812:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 73813:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 73814:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 73815:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 73816:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 73817:20]
  assign io_z = ~x72; // @[Snxn100k.scala 73818:16]
endmodule
module SnxnLv4Inst33(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 74227:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 74228:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 74229:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 74230:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 74231:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 74232:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 74233:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 74234:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 74235:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 74236:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 74237:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 74238:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 74239:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 74240:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 74241:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 74242:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 74243:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 74244:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 74245:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 74246:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 74247:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 74248:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 74249:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 74250:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 74251:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 74252:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 74253:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 74254:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 74255:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 74256:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 74257:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 74258:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 74259:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 74260:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 74261:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 74262:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 74263:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 74264:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 74265:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 74266:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 74267:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 74268:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 74269:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 74270:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 74271:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 74272:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 74273:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 74274:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 74275:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 74276:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 74277:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 74278:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 74279:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 74280:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 74281:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 74282:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 74283:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 74284:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 74285:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 74286:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 74287:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 74288:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 74289:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 74290:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 74291:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 74292:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 74293:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 74294:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 74295:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 74296:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 74297:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 74298:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 74299:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 74300:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 74301:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 74302:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 74303:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 74304:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 74305:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 74306:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 74307:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 74308:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 74309:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 74310:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 74311:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 74312:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 74313:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 74314:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 74315:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 74316:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 74317:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 74318:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 74319:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 74320:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 74321:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 74322:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 74323:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 74324:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 74325:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 74326:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 74327:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 74328:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 74329:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 74330:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 74331:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 74332:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 74333:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 74334:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 74335:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 74336:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 74337:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 74338:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 74339:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 74340:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 74341:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 74342:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 74343:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 74344:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 74345:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 74346:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 74347:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 74348:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 74349:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 74350:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 74351:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 74352:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 74353:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 74354:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 74355:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 74356:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 74357:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 74358:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 74359:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 74360:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 74361:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 74362:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 74363:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 74364:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 74365:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 74366:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 74367:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 74368:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 74369:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 74370:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 74371:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 74372:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 74373:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 74374:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 74375:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 74376:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 74377:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 74378:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 74379:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 74380:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 74381:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 74382:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 74383:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 74384:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 74385:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 74386:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 74387:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 74388:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 74389:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 74390:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 74391:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 74392:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 74393:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 74394:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 74395:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 74396:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 74397:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 74398:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 74399:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 74400:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 74401:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 74402:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 74403:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 74404:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 74405:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 74406:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 74407:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 74408:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 74409:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 74410:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 74411:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 74412:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 74413:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 74414:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 74415:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 74416:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 74417:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 74418:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 74419:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 74420:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 74421:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 74422:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 74423:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 74424:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 74425:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 74426:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 74427:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 74428:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 74429:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 74430:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 74431:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 74432:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 74433:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 74434:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 74435:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 74436:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 74437:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 74438:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 74439:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 74440:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 74441:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 74442:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 74443:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 74444:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 74445:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 74446:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 74447:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 74448:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 74449:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 74450:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 74451:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 74452:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 74453:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 74454:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 74455:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 74456:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 74457:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 74458:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 74459:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 74460:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 74461:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 74462:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 74463:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 74464:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 74465:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 74466:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 74467:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 74468:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 74469:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 74470:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 74471:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 74472:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 74473:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 74474:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 74475:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 74476:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 74477:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 74478:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 74479:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 74480:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 74481:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 74482:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 74483:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 74484:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 74485:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 74486:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 74487:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 74488:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 74489:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 74490:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 74491:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 74492:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 74493:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 74494:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 74495:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 74496:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 74497:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 74498:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 74499:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 74500:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 74501:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 74502:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 74503:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 74504:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 74505:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 74506:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 74507:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 74508:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 74509:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 74510:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 74511:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 74512:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 74513:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 74514:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 74515:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 74516:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 74517:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 74518:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 74519:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 74520:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 74521:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 74522:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 74523:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 74524:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 74525:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 74526:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 74527:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 74528:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 74529:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 74530:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 74531:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 74532:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 74533:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 74534:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 74535:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 74536:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 74537:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 74538:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 74539:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 74540:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 74541:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 74542:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 74543:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 74544:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 74545:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 74546:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 74547:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 74548:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 74549:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 74550:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 74551:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 74552:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 74553:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 74554:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 74555:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 74556:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 74557:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 74558:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 74559:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 74560:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 74561:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 74562:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 74563:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 74564:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 74565:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 74566:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 74567:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 74568:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 74569:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 74570:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 74571:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 74572:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 74573:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 74574:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 74575:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 74576:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 74577:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 74578:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 74579:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 74580:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 74581:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 74582:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 74583:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 74584:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 74585:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 74586:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 74587:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 74588:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 74589:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 74590:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 74591:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 74592:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 74593:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 74594:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 74595:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 74596:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 74597:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 74598:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 74599:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 74600:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 74601:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 74602:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 74603:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 74604:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 74605:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 74606:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 74607:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 74608:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 74609:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 74610:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 74611:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 74612:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 74613:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 74614:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 74615:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 74616:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 74617:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 74618:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 74619:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 74620:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 74621:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 74622:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 74623:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 74624:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 74625:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 74626:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 74627:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 74628:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 74629:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 74630:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 74631:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 74632:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 74633:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 74634:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 74635:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 74636:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 74637:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 74638:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 74639:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 74640:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 74641:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 74642:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 74643:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 74644:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 74645:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 74646:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 74647:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 74648:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 74649:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 74650:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 74651:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 74652:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 74653:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 74654:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 74655:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 74656:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 74657:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 74658:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 74659:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 74660:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 74661:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 74662:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 74663:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 74664:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 74665:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 74666:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 74667:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 74668:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 74669:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 74670:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 74671:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 74672:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 74673:22]
  assign io_z = ~x111; // @[Snxn100k.scala 74674:17]
endmodule
module SnxnLv4Inst34(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 74685:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 74686:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 74687:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 74688:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 74689:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 74690:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 74691:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 74692:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 74693:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 74694:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 74695:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 74696:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 74697:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 74698:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 74699:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 74700:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 74701:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 74702:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 74703:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 74704:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 74705:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 74706:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 74707:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 74708:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 74709:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 74710:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 74711:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 74712:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 74713:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 74714:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 74715:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 74716:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 74717:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 74718:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 74719:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 74720:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 74721:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 74722:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 74723:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 74724:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 74725:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 74726:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 74727:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 74728:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 74729:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 74730:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 74731:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 74732:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 74733:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 74734:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 74735:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 74736:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 74737:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 74738:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 74739:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 74740:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 74741:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 74742:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 74743:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 74744:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 74745:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 74746:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 74747:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 74748:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 74749:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 74750:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 74751:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 74752:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 74753:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 74754:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 74755:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 74756:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 74757:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 74758:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 74759:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 74760:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 74761:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 74762:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 74763:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 74764:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 74765:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 74766:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 74767:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 74768:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 74769:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 74770:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 74771:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 74772:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 74773:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 74774:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 74775:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 74776:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 74777:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 74778:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 74779:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 74780:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 74781:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 74782:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 74783:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 74784:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 74785:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 74786:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 74787:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 74788:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 74789:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 74790:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 74791:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 74792:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 74793:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 74794:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 74795:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 74796:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 74797:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 74798:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 74799:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 74800:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 74801:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 74802:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 74803:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 74804:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 74805:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 74806:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 74807:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 74808:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 74809:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 74810:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 74811:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 74812:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 74813:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 74814:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 74815:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 74816:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 74817:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 74818:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 74819:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 74820:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 74821:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 74822:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 74823:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 74824:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 74825:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 74826:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 74827:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 74828:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 74829:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 74830:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 74831:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 74832:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 74833:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 74834:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 74835:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 74836:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 74837:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 74838:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 74839:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 74840:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 74841:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 74842:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 74843:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 74844:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 74845:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 74846:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 74847:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 74848:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 74849:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 74850:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 74851:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 74852:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 74853:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 74854:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 74855:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 74856:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 74857:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 74858:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 74859:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 74860:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 74861:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 74862:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 74863:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 74864:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 74865:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 74866:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 74867:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 74868:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 74869:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 74870:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 74871:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 74872:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 74873:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 74874:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 74875:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 74876:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 74877:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 74878:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 74879:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 74880:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 74881:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 74882:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 74883:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 74884:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 74885:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 74886:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 74887:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 74888:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 74889:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 74890:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 74891:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 74892:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 74893:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 74894:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 74895:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 74896:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 74897:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 74898:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 74899:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 74900:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 74901:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 74902:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 74903:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 74904:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 74905:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 74906:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 74907:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 74908:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 74909:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 74910:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 74911:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 74912:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 74913:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 74914:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 74915:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 74916:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 74917:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 74918:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 74919:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 74920:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 74921:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 74922:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 74923:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 74924:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 74925:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 74926:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 74927:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 74928:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 74929:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 74930:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 74931:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 74932:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 74933:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 74934:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 74935:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 74936:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 74937:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 74938:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 74939:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 74940:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 74941:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 74942:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 74943:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 74944:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 74945:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 74946:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 74947:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 74948:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 74949:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 74950:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 74951:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 74952:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 74953:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 74954:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 74955:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 74956:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 74957:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 74958:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 74959:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 74960:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 74961:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 74962:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 74963:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 74964:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 74965:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 74966:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 74967:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 74968:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 74969:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 74970:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 74971:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 74972:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 74973:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 74974:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 74975:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 74976:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 74977:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 74978:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 74979:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 74980:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 74981:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 74982:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 74983:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 74984:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 74985:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 74986:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 74987:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 74988:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 74989:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 74990:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 74991:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 74992:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 74993:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 74994:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 74995:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 74996:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 74997:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 74998:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 74999:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 75000:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 75001:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 75002:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 75003:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 75004:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 75005:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 75006:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 75007:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 75008:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 75009:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 75010:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 75011:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 75012:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 75013:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 75014:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 75015:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 75016:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 75017:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 75018:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 75019:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 75020:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 75021:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 75022:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 75023:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 75024:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 75025:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 75026:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 75027:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 75028:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 75029:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 75030:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 75031:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 75032:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 75033:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 75034:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 75035:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 75036:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 75037:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 75038:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 75039:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 75040:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 75041:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 75042:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 75043:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 75044:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 75045:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 75046:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 75047:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 75048:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 75049:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 75050:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 75051:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 75052:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 75053:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 75054:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 75055:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 75056:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 75057:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 75058:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 75059:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 75060:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 75061:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 75062:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 75063:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 75064:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 75065:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 75066:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 75067:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 75068:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 75069:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 75070:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 75071:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 75072:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 75073:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 75074:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 75075:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 75076:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 75077:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 75078:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 75079:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 75080:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 75081:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 75082:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 75083:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 75084:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 75085:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 75086:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 75087:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 75088:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 75089:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 75090:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 75091:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 75092:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 75093:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 75094:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 75095:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 75096:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 75097:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 75098:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 75099:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 75100:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 75101:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 75102:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 75103:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 75104:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 75105:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 75106:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 75107:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 75108:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 75109:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 75110:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 75111:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 75112:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 75113:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 75114:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 75115:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 75116:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 75117:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 75118:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 75119:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 75120:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 75121:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 75122:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 75123:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 75124:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 75125:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 75126:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 75127:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 75128:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 75129:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 75130:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 75131:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 75132:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 75133:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 75134:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 75135:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 75136:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 75137:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 75138:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 75139:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 75140:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 75141:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 75142:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 75143:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 75144:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 75145:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 75146:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 75147:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 75148:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 75149:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 75150:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 75151:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 75152:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 75153:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 75154:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 75155:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 75156:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 75157:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 75158:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 75159:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 75160:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 75161:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 75162:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 75163:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 75164:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 75165:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 75166:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 75167:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 75168:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 75169:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 75170:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 75171:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 75172:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 75173:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 75174:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 75175:22]
  assign io_z = ~x122; // @[Snxn100k.scala 75176:17]
endmodule
module SnxnLv3Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst32_io_a; // @[Snxn100k.scala 23202:34]
  wire  inst_SnxnLv4Inst32_io_b; // @[Snxn100k.scala 23202:34]
  wire  inst_SnxnLv4Inst32_io_z; // @[Snxn100k.scala 23202:34]
  wire  inst_SnxnLv4Inst33_io_a; // @[Snxn100k.scala 23206:34]
  wire  inst_SnxnLv4Inst33_io_b; // @[Snxn100k.scala 23206:34]
  wire  inst_SnxnLv4Inst33_io_z; // @[Snxn100k.scala 23206:34]
  wire  inst_SnxnLv4Inst34_io_a; // @[Snxn100k.scala 23210:34]
  wire  inst_SnxnLv4Inst34_io_b; // @[Snxn100k.scala 23210:34]
  wire  inst_SnxnLv4Inst34_io_z; // @[Snxn100k.scala 23210:34]
  wire  inst_SnxnLv4Inst35_io_a; // @[Snxn100k.scala 23214:34]
  wire  inst_SnxnLv4Inst35_io_b; // @[Snxn100k.scala 23214:34]
  wire  inst_SnxnLv4Inst35_io_z; // @[Snxn100k.scala 23214:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst32_io_z + inst_SnxnLv4Inst33_io_z; // @[Snxn100k.scala 23218:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst34_io_z; // @[Snxn100k.scala 23218:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst35_io_z; // @[Snxn100k.scala 23218:89]
  SnxnLv4Inst32 inst_SnxnLv4Inst32 ( // @[Snxn100k.scala 23202:34]
    .io_a(inst_SnxnLv4Inst32_io_a),
    .io_b(inst_SnxnLv4Inst32_io_b),
    .io_z(inst_SnxnLv4Inst32_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst33 ( // @[Snxn100k.scala 23206:34]
    .io_a(inst_SnxnLv4Inst33_io_a),
    .io_b(inst_SnxnLv4Inst33_io_b),
    .io_z(inst_SnxnLv4Inst33_io_z)
  );
  SnxnLv4Inst34 inst_SnxnLv4Inst34 ( // @[Snxn100k.scala 23210:34]
    .io_a(inst_SnxnLv4Inst34_io_a),
    .io_b(inst_SnxnLv4Inst34_io_b),
    .io_z(inst_SnxnLv4Inst34_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst35 ( // @[Snxn100k.scala 23214:34]
    .io_a(inst_SnxnLv4Inst35_io_a),
    .io_b(inst_SnxnLv4Inst35_io_b),
    .io_z(inst_SnxnLv4Inst35_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23219:15]
  assign inst_SnxnLv4Inst32_io_a = io_a; // @[Snxn100k.scala 23203:27]
  assign inst_SnxnLv4Inst32_io_b = io_b; // @[Snxn100k.scala 23204:27]
  assign inst_SnxnLv4Inst33_io_a = io_a; // @[Snxn100k.scala 23207:27]
  assign inst_SnxnLv4Inst33_io_b = io_b; // @[Snxn100k.scala 23208:27]
  assign inst_SnxnLv4Inst34_io_a = io_a; // @[Snxn100k.scala 23211:27]
  assign inst_SnxnLv4Inst34_io_b = io_b; // @[Snxn100k.scala 23212:27]
  assign inst_SnxnLv4Inst35_io_a = io_a; // @[Snxn100k.scala 23215:27]
  assign inst_SnxnLv4Inst35_io_b = io_b; // @[Snxn100k.scala 23216:27]
endmodule
module SnxnLv4Inst36(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 76539:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 76540:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 76541:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 76542:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 76543:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 76544:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 76545:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 76546:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 76547:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 76548:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 76549:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 76550:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 76551:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 76552:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 76553:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 76554:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 76555:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 76556:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 76557:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 76558:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 76559:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 76560:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 76561:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 76562:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 76563:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 76564:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 76565:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 76566:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 76567:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 76568:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 76569:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 76570:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 76571:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 76572:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 76573:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 76574:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 76575:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 76576:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 76577:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 76578:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 76579:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 76580:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 76581:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 76582:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 76583:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 76584:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 76585:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 76586:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 76587:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 76588:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 76589:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 76590:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 76591:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 76592:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 76593:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 76594:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 76595:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 76596:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 76597:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 76598:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 76599:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 76600:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 76601:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 76602:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 76603:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 76604:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 76605:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 76606:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 76607:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 76608:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 76609:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 76610:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 76611:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 76612:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 76613:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 76614:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 76615:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 76616:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 76617:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 76618:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 76619:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 76620:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 76621:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 76622:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 76623:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 76624:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 76625:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 76626:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 76627:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 76628:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 76629:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 76630:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 76631:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 76632:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 76633:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 76634:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 76635:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 76636:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 76637:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 76638:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 76639:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 76640:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 76641:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 76642:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 76643:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 76644:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 76645:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 76646:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 76647:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 76648:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 76649:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 76650:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 76651:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 76652:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 76653:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 76654:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 76655:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 76656:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 76657:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 76658:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 76659:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 76660:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 76661:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 76662:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 76663:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 76664:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 76665:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 76666:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 76667:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 76668:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 76669:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 76670:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 76671:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 76672:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 76673:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 76674:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 76675:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 76676:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 76677:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 76678:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 76679:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 76680:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 76681:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 76682:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 76683:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 76684:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 76685:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 76686:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 76687:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 76688:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 76689:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 76690:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 76691:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 76692:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 76693:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 76694:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 76695:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 76696:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 76697:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 76698:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 76699:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 76700:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 76701:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 76702:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 76703:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 76704:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 76705:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 76706:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 76707:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 76708:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 76709:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 76710:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 76711:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 76712:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 76713:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 76714:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 76715:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 76716:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 76717:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 76718:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 76719:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 76720:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 76721:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 76722:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 76723:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 76724:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 76725:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 76726:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 76727:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 76728:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 76729:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 76730:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 76731:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 76732:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 76733:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 76734:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 76735:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 76736:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 76737:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 76738:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 76739:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 76740:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 76741:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 76742:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 76743:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 76744:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 76745:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 76746:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 76747:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 76748:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 76749:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 76750:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 76751:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 76752:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 76753:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 76754:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 76755:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 76756:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 76757:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 76758:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 76759:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 76760:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 76761:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 76762:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 76763:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 76764:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 76765:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 76766:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 76767:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 76768:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 76769:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 76770:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 76771:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 76772:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 76773:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 76774:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 76775:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 76776:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 76777:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 76778:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 76779:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 76780:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 76781:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 76782:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 76783:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 76784:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 76785:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 76786:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 76787:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 76788:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 76789:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 76790:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 76791:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 76792:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 76793:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 76794:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 76795:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 76796:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 76797:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 76798:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 76799:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 76800:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 76801:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 76802:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 76803:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 76804:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 76805:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 76806:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 76807:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 76808:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 76809:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 76810:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 76811:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 76812:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 76813:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 76814:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 76815:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 76816:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 76817:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 76818:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 76819:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 76820:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 76821:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 76822:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 76823:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 76824:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 76825:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 76826:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 76827:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 76828:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 76829:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 76830:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 76831:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 76832:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 76833:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 76834:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 76835:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 76836:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 76837:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 76838:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 76839:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 76840:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 76841:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 76842:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 76843:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 76844:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 76845:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 76846:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 76847:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 76848:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 76849:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 76850:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 76851:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 76852:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 76853:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 76854:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 76855:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 76856:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 76857:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 76858:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 76859:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 76860:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 76861:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 76862:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 76863:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 76864:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 76865:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 76866:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 76867:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 76868:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 76869:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 76870:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 76871:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 76872:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 76873:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 76874:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 76875:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 76876:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 76877:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 76878:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 76879:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 76880:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 76881:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 76882:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 76883:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 76884:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 76885:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 76886:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 76887:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 76888:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 76889:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 76890:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 76891:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 76892:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 76893:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 76894:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 76895:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 76896:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 76897:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 76898:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 76899:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 76900:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 76901:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 76902:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 76903:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 76904:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 76905:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 76906:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 76907:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 76908:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 76909:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 76910:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 76911:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 76912:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 76913:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 76914:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 76915:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 76916:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 76917:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 76918:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 76919:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 76920:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 76921:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 76922:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 76923:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 76924:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 76925:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 76926:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 76927:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 76928:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 76929:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 76930:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 76931:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 76932:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 76933:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 76934:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 76935:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 76936:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 76937:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 76938:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 76939:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 76940:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 76941:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 76942:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 76943:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 76944:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 76945:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 76946:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 76947:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 76948:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 76949:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 76950:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 76951:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 76952:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 76953:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 76954:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 76955:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 76956:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 76957:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 76958:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 76959:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 76960:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 76961:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 76962:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 76963:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 76964:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 76965:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 76966:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 76967:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 76968:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 76969:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 76970:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 76971:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 76972:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 76973:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 76974:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 76975:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 76976:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 76977:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 76978:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 76979:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 76980:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 76981:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 76982:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 76983:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 76984:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 76985:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 76986:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 76987:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 76988:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 76989:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 76990:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 76991:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 76992:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 76993:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 76994:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 76995:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 76996:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 76997:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 76998:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 76999:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 77000:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 77001:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 77002:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 77003:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 77004:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 77005:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 77006:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 77007:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 77008:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 77009:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 77010:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 77011:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 77012:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 77013:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 77014:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 77015:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 77016:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 77017:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 77018:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 77019:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 77020:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 77021:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 77022:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 77023:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 77024:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 77025:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 77026:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 77027:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 77028:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 77029:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 77030:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 77031:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 77032:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 77033:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 77034:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 77035:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 77036:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 77037:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 77038:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 77039:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 77040:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 77041:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 77042:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 77043:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 77044:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 77045:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 77046:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 77047:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 77048:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 77049:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 77050:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 77051:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 77052:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 77053:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 77054:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 77055:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 77056:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 77057:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 77058:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 77059:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 77060:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 77061:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 77062:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 77063:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 77064:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 77065:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 77066:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 77067:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 77068:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 77069:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 77070:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 77071:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 77072:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 77073:22]
  assign io_z = ~x133; // @[Snxn100k.scala 77074:17]
endmodule
module SnxnLv4Inst38(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75967:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75968:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75969:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75970:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75971:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75972:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75973:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75974:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75975:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75976:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75977:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75978:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75979:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75980:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75981:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75982:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75983:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75984:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75985:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75986:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75987:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75988:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75989:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75990:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75991:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75992:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75993:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75994:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75995:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75996:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75997:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75998:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75999:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 76000:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 76001:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 76002:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 76003:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 76004:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 76005:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 76006:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 76007:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 76008:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 76009:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 76010:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 76011:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 76012:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 76013:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 76014:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 76015:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 76016:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 76017:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 76018:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 76019:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 76020:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 76021:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 76022:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 76023:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 76024:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 76025:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 76026:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 76027:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 76028:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 76029:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 76030:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 76031:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 76032:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 76033:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 76034:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 76035:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 76036:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 76037:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 76038:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 76039:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 76040:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 76041:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 76042:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 76043:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 76044:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 76045:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 76046:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 76047:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 76048:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 76049:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 76050:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 76051:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 76052:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 76053:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 76054:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 76055:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 76056:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 76057:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 76058:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 76059:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 76060:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 76061:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 76062:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 76063:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 76064:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 76065:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 76066:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 76067:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 76068:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 76069:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 76070:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 76071:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 76072:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 76073:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 76074:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 76075:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 76076:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 76077:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 76078:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 76079:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 76080:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 76081:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 76082:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 76083:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 76084:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 76085:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 76086:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 76087:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 76088:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 76089:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 76090:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 76091:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 76092:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 76093:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 76094:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 76095:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 76096:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 76097:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 76098:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 76099:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 76100:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 76101:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 76102:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 76103:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 76104:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 76105:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 76106:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 76107:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 76108:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 76109:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 76110:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 76111:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 76112:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 76113:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 76114:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 76115:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 76116:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 76117:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 76118:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 76119:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 76120:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 76121:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 76122:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 76123:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 76124:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 76125:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 76126:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 76127:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 76128:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 76129:20]
  assign io_z = ~x40; // @[Snxn100k.scala 76130:16]
endmodule
module SnxnLv3Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst36_io_a; // @[Snxn100k.scala 23572:34]
  wire  inst_SnxnLv4Inst36_io_b; // @[Snxn100k.scala 23572:34]
  wire  inst_SnxnLv4Inst36_io_z; // @[Snxn100k.scala 23572:34]
  wire  inst_SnxnLv4Inst37_io_a; // @[Snxn100k.scala 23576:34]
  wire  inst_SnxnLv4Inst37_io_b; // @[Snxn100k.scala 23576:34]
  wire  inst_SnxnLv4Inst37_io_z; // @[Snxn100k.scala 23576:34]
  wire  inst_SnxnLv4Inst38_io_a; // @[Snxn100k.scala 23580:34]
  wire  inst_SnxnLv4Inst38_io_b; // @[Snxn100k.scala 23580:34]
  wire  inst_SnxnLv4Inst38_io_z; // @[Snxn100k.scala 23580:34]
  wire  inst_SnxnLv4Inst39_io_a; // @[Snxn100k.scala 23584:34]
  wire  inst_SnxnLv4Inst39_io_b; // @[Snxn100k.scala 23584:34]
  wire  inst_SnxnLv4Inst39_io_z; // @[Snxn100k.scala 23584:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst36_io_z + inst_SnxnLv4Inst37_io_z; // @[Snxn100k.scala 23588:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst38_io_z; // @[Snxn100k.scala 23588:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst39_io_z; // @[Snxn100k.scala 23588:89]
  SnxnLv4Inst36 inst_SnxnLv4Inst36 ( // @[Snxn100k.scala 23572:34]
    .io_a(inst_SnxnLv4Inst36_io_a),
    .io_b(inst_SnxnLv4Inst36_io_b),
    .io_z(inst_SnxnLv4Inst36_io_z)
  );
  SnxnLv4Inst36 inst_SnxnLv4Inst37 ( // @[Snxn100k.scala 23576:34]
    .io_a(inst_SnxnLv4Inst37_io_a),
    .io_b(inst_SnxnLv4Inst37_io_b),
    .io_z(inst_SnxnLv4Inst37_io_z)
  );
  SnxnLv4Inst38 inst_SnxnLv4Inst38 ( // @[Snxn100k.scala 23580:34]
    .io_a(inst_SnxnLv4Inst38_io_a),
    .io_b(inst_SnxnLv4Inst38_io_b),
    .io_z(inst_SnxnLv4Inst38_io_z)
  );
  SnxnLv4Inst22 inst_SnxnLv4Inst39 ( // @[Snxn100k.scala 23584:34]
    .io_a(inst_SnxnLv4Inst39_io_a),
    .io_b(inst_SnxnLv4Inst39_io_b),
    .io_z(inst_SnxnLv4Inst39_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23589:15]
  assign inst_SnxnLv4Inst36_io_a = io_a; // @[Snxn100k.scala 23573:27]
  assign inst_SnxnLv4Inst36_io_b = io_b; // @[Snxn100k.scala 23574:27]
  assign inst_SnxnLv4Inst37_io_a = io_a; // @[Snxn100k.scala 23577:27]
  assign inst_SnxnLv4Inst37_io_b = io_b; // @[Snxn100k.scala 23578:27]
  assign inst_SnxnLv4Inst38_io_a = io_a; // @[Snxn100k.scala 23581:27]
  assign inst_SnxnLv4Inst38_io_b = io_b; // @[Snxn100k.scala 23582:27]
  assign inst_SnxnLv4Inst39_io_a = io_a; // @[Snxn100k.scala 23585:27]
  assign inst_SnxnLv4Inst39_io_b = io_b; // @[Snxn100k.scala 23586:27]
endmodule
module SnxnLv4Inst40(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75855:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75856:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75857:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75858:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75859:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75860:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75861:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75862:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75863:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75864:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75865:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75866:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75867:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75868:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75869:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75870:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75871:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75872:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75873:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75874:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75875:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75876:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75877:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75878:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75879:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75880:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75881:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75882:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75883:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75884:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75885:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75886:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75887:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 75888:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 75889:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 75890:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 75891:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 75892:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 75893:18]
  assign io_z = ~x9; // @[Snxn100k.scala 75894:15]
endmodule
module SnxnLv4Inst41(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75187:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75188:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75189:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75190:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75191:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75192:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75193:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75194:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75195:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75196:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75197:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75198:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75199:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75200:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75201:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75202:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75203:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75204:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75205:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75206:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75207:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75208:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75209:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75210:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75211:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75212:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75213:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75214:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75215:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75216:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75217:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75218:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75219:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 75220:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 75221:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 75222:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 75223:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 75224:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 75225:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 75226:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 75227:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 75228:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 75229:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 75230:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 75231:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 75232:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 75233:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 75234:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 75235:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 75236:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 75237:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 75238:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 75239:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 75240:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 75241:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 75242:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 75243:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 75244:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 75245:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 75246:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 75247:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 75248:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 75249:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 75250:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 75251:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 75252:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 75253:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 75254:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 75255:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 75256:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 75257:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 75258:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 75259:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 75260:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 75261:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 75262:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 75263:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 75264:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 75265:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 75266:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 75267:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 75268:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 75269:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 75270:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 75271:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 75272:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 75273:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 75274:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 75275:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 75276:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 75277:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 75278:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 75279:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 75280:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 75281:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 75282:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 75283:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 75284:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 75285:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 75286:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 75287:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 75288:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 75289:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 75290:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 75291:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 75292:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 75293:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 75294:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 75295:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 75296:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 75297:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 75298:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 75299:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 75300:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 75301:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 75302:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 75303:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 75304:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 75305:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 75306:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 75307:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 75308:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 75309:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 75310:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 75311:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 75312:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 75313:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 75314:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 75315:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 75316:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 75317:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 75318:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 75319:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 75320:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 75321:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 75322:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 75323:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 75324:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 75325:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 75326:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 75327:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 75328:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 75329:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 75330:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 75331:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 75332:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 75333:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 75334:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 75335:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 75336:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 75337:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 75338:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 75339:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 75340:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 75341:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 75342:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 75343:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 75344:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 75345:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 75346:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 75347:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 75348:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 75349:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 75350:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 75351:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 75352:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 75353:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 75354:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 75355:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 75356:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 75357:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 75358:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 75359:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 75360:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 75361:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 75362:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 75363:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 75364:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 75365:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 75366:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 75367:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 75368:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 75369:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 75370:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 75371:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 75372:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 75373:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 75374:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 75375:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 75376:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 75377:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 75378:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 75379:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 75380:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 75381:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 75382:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 75383:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 75384:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 75385:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 75386:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 75387:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 75388:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 75389:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 75390:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 75391:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 75392:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 75393:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 75394:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 75395:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 75396:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 75397:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 75398:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 75399:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 75400:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 75401:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 75402:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 75403:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 75404:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 75405:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 75406:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 75407:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 75408:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 75409:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 75410:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 75411:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 75412:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 75413:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 75414:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 75415:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 75416:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 75417:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 75418:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 75419:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 75420:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 75421:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 75422:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 75423:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 75424:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 75425:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 75426:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 75427:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 75428:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 75429:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 75430:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 75431:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 75432:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 75433:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 75434:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 75435:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 75436:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 75437:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 75438:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 75439:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 75440:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 75441:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 75442:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 75443:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 75444:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 75445:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 75446:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 75447:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 75448:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 75449:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 75450:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 75451:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 75452:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 75453:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 75454:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 75455:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 75456:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 75457:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 75458:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 75459:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 75460:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 75461:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 75462:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 75463:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 75464:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 75465:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 75466:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 75467:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 75468:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 75469:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 75470:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 75471:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 75472:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 75473:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 75474:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 75475:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 75476:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 75477:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 75478:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 75479:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 75480:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 75481:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 75482:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 75483:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 75484:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 75485:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 75486:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 75487:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 75488:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 75489:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 75490:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 75491:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 75492:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 75493:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 75494:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 75495:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 75496:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 75497:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 75498:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 75499:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 75500:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 75501:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 75502:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 75503:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 75504:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 75505:20]
  assign io_z = ~x79; // @[Snxn100k.scala 75506:16]
endmodule
module SnxnLv4Inst42(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75905:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75906:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75907:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75908:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75909:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75910:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75911:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75912:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75913:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75914:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75915:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75916:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75917:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75918:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75919:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75920:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75921:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75922:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75923:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75924:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75925:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75926:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75927:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75928:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75929:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75930:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75931:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75932:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75933:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75934:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75935:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75936:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75937:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 75938:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 75939:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 75940:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 75941:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 75942:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 75943:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 75944:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 75945:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 75946:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 75947:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 75948:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 75949:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 75950:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 75951:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 75952:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 75953:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 75954:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 75955:20]
  assign io_z = ~x12; // @[Snxn100k.scala 75956:16]
endmodule
module SnxnLv4Inst43(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 75517:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 75518:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 75519:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 75520:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 75521:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 75522:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 75523:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 75524:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 75525:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 75526:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 75527:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 75528:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 75529:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 75530:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 75531:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 75532:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 75533:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 75534:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 75535:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 75536:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 75537:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 75538:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 75539:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 75540:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 75541:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 75542:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 75543:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 75544:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 75545:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 75546:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 75547:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 75548:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 75549:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 75550:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 75551:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 75552:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 75553:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 75554:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 75555:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 75556:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 75557:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 75558:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 75559:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 75560:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 75561:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 75562:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 75563:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 75564:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 75565:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 75566:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 75567:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 75568:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 75569:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 75570:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 75571:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 75572:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 75573:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 75574:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 75575:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 75576:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 75577:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 75578:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 75579:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 75580:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 75581:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 75582:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 75583:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 75584:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 75585:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 75586:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 75587:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 75588:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 75589:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 75590:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 75591:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 75592:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 75593:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 75594:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 75595:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 75596:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 75597:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 75598:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 75599:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 75600:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 75601:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 75602:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 75603:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 75604:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 75605:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 75606:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 75607:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 75608:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 75609:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 75610:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 75611:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 75612:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 75613:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 75614:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 75615:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 75616:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 75617:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 75618:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 75619:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 75620:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 75621:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 75622:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 75623:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 75624:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 75625:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 75626:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 75627:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 75628:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 75629:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 75630:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 75631:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 75632:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 75633:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 75634:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 75635:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 75636:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 75637:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 75638:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 75639:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 75640:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 75641:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 75642:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 75643:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 75644:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 75645:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 75646:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 75647:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 75648:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 75649:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 75650:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 75651:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 75652:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 75653:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 75654:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 75655:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 75656:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 75657:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 75658:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 75659:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 75660:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 75661:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 75662:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 75663:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 75664:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 75665:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 75666:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 75667:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 75668:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 75669:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 75670:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 75671:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 75672:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 75673:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 75674:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 75675:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 75676:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 75677:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 75678:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 75679:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 75680:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 75681:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 75682:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 75683:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 75684:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 75685:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 75686:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 75687:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 75688:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 75689:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 75690:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 75691:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 75692:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 75693:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 75694:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 75695:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 75696:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 75697:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 75698:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 75699:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 75700:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 75701:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 75702:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 75703:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 75704:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 75705:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 75706:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 75707:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 75708:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 75709:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 75710:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 75711:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 75712:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 75713:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 75714:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 75715:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 75716:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 75717:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 75718:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 75719:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 75720:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 75721:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 75722:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 75723:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 75724:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 75725:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 75726:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 75727:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 75728:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 75729:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 75730:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 75731:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 75732:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 75733:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 75734:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 75735:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 75736:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 75737:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 75738:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 75739:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 75740:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 75741:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 75742:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 75743:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 75744:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 75745:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 75746:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 75747:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 75748:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 75749:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 75750:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 75751:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 75752:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 75753:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 75754:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 75755:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 75756:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 75757:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 75758:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 75759:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 75760:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 75761:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 75762:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 75763:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 75764:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 75765:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 75766:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 75767:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 75768:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 75769:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 75770:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 75771:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 75772:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 75773:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 75774:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 75775:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 75776:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 75777:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 75778:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 75779:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 75780:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 75781:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 75782:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 75783:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 75784:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 75785:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 75786:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 75787:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 75788:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 75789:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 75790:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 75791:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 75792:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 75793:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 75794:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 75795:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 75796:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 75797:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 75798:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 75799:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 75800:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 75801:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 75802:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 75803:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 75804:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 75805:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 75806:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 75807:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 75808:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 75809:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 75810:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 75811:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 75812:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 75813:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 75814:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 75815:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 75816:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 75817:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 75818:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 75819:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 75820:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 75821:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 75822:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 75823:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 75824:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 75825:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 75826:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 75827:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 75828:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 75829:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 75830:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 75831:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 75832:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 75833:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 75834:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 75835:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 75836:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 75837:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 75838:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 75839:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 75840:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 75841:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 75842:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 75843:20]
  assign io_z = ~x81; // @[Snxn100k.scala 75844:16]
endmodule
module SnxnLv3Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst40_io_a; // @[Snxn100k.scala 23513:34]
  wire  inst_SnxnLv4Inst40_io_b; // @[Snxn100k.scala 23513:34]
  wire  inst_SnxnLv4Inst40_io_z; // @[Snxn100k.scala 23513:34]
  wire  inst_SnxnLv4Inst41_io_a; // @[Snxn100k.scala 23517:34]
  wire  inst_SnxnLv4Inst41_io_b; // @[Snxn100k.scala 23517:34]
  wire  inst_SnxnLv4Inst41_io_z; // @[Snxn100k.scala 23517:34]
  wire  inst_SnxnLv4Inst42_io_a; // @[Snxn100k.scala 23521:34]
  wire  inst_SnxnLv4Inst42_io_b; // @[Snxn100k.scala 23521:34]
  wire  inst_SnxnLv4Inst42_io_z; // @[Snxn100k.scala 23521:34]
  wire  inst_SnxnLv4Inst43_io_a; // @[Snxn100k.scala 23525:34]
  wire  inst_SnxnLv4Inst43_io_b; // @[Snxn100k.scala 23525:34]
  wire  inst_SnxnLv4Inst43_io_z; // @[Snxn100k.scala 23525:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst40_io_z + inst_SnxnLv4Inst41_io_z; // @[Snxn100k.scala 23529:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst42_io_z; // @[Snxn100k.scala 23529:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst43_io_z; // @[Snxn100k.scala 23529:89]
  SnxnLv4Inst40 inst_SnxnLv4Inst40 ( // @[Snxn100k.scala 23513:34]
    .io_a(inst_SnxnLv4Inst40_io_a),
    .io_b(inst_SnxnLv4Inst40_io_b),
    .io_z(inst_SnxnLv4Inst40_io_z)
  );
  SnxnLv4Inst41 inst_SnxnLv4Inst41 ( // @[Snxn100k.scala 23517:34]
    .io_a(inst_SnxnLv4Inst41_io_a),
    .io_b(inst_SnxnLv4Inst41_io_b),
    .io_z(inst_SnxnLv4Inst41_io_z)
  );
  SnxnLv4Inst42 inst_SnxnLv4Inst42 ( // @[Snxn100k.scala 23521:34]
    .io_a(inst_SnxnLv4Inst42_io_a),
    .io_b(inst_SnxnLv4Inst42_io_b),
    .io_z(inst_SnxnLv4Inst42_io_z)
  );
  SnxnLv4Inst43 inst_SnxnLv4Inst43 ( // @[Snxn100k.scala 23525:34]
    .io_a(inst_SnxnLv4Inst43_io_a),
    .io_b(inst_SnxnLv4Inst43_io_b),
    .io_z(inst_SnxnLv4Inst43_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 23530:15]
  assign inst_SnxnLv4Inst40_io_a = io_a; // @[Snxn100k.scala 23514:27]
  assign inst_SnxnLv4Inst40_io_b = io_b; // @[Snxn100k.scala 23515:27]
  assign inst_SnxnLv4Inst41_io_a = io_a; // @[Snxn100k.scala 23518:27]
  assign inst_SnxnLv4Inst41_io_b = io_b; // @[Snxn100k.scala 23519:27]
  assign inst_SnxnLv4Inst42_io_a = io_a; // @[Snxn100k.scala 23522:27]
  assign inst_SnxnLv4Inst42_io_b = io_b; // @[Snxn100k.scala 23523:27]
  assign inst_SnxnLv4Inst43_io_a = io_a; // @[Snxn100k.scala 23526:27]
  assign inst_SnxnLv4Inst43_io_b = io_b; // @[Snxn100k.scala 23527:27]
endmodule
module SnxnLv4Inst44(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78337:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78338:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78339:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78340:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78341:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78342:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78343:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78344:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78345:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78346:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78347:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78348:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78349:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78350:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78351:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78352:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78353:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78354:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78355:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78356:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78357:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78358:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78359:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78360:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78361:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78362:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78363:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78364:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78365:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78366:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78367:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78368:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78369:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78370:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78371:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78372:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78373:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78374:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78375:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78376:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78377:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78378:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78379:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78380:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78381:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78382:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78383:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78384:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78385:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78386:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78387:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78388:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78389:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78390:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78391:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78392:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78393:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78394:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78395:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78396:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78397:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78398:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78399:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78400:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78401:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78402:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78403:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78404:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78405:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78406:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78407:20]
  assign io_z = ~x17; // @[Snxn100k.scala 78408:16]
endmodule
module SnxnLv4Inst46(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 78051:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 78052:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 78053:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 78054:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 78055:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 78056:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 78057:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 78058:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 78059:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 78060:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 78061:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 78062:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 78063:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 78064:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 78065:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 78066:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 78067:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 78068:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 78069:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 78070:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 78071:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 78072:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 78073:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 78074:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 78075:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 78076:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 78077:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 78078:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 78079:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 78080:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 78081:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 78082:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 78083:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 78084:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 78085:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 78086:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 78087:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 78088:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 78089:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 78090:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 78091:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 78092:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 78093:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 78094:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 78095:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 78096:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 78097:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 78098:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 78099:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 78100:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 78101:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 78102:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 78103:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 78104:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 78105:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 78106:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 78107:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 78108:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 78109:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 78110:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 78111:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 78112:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 78113:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 78114:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 78115:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 78116:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 78117:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 78118:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 78119:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 78120:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 78121:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 78122:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 78123:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 78124:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 78125:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 78126:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 78127:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 78128:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 78129:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 78130:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 78131:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 78132:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 78133:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 78134:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 78135:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 78136:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 78137:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 78138:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 78139:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 78140:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 78141:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 78142:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 78143:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 78144:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 78145:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 78146:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 78147:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 78148:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 78149:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 78150:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 78151:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 78152:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 78153:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 78154:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 78155:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 78156:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 78157:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 78158:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 78159:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 78160:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 78161:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 78162:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 78163:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 78164:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 78165:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 78166:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 78167:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 78168:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 78169:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 78170:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 78171:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 78172:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 78173:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 78174:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 78175:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 78176:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 78177:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 78178:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 78179:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 78180:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 78181:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 78182:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 78183:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 78184:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 78185:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 78186:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 78187:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 78188:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 78189:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 78190:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 78191:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 78192:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 78193:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 78194:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 78195:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 78196:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 78197:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 78198:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 78199:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 78200:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 78201:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 78202:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 78203:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 78204:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 78205:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 78206:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 78207:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 78208:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 78209:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 78210:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 78211:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 78212:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 78213:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 78214:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 78215:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 78216:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 78217:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 78218:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 78219:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 78220:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 78221:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 78222:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 78223:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 78224:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 78225:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 78226:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 78227:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 78228:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 78229:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 78230:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 78231:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 78232:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 78233:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 78234:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 78235:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 78236:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 78237:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 78238:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 78239:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 78240:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 78241:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 78242:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 78243:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 78244:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 78245:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 78246:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 78247:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 78248:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 78249:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 78250:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 78251:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 78252:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 78253:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 78254:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 78255:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 78256:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 78257:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 78258:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 78259:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 78260:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 78261:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 78262:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 78263:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 78264:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 78265:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 78266:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 78267:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 78268:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 78269:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 78270:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 78271:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 78272:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 78273:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 78274:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 78275:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 78276:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 78277:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 78278:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 78279:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 78280:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 78281:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 78282:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 78283:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 78284:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 78285:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 78286:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 78287:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 78288:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 78289:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 78290:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 78291:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 78292:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 78293:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 78294:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 78295:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 78296:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 78297:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 78298:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 78299:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 78300:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 78301:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 78302:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 78303:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 78304:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 78305:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 78306:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 78307:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 78308:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 78309:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 78310:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 78311:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 78312:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 78313:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 78314:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 78315:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 78316:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 78317:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 78318:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 78319:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 78320:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 78321:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 78322:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 78323:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 78324:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 78325:20]
  assign io_z = ~x68; // @[Snxn100k.scala 78326:16]
endmodule
module SnxnLv4Inst47(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 77821:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 77822:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 77823:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 77824:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 77825:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 77826:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 77827:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 77828:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 77829:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 77830:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 77831:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 77832:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 77833:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 77834:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 77835:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 77836:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 77837:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 77838:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 77839:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 77840:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 77841:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 77842:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 77843:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 77844:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 77845:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 77846:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 77847:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 77848:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 77849:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 77850:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 77851:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 77852:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 77853:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 77854:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 77855:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 77856:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 77857:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 77858:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 77859:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 77860:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 77861:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 77862:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 77863:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 77864:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 77865:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 77866:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 77867:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 77868:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 77869:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 77870:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 77871:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 77872:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 77873:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 77874:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 77875:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 77876:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 77877:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 77878:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 77879:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 77880:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 77881:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 77882:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 77883:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 77884:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 77885:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 77886:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 77887:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 77888:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 77889:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 77890:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 77891:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 77892:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 77893:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 77894:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 77895:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 77896:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 77897:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 77898:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 77899:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 77900:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 77901:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 77902:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 77903:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 77904:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 77905:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 77906:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 77907:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 77908:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 77909:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 77910:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 77911:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 77912:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 77913:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 77914:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 77915:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 77916:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 77917:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 77918:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 77919:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 77920:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 77921:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 77922:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 77923:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 77924:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 77925:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 77926:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 77927:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 77928:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 77929:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 77930:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 77931:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 77932:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 77933:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 77934:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 77935:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 77936:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 77937:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 77938:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 77939:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 77940:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 77941:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 77942:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 77943:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 77944:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 77945:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 77946:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 77947:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 77948:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 77949:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 77950:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 77951:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 77952:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 77953:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 77954:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 77955:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 77956:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 77957:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 77958:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 77959:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 77960:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 77961:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 77962:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 77963:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 77964:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 77965:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 77966:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 77967:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 77968:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 77969:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 77970:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 77971:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 77972:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 77973:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 77974:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 77975:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 77976:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 77977:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 77978:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 77979:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 77980:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 77981:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 77982:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 77983:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 77984:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 77985:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 77986:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 77987:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 77988:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 77989:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 77990:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 77991:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 77992:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 77993:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 77994:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 77995:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 77996:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 77997:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 77998:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 77999:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 78000:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 78001:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 78002:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 78003:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 78004:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 78005:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 78006:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 78007:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 78008:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 78009:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 78010:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 78011:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 78012:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 78013:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 78014:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 78015:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 78016:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 78017:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 78018:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 78019:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 78020:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 78021:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 78022:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 78023:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 78024:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 78025:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 78026:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 78027:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 78028:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 78029:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 78030:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 78031:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 78032:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 78033:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 78034:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 78035:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 78036:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 78037:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 78038:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 78039:20]
  assign io_z = ~x54; // @[Snxn100k.scala 78040:16]
endmodule
module SnxnLv3Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst44_io_a; // @[Snxn100k.scala 24007:34]
  wire  inst_SnxnLv4Inst44_io_b; // @[Snxn100k.scala 24007:34]
  wire  inst_SnxnLv4Inst44_io_z; // @[Snxn100k.scala 24007:34]
  wire  inst_SnxnLv4Inst45_io_a; // @[Snxn100k.scala 24011:34]
  wire  inst_SnxnLv4Inst45_io_b; // @[Snxn100k.scala 24011:34]
  wire  inst_SnxnLv4Inst45_io_z; // @[Snxn100k.scala 24011:34]
  wire  inst_SnxnLv4Inst46_io_a; // @[Snxn100k.scala 24015:34]
  wire  inst_SnxnLv4Inst46_io_b; // @[Snxn100k.scala 24015:34]
  wire  inst_SnxnLv4Inst46_io_z; // @[Snxn100k.scala 24015:34]
  wire  inst_SnxnLv4Inst47_io_a; // @[Snxn100k.scala 24019:34]
  wire  inst_SnxnLv4Inst47_io_b; // @[Snxn100k.scala 24019:34]
  wire  inst_SnxnLv4Inst47_io_z; // @[Snxn100k.scala 24019:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst44_io_z + inst_SnxnLv4Inst45_io_z; // @[Snxn100k.scala 24023:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst46_io_z; // @[Snxn100k.scala 24023:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst47_io_z; // @[Snxn100k.scala 24023:89]
  SnxnLv4Inst44 inst_SnxnLv4Inst44 ( // @[Snxn100k.scala 24007:34]
    .io_a(inst_SnxnLv4Inst44_io_a),
    .io_b(inst_SnxnLv4Inst44_io_b),
    .io_z(inst_SnxnLv4Inst44_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst45 ( // @[Snxn100k.scala 24011:34]
    .io_a(inst_SnxnLv4Inst45_io_a),
    .io_b(inst_SnxnLv4Inst45_io_b),
    .io_z(inst_SnxnLv4Inst45_io_z)
  );
  SnxnLv4Inst46 inst_SnxnLv4Inst46 ( // @[Snxn100k.scala 24015:34]
    .io_a(inst_SnxnLv4Inst46_io_a),
    .io_b(inst_SnxnLv4Inst46_io_b),
    .io_z(inst_SnxnLv4Inst46_io_z)
  );
  SnxnLv4Inst47 inst_SnxnLv4Inst47 ( // @[Snxn100k.scala 24019:34]
    .io_a(inst_SnxnLv4Inst47_io_a),
    .io_b(inst_SnxnLv4Inst47_io_b),
    .io_z(inst_SnxnLv4Inst47_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 24024:15]
  assign inst_SnxnLv4Inst44_io_a = io_a; // @[Snxn100k.scala 24008:27]
  assign inst_SnxnLv4Inst44_io_b = io_b; // @[Snxn100k.scala 24009:27]
  assign inst_SnxnLv4Inst45_io_a = io_a; // @[Snxn100k.scala 24012:27]
  assign inst_SnxnLv4Inst45_io_b = io_b; // @[Snxn100k.scala 24013:27]
  assign inst_SnxnLv4Inst46_io_a = io_a; // @[Snxn100k.scala 24016:27]
  assign inst_SnxnLv4Inst46_io_b = io_b; // @[Snxn100k.scala 24017:27]
  assign inst_SnxnLv4Inst47_io_a = io_a; // @[Snxn100k.scala 24020:27]
  assign inst_SnxnLv4Inst47_io_b = io_b; // @[Snxn100k.scala 24021:27]
endmodule
module SnxnLv2Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst8_io_a; // @[Snxn100k.scala 7098:33]
  wire  inst_SnxnLv3Inst8_io_b; // @[Snxn100k.scala 7098:33]
  wire  inst_SnxnLv3Inst8_io_z; // @[Snxn100k.scala 7098:33]
  wire  inst_SnxnLv3Inst9_io_a; // @[Snxn100k.scala 7102:33]
  wire  inst_SnxnLv3Inst9_io_b; // @[Snxn100k.scala 7102:33]
  wire  inst_SnxnLv3Inst9_io_z; // @[Snxn100k.scala 7102:33]
  wire  inst_SnxnLv3Inst10_io_a; // @[Snxn100k.scala 7106:34]
  wire  inst_SnxnLv3Inst10_io_b; // @[Snxn100k.scala 7106:34]
  wire  inst_SnxnLv3Inst10_io_z; // @[Snxn100k.scala 7106:34]
  wire  inst_SnxnLv3Inst11_io_a; // @[Snxn100k.scala 7110:34]
  wire  inst_SnxnLv3Inst11_io_b; // @[Snxn100k.scala 7110:34]
  wire  inst_SnxnLv3Inst11_io_z; // @[Snxn100k.scala 7110:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst8_io_z + inst_SnxnLv3Inst9_io_z; // @[Snxn100k.scala 7114:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst10_io_z; // @[Snxn100k.scala 7114:61]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst11_io_z; // @[Snxn100k.scala 7114:87]
  SnxnLv3Inst8 inst_SnxnLv3Inst8 ( // @[Snxn100k.scala 7098:33]
    .io_a(inst_SnxnLv3Inst8_io_a),
    .io_b(inst_SnxnLv3Inst8_io_b),
    .io_z(inst_SnxnLv3Inst8_io_z)
  );
  SnxnLv3Inst9 inst_SnxnLv3Inst9 ( // @[Snxn100k.scala 7102:33]
    .io_a(inst_SnxnLv3Inst9_io_a),
    .io_b(inst_SnxnLv3Inst9_io_b),
    .io_z(inst_SnxnLv3Inst9_io_z)
  );
  SnxnLv3Inst10 inst_SnxnLv3Inst10 ( // @[Snxn100k.scala 7106:34]
    .io_a(inst_SnxnLv3Inst10_io_a),
    .io_b(inst_SnxnLv3Inst10_io_b),
    .io_z(inst_SnxnLv3Inst10_io_z)
  );
  SnxnLv3Inst11 inst_SnxnLv3Inst11 ( // @[Snxn100k.scala 7110:34]
    .io_a(inst_SnxnLv3Inst11_io_a),
    .io_b(inst_SnxnLv3Inst11_io_b),
    .io_z(inst_SnxnLv3Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7115:15]
  assign inst_SnxnLv3Inst8_io_a = io_a; // @[Snxn100k.scala 7099:26]
  assign inst_SnxnLv3Inst8_io_b = io_b; // @[Snxn100k.scala 7100:26]
  assign inst_SnxnLv3Inst9_io_a = io_a; // @[Snxn100k.scala 7103:26]
  assign inst_SnxnLv3Inst9_io_b = io_b; // @[Snxn100k.scala 7104:26]
  assign inst_SnxnLv3Inst10_io_a = io_a; // @[Snxn100k.scala 7107:27]
  assign inst_SnxnLv3Inst10_io_b = io_b; // @[Snxn100k.scala 7108:27]
  assign inst_SnxnLv3Inst11_io_a = io_a; // @[Snxn100k.scala 7111:27]
  assign inst_SnxnLv3Inst11_io_b = io_b; // @[Snxn100k.scala 7112:27]
endmodule
module SnxnLv4Inst48(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 67397:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 67398:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 67399:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 67400:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 67401:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 67402:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 67403:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 67404:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 67405:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 67406:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 67407:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 67408:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 67409:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 67410:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 67411:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 67412:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 67413:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 67414:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 67415:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 67416:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 67417:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 67418:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 67419:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 67420:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 67421:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 67422:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 67423:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 67424:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 67425:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 67426:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 67427:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 67428:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 67429:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 67430:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 67431:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 67432:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 67433:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 67434:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 67435:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 67436:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 67437:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 67438:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 67439:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 67440:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 67441:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 67442:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 67443:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 67444:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 67445:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 67446:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 67447:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 67448:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 67449:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 67450:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 67451:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 67452:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 67453:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 67454:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 67455:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 67456:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 67457:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 67458:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 67459:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 67460:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 67461:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 67462:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 67463:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 67464:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 67465:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 67466:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 67467:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 67468:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 67469:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 67470:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 67471:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 67472:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 67473:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 67474:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 67475:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 67476:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 67477:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 67478:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 67479:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 67480:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 67481:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 67482:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 67483:20]
  assign io_z = ~x21; // @[Snxn100k.scala 67484:16]
endmodule
module SnxnLv4Inst49(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 66843:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 66844:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 66845:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 66846:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 66847:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 66848:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 66849:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 66850:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 66851:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 66852:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 66853:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 66854:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 66855:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 66856:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 66857:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 66858:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 66859:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 66860:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 66861:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 66862:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 66863:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 66864:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 66865:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 66866:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 66867:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 66868:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 66869:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 66870:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 66871:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 66872:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 66873:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 66874:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 66875:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 66876:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 66877:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 66878:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 66879:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 66880:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 66881:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 66882:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 66883:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 66884:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 66885:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 66886:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 66887:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 66888:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 66889:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 66890:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 66891:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 66892:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 66893:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 66894:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 66895:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 66896:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 66897:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 66898:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 66899:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 66900:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 66901:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 66902:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 66903:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 66904:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 66905:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 66906:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 66907:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 66908:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 66909:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 66910:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 66911:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 66912:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 66913:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 66914:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 66915:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 66916:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 66917:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 66918:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 66919:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 66920:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 66921:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 66922:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 66923:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 66924:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 66925:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 66926:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 66927:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 66928:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 66929:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 66930:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 66931:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 66932:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 66933:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 66934:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 66935:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 66936:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 66937:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 66938:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 66939:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 66940:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 66941:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 66942:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 66943:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 66944:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 66945:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 66946:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 66947:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 66948:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 66949:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 66950:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 66951:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 66952:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 66953:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 66954:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 66955:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 66956:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 66957:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 66958:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 66959:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 66960:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 66961:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 66962:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 66963:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 66964:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 66965:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 66966:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 66967:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 66968:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 66969:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 66970:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 66971:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 66972:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 66973:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 66974:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 66975:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 66976:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 66977:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 66978:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 66979:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 66980:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 66981:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 66982:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 66983:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 66984:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 66985:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 66986:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 66987:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 66988:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 66989:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 66990:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 66991:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 66992:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 66993:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 66994:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 66995:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 66996:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 66997:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 66998:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 66999:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 67000:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 67001:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 67002:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 67003:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 67004:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 67005:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 67006:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 67007:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 67008:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 67009:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 67010:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 67011:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 67012:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 67013:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 67014:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 67015:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 67016:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 67017:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 67018:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 67019:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 67020:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 67021:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 67022:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 67023:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 67024:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 67025:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 67026:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 67027:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 67028:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 67029:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 67030:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 67031:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 67032:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 67033:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 67034:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 67035:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 67036:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 67037:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 67038:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 67039:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 67040:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 67041:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 67042:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 67043:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 67044:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 67045:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 67046:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 67047:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 67048:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 67049:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 67050:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 67051:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 67052:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 67053:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 67054:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 67055:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 67056:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 67057:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 67058:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 67059:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 67060:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 67061:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 67062:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 67063:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 67064:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 67065:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 67066:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 67067:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 67068:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 67069:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 67070:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 67071:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 67072:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 67073:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 67074:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 67075:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 67076:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 67077:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 67078:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 67079:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 67080:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 67081:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 67082:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 67083:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 67084:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 67085:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 67086:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 67087:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 67088:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 67089:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 67090:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 67091:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 67092:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 67093:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 67094:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 67095:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 67096:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 67097:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 67098:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 67099:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 67100:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 67101:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 67102:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 67103:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 67104:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 67105:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 67106:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 67107:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 67108:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 67109:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 67110:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 67111:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 67112:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 67113:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 67114:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 67115:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 67116:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 67117:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 67118:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 67119:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 67120:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 67121:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 67122:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 67123:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 67124:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 67125:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 67126:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 67127:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 67128:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 67129:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 67130:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 67131:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 67132:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 67133:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 67134:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 67135:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 67136:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 67137:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 67138:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 67139:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 67140:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 67141:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 67142:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 67143:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 67144:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 67145:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 67146:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 67147:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 67148:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 67149:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 67150:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 67151:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 67152:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 67153:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 67154:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 67155:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 67156:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 67157:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 67158:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 67159:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 67160:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 67161:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 67162:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 67163:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 67164:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 67165:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 67166:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 67167:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 67168:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 67169:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 67170:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 67171:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 67172:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 67173:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 67174:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 67175:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 67176:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 67177:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 67178:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 67179:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 67180:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 67181:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 67182:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 67183:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 67184:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 67185:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 67186:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 67187:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 67188:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 67189:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 67190:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 67191:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 67192:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 67193:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 67194:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 67195:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 67196:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 67197:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 67198:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 67199:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 67200:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 67201:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 67202:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 67203:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 67204:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 67205:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 67206:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 67207:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 67208:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 67209:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 67210:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 67211:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 67212:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 67213:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 67214:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 67215:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 67216:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 67217:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 67218:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 67219:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 67220:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 67221:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 67222:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 67223:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 67224:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 67225:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 67226:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 67227:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 67228:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 67229:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 67230:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 67231:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 67232:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 67233:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 67234:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 67235:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 67236:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 67237:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 67238:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 67239:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 67240:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 67241:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 67242:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 67243:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 67244:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 67245:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 67246:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 67247:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 67248:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 67249:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 67250:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 67251:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 67252:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 67253:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 67254:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 67255:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 67256:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 67257:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 67258:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 67259:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 67260:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 67261:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 67262:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 67263:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 67264:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 67265:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 67266:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 67267:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 67268:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 67269:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 67270:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 67271:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 67272:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 67273:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 67274:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 67275:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 67276:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 67277:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 67278:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 67279:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 67280:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 67281:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 67282:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 67283:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 67284:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 67285:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 67286:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 67287:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 67288:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 67289:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 67290:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 67291:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 67292:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 67293:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 67294:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 67295:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 67296:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 67297:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 67298:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 67299:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 67300:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 67301:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 67302:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 67303:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 67304:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 67305:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 67306:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 67307:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 67308:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 67309:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 67310:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 67311:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 67312:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 67313:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 67314:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 67315:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 67316:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 67317:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 67318:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 67319:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 67320:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 67321:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 67322:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 67323:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 67324:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 67325:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 67326:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 67327:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 67328:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 67329:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 67330:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 67331:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 67332:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 67333:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 67334:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 67335:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 67336:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 67337:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 67338:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 67339:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 67340:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 67341:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 67342:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 67343:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 67344:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 67345:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 67346:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 67347:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 67348:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 67349:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 67350:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 67351:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 67352:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 67353:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 67354:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 67355:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 67356:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 67357:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 67358:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 67359:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 67360:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 67361:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 67362:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 67363:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 67364:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 67365:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 67366:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 67367:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 67368:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 67369:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 67370:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 67371:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 67372:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 67373:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 67374:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 67375:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 67376:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 67377:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 67378:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 67379:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 67380:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 67381:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 67382:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 67383:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 67384:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 67385:22]
  assign io_z = ~x135; // @[Snxn100k.scala 67386:17]
endmodule
module SnxnLv4Inst51(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 66329:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 66330:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 66331:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 66332:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 66333:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 66334:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 66335:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 66336:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 66337:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 66338:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 66339:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 66340:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 66341:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 66342:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 66343:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 66344:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 66345:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 66346:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 66347:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 66348:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 66349:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 66350:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 66351:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 66352:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 66353:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 66354:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 66355:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 66356:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 66357:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 66358:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 66359:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 66360:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 66361:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 66362:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 66363:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 66364:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 66365:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 66366:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 66367:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 66368:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 66369:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 66370:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 66371:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 66372:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 66373:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 66374:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 66375:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 66376:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 66377:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 66378:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 66379:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 66380:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 66381:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 66382:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 66383:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 66384:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 66385:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 66386:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 66387:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 66388:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 66389:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 66390:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 66391:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 66392:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 66393:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 66394:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 66395:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 66396:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 66397:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 66398:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 66399:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 66400:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 66401:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 66402:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 66403:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 66404:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 66405:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 66406:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 66407:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 66408:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 66409:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 66410:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 66411:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 66412:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 66413:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 66414:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 66415:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 66416:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 66417:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 66418:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 66419:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 66420:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 66421:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 66422:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 66423:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 66424:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 66425:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 66426:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 66427:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 66428:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 66429:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 66430:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 66431:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 66432:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 66433:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 66434:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 66435:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 66436:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 66437:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 66438:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 66439:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 66440:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 66441:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 66442:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 66443:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 66444:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 66445:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 66446:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 66447:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 66448:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 66449:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 66450:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 66451:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 66452:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 66453:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 66454:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 66455:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 66456:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 66457:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 66458:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 66459:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 66460:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 66461:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 66462:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 66463:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 66464:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 66465:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 66466:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 66467:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 66468:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 66469:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 66470:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 66471:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 66472:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 66473:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 66474:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 66475:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 66476:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 66477:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 66478:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 66479:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 66480:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 66481:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 66482:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 66483:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 66484:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 66485:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 66486:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 66487:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 66488:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 66489:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 66490:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 66491:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 66492:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 66493:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 66494:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 66495:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 66496:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 66497:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 66498:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 66499:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 66500:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 66501:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 66502:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 66503:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 66504:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 66505:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 66506:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 66507:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 66508:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 66509:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 66510:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 66511:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 66512:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 66513:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 66514:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 66515:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 66516:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 66517:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 66518:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 66519:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 66520:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 66521:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 66522:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 66523:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 66524:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 66525:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 66526:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 66527:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 66528:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 66529:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 66530:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 66531:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 66532:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 66533:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 66534:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 66535:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 66536:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 66537:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 66538:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 66539:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 66540:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 66541:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 66542:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 66543:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 66544:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 66545:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 66546:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 66547:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 66548:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 66549:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 66550:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 66551:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 66552:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 66553:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 66554:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 66555:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 66556:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 66557:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 66558:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 66559:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 66560:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 66561:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 66562:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 66563:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 66564:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 66565:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 66566:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 66567:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 66568:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 66569:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 66570:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 66571:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 66572:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 66573:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 66574:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 66575:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 66576:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 66577:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 66578:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 66579:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 66580:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 66581:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 66582:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 66583:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 66584:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 66585:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 66586:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 66587:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 66588:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 66589:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 66590:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 66591:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 66592:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 66593:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 66594:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 66595:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 66596:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 66597:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 66598:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 66599:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 66600:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 66601:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 66602:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 66603:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 66604:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 66605:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 66606:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 66607:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 66608:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 66609:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 66610:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 66611:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 66612:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 66613:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 66614:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 66615:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 66616:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 66617:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 66618:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 66619:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 66620:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 66621:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 66622:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 66623:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 66624:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 66625:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 66626:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 66627:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 66628:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 66629:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 66630:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 66631:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 66632:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 66633:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 66634:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 66635:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 66636:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 66637:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 66638:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 66639:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 66640:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 66641:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 66642:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 66643:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 66644:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 66645:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 66646:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 66647:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 66648:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 66649:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 66650:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 66651:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 66652:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 66653:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 66654:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 66655:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 66656:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 66657:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 66658:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 66659:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 66660:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 66661:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 66662:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 66663:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 66664:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 66665:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 66666:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 66667:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 66668:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 66669:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 66670:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 66671:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 66672:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 66673:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 66674:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 66675:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 66676:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 66677:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 66678:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 66679:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 66680:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 66681:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 66682:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 66683:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 66684:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 66685:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 66686:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 66687:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 66688:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 66689:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 66690:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 66691:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 66692:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 66693:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 66694:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 66695:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 66696:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 66697:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 66698:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 66699:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 66700:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 66701:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 66702:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 66703:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 66704:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 66705:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 66706:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 66707:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 66708:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 66709:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 66710:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 66711:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 66712:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 66713:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 66714:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 66715:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 66716:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 66717:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 66718:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 66719:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 66720:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 66721:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 66722:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 66723:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 66724:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 66725:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 66726:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 66727:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 66728:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 66729:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 66730:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 66731:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 66732:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 66733:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 66734:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 66735:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 66736:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 66737:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 66738:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 66739:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 66740:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 66741:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 66742:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 66743:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 66744:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 66745:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 66746:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 66747:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 66748:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 66749:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 66750:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 66751:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 66752:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 66753:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 66754:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 66755:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 66756:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 66757:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 66758:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 66759:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 66760:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 66761:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 66762:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 66763:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 66764:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 66765:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 66766:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 66767:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 66768:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 66769:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 66770:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 66771:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 66772:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 66773:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 66774:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 66775:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 66776:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 66777:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 66778:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 66779:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 66780:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 66781:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 66782:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 66783:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 66784:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 66785:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 66786:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 66787:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 66788:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 66789:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 66790:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 66791:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 66792:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 66793:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 66794:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 66795:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 66796:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 66797:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 66798:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 66799:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 66800:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 66801:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 66802:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 66803:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 66804:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 66805:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 66806:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 66807:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 66808:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 66809:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 66810:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 66811:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 66812:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 66813:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 66814:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 66815:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 66816:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 66817:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 66818:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 66819:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 66820:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 66821:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 66822:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 66823:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 66824:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 66825:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 66826:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 66827:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 66828:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 66829:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 66830:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 66831:22]
  assign io_z = ~x125; // @[Snxn100k.scala 66832:17]
endmodule
module SnxnLv3Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst48_io_a; // @[Snxn100k.scala 21552:34]
  wire  inst_SnxnLv4Inst48_io_b; // @[Snxn100k.scala 21552:34]
  wire  inst_SnxnLv4Inst48_io_z; // @[Snxn100k.scala 21552:34]
  wire  inst_SnxnLv4Inst49_io_a; // @[Snxn100k.scala 21556:34]
  wire  inst_SnxnLv4Inst49_io_b; // @[Snxn100k.scala 21556:34]
  wire  inst_SnxnLv4Inst49_io_z; // @[Snxn100k.scala 21556:34]
  wire  inst_SnxnLv4Inst50_io_a; // @[Snxn100k.scala 21560:34]
  wire  inst_SnxnLv4Inst50_io_b; // @[Snxn100k.scala 21560:34]
  wire  inst_SnxnLv4Inst50_io_z; // @[Snxn100k.scala 21560:34]
  wire  inst_SnxnLv4Inst51_io_a; // @[Snxn100k.scala 21564:34]
  wire  inst_SnxnLv4Inst51_io_b; // @[Snxn100k.scala 21564:34]
  wire  inst_SnxnLv4Inst51_io_z; // @[Snxn100k.scala 21564:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst48_io_z + inst_SnxnLv4Inst49_io_z; // @[Snxn100k.scala 21568:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst50_io_z; // @[Snxn100k.scala 21568:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst51_io_z; // @[Snxn100k.scala 21568:89]
  SnxnLv4Inst48 inst_SnxnLv4Inst48 ( // @[Snxn100k.scala 21552:34]
    .io_a(inst_SnxnLv4Inst48_io_a),
    .io_b(inst_SnxnLv4Inst48_io_b),
    .io_z(inst_SnxnLv4Inst48_io_z)
  );
  SnxnLv4Inst49 inst_SnxnLv4Inst49 ( // @[Snxn100k.scala 21556:34]
    .io_a(inst_SnxnLv4Inst49_io_a),
    .io_b(inst_SnxnLv4Inst49_io_b),
    .io_z(inst_SnxnLv4Inst49_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst50 ( // @[Snxn100k.scala 21560:34]
    .io_a(inst_SnxnLv4Inst50_io_a),
    .io_b(inst_SnxnLv4Inst50_io_b),
    .io_z(inst_SnxnLv4Inst50_io_z)
  );
  SnxnLv4Inst51 inst_SnxnLv4Inst51 ( // @[Snxn100k.scala 21564:34]
    .io_a(inst_SnxnLv4Inst51_io_a),
    .io_b(inst_SnxnLv4Inst51_io_b),
    .io_z(inst_SnxnLv4Inst51_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21569:15]
  assign inst_SnxnLv4Inst48_io_a = io_a; // @[Snxn100k.scala 21553:27]
  assign inst_SnxnLv4Inst48_io_b = io_b; // @[Snxn100k.scala 21554:27]
  assign inst_SnxnLv4Inst49_io_a = io_a; // @[Snxn100k.scala 21557:27]
  assign inst_SnxnLv4Inst49_io_b = io_b; // @[Snxn100k.scala 21558:27]
  assign inst_SnxnLv4Inst50_io_a = io_a; // @[Snxn100k.scala 21561:27]
  assign inst_SnxnLv4Inst50_io_b = io_b; // @[Snxn100k.scala 21562:27]
  assign inst_SnxnLv4Inst51_io_a = io_a; // @[Snxn100k.scala 21565:27]
  assign inst_SnxnLv4Inst51_io_b = io_b; // @[Snxn100k.scala 21566:27]
endmodule
module SnxnLv4Inst52(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 65159:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 65160:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 65161:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 65162:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 65163:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 65164:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 65165:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 65166:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 65167:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 65168:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 65169:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 65170:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 65171:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 65172:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 65173:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 65174:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 65175:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 65176:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 65177:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 65178:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 65179:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 65180:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 65181:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 65182:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 65183:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 65184:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 65185:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 65186:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 65187:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 65188:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 65189:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 65190:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 65191:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 65192:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 65193:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 65194:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 65195:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 65196:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 65197:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 65198:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 65199:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 65200:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 65201:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 65202:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 65203:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 65204:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 65205:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 65206:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 65207:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 65208:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 65209:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 65210:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 65211:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 65212:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 65213:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 65214:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 65215:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 65216:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 65217:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 65218:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 65219:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 65220:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 65221:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 65222:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 65223:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 65224:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 65225:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 65226:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 65227:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 65228:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 65229:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 65230:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 65231:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 65232:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 65233:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 65234:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 65235:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 65236:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 65237:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 65238:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 65239:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 65240:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 65241:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 65242:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 65243:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 65244:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 65245:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 65246:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 65247:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 65248:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 65249:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 65250:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 65251:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 65252:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 65253:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 65254:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 65255:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 65256:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 65257:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 65258:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 65259:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 65260:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 65261:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 65262:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 65263:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 65264:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 65265:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 65266:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 65267:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 65268:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 65269:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 65270:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 65271:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 65272:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 65273:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 65274:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 65275:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 65276:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 65277:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 65278:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 65279:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 65280:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 65281:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 65282:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 65283:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 65284:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 65285:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 65286:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 65287:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 65288:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 65289:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 65290:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 65291:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 65292:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 65293:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 65294:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 65295:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 65296:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 65297:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 65298:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 65299:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 65300:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 65301:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 65302:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 65303:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 65304:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 65305:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 65306:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 65307:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 65308:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 65309:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 65310:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 65311:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 65312:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 65313:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 65314:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 65315:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 65316:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 65317:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 65318:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 65319:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 65320:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 65321:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 65322:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 65323:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 65324:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 65325:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 65326:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 65327:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 65328:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 65329:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 65330:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 65331:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 65332:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 65333:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 65334:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 65335:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 65336:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 65337:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 65338:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 65339:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 65340:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 65341:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 65342:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 65343:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 65344:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 65345:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 65346:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 65347:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 65348:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 65349:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 65350:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 65351:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 65352:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 65353:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 65354:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 65355:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 65356:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 65357:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 65358:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 65359:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 65360:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 65361:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 65362:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 65363:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 65364:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 65365:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 65366:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 65367:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 65368:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 65369:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 65370:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 65371:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 65372:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 65373:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 65374:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 65375:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 65376:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 65377:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 65378:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 65379:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 65380:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 65381:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 65382:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 65383:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 65384:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 65385:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 65386:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 65387:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 65388:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 65389:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 65390:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 65391:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 65392:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 65393:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 65394:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 65395:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 65396:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 65397:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 65398:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 65399:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 65400:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 65401:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 65402:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 65403:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 65404:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 65405:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 65406:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 65407:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 65408:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 65409:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 65410:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 65411:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 65412:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 65413:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 65414:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 65415:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 65416:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 65417:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 65418:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 65419:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 65420:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 65421:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 65422:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 65423:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 65424:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 65425:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 65426:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 65427:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 65428:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 65429:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 65430:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 65431:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 65432:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 65433:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 65434:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 65435:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 65436:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 65437:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 65438:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 65439:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 65440:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 65441:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 65442:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 65443:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 65444:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 65445:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 65446:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 65447:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 65448:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 65449:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 65450:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 65451:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 65452:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 65453:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 65454:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 65455:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 65456:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 65457:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 65458:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 65459:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 65460:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 65461:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 65462:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 65463:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 65464:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 65465:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 65466:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 65467:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 65468:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 65469:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 65470:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 65471:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 65472:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 65473:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 65474:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 65475:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 65476:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 65477:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 65478:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 65479:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 65480:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 65481:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 65482:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 65483:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 65484:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 65485:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 65486:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 65487:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 65488:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 65489:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 65490:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 65491:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 65492:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 65493:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 65494:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 65495:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 65496:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 65497:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 65498:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 65499:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 65500:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 65501:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 65502:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 65503:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 65504:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 65505:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 65506:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 65507:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 65508:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 65509:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 65510:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 65511:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 65512:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 65513:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 65514:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 65515:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 65516:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 65517:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 65518:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 65519:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 65520:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 65521:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 65522:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 65523:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 65524:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 65525:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 65526:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 65527:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 65528:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 65529:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 65530:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 65531:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 65532:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 65533:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 65534:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 65535:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 65536:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 65537:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 65538:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 65539:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 65540:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 65541:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 65542:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 65543:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 65544:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 65545:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 65546:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 65547:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 65548:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 65549:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 65550:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 65551:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 65552:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 65553:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 65554:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 65555:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 65556:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 65557:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 65558:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 65559:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 65560:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 65561:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 65562:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 65563:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 65564:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 65565:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 65566:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 65567:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 65568:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 65569:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 65570:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 65571:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 65572:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 65573:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 65574:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 65575:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 65576:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 65577:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 65578:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 65579:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 65580:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 65581:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 65582:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 65583:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 65584:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 65585:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 65586:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 65587:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 65588:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 65589:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 65590:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 65591:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 65592:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 65593:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 65594:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 65595:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 65596:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 65597:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 65598:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 65599:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 65600:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 65601:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 65602:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 65603:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 65604:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 65605:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 65606:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 65607:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 65608:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 65609:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 65610:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 65611:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 65612:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 65613:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 65614:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 65615:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 65616:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 65617:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 65618:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 65619:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 65620:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 65621:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 65622:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 65623:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 65624:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 65625:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 65626:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 65627:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 65628:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 65629:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 65630:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 65631:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 65632:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 65633:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 65634:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 65635:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 65636:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 65637:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 65638:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 65639:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 65640:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 65641:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 65642:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 65643:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 65644:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 65645:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 65646:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 65647:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 65648:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 65649:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 65650:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 65651:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 65652:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 65653:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 65654:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 65655:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 65656:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 65657:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 65658:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 65659:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 65660:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 65661:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 65662:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 65663:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 65664:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 65665:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 65666:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 65667:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 65668:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 65669:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 65670:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 65671:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 65672:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 65673:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 65674:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 65675:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 65676:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 65677:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 65678:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 65679:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 65680:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 65681:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 65682:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 65683:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 65684:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 65685:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 65686:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 65687:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 65688:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 65689:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 65690:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 65691:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 65692:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 65693:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 65694:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 65695:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 65696:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 65697:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 65698:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 65699:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 65700:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 65701:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 65702:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 65703:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 65704:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 65705:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 65706:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 65707:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 65708:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 65709:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 65710:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 65711:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 65712:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 65713:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 65714:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 65715:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 65716:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 65717:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 65718:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 65719:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 65720:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 65721:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 65722:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 65723:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 65724:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 65725:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 65726:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 65727:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 65728:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 65729:22]
  wire  invx142 = ~x142; // @[Snxn100k.scala 65730:17]
  wire  t143 = x142 + invx142; // @[Snxn100k.scala 65731:22]
  wire  inv143 = ~t143; // @[Snxn100k.scala 65732:17]
  wire  x143 = t143 ^ inv143; // @[Snxn100k.scala 65733:22]
  wire  invx143 = ~x143; // @[Snxn100k.scala 65734:17]
  wire  t144 = x143 + invx143; // @[Snxn100k.scala 65735:22]
  wire  inv144 = ~t144; // @[Snxn100k.scala 65736:17]
  wire  x144 = t144 ^ inv144; // @[Snxn100k.scala 65737:22]
  assign io_z = ~x144; // @[Snxn100k.scala 65738:17]
endmodule
module SnxnLv4Inst54(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 64725:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 64726:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 64727:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 64728:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 64729:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 64730:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 64731:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 64732:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 64733:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 64734:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 64735:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 64736:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 64737:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 64738:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 64739:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 64740:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 64741:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 64742:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 64743:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 64744:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 64745:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 64746:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 64747:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 64748:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 64749:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 64750:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 64751:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 64752:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 64753:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 64754:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 64755:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 64756:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 64757:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 64758:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 64759:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 64760:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 64761:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 64762:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 64763:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 64764:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 64765:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 64766:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 64767:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 64768:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 64769:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 64770:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 64771:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 64772:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 64773:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 64774:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 64775:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 64776:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 64777:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 64778:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 64779:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 64780:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 64781:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 64782:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 64783:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 64784:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 64785:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 64786:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 64787:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 64788:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 64789:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 64790:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 64791:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 64792:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 64793:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 64794:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 64795:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 64796:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 64797:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 64798:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 64799:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 64800:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 64801:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 64802:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 64803:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 64804:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 64805:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 64806:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 64807:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 64808:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 64809:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 64810:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 64811:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 64812:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 64813:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 64814:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 64815:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 64816:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 64817:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 64818:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 64819:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 64820:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 64821:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 64822:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 64823:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 64824:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 64825:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 64826:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 64827:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 64828:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 64829:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 64830:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 64831:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 64832:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 64833:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 64834:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 64835:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 64836:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 64837:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 64838:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 64839:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 64840:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 64841:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 64842:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 64843:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 64844:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 64845:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 64846:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 64847:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 64848:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 64849:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 64850:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 64851:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 64852:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 64853:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 64854:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 64855:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 64856:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 64857:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 64858:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 64859:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 64860:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 64861:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 64862:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 64863:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 64864:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 64865:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 64866:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 64867:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 64868:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 64869:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 64870:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 64871:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 64872:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 64873:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 64874:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 64875:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 64876:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 64877:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 64878:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 64879:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 64880:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 64881:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 64882:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 64883:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 64884:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 64885:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 64886:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 64887:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 64888:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 64889:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 64890:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 64891:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 64892:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 64893:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 64894:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 64895:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 64896:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 64897:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 64898:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 64899:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 64900:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 64901:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 64902:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 64903:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 64904:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 64905:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 64906:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 64907:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 64908:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 64909:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 64910:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 64911:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 64912:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 64913:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 64914:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 64915:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 64916:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 64917:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 64918:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 64919:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 64920:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 64921:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 64922:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 64923:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 64924:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 64925:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 64926:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 64927:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 64928:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 64929:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 64930:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 64931:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 64932:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 64933:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 64934:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 64935:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 64936:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 64937:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 64938:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 64939:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 64940:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 64941:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 64942:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 64943:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 64944:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 64945:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 64946:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 64947:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 64948:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 64949:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 64950:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 64951:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 64952:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 64953:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 64954:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 64955:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 64956:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 64957:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 64958:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 64959:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 64960:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 64961:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 64962:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 64963:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 64964:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 64965:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 64966:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 64967:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 64968:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 64969:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 64970:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 64971:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 64972:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 64973:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 64974:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 64975:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 64976:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 64977:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 64978:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 64979:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 64980:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 64981:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 64982:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 64983:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 64984:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 64985:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 64986:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 64987:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 64988:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 64989:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 64990:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 64991:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 64992:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 64993:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 64994:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 64995:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 64996:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 64997:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 64998:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 64999:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 65000:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 65001:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 65002:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 65003:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 65004:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 65005:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 65006:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 65007:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 65008:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 65009:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 65010:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 65011:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 65012:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 65013:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 65014:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 65015:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 65016:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 65017:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 65018:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 65019:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 65020:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 65021:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 65022:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 65023:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 65024:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 65025:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 65026:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 65027:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 65028:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 65029:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 65030:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 65031:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 65032:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 65033:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 65034:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 65035:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 65036:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 65037:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 65038:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 65039:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 65040:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 65041:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 65042:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 65043:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 65044:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 65045:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 65046:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 65047:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 65048:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 65049:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 65050:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 65051:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 65052:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 65053:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 65054:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 65055:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 65056:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 65057:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 65058:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 65059:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 65060:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 65061:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 65062:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 65063:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 65064:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 65065:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 65066:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 65067:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 65068:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 65069:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 65070:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 65071:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 65072:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 65073:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 65074:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 65075:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 65076:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 65077:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 65078:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 65079:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 65080:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 65081:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 65082:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 65083:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 65084:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 65085:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 65086:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 65087:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 65088:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 65089:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 65090:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 65091:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 65092:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 65093:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 65094:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 65095:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 65096:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 65097:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 65098:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 65099:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 65100:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 65101:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 65102:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 65103:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 65104:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 65105:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 65106:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 65107:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 65108:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 65109:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 65110:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 65111:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 65112:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 65113:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 65114:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 65115:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 65116:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 65117:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 65118:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 65119:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 65120:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 65121:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 65122:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 65123:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 65124:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 65125:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 65126:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 65127:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 65128:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 65129:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 65130:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 65131:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 65132:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 65133:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 65134:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 65135:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 65136:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 65137:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 65138:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 65139:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 65140:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 65141:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 65142:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 65143:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 65144:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 65145:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 65146:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 65147:22]
  assign io_z = ~x105; // @[Snxn100k.scala 65148:17]
endmodule
module SnxnLv4Inst55(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 65749:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 65750:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 65751:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 65752:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 65753:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 65754:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 65755:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 65756:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 65757:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 65758:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 65759:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 65760:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 65761:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 65762:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 65763:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 65764:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 65765:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 65766:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 65767:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 65768:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 65769:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 65770:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 65771:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 65772:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 65773:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 65774:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 65775:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 65776:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 65777:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 65778:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 65779:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 65780:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 65781:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 65782:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 65783:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 65784:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 65785:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 65786:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 65787:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 65788:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 65789:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 65790:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 65791:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 65792:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 65793:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 65794:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 65795:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 65796:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 65797:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 65798:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 65799:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 65800:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 65801:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 65802:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 65803:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 65804:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 65805:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 65806:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 65807:20]
  assign io_z = ~x14; // @[Snxn100k.scala 65808:16]
endmodule
module SnxnLv3Inst13(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst52_io_a; // @[Snxn100k.scala 21269:34]
  wire  inst_SnxnLv4Inst52_io_b; // @[Snxn100k.scala 21269:34]
  wire  inst_SnxnLv4Inst52_io_z; // @[Snxn100k.scala 21269:34]
  wire  inst_SnxnLv4Inst53_io_a; // @[Snxn100k.scala 21273:34]
  wire  inst_SnxnLv4Inst53_io_b; // @[Snxn100k.scala 21273:34]
  wire  inst_SnxnLv4Inst53_io_z; // @[Snxn100k.scala 21273:34]
  wire  inst_SnxnLv4Inst54_io_a; // @[Snxn100k.scala 21277:34]
  wire  inst_SnxnLv4Inst54_io_b; // @[Snxn100k.scala 21277:34]
  wire  inst_SnxnLv4Inst54_io_z; // @[Snxn100k.scala 21277:34]
  wire  inst_SnxnLv4Inst55_io_a; // @[Snxn100k.scala 21281:34]
  wire  inst_SnxnLv4Inst55_io_b; // @[Snxn100k.scala 21281:34]
  wire  inst_SnxnLv4Inst55_io_z; // @[Snxn100k.scala 21281:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst52_io_z + inst_SnxnLv4Inst53_io_z; // @[Snxn100k.scala 21285:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst54_io_z; // @[Snxn100k.scala 21285:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst55_io_z; // @[Snxn100k.scala 21285:89]
  SnxnLv4Inst52 inst_SnxnLv4Inst52 ( // @[Snxn100k.scala 21269:34]
    .io_a(inst_SnxnLv4Inst52_io_a),
    .io_b(inst_SnxnLv4Inst52_io_b),
    .io_z(inst_SnxnLv4Inst52_io_z)
  );
  SnxnLv4Inst38 inst_SnxnLv4Inst53 ( // @[Snxn100k.scala 21273:34]
    .io_a(inst_SnxnLv4Inst53_io_a),
    .io_b(inst_SnxnLv4Inst53_io_b),
    .io_z(inst_SnxnLv4Inst53_io_z)
  );
  SnxnLv4Inst54 inst_SnxnLv4Inst54 ( // @[Snxn100k.scala 21277:34]
    .io_a(inst_SnxnLv4Inst54_io_a),
    .io_b(inst_SnxnLv4Inst54_io_b),
    .io_z(inst_SnxnLv4Inst54_io_z)
  );
  SnxnLv4Inst55 inst_SnxnLv4Inst55 ( // @[Snxn100k.scala 21281:34]
    .io_a(inst_SnxnLv4Inst55_io_a),
    .io_b(inst_SnxnLv4Inst55_io_b),
    .io_z(inst_SnxnLv4Inst55_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21286:15]
  assign inst_SnxnLv4Inst52_io_a = io_a; // @[Snxn100k.scala 21270:27]
  assign inst_SnxnLv4Inst52_io_b = io_b; // @[Snxn100k.scala 21271:27]
  assign inst_SnxnLv4Inst53_io_a = io_a; // @[Snxn100k.scala 21274:27]
  assign inst_SnxnLv4Inst53_io_b = io_b; // @[Snxn100k.scala 21275:27]
  assign inst_SnxnLv4Inst54_io_a = io_a; // @[Snxn100k.scala 21278:27]
  assign inst_SnxnLv4Inst54_io_b = io_b; // @[Snxn100k.scala 21279:27]
  assign inst_SnxnLv4Inst55_io_a = io_a; // @[Snxn100k.scala 21282:27]
  assign inst_SnxnLv4Inst55_io_b = io_b; // @[Snxn100k.scala 21283:27]
endmodule
module SnxnLv4Inst56(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 63383:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 63384:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 63385:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 63386:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 63387:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 63388:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 63389:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 63390:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 63391:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 63392:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 63393:18]
  assign io_z = ~x2; // @[Snxn100k.scala 63394:15]
endmodule
module SnxnLv4Inst58(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 64013:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 64014:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 64015:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 64016:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 64017:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 64018:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 64019:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 64020:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 64021:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 64022:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 64023:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 64024:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 64025:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 64026:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 64027:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 64028:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 64029:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 64030:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 64031:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 64032:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 64033:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 64034:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 64035:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 64036:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 64037:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 64038:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 64039:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 64040:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 64041:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 64042:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 64043:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 64044:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 64045:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 64046:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 64047:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 64048:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 64049:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 64050:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 64051:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 64052:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 64053:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 64054:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 64055:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 64056:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 64057:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 64058:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 64059:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 64060:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 64061:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 64062:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 64063:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 64064:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 64065:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 64066:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 64067:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 64068:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 64069:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 64070:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 64071:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 64072:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 64073:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 64074:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 64075:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 64076:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 64077:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 64078:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 64079:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 64080:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 64081:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 64082:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 64083:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 64084:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 64085:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 64086:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 64087:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 64088:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 64089:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 64090:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 64091:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 64092:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 64093:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 64094:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 64095:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 64096:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 64097:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 64098:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 64099:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 64100:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 64101:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 64102:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 64103:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 64104:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 64105:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 64106:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 64107:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 64108:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 64109:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 64110:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 64111:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 64112:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 64113:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 64114:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 64115:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 64116:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 64117:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 64118:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 64119:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 64120:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 64121:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 64122:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 64123:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 64124:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 64125:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 64126:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 64127:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 64128:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 64129:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 64130:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 64131:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 64132:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 64133:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 64134:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 64135:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 64136:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 64137:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 64138:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 64139:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 64140:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 64141:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 64142:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 64143:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 64144:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 64145:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 64146:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 64147:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 64148:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 64149:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 64150:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 64151:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 64152:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 64153:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 64154:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 64155:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 64156:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 64157:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 64158:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 64159:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 64160:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 64161:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 64162:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 64163:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 64164:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 64165:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 64166:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 64167:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 64168:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 64169:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 64170:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 64171:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 64172:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 64173:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 64174:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 64175:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 64176:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 64177:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 64178:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 64179:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 64180:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 64181:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 64182:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 64183:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 64184:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 64185:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 64186:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 64187:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 64188:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 64189:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 64190:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 64191:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 64192:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 64193:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 64194:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 64195:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 64196:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 64197:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 64198:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 64199:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 64200:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 64201:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 64202:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 64203:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 64204:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 64205:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 64206:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 64207:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 64208:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 64209:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 64210:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 64211:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 64212:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 64213:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 64214:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 64215:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 64216:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 64217:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 64218:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 64219:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 64220:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 64221:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 64222:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 64223:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 64224:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 64225:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 64226:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 64227:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 64228:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 64229:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 64230:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 64231:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 64232:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 64233:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 64234:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 64235:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 64236:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 64237:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 64238:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 64239:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 64240:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 64241:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 64242:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 64243:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 64244:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 64245:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 64246:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 64247:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 64248:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 64249:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 64250:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 64251:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 64252:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 64253:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 64254:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 64255:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 64256:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 64257:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 64258:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 64259:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 64260:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 64261:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 64262:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 64263:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 64264:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 64265:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 64266:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 64267:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 64268:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 64269:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 64270:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 64271:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 64272:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 64273:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 64274:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 64275:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 64276:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 64277:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 64278:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 64279:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 64280:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 64281:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 64282:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 64283:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 64284:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 64285:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 64286:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 64287:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 64288:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 64289:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 64290:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 64291:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 64292:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 64293:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 64294:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 64295:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 64296:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 64297:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 64298:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 64299:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 64300:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 64301:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 64302:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 64303:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 64304:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 64305:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 64306:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 64307:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 64308:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 64309:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 64310:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 64311:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 64312:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 64313:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 64314:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 64315:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 64316:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 64317:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 64318:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 64319:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 64320:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 64321:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 64322:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 64323:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 64324:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 64325:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 64326:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 64327:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 64328:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 64329:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 64330:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 64331:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 64332:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 64333:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 64334:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 64335:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 64336:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 64337:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 64338:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 64339:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 64340:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 64341:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 64342:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 64343:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 64344:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 64345:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 64346:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 64347:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 64348:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 64349:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 64350:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 64351:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 64352:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 64353:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 64354:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 64355:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 64356:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 64357:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 64358:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 64359:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 64360:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 64361:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 64362:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 64363:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 64364:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 64365:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 64366:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 64367:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 64368:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 64369:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 64370:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 64371:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 64372:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 64373:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 64374:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 64375:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 64376:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 64377:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 64378:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 64379:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 64380:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 64381:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 64382:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 64383:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 64384:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 64385:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 64386:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 64387:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 64388:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 64389:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 64390:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 64391:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 64392:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 64393:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 64394:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 64395:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 64396:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 64397:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 64398:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 64399:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 64400:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 64401:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 64402:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 64403:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 64404:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 64405:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 64406:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 64407:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 64408:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 64409:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 64410:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 64411:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 64412:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 64413:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 64414:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 64415:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 64416:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 64417:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 64418:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 64419:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 64420:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 64421:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 64422:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 64423:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 64424:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 64425:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 64426:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 64427:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 64428:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 64429:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 64430:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 64431:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 64432:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 64433:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 64434:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 64435:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 64436:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 64437:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 64438:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 64439:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 64440:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 64441:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 64442:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 64443:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 64444:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 64445:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 64446:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 64447:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 64448:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 64449:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 64450:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 64451:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 64452:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 64453:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 64454:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 64455:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 64456:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 64457:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 64458:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 64459:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 64460:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 64461:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 64462:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 64463:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 64464:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 64465:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 64466:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 64467:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 64468:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 64469:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 64470:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 64471:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 64472:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 64473:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 64474:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 64475:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 64476:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 64477:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 64478:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 64479:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 64480:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 64481:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 64482:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 64483:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 64484:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 64485:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 64486:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 64487:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 64488:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 64489:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 64490:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 64491:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 64492:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 64493:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 64494:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 64495:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 64496:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 64497:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 64498:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 64499:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 64500:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 64501:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 64502:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 64503:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 64504:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 64505:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 64506:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 64507:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 64508:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 64509:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 64510:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 64511:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 64512:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 64513:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 64514:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 64515:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 64516:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 64517:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 64518:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 64519:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 64520:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 64521:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 64522:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 64523:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 64524:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 64525:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 64526:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 64527:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 64528:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 64529:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 64530:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 64531:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 64532:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 64533:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 64534:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 64535:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 64536:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 64537:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 64538:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 64539:22]
  assign io_z = ~x131; // @[Snxn100k.scala 64540:17]
endmodule
module SnxnLv4Inst59(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 63405:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 63406:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 63407:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 63408:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 63409:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 63410:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 63411:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 63412:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 63413:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 63414:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 63415:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 63416:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 63417:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 63418:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 63419:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 63420:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 63421:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 63422:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 63423:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 63424:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 63425:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 63426:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 63427:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 63428:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 63429:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 63430:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 63431:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 63432:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 63433:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 63434:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 63435:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 63436:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 63437:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 63438:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 63439:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 63440:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 63441:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 63442:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 63443:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 63444:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 63445:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 63446:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 63447:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 63448:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 63449:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 63450:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 63451:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 63452:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 63453:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 63454:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 63455:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 63456:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 63457:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 63458:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 63459:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 63460:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 63461:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 63462:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 63463:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 63464:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 63465:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 63466:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 63467:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 63468:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 63469:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 63470:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 63471:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 63472:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 63473:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 63474:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 63475:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 63476:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 63477:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 63478:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 63479:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 63480:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 63481:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 63482:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 63483:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 63484:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 63485:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 63486:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 63487:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 63488:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 63489:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 63490:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 63491:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 63492:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 63493:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 63494:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 63495:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 63496:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 63497:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 63498:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 63499:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 63500:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 63501:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 63502:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 63503:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 63504:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 63505:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 63506:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 63507:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 63508:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 63509:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 63510:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 63511:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 63512:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 63513:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 63514:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 63515:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 63516:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 63517:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 63518:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 63519:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 63520:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 63521:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 63522:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 63523:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 63524:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 63525:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 63526:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 63527:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 63528:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 63529:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 63530:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 63531:20]
  assign io_z = ~x31; // @[Snxn100k.scala 63532:16]
endmodule
module SnxnLv3Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst56_io_a; // @[Snxn100k.scala 21026:34]
  wire  inst_SnxnLv4Inst56_io_b; // @[Snxn100k.scala 21026:34]
  wire  inst_SnxnLv4Inst56_io_z; // @[Snxn100k.scala 21026:34]
  wire  inst_SnxnLv4Inst57_io_a; // @[Snxn100k.scala 21030:34]
  wire  inst_SnxnLv4Inst57_io_b; // @[Snxn100k.scala 21030:34]
  wire  inst_SnxnLv4Inst57_io_z; // @[Snxn100k.scala 21030:34]
  wire  inst_SnxnLv4Inst58_io_a; // @[Snxn100k.scala 21034:34]
  wire  inst_SnxnLv4Inst58_io_b; // @[Snxn100k.scala 21034:34]
  wire  inst_SnxnLv4Inst58_io_z; // @[Snxn100k.scala 21034:34]
  wire  inst_SnxnLv4Inst59_io_a; // @[Snxn100k.scala 21038:34]
  wire  inst_SnxnLv4Inst59_io_b; // @[Snxn100k.scala 21038:34]
  wire  inst_SnxnLv4Inst59_io_z; // @[Snxn100k.scala 21038:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst56_io_z + inst_SnxnLv4Inst57_io_z; // @[Snxn100k.scala 21042:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst58_io_z; // @[Snxn100k.scala 21042:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst59_io_z; // @[Snxn100k.scala 21042:89]
  SnxnLv4Inst56 inst_SnxnLv4Inst56 ( // @[Snxn100k.scala 21026:34]
    .io_a(inst_SnxnLv4Inst56_io_a),
    .io_b(inst_SnxnLv4Inst56_io_b),
    .io_z(inst_SnxnLv4Inst56_io_z)
  );
  SnxnLv4Inst8 inst_SnxnLv4Inst57 ( // @[Snxn100k.scala 21030:34]
    .io_a(inst_SnxnLv4Inst57_io_a),
    .io_b(inst_SnxnLv4Inst57_io_b),
    .io_z(inst_SnxnLv4Inst57_io_z)
  );
  SnxnLv4Inst58 inst_SnxnLv4Inst58 ( // @[Snxn100k.scala 21034:34]
    .io_a(inst_SnxnLv4Inst58_io_a),
    .io_b(inst_SnxnLv4Inst58_io_b),
    .io_z(inst_SnxnLv4Inst58_io_z)
  );
  SnxnLv4Inst59 inst_SnxnLv4Inst59 ( // @[Snxn100k.scala 21038:34]
    .io_a(inst_SnxnLv4Inst59_io_a),
    .io_b(inst_SnxnLv4Inst59_io_b),
    .io_z(inst_SnxnLv4Inst59_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21043:15]
  assign inst_SnxnLv4Inst56_io_a = io_a; // @[Snxn100k.scala 21027:27]
  assign inst_SnxnLv4Inst56_io_b = io_b; // @[Snxn100k.scala 21028:27]
  assign inst_SnxnLv4Inst57_io_a = io_a; // @[Snxn100k.scala 21031:27]
  assign inst_SnxnLv4Inst57_io_b = io_b; // @[Snxn100k.scala 21032:27]
  assign inst_SnxnLv4Inst58_io_a = io_a; // @[Snxn100k.scala 21035:27]
  assign inst_SnxnLv4Inst58_io_b = io_b; // @[Snxn100k.scala 21036:27]
  assign inst_SnxnLv4Inst59_io_a = io_a; // @[Snxn100k.scala 21039:27]
  assign inst_SnxnLv4Inst59_io_b = io_b; // @[Snxn100k.scala 21040:27]
endmodule
module SnxnLv4Inst61(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 67521:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 67522:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 67523:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 67524:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 67525:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 67526:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 67527:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 67528:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 67529:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 67530:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 67531:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 67532:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 67533:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 67534:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 67535:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 67536:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 67537:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 67538:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 67539:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 67540:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 67541:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 67542:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 67543:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 67544:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 67545:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 67546:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 67547:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 67548:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 67549:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 67550:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 67551:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 67552:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 67553:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 67554:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 67555:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 67556:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 67557:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 67558:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 67559:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 67560:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 67561:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 67562:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 67563:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 67564:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 67565:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 67566:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 67567:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 67568:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 67569:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 67570:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 67571:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 67572:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 67573:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 67574:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 67575:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 67576:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 67577:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 67578:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 67579:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 67580:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 67581:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 67582:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 67583:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 67584:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 67585:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 67586:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 67587:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 67588:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 67589:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 67590:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 67591:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 67592:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 67593:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 67594:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 67595:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 67596:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 67597:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 67598:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 67599:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 67600:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 67601:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 67602:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 67603:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 67604:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 67605:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 67606:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 67607:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 67608:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 67609:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 67610:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 67611:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 67612:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 67613:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 67614:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 67615:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 67616:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 67617:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 67618:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 67619:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 67620:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 67621:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 67622:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 67623:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 67624:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 67625:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 67626:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 67627:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 67628:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 67629:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 67630:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 67631:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 67632:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 67633:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 67634:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 67635:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 67636:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 67637:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 67638:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 67639:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 67640:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 67641:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 67642:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 67643:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 67644:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 67645:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 67646:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 67647:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 67648:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 67649:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 67650:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 67651:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 67652:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 67653:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 67654:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 67655:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 67656:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 67657:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 67658:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 67659:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 67660:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 67661:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 67662:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 67663:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 67664:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 67665:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 67666:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 67667:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 67668:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 67669:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 67670:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 67671:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 67672:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 67673:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 67674:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 67675:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 67676:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 67677:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 67678:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 67679:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 67680:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 67681:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 67682:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 67683:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 67684:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 67685:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 67686:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 67687:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 67688:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 67689:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 67690:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 67691:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 67692:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 67693:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 67694:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 67695:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 67696:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 67697:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 67698:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 67699:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 67700:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 67701:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 67702:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 67703:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 67704:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 67705:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 67706:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 67707:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 67708:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 67709:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 67710:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 67711:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 67712:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 67713:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 67714:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 67715:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 67716:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 67717:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 67718:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 67719:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 67720:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 67721:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 67722:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 67723:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 67724:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 67725:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 67726:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 67727:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 67728:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 67729:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 67730:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 67731:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 67732:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 67733:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 67734:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 67735:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 67736:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 67737:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 67738:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 67739:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 67740:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 67741:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 67742:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 67743:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 67744:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 67745:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 67746:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 67747:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 67748:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 67749:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 67750:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 67751:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 67752:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 67753:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 67754:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 67755:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 67756:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 67757:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 67758:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 67759:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 67760:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 67761:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 67762:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 67763:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 67764:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 67765:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 67766:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 67767:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 67768:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 67769:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 67770:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 67771:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 67772:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 67773:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 67774:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 67775:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 67776:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 67777:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 67778:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 67779:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 67780:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 67781:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 67782:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 67783:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 67784:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 67785:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 67786:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 67787:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 67788:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 67789:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 67790:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 67791:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 67792:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 67793:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 67794:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 67795:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 67796:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 67797:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 67798:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 67799:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 67800:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 67801:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 67802:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 67803:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 67804:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 67805:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 67806:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 67807:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 67808:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 67809:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 67810:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 67811:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 67812:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 67813:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 67814:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 67815:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 67816:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 67817:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 67818:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 67819:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 67820:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 67821:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 67822:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 67823:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 67824:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 67825:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 67826:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 67827:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 67828:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 67829:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 67830:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 67831:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 67832:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 67833:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 67834:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 67835:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 67836:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 67837:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 67838:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 67839:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 67840:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 67841:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 67842:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 67843:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 67844:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 67845:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 67846:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 67847:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 67848:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 67849:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 67850:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 67851:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 67852:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 67853:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 67854:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 67855:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 67856:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 67857:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 67858:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 67859:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 67860:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 67861:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 67862:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 67863:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 67864:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 67865:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 67866:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 67867:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 67868:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 67869:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 67870:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 67871:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 67872:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 67873:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 67874:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 67875:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 67876:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 67877:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 67878:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 67879:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 67880:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 67881:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 67882:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 67883:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 67884:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 67885:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 67886:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 67887:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 67888:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 67889:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 67890:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 67891:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 67892:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 67893:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 67894:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 67895:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 67896:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 67897:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 67898:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 67899:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 67900:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 67901:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 67902:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 67903:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 67904:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 67905:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 67906:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 67907:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 67908:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 67909:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 67910:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 67911:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 67912:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 67913:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 67914:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 67915:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 67916:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 67917:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 67918:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 67919:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 67920:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 67921:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 67922:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 67923:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 67924:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 67925:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 67926:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 67927:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 67928:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 67929:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 67930:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 67931:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 67932:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 67933:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 67934:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 67935:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 67936:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 67937:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 67938:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 67939:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 67940:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 67941:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 67942:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 67943:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 67944:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 67945:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 67946:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 67947:22]
  assign io_z = ~x106; // @[Snxn100k.scala 67948:17]
endmodule
module SnxnLv4Inst63(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 67495:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 67496:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 67497:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 67498:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 67499:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 67500:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 67501:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 67502:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 67503:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 67504:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 67505:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 67506:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 67507:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 67508:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 67509:18]
  assign io_z = ~x3; // @[Snxn100k.scala 67510:15]
endmodule
module SnxnLv3Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst60_io_a; // @[Snxn100k.scala 21887:34]
  wire  inst_SnxnLv4Inst60_io_b; // @[Snxn100k.scala 21887:34]
  wire  inst_SnxnLv4Inst60_io_z; // @[Snxn100k.scala 21887:34]
  wire  inst_SnxnLv4Inst61_io_a; // @[Snxn100k.scala 21891:34]
  wire  inst_SnxnLv4Inst61_io_b; // @[Snxn100k.scala 21891:34]
  wire  inst_SnxnLv4Inst61_io_z; // @[Snxn100k.scala 21891:34]
  wire  inst_SnxnLv4Inst62_io_a; // @[Snxn100k.scala 21895:34]
  wire  inst_SnxnLv4Inst62_io_b; // @[Snxn100k.scala 21895:34]
  wire  inst_SnxnLv4Inst62_io_z; // @[Snxn100k.scala 21895:34]
  wire  inst_SnxnLv4Inst63_io_a; // @[Snxn100k.scala 21899:34]
  wire  inst_SnxnLv4Inst63_io_b; // @[Snxn100k.scala 21899:34]
  wire  inst_SnxnLv4Inst63_io_z; // @[Snxn100k.scala 21899:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst60_io_z + inst_SnxnLv4Inst61_io_z; // @[Snxn100k.scala 21903:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst62_io_z; // @[Snxn100k.scala 21903:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst63_io_z; // @[Snxn100k.scala 21903:89]
  SnxnLv4Inst24 inst_SnxnLv4Inst60 ( // @[Snxn100k.scala 21887:34]
    .io_a(inst_SnxnLv4Inst60_io_a),
    .io_b(inst_SnxnLv4Inst60_io_b),
    .io_z(inst_SnxnLv4Inst60_io_z)
  );
  SnxnLv4Inst61 inst_SnxnLv4Inst61 ( // @[Snxn100k.scala 21891:34]
    .io_a(inst_SnxnLv4Inst61_io_a),
    .io_b(inst_SnxnLv4Inst61_io_b),
    .io_z(inst_SnxnLv4Inst61_io_z)
  );
  SnxnLv4Inst61 inst_SnxnLv4Inst62 ( // @[Snxn100k.scala 21895:34]
    .io_a(inst_SnxnLv4Inst62_io_a),
    .io_b(inst_SnxnLv4Inst62_io_b),
    .io_z(inst_SnxnLv4Inst62_io_z)
  );
  SnxnLv4Inst63 inst_SnxnLv4Inst63 ( // @[Snxn100k.scala 21899:34]
    .io_a(inst_SnxnLv4Inst63_io_a),
    .io_b(inst_SnxnLv4Inst63_io_b),
    .io_z(inst_SnxnLv4Inst63_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 21904:15]
  assign inst_SnxnLv4Inst60_io_a = io_a; // @[Snxn100k.scala 21888:27]
  assign inst_SnxnLv4Inst60_io_b = io_b; // @[Snxn100k.scala 21889:27]
  assign inst_SnxnLv4Inst61_io_a = io_a; // @[Snxn100k.scala 21892:27]
  assign inst_SnxnLv4Inst61_io_b = io_b; // @[Snxn100k.scala 21893:27]
  assign inst_SnxnLv4Inst62_io_a = io_a; // @[Snxn100k.scala 21896:27]
  assign inst_SnxnLv4Inst62_io_b = io_b; // @[Snxn100k.scala 21897:27]
  assign inst_SnxnLv4Inst63_io_a = io_a; // @[Snxn100k.scala 21900:27]
  assign inst_SnxnLv4Inst63_io_b = io_b; // @[Snxn100k.scala 21901:27]
endmodule
module SnxnLv2Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst12_io_a; // @[Snxn100k.scala 5880:34]
  wire  inst_SnxnLv3Inst12_io_b; // @[Snxn100k.scala 5880:34]
  wire  inst_SnxnLv3Inst12_io_z; // @[Snxn100k.scala 5880:34]
  wire  inst_SnxnLv3Inst13_io_a; // @[Snxn100k.scala 5884:34]
  wire  inst_SnxnLv3Inst13_io_b; // @[Snxn100k.scala 5884:34]
  wire  inst_SnxnLv3Inst13_io_z; // @[Snxn100k.scala 5884:34]
  wire  inst_SnxnLv3Inst14_io_a; // @[Snxn100k.scala 5888:34]
  wire  inst_SnxnLv3Inst14_io_b; // @[Snxn100k.scala 5888:34]
  wire  inst_SnxnLv3Inst14_io_z; // @[Snxn100k.scala 5888:34]
  wire  inst_SnxnLv3Inst15_io_a; // @[Snxn100k.scala 5892:34]
  wire  inst_SnxnLv3Inst15_io_b; // @[Snxn100k.scala 5892:34]
  wire  inst_SnxnLv3Inst15_io_z; // @[Snxn100k.scala 5892:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst12_io_z + inst_SnxnLv3Inst13_io_z; // @[Snxn100k.scala 5896:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst14_io_z; // @[Snxn100k.scala 5896:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst15_io_z; // @[Snxn100k.scala 5896:89]
  SnxnLv3Inst12 inst_SnxnLv3Inst12 ( // @[Snxn100k.scala 5880:34]
    .io_a(inst_SnxnLv3Inst12_io_a),
    .io_b(inst_SnxnLv3Inst12_io_b),
    .io_z(inst_SnxnLv3Inst12_io_z)
  );
  SnxnLv3Inst13 inst_SnxnLv3Inst13 ( // @[Snxn100k.scala 5884:34]
    .io_a(inst_SnxnLv3Inst13_io_a),
    .io_b(inst_SnxnLv3Inst13_io_b),
    .io_z(inst_SnxnLv3Inst13_io_z)
  );
  SnxnLv3Inst14 inst_SnxnLv3Inst14 ( // @[Snxn100k.scala 5888:34]
    .io_a(inst_SnxnLv3Inst14_io_a),
    .io_b(inst_SnxnLv3Inst14_io_b),
    .io_z(inst_SnxnLv3Inst14_io_z)
  );
  SnxnLv3Inst15 inst_SnxnLv3Inst15 ( // @[Snxn100k.scala 5892:34]
    .io_a(inst_SnxnLv3Inst15_io_a),
    .io_b(inst_SnxnLv3Inst15_io_b),
    .io_z(inst_SnxnLv3Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 5897:15]
  assign inst_SnxnLv3Inst12_io_a = io_a; // @[Snxn100k.scala 5881:27]
  assign inst_SnxnLv3Inst12_io_b = io_b; // @[Snxn100k.scala 5882:27]
  assign inst_SnxnLv3Inst13_io_a = io_a; // @[Snxn100k.scala 5885:27]
  assign inst_SnxnLv3Inst13_io_b = io_b; // @[Snxn100k.scala 5886:27]
  assign inst_SnxnLv3Inst14_io_a = io_a; // @[Snxn100k.scala 5889:27]
  assign inst_SnxnLv3Inst14_io_b = io_b; // @[Snxn100k.scala 5890:27]
  assign inst_SnxnLv3Inst15_io_a = io_a; // @[Snxn100k.scala 5893:27]
  assign inst_SnxnLv3Inst15_io_b = io_b; // @[Snxn100k.scala 5894:27]
endmodule
module SnxnLv1Inst0(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst0_io_a; // @[Snxn100k.scala 1038:33]
  wire  inst_SnxnLv2Inst0_io_b; // @[Snxn100k.scala 1038:33]
  wire  inst_SnxnLv2Inst0_io_z; // @[Snxn100k.scala 1038:33]
  wire  inst_SnxnLv2Inst1_io_a; // @[Snxn100k.scala 1042:33]
  wire  inst_SnxnLv2Inst1_io_b; // @[Snxn100k.scala 1042:33]
  wire  inst_SnxnLv2Inst1_io_z; // @[Snxn100k.scala 1042:33]
  wire  inst_SnxnLv2Inst2_io_a; // @[Snxn100k.scala 1046:33]
  wire  inst_SnxnLv2Inst2_io_b; // @[Snxn100k.scala 1046:33]
  wire  inst_SnxnLv2Inst2_io_z; // @[Snxn100k.scala 1046:33]
  wire  inst_SnxnLv2Inst3_io_a; // @[Snxn100k.scala 1050:33]
  wire  inst_SnxnLv2Inst3_io_b; // @[Snxn100k.scala 1050:33]
  wire  inst_SnxnLv2Inst3_io_z; // @[Snxn100k.scala 1050:33]
  wire  _sum_T_1 = inst_SnxnLv2Inst0_io_z + inst_SnxnLv2Inst1_io_z; // @[Snxn100k.scala 1054:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst2_io_z; // @[Snxn100k.scala 1054:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst3_io_z; // @[Snxn100k.scala 1054:86]
  SnxnLv2Inst0 inst_SnxnLv2Inst0 ( // @[Snxn100k.scala 1038:33]
    .io_a(inst_SnxnLv2Inst0_io_a),
    .io_b(inst_SnxnLv2Inst0_io_b),
    .io_z(inst_SnxnLv2Inst0_io_z)
  );
  SnxnLv2Inst1 inst_SnxnLv2Inst1 ( // @[Snxn100k.scala 1042:33]
    .io_a(inst_SnxnLv2Inst1_io_a),
    .io_b(inst_SnxnLv2Inst1_io_b),
    .io_z(inst_SnxnLv2Inst1_io_z)
  );
  SnxnLv2Inst2 inst_SnxnLv2Inst2 ( // @[Snxn100k.scala 1046:33]
    .io_a(inst_SnxnLv2Inst2_io_a),
    .io_b(inst_SnxnLv2Inst2_io_b),
    .io_z(inst_SnxnLv2Inst2_io_z)
  );
  SnxnLv2Inst3 inst_SnxnLv2Inst3 ( // @[Snxn100k.scala 1050:33]
    .io_a(inst_SnxnLv2Inst3_io_a),
    .io_b(inst_SnxnLv2Inst3_io_b),
    .io_z(inst_SnxnLv2Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1055:15]
  assign inst_SnxnLv2Inst0_io_a = io_a; // @[Snxn100k.scala 1039:26]
  assign inst_SnxnLv2Inst0_io_b = io_b; // @[Snxn100k.scala 1040:26]
  assign inst_SnxnLv2Inst1_io_a = io_a; // @[Snxn100k.scala 1043:26]
  assign inst_SnxnLv2Inst1_io_b = io_b; // @[Snxn100k.scala 1044:26]
  assign inst_SnxnLv2Inst2_io_a = io_a; // @[Snxn100k.scala 1047:26]
  assign inst_SnxnLv2Inst2_io_b = io_b; // @[Snxn100k.scala 1048:26]
  assign inst_SnxnLv2Inst3_io_a = io_a; // @[Snxn100k.scala 1051:26]
  assign inst_SnxnLv2Inst3_io_b = io_b; // @[Snxn100k.scala 1052:26]
endmodule
module SnxnLv4Inst64(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 42331:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 42332:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 42333:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 42334:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 42335:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 42336:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 42337:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 42338:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 42339:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 42340:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 42341:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 42342:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 42343:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 42344:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 42345:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 42346:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 42347:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 42348:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 42349:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 42350:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 42351:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 42352:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 42353:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 42354:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 42355:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 42356:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 42357:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 42358:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 42359:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 42360:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 42361:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 42362:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 42363:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 42364:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 42365:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 42366:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 42367:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 42368:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 42369:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 42370:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 42371:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 42372:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 42373:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 42374:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 42375:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 42376:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 42377:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 42378:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 42379:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 42380:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 42381:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 42382:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 42383:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 42384:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 42385:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 42386:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 42387:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 42388:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 42389:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 42390:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 42391:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 42392:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 42393:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 42394:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 42395:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 42396:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 42397:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 42398:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 42399:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 42400:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 42401:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 42402:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 42403:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 42404:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 42405:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 42406:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 42407:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 42408:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 42409:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 42410:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 42411:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 42412:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 42413:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 42414:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 42415:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 42416:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 42417:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 42418:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 42419:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 42420:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 42421:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 42422:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 42423:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 42424:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 42425:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 42426:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 42427:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 42428:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 42429:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 42430:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 42431:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 42432:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 42433:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 42434:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 42435:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 42436:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 42437:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 42438:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 42439:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 42440:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 42441:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 42442:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 42443:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 42444:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 42445:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 42446:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 42447:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 42448:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 42449:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 42450:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 42451:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 42452:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 42453:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 42454:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 42455:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 42456:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 42457:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 42458:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 42459:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 42460:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 42461:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 42462:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 42463:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 42464:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 42465:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 42466:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 42467:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 42468:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 42469:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 42470:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 42471:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 42472:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 42473:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 42474:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 42475:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 42476:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 42477:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 42478:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 42479:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 42480:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 42481:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 42482:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 42483:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 42484:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 42485:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 42486:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 42487:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 42488:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 42489:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 42490:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 42491:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 42492:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 42493:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 42494:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 42495:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 42496:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 42497:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 42498:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 42499:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 42500:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 42501:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 42502:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 42503:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 42504:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 42505:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 42506:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 42507:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 42508:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 42509:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 42510:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 42511:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 42512:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 42513:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 42514:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 42515:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 42516:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 42517:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 42518:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 42519:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 42520:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 42521:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 42522:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 42523:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 42524:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 42525:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 42526:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 42527:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 42528:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 42529:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 42530:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 42531:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 42532:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 42533:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 42534:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 42535:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 42536:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 42537:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 42538:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 42539:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 42540:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 42541:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 42542:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 42543:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 42544:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 42545:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 42546:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 42547:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 42548:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 42549:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 42550:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 42551:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 42552:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 42553:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 42554:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 42555:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 42556:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 42557:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 42558:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 42559:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 42560:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 42561:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 42562:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 42563:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 42564:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 42565:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 42566:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 42567:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 42568:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 42569:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 42570:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 42571:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 42572:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 42573:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 42574:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 42575:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 42576:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 42577:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 42578:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 42579:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 42580:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 42581:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 42582:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 42583:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 42584:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 42585:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 42586:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 42587:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 42588:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 42589:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 42590:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 42591:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 42592:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 42593:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 42594:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 42595:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 42596:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 42597:20]
  assign io_z = ~x66; // @[Snxn100k.scala 42598:16]
endmodule
module SnxnLv4Inst65(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 42161:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 42162:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 42163:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 42164:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 42165:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 42166:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 42167:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 42168:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 42169:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 42170:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 42171:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 42172:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 42173:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 42174:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 42175:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 42176:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 42177:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 42178:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 42179:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 42180:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 42181:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 42182:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 42183:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 42184:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 42185:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 42186:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 42187:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 42188:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 42189:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 42190:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 42191:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 42192:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 42193:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 42194:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 42195:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 42196:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 42197:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 42198:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 42199:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 42200:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 42201:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 42202:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 42203:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 42204:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 42205:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 42206:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 42207:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 42208:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 42209:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 42210:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 42211:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 42212:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 42213:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 42214:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 42215:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 42216:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 42217:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 42218:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 42219:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 42220:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 42221:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 42222:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 42223:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 42224:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 42225:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 42226:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 42227:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 42228:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 42229:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 42230:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 42231:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 42232:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 42233:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 42234:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 42235:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 42236:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 42237:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 42238:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 42239:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 42240:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 42241:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 42242:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 42243:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 42244:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 42245:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 42246:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 42247:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 42248:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 42249:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 42250:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 42251:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 42252:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 42253:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 42254:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 42255:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 42256:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 42257:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 42258:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 42259:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 42260:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 42261:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 42262:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 42263:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 42264:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 42265:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 42266:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 42267:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 42268:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 42269:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 42270:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 42271:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 42272:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 42273:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 42274:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 42275:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 42276:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 42277:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 42278:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 42279:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 42280:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 42281:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 42282:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 42283:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 42284:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 42285:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 42286:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 42287:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 42288:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 42289:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 42290:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 42291:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 42292:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 42293:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 42294:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 42295:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 42296:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 42297:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 42298:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 42299:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 42300:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 42301:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 42302:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 42303:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 42304:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 42305:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 42306:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 42307:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 42308:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 42309:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 42310:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 42311:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 42312:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 42313:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 42314:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 42315:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 42316:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 42317:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 42318:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 42319:20]
  assign io_z = ~x39; // @[Snxn100k.scala 42320:16]
endmodule
module SnxnLv4Inst67(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 42609:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 42610:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 42611:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 42612:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 42613:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 42614:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 42615:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 42616:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 42617:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 42618:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 42619:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 42620:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 42621:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 42622:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 42623:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 42624:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 42625:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 42626:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 42627:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 42628:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 42629:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 42630:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 42631:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 42632:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 42633:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 42634:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 42635:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 42636:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 42637:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 42638:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 42639:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 42640:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 42641:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 42642:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 42643:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 42644:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 42645:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 42646:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 42647:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 42648:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 42649:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 42650:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 42651:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 42652:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 42653:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 42654:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 42655:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 42656:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 42657:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 42658:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 42659:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 42660:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 42661:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 42662:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 42663:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 42664:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 42665:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 42666:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 42667:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 42668:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 42669:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 42670:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 42671:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 42672:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 42673:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 42674:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 42675:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 42676:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 42677:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 42678:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 42679:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 42680:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 42681:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 42682:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 42683:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 42684:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 42685:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 42686:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 42687:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 42688:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 42689:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 42690:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 42691:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 42692:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 42693:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 42694:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 42695:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 42696:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 42697:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 42698:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 42699:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 42700:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 42701:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 42702:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 42703:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 42704:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 42705:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 42706:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 42707:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 42708:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 42709:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 42710:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 42711:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 42712:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 42713:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 42714:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 42715:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 42716:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 42717:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 42718:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 42719:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 42720:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 42721:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 42722:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 42723:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 42724:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 42725:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 42726:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 42727:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 42728:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 42729:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 42730:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 42731:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 42732:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 42733:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 42734:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 42735:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 42736:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 42737:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 42738:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 42739:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 42740:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 42741:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 42742:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 42743:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 42744:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 42745:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 42746:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 42747:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 42748:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 42749:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 42750:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 42751:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 42752:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 42753:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 42754:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 42755:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 42756:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 42757:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 42758:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 42759:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 42760:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 42761:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 42762:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 42763:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 42764:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 42765:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 42766:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 42767:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 42768:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 42769:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 42770:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 42771:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 42772:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 42773:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 42774:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 42775:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 42776:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 42777:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 42778:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 42779:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 42780:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 42781:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 42782:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 42783:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 42784:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 42785:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 42786:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 42787:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 42788:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 42789:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 42790:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 42791:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 42792:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 42793:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 42794:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 42795:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 42796:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 42797:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 42798:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 42799:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 42800:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 42801:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 42802:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 42803:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 42804:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 42805:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 42806:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 42807:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 42808:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 42809:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 42810:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 42811:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 42812:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 42813:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 42814:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 42815:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 42816:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 42817:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 42818:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 42819:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 42820:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 42821:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 42822:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 42823:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 42824:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 42825:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 42826:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 42827:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 42828:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 42829:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 42830:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 42831:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 42832:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 42833:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 42834:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 42835:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 42836:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 42837:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 42838:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 42839:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 42840:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 42841:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 42842:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 42843:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 42844:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 42845:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 42846:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 42847:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 42848:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 42849:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 42850:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 42851:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 42852:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 42853:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 42854:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 42855:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 42856:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 42857:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 42858:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 42859:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 42860:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 42861:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 42862:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 42863:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 42864:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 42865:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 42866:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 42867:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 42868:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 42869:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 42870:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 42871:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 42872:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 42873:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 42874:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 42875:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 42876:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 42877:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 42878:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 42879:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 42880:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 42881:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 42882:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 42883:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 42884:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 42885:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 42886:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 42887:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 42888:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 42889:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 42890:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 42891:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 42892:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 42893:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 42894:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 42895:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 42896:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 42897:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 42898:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 42899:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 42900:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 42901:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 42902:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 42903:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 42904:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 42905:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 42906:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 42907:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 42908:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 42909:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 42910:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 42911:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 42912:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 42913:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 42914:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 42915:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 42916:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 42917:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 42918:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 42919:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 42920:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 42921:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 42922:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 42923:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 42924:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 42925:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 42926:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 42927:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 42928:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 42929:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 42930:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 42931:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 42932:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 42933:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 42934:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 42935:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 42936:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 42937:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 42938:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 42939:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 42940:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 42941:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 42942:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 42943:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 42944:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 42945:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 42946:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 42947:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 42948:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 42949:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 42950:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 42951:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 42952:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 42953:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 42954:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 42955:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 42956:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 42957:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 42958:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 42959:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 42960:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 42961:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 42962:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 42963:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 42964:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 42965:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 42966:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 42967:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 42968:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 42969:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 42970:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 42971:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 42972:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 42973:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 42974:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 42975:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 42976:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 42977:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 42978:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 42979:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 42980:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 42981:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 42982:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 42983:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 42984:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 42985:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 42986:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 42987:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 42988:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 42989:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 42990:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 42991:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 42992:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 42993:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 42994:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 42995:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 42996:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 42997:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 42998:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 42999:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 43000:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 43001:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 43002:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 43003:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 43004:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 43005:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 43006:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 43007:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 43008:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 43009:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 43010:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 43011:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 43012:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 43013:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 43014:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 43015:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 43016:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 43017:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 43018:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 43019:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 43020:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 43021:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 43022:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 43023:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 43024:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 43025:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 43026:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 43027:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 43028:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 43029:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 43030:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 43031:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 43032:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 43033:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 43034:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 43035:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 43036:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 43037:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 43038:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 43039:22]
  assign io_z = ~x107; // @[Snxn100k.scala 43040:17]
endmodule
module SnxnLv3Inst16(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst64_io_a; // @[Snxn100k.scala 12426:34]
  wire  inst_SnxnLv4Inst64_io_b; // @[Snxn100k.scala 12426:34]
  wire  inst_SnxnLv4Inst64_io_z; // @[Snxn100k.scala 12426:34]
  wire  inst_SnxnLv4Inst65_io_a; // @[Snxn100k.scala 12430:34]
  wire  inst_SnxnLv4Inst65_io_b; // @[Snxn100k.scala 12430:34]
  wire  inst_SnxnLv4Inst65_io_z; // @[Snxn100k.scala 12430:34]
  wire  inst_SnxnLv4Inst66_io_a; // @[Snxn100k.scala 12434:34]
  wire  inst_SnxnLv4Inst66_io_b; // @[Snxn100k.scala 12434:34]
  wire  inst_SnxnLv4Inst66_io_z; // @[Snxn100k.scala 12434:34]
  wire  inst_SnxnLv4Inst67_io_a; // @[Snxn100k.scala 12438:34]
  wire  inst_SnxnLv4Inst67_io_b; // @[Snxn100k.scala 12438:34]
  wire  inst_SnxnLv4Inst67_io_z; // @[Snxn100k.scala 12438:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst64_io_z + inst_SnxnLv4Inst65_io_z; // @[Snxn100k.scala 12442:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst66_io_z; // @[Snxn100k.scala 12442:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst67_io_z; // @[Snxn100k.scala 12442:89]
  SnxnLv4Inst64 inst_SnxnLv4Inst64 ( // @[Snxn100k.scala 12426:34]
    .io_a(inst_SnxnLv4Inst64_io_a),
    .io_b(inst_SnxnLv4Inst64_io_b),
    .io_z(inst_SnxnLv4Inst64_io_z)
  );
  SnxnLv4Inst65 inst_SnxnLv4Inst65 ( // @[Snxn100k.scala 12430:34]
    .io_a(inst_SnxnLv4Inst65_io_a),
    .io_b(inst_SnxnLv4Inst65_io_b),
    .io_z(inst_SnxnLv4Inst65_io_z)
  );
  SnxnLv4Inst14 inst_SnxnLv4Inst66 ( // @[Snxn100k.scala 12434:34]
    .io_a(inst_SnxnLv4Inst66_io_a),
    .io_b(inst_SnxnLv4Inst66_io_b),
    .io_z(inst_SnxnLv4Inst66_io_z)
  );
  SnxnLv4Inst67 inst_SnxnLv4Inst67 ( // @[Snxn100k.scala 12438:34]
    .io_a(inst_SnxnLv4Inst67_io_a),
    .io_b(inst_SnxnLv4Inst67_io_b),
    .io_z(inst_SnxnLv4Inst67_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 12443:15]
  assign inst_SnxnLv4Inst64_io_a = io_a; // @[Snxn100k.scala 12427:27]
  assign inst_SnxnLv4Inst64_io_b = io_b; // @[Snxn100k.scala 12428:27]
  assign inst_SnxnLv4Inst65_io_a = io_a; // @[Snxn100k.scala 12431:27]
  assign inst_SnxnLv4Inst65_io_b = io_b; // @[Snxn100k.scala 12432:27]
  assign inst_SnxnLv4Inst66_io_a = io_a; // @[Snxn100k.scala 12435:27]
  assign inst_SnxnLv4Inst66_io_b = io_b; // @[Snxn100k.scala 12436:27]
  assign inst_SnxnLv4Inst67_io_a = io_a; // @[Snxn100k.scala 12439:27]
  assign inst_SnxnLv4Inst67_io_b = io_b; // @[Snxn100k.scala 12440:27]
endmodule
module SnxnLv4Inst69(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 39335:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 39336:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 39337:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 39338:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 39339:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 39340:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 39341:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 39342:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 39343:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 39344:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 39345:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 39346:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 39347:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 39348:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 39349:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 39350:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 39351:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 39352:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 39353:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 39354:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 39355:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 39356:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 39357:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 39358:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 39359:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 39360:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 39361:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 39362:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 39363:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 39364:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 39365:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 39366:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 39367:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 39368:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 39369:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 39370:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 39371:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 39372:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 39373:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 39374:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 39375:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 39376:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 39377:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 39378:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 39379:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 39380:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 39381:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 39382:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 39383:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 39384:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 39385:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 39386:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 39387:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 39388:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 39389:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 39390:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 39391:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 39392:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 39393:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 39394:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 39395:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 39396:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 39397:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 39398:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 39399:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 39400:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 39401:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 39402:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 39403:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 39404:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 39405:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 39406:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 39407:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 39408:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 39409:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 39410:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 39411:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 39412:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 39413:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 39414:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 39415:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 39416:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 39417:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 39418:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 39419:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 39420:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 39421:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 39422:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 39423:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 39424:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 39425:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 39426:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 39427:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 39428:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 39429:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 39430:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 39431:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 39432:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 39433:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 39434:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 39435:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 39436:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 39437:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 39438:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 39439:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 39440:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 39441:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 39442:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 39443:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 39444:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 39445:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 39446:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 39447:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 39448:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 39449:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 39450:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 39451:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 39452:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 39453:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 39454:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 39455:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 39456:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 39457:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 39458:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 39459:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 39460:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 39461:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 39462:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 39463:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 39464:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 39465:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 39466:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 39467:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 39468:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 39469:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 39470:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 39471:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 39472:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 39473:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 39474:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 39475:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 39476:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 39477:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 39478:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 39479:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 39480:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 39481:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 39482:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 39483:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 39484:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 39485:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 39486:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 39487:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 39488:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 39489:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 39490:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 39491:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 39492:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 39493:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 39494:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 39495:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 39496:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 39497:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 39498:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 39499:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 39500:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 39501:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 39502:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 39503:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 39504:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 39505:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 39506:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 39507:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 39508:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 39509:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 39510:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 39511:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 39512:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 39513:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 39514:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 39515:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 39516:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 39517:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 39518:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 39519:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 39520:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 39521:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 39522:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 39523:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 39524:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 39525:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 39526:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 39527:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 39528:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 39529:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 39530:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 39531:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 39532:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 39533:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 39534:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 39535:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 39536:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 39537:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 39538:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 39539:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 39540:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 39541:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 39542:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 39543:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 39544:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 39545:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 39546:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 39547:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 39548:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 39549:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 39550:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 39551:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 39552:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 39553:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 39554:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 39555:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 39556:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 39557:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 39558:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 39559:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 39560:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 39561:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 39562:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 39563:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 39564:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 39565:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 39566:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 39567:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 39568:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 39569:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 39570:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 39571:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 39572:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 39573:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 39574:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 39575:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 39576:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 39577:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 39578:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 39579:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 39580:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 39581:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 39582:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 39583:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 39584:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 39585:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 39586:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 39587:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 39588:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 39589:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 39590:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 39591:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 39592:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 39593:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 39594:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 39595:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 39596:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 39597:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 39598:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 39599:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 39600:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 39601:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 39602:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 39603:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 39604:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 39605:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 39606:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 39607:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 39608:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 39609:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 39610:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 39611:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 39612:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 39613:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 39614:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 39615:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 39616:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 39617:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 39618:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 39619:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 39620:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 39621:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 39622:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 39623:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 39624:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 39625:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 39626:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 39627:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 39628:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 39629:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 39630:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 39631:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 39632:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 39633:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 39634:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 39635:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 39636:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 39637:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 39638:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 39639:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 39640:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 39641:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 39642:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 39643:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 39644:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 39645:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 39646:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 39647:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 39648:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 39649:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 39650:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 39651:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 39652:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 39653:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 39654:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 39655:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 39656:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 39657:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 39658:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 39659:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 39660:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 39661:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 39662:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 39663:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 39664:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 39665:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 39666:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 39667:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 39668:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 39669:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 39670:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 39671:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 39672:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 39673:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 39674:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 39675:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 39676:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 39677:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 39678:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 39679:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 39680:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 39681:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 39682:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 39683:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 39684:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 39685:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 39686:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 39687:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 39688:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 39689:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 39690:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 39691:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 39692:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 39693:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 39694:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 39695:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 39696:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 39697:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 39698:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 39699:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 39700:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 39701:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 39702:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 39703:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 39704:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 39705:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 39706:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 39707:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 39708:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 39709:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 39710:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 39711:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 39712:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 39713:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 39714:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 39715:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 39716:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 39717:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 39718:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 39719:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 39720:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 39721:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 39722:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 39723:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 39724:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 39725:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 39726:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 39727:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 39728:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 39729:20]
  assign io_z = ~x98; // @[Snxn100k.scala 39730:16]
endmodule
module SnxnLv4Inst71(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 40199:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 40200:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 40201:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 40202:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 40203:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 40204:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 40205:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 40206:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 40207:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 40208:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 40209:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 40210:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 40211:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 40212:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 40213:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 40214:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 40215:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 40216:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 40217:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 40218:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 40219:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 40220:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 40221:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 40222:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 40223:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 40224:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 40225:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 40226:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 40227:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 40228:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 40229:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 40230:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 40231:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 40232:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 40233:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 40234:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 40235:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 40236:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 40237:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 40238:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 40239:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 40240:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 40241:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 40242:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 40243:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 40244:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 40245:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 40246:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 40247:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 40248:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 40249:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 40250:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 40251:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 40252:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 40253:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 40254:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 40255:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 40256:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 40257:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 40258:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 40259:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 40260:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 40261:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 40262:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 40263:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 40264:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 40265:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 40266:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 40267:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 40268:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 40269:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 40270:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 40271:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 40272:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 40273:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 40274:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 40275:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 40276:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 40277:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 40278:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 40279:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 40280:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 40281:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 40282:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 40283:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 40284:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 40285:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 40286:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 40287:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 40288:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 40289:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 40290:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 40291:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 40292:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 40293:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 40294:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 40295:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 40296:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 40297:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 40298:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 40299:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 40300:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 40301:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 40302:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 40303:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 40304:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 40305:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 40306:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 40307:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 40308:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 40309:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 40310:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 40311:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 40312:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 40313:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 40314:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 40315:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 40316:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 40317:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 40318:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 40319:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 40320:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 40321:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 40322:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 40323:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 40324:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 40325:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 40326:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 40327:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 40328:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 40329:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 40330:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 40331:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 40332:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 40333:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 40334:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 40335:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 40336:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 40337:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 40338:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 40339:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 40340:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 40341:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 40342:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 40343:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 40344:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 40345:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 40346:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 40347:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 40348:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 40349:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 40350:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 40351:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 40352:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 40353:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 40354:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 40355:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 40356:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 40357:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 40358:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 40359:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 40360:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 40361:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 40362:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 40363:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 40364:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 40365:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 40366:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 40367:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 40368:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 40369:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 40370:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 40371:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 40372:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 40373:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 40374:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 40375:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 40376:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 40377:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 40378:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 40379:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 40380:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 40381:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 40382:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 40383:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 40384:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 40385:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 40386:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 40387:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 40388:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 40389:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 40390:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 40391:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 40392:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 40393:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 40394:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 40395:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 40396:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 40397:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 40398:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 40399:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 40400:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 40401:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 40402:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 40403:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 40404:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 40405:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 40406:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 40407:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 40408:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 40409:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 40410:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 40411:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 40412:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 40413:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 40414:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 40415:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 40416:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 40417:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 40418:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 40419:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 40420:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 40421:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 40422:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 40423:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 40424:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 40425:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 40426:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 40427:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 40428:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 40429:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 40430:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 40431:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 40432:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 40433:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 40434:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 40435:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 40436:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 40437:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 40438:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 40439:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 40440:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 40441:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 40442:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 40443:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 40444:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 40445:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 40446:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 40447:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 40448:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 40449:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 40450:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 40451:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 40452:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 40453:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 40454:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 40455:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 40456:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 40457:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 40458:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 40459:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 40460:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 40461:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 40462:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 40463:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 40464:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 40465:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 40466:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 40467:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 40468:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 40469:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 40470:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 40471:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 40472:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 40473:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 40474:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 40475:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 40476:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 40477:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 40478:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 40479:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 40480:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 40481:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 40482:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 40483:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 40484:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 40485:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 40486:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 40487:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 40488:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 40489:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 40490:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 40491:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 40492:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 40493:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 40494:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 40495:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 40496:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 40497:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 40498:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 40499:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 40500:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 40501:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 40502:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 40503:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 40504:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 40505:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 40506:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 40507:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 40508:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 40509:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 40510:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 40511:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 40512:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 40513:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 40514:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 40515:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 40516:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 40517:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 40518:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 40519:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 40520:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 40521:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 40522:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 40523:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 40524:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 40525:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 40526:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 40527:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 40528:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 40529:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 40530:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 40531:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 40532:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 40533:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 40534:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 40535:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 40536:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 40537:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 40538:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 40539:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 40540:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 40541:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 40542:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 40543:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 40544:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 40545:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 40546:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 40547:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 40548:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 40549:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 40550:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 40551:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 40552:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 40553:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 40554:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 40555:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 40556:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 40557:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 40558:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 40559:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 40560:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 40561:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 40562:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 40563:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 40564:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 40565:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 40566:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 40567:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 40568:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 40569:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 40570:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 40571:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 40572:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 40573:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 40574:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 40575:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 40576:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 40577:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 40578:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 40579:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 40580:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 40581:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 40582:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 40583:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 40584:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 40585:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 40586:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 40587:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 40588:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 40589:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 40590:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 40591:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 40592:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 40593:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 40594:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 40595:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 40596:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 40597:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 40598:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 40599:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 40600:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 40601:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 40602:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 40603:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 40604:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 40605:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 40606:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 40607:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 40608:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 40609:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 40610:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 40611:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 40612:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 40613:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 40614:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 40615:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 40616:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 40617:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 40618:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 40619:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 40620:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 40621:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 40622:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 40623:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 40624:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 40625:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 40626:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 40627:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 40628:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 40629:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 40630:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 40631:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 40632:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 40633:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 40634:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 40635:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 40636:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 40637:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 40638:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 40639:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 40640:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 40641:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 40642:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 40643:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 40644:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 40645:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 40646:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 40647:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 40648:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 40649:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 40650:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 40651:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 40652:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 40653:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 40654:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 40655:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 40656:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 40657:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 40658:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 40659:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 40660:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 40661:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 40662:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 40663:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 40664:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 40665:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 40666:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 40667:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 40668:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 40669:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 40670:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 40671:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 40672:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 40673:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 40674:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 40675:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 40676:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 40677:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 40678:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 40679:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 40680:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 40681:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 40682:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 40683:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 40684:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 40685:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 40686:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 40687:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 40688:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 40689:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 40690:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 40691:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 40692:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 40693:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 40694:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 40695:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 40696:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 40697:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 40698:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 40699:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 40700:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 40701:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 40702:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 40703:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 40704:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 40705:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 40706:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 40707:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 40708:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 40709:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 40710:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 40711:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 40712:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 40713:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 40714:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 40715:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 40716:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 40717:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 40718:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 40719:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 40720:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 40721:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 40722:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 40723:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 40724:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 40725:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 40726:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 40727:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 40728:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 40729:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 40730:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 40731:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 40732:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 40733:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 40734:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 40735:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 40736:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 40737:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 40738:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 40739:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 40740:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 40741:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 40742:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 40743:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 40744:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 40745:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 40746:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 40747:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 40748:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 40749:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 40750:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 40751:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 40752:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 40753:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 40754:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 40755:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 40756:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 40757:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 40758:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 40759:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 40760:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 40761:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 40762:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 40763:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 40764:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 40765:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 40766:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 40767:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 40768:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 40769:22]
  wire  invx142 = ~x142; // @[Snxn100k.scala 40770:17]
  wire  t143 = x142 + invx142; // @[Snxn100k.scala 40771:22]
  wire  inv143 = ~t143; // @[Snxn100k.scala 40772:17]
  wire  x143 = t143 ^ inv143; // @[Snxn100k.scala 40773:22]
  wire  invx143 = ~x143; // @[Snxn100k.scala 40774:17]
  wire  t144 = x143 + invx143; // @[Snxn100k.scala 40775:22]
  wire  inv144 = ~t144; // @[Snxn100k.scala 40776:17]
  wire  x144 = t144 ^ inv144; // @[Snxn100k.scala 40777:22]
  wire  invx144 = ~x144; // @[Snxn100k.scala 40778:17]
  wire  t145 = x144 + invx144; // @[Snxn100k.scala 40779:22]
  wire  inv145 = ~t145; // @[Snxn100k.scala 40780:17]
  wire  x145 = t145 ^ inv145; // @[Snxn100k.scala 40781:22]
  wire  invx145 = ~x145; // @[Snxn100k.scala 40782:17]
  wire  t146 = x145 + invx145; // @[Snxn100k.scala 40783:22]
  wire  inv146 = ~t146; // @[Snxn100k.scala 40784:17]
  wire  x146 = t146 ^ inv146; // @[Snxn100k.scala 40785:22]
  wire  invx146 = ~x146; // @[Snxn100k.scala 40786:17]
  wire  t147 = x146 + invx146; // @[Snxn100k.scala 40787:22]
  wire  inv147 = ~t147; // @[Snxn100k.scala 40788:17]
  wire  x147 = t147 ^ inv147; // @[Snxn100k.scala 40789:22]
  wire  invx147 = ~x147; // @[Snxn100k.scala 40790:17]
  wire  t148 = x147 + invx147; // @[Snxn100k.scala 40791:22]
  wire  inv148 = ~t148; // @[Snxn100k.scala 40792:17]
  wire  x148 = t148 ^ inv148; // @[Snxn100k.scala 40793:22]
  assign io_z = ~x148; // @[Snxn100k.scala 40794:17]
endmodule
module SnxnLv3Inst17(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst68_io_a; // @[Snxn100k.scala 11552:34]
  wire  inst_SnxnLv4Inst68_io_b; // @[Snxn100k.scala 11552:34]
  wire  inst_SnxnLv4Inst68_io_z; // @[Snxn100k.scala 11552:34]
  wire  inst_SnxnLv4Inst69_io_a; // @[Snxn100k.scala 11556:34]
  wire  inst_SnxnLv4Inst69_io_b; // @[Snxn100k.scala 11556:34]
  wire  inst_SnxnLv4Inst69_io_z; // @[Snxn100k.scala 11556:34]
  wire  inst_SnxnLv4Inst70_io_a; // @[Snxn100k.scala 11560:34]
  wire  inst_SnxnLv4Inst70_io_b; // @[Snxn100k.scala 11560:34]
  wire  inst_SnxnLv4Inst70_io_z; // @[Snxn100k.scala 11560:34]
  wire  inst_SnxnLv4Inst71_io_a; // @[Snxn100k.scala 11564:34]
  wire  inst_SnxnLv4Inst71_io_b; // @[Snxn100k.scala 11564:34]
  wire  inst_SnxnLv4Inst71_io_z; // @[Snxn100k.scala 11564:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst68_io_z + inst_SnxnLv4Inst69_io_z; // @[Snxn100k.scala 11568:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst70_io_z; // @[Snxn100k.scala 11568:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst71_io_z; // @[Snxn100k.scala 11568:89]
  SnxnLv4Inst6 inst_SnxnLv4Inst68 ( // @[Snxn100k.scala 11552:34]
    .io_a(inst_SnxnLv4Inst68_io_a),
    .io_b(inst_SnxnLv4Inst68_io_b),
    .io_z(inst_SnxnLv4Inst68_io_z)
  );
  SnxnLv4Inst69 inst_SnxnLv4Inst69 ( // @[Snxn100k.scala 11556:34]
    .io_a(inst_SnxnLv4Inst69_io_a),
    .io_b(inst_SnxnLv4Inst69_io_b),
    .io_z(inst_SnxnLv4Inst69_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst70 ( // @[Snxn100k.scala 11560:34]
    .io_a(inst_SnxnLv4Inst70_io_a),
    .io_b(inst_SnxnLv4Inst70_io_b),
    .io_z(inst_SnxnLv4Inst70_io_z)
  );
  SnxnLv4Inst71 inst_SnxnLv4Inst71 ( // @[Snxn100k.scala 11564:34]
    .io_a(inst_SnxnLv4Inst71_io_a),
    .io_b(inst_SnxnLv4Inst71_io_b),
    .io_z(inst_SnxnLv4Inst71_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11569:15]
  assign inst_SnxnLv4Inst68_io_a = io_a; // @[Snxn100k.scala 11553:27]
  assign inst_SnxnLv4Inst68_io_b = io_b; // @[Snxn100k.scala 11554:27]
  assign inst_SnxnLv4Inst69_io_a = io_a; // @[Snxn100k.scala 11557:27]
  assign inst_SnxnLv4Inst69_io_b = io_b; // @[Snxn100k.scala 11558:27]
  assign inst_SnxnLv4Inst70_io_a = io_a; // @[Snxn100k.scala 11561:27]
  assign inst_SnxnLv4Inst70_io_b = io_b; // @[Snxn100k.scala 11562:27]
  assign inst_SnxnLv4Inst71_io_a = io_a; // @[Snxn100k.scala 11565:27]
  assign inst_SnxnLv4Inst71_io_b = io_b; // @[Snxn100k.scala 11566:27]
endmodule
module SnxnLv4Inst72(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 41217:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 41218:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 41219:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 41220:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 41221:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 41222:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 41223:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 41224:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 41225:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 41226:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 41227:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 41228:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 41229:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 41230:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 41231:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 41232:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 41233:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 41234:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 41235:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 41236:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 41237:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 41238:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 41239:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 41240:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 41241:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 41242:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 41243:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 41244:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 41245:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 41246:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 41247:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 41248:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 41249:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 41250:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 41251:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 41252:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 41253:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 41254:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 41255:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 41256:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 41257:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 41258:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 41259:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 41260:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 41261:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 41262:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 41263:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 41264:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 41265:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 41266:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 41267:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 41268:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 41269:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 41270:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 41271:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 41272:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 41273:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 41274:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 41275:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 41276:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 41277:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 41278:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 41279:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 41280:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 41281:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 41282:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 41283:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 41284:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 41285:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 41286:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 41287:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 41288:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 41289:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 41290:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 41291:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 41292:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 41293:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 41294:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 41295:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 41296:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 41297:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 41298:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 41299:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 41300:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 41301:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 41302:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 41303:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 41304:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 41305:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 41306:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 41307:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 41308:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 41309:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 41310:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 41311:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 41312:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 41313:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 41314:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 41315:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 41316:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 41317:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 41318:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 41319:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 41320:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 41321:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 41322:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 41323:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 41324:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 41325:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 41326:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 41327:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 41328:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 41329:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 41330:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 41331:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 41332:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 41333:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 41334:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 41335:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 41336:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 41337:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 41338:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 41339:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 41340:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 41341:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 41342:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 41343:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 41344:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 41345:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 41346:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 41347:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 41348:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 41349:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 41350:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 41351:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 41352:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 41353:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 41354:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 41355:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 41356:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 41357:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 41358:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 41359:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 41360:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 41361:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 41362:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 41363:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 41364:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 41365:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 41366:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 41367:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 41368:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 41369:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 41370:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 41371:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 41372:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 41373:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 41374:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 41375:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 41376:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 41377:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 41378:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 41379:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 41380:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 41381:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 41382:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 41383:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 41384:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 41385:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 41386:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 41387:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 41388:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 41389:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 41390:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 41391:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 41392:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 41393:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 41394:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 41395:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 41396:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 41397:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 41398:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 41399:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 41400:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 41401:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 41402:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 41403:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 41404:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 41405:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 41406:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 41407:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 41408:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 41409:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 41410:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 41411:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 41412:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 41413:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 41414:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 41415:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 41416:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 41417:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 41418:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 41419:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 41420:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 41421:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 41422:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 41423:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 41424:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 41425:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 41426:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 41427:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 41428:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 41429:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 41430:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 41431:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 41432:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 41433:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 41434:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 41435:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 41436:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 41437:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 41438:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 41439:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 41440:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 41441:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 41442:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 41443:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 41444:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 41445:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 41446:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 41447:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 41448:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 41449:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 41450:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 41451:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 41452:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 41453:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 41454:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 41455:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 41456:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 41457:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 41458:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 41459:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 41460:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 41461:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 41462:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 41463:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 41464:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 41465:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 41466:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 41467:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 41468:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 41469:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 41470:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 41471:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 41472:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 41473:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 41474:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 41475:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 41476:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 41477:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 41478:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 41479:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 41480:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 41481:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 41482:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 41483:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 41484:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 41485:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 41486:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 41487:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 41488:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 41489:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 41490:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 41491:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 41492:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 41493:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 41494:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 41495:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 41496:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 41497:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 41498:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 41499:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 41500:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 41501:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 41502:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 41503:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 41504:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 41505:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 41506:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 41507:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 41508:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 41509:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 41510:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 41511:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 41512:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 41513:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 41514:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 41515:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 41516:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 41517:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 41518:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 41519:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 41520:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 41521:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 41522:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 41523:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 41524:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 41525:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 41526:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 41527:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 41528:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 41529:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 41530:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 41531:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 41532:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 41533:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 41534:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 41535:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 41536:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 41537:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 41538:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 41539:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 41540:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 41541:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 41542:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 41543:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 41544:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 41545:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 41546:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 41547:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 41548:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 41549:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 41550:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 41551:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 41552:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 41553:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 41554:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 41555:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 41556:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 41557:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 41558:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 41559:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 41560:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 41561:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 41562:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 41563:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 41564:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 41565:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 41566:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 41567:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 41568:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 41569:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 41570:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 41571:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 41572:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 41573:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 41574:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 41575:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 41576:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 41577:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 41578:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 41579:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 41580:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 41581:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 41582:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 41583:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 41584:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 41585:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 41586:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 41587:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 41588:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 41589:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 41590:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 41591:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 41592:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 41593:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 41594:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 41595:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 41596:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 41597:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 41598:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 41599:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 41600:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 41601:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 41602:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 41603:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 41604:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 41605:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 41606:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 41607:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 41608:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 41609:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 41610:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 41611:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 41612:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 41613:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 41614:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 41615:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 41616:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 41617:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 41618:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 41619:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 41620:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 41621:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 41622:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 41623:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 41624:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 41625:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 41626:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 41627:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 41628:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 41629:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 41630:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 41631:22]
  assign io_z = ~x103; // @[Snxn100k.scala 41632:17]
endmodule
module SnxnLv4Inst74(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 40805:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 40806:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 40807:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 40808:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 40809:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 40810:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 40811:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 40812:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 40813:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 40814:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 40815:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 40816:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 40817:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 40818:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 40819:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 40820:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 40821:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 40822:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 40823:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 40824:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 40825:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 40826:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 40827:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 40828:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 40829:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 40830:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 40831:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 40832:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 40833:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 40834:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 40835:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 40836:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 40837:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 40838:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 40839:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 40840:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 40841:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 40842:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 40843:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 40844:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 40845:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 40846:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 40847:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 40848:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 40849:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 40850:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 40851:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 40852:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 40853:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 40854:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 40855:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 40856:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 40857:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 40858:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 40859:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 40860:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 40861:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 40862:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 40863:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 40864:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 40865:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 40866:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 40867:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 40868:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 40869:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 40870:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 40871:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 40872:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 40873:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 40874:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 40875:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 40876:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 40877:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 40878:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 40879:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 40880:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 40881:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 40882:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 40883:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 40884:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 40885:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 40886:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 40887:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 40888:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 40889:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 40890:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 40891:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 40892:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 40893:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 40894:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 40895:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 40896:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 40897:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 40898:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 40899:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 40900:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 40901:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 40902:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 40903:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 40904:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 40905:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 40906:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 40907:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 40908:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 40909:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 40910:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 40911:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 40912:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 40913:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 40914:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 40915:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 40916:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 40917:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 40918:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 40919:20]
  assign io_z = ~x28; // @[Snxn100k.scala 40920:16]
endmodule
module SnxnLv3Inst18(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst72_io_a; // @[Snxn100k.scala 11939:34]
  wire  inst_SnxnLv4Inst72_io_b; // @[Snxn100k.scala 11939:34]
  wire  inst_SnxnLv4Inst72_io_z; // @[Snxn100k.scala 11939:34]
  wire  inst_SnxnLv4Inst73_io_a; // @[Snxn100k.scala 11943:34]
  wire  inst_SnxnLv4Inst73_io_b; // @[Snxn100k.scala 11943:34]
  wire  inst_SnxnLv4Inst73_io_z; // @[Snxn100k.scala 11943:34]
  wire  inst_SnxnLv4Inst74_io_a; // @[Snxn100k.scala 11947:34]
  wire  inst_SnxnLv4Inst74_io_b; // @[Snxn100k.scala 11947:34]
  wire  inst_SnxnLv4Inst74_io_z; // @[Snxn100k.scala 11947:34]
  wire  inst_SnxnLv4Inst75_io_a; // @[Snxn100k.scala 11951:34]
  wire  inst_SnxnLv4Inst75_io_b; // @[Snxn100k.scala 11951:34]
  wire  inst_SnxnLv4Inst75_io_z; // @[Snxn100k.scala 11951:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst72_io_z + inst_SnxnLv4Inst73_io_z; // @[Snxn100k.scala 11955:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst74_io_z; // @[Snxn100k.scala 11955:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst75_io_z; // @[Snxn100k.scala 11955:89]
  SnxnLv4Inst72 inst_SnxnLv4Inst72 ( // @[Snxn100k.scala 11939:34]
    .io_a(inst_SnxnLv4Inst72_io_a),
    .io_b(inst_SnxnLv4Inst72_io_b),
    .io_z(inst_SnxnLv4Inst72_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst73 ( // @[Snxn100k.scala 11943:34]
    .io_a(inst_SnxnLv4Inst73_io_a),
    .io_b(inst_SnxnLv4Inst73_io_b),
    .io_z(inst_SnxnLv4Inst73_io_z)
  );
  SnxnLv4Inst74 inst_SnxnLv4Inst74 ( // @[Snxn100k.scala 11947:34]
    .io_a(inst_SnxnLv4Inst74_io_a),
    .io_b(inst_SnxnLv4Inst74_io_b),
    .io_z(inst_SnxnLv4Inst74_io_z)
  );
  SnxnLv4Inst46 inst_SnxnLv4Inst75 ( // @[Snxn100k.scala 11951:34]
    .io_a(inst_SnxnLv4Inst75_io_a),
    .io_b(inst_SnxnLv4Inst75_io_b),
    .io_z(inst_SnxnLv4Inst75_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11956:15]
  assign inst_SnxnLv4Inst72_io_a = io_a; // @[Snxn100k.scala 11940:27]
  assign inst_SnxnLv4Inst72_io_b = io_b; // @[Snxn100k.scala 11941:27]
  assign inst_SnxnLv4Inst73_io_a = io_a; // @[Snxn100k.scala 11944:27]
  assign inst_SnxnLv4Inst73_io_b = io_b; // @[Snxn100k.scala 11945:27]
  assign inst_SnxnLv4Inst74_io_a = io_a; // @[Snxn100k.scala 11948:27]
  assign inst_SnxnLv4Inst74_io_b = io_b; // @[Snxn100k.scala 11949:27]
  assign inst_SnxnLv4Inst75_io_a = io_a; // @[Snxn100k.scala 11952:27]
  assign inst_SnxnLv4Inst75_io_b = io_b; // @[Snxn100k.scala 11953:27]
endmodule
module SnxnLv4Inst76(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 44023:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 44024:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 44025:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 44026:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 44027:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 44028:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 44029:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 44030:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 44031:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 44032:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 44033:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 44034:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 44035:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 44036:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 44037:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 44038:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 44039:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 44040:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 44041:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 44042:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 44043:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 44044:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 44045:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 44046:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 44047:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 44048:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 44049:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 44050:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 44051:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 44052:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 44053:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 44054:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 44055:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 44056:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 44057:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 44058:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 44059:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 44060:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 44061:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 44062:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 44063:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 44064:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 44065:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 44066:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 44067:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 44068:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 44069:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 44070:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 44071:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 44072:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 44073:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 44074:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 44075:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 44076:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 44077:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 44078:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 44079:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 44080:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 44081:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 44082:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 44083:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 44084:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 44085:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 44086:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 44087:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 44088:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 44089:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 44090:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 44091:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 44092:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 44093:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 44094:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 44095:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 44096:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 44097:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 44098:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 44099:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 44100:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 44101:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 44102:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 44103:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 44104:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 44105:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 44106:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 44107:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 44108:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 44109:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 44110:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 44111:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 44112:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 44113:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 44114:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 44115:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 44116:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 44117:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 44118:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 44119:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 44120:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 44121:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 44122:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 44123:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 44124:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 44125:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 44126:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 44127:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 44128:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 44129:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 44130:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 44131:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 44132:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 44133:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 44134:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 44135:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 44136:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 44137:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 44138:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 44139:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 44140:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 44141:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 44142:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 44143:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 44144:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 44145:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 44146:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 44147:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 44148:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 44149:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 44150:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 44151:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 44152:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 44153:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 44154:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 44155:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 44156:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 44157:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 44158:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 44159:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 44160:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 44161:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 44162:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 44163:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 44164:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 44165:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 44166:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 44167:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 44168:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 44169:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 44170:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 44171:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 44172:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 44173:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 44174:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 44175:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 44176:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 44177:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 44178:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 44179:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 44180:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 44181:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 44182:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 44183:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 44184:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 44185:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 44186:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 44187:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 44188:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 44189:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 44190:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 44191:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 44192:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 44193:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 44194:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 44195:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 44196:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 44197:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 44198:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 44199:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 44200:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 44201:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 44202:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 44203:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 44204:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 44205:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 44206:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 44207:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 44208:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 44209:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 44210:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 44211:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 44212:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 44213:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 44214:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 44215:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 44216:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 44217:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 44218:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 44219:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 44220:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 44221:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 44222:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 44223:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 44224:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 44225:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 44226:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 44227:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 44228:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 44229:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 44230:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 44231:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 44232:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 44233:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 44234:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 44235:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 44236:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 44237:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 44238:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 44239:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 44240:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 44241:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 44242:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 44243:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 44244:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 44245:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 44246:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 44247:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 44248:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 44249:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 44250:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 44251:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 44252:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 44253:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 44254:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 44255:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 44256:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 44257:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 44258:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 44259:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 44260:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 44261:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 44262:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 44263:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 44264:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 44265:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 44266:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 44267:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 44268:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 44269:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 44270:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 44271:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 44272:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 44273:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 44274:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 44275:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 44276:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 44277:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 44278:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 44279:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 44280:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 44281:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 44282:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 44283:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 44284:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 44285:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 44286:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 44287:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 44288:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 44289:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 44290:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 44291:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 44292:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 44293:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 44294:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 44295:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 44296:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 44297:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 44298:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 44299:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 44300:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 44301:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 44302:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 44303:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 44304:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 44305:20]
  assign io_z = ~x70; // @[Snxn100k.scala 44306:16]
endmodule
module SnxnLv4Inst77(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 43821:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 43822:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 43823:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 43824:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 43825:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 43826:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 43827:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 43828:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 43829:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 43830:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 43831:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 43832:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 43833:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 43834:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 43835:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 43836:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 43837:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 43838:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 43839:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 43840:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 43841:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 43842:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 43843:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 43844:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 43845:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 43846:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 43847:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 43848:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 43849:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 43850:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 43851:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 43852:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 43853:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 43854:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 43855:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 43856:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 43857:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 43858:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 43859:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 43860:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 43861:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 43862:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 43863:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 43864:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 43865:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 43866:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 43867:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 43868:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 43869:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 43870:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 43871:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 43872:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 43873:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 43874:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 43875:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 43876:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 43877:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 43878:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 43879:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 43880:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 43881:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 43882:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 43883:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 43884:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 43885:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 43886:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 43887:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 43888:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 43889:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 43890:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 43891:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 43892:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 43893:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 43894:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 43895:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 43896:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 43897:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 43898:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 43899:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 43900:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 43901:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 43902:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 43903:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 43904:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 43905:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 43906:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 43907:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 43908:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 43909:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 43910:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 43911:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 43912:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 43913:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 43914:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 43915:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 43916:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 43917:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 43918:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 43919:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 43920:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 43921:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 43922:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 43923:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 43924:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 43925:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 43926:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 43927:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 43928:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 43929:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 43930:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 43931:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 43932:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 43933:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 43934:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 43935:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 43936:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 43937:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 43938:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 43939:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 43940:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 43941:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 43942:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 43943:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 43944:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 43945:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 43946:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 43947:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 43948:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 43949:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 43950:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 43951:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 43952:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 43953:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 43954:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 43955:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 43956:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 43957:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 43958:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 43959:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 43960:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 43961:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 43962:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 43963:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 43964:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 43965:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 43966:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 43967:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 43968:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 43969:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 43970:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 43971:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 43972:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 43973:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 43974:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 43975:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 43976:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 43977:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 43978:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 43979:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 43980:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 43981:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 43982:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 43983:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 43984:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 43985:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 43986:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 43987:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 43988:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 43989:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 43990:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 43991:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 43992:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 43993:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 43994:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 43995:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 43996:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 43997:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 43998:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 43999:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 44000:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 44001:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 44002:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 44003:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 44004:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 44005:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 44006:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 44007:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 44008:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 44009:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 44010:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 44011:20]
  assign io_z = ~x47; // @[Snxn100k.scala 44012:16]
endmodule
module SnxnLv4Inst78(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 43643:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 43644:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 43645:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 43646:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 43647:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 43648:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 43649:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 43650:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 43651:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 43652:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 43653:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 43654:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 43655:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 43656:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 43657:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 43658:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 43659:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 43660:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 43661:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 43662:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 43663:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 43664:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 43665:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 43666:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 43667:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 43668:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 43669:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 43670:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 43671:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 43672:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 43673:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 43674:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 43675:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 43676:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 43677:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 43678:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 43679:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 43680:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 43681:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 43682:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 43683:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 43684:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 43685:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 43686:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 43687:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 43688:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 43689:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 43690:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 43691:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 43692:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 43693:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 43694:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 43695:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 43696:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 43697:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 43698:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 43699:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 43700:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 43701:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 43702:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 43703:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 43704:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 43705:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 43706:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 43707:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 43708:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 43709:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 43710:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 43711:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 43712:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 43713:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 43714:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 43715:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 43716:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 43717:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 43718:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 43719:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 43720:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 43721:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 43722:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 43723:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 43724:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 43725:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 43726:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 43727:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 43728:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 43729:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 43730:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 43731:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 43732:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 43733:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 43734:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 43735:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 43736:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 43737:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 43738:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 43739:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 43740:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 43741:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 43742:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 43743:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 43744:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 43745:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 43746:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 43747:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 43748:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 43749:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 43750:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 43751:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 43752:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 43753:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 43754:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 43755:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 43756:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 43757:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 43758:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 43759:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 43760:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 43761:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 43762:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 43763:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 43764:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 43765:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 43766:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 43767:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 43768:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 43769:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 43770:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 43771:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 43772:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 43773:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 43774:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 43775:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 43776:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 43777:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 43778:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 43779:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 43780:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 43781:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 43782:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 43783:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 43784:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 43785:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 43786:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 43787:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 43788:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 43789:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 43790:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 43791:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 43792:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 43793:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 43794:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 43795:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 43796:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 43797:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 43798:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 43799:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 43800:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 43801:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 43802:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 43803:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 43804:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 43805:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 43806:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 43807:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 43808:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 43809:20]
  assign io_z = ~x41; // @[Snxn100k.scala 43810:16]
endmodule
module SnxnLv3Inst19(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst76_io_a; // @[Snxn100k.scala 12917:34]
  wire  inst_SnxnLv4Inst76_io_b; // @[Snxn100k.scala 12917:34]
  wire  inst_SnxnLv4Inst76_io_z; // @[Snxn100k.scala 12917:34]
  wire  inst_SnxnLv4Inst77_io_a; // @[Snxn100k.scala 12921:34]
  wire  inst_SnxnLv4Inst77_io_b; // @[Snxn100k.scala 12921:34]
  wire  inst_SnxnLv4Inst77_io_z; // @[Snxn100k.scala 12921:34]
  wire  inst_SnxnLv4Inst78_io_a; // @[Snxn100k.scala 12925:34]
  wire  inst_SnxnLv4Inst78_io_b; // @[Snxn100k.scala 12925:34]
  wire  inst_SnxnLv4Inst78_io_z; // @[Snxn100k.scala 12925:34]
  wire  inst_SnxnLv4Inst79_io_a; // @[Snxn100k.scala 12929:34]
  wire  inst_SnxnLv4Inst79_io_b; // @[Snxn100k.scala 12929:34]
  wire  inst_SnxnLv4Inst79_io_z; // @[Snxn100k.scala 12929:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst76_io_z + inst_SnxnLv4Inst77_io_z; // @[Snxn100k.scala 12933:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst78_io_z; // @[Snxn100k.scala 12933:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst79_io_z; // @[Snxn100k.scala 12933:89]
  SnxnLv4Inst76 inst_SnxnLv4Inst76 ( // @[Snxn100k.scala 12917:34]
    .io_a(inst_SnxnLv4Inst76_io_a),
    .io_b(inst_SnxnLv4Inst76_io_b),
    .io_z(inst_SnxnLv4Inst76_io_z)
  );
  SnxnLv4Inst77 inst_SnxnLv4Inst77 ( // @[Snxn100k.scala 12921:34]
    .io_a(inst_SnxnLv4Inst77_io_a),
    .io_b(inst_SnxnLv4Inst77_io_b),
    .io_z(inst_SnxnLv4Inst77_io_z)
  );
  SnxnLv4Inst78 inst_SnxnLv4Inst78 ( // @[Snxn100k.scala 12925:34]
    .io_a(inst_SnxnLv4Inst78_io_a),
    .io_b(inst_SnxnLv4Inst78_io_b),
    .io_z(inst_SnxnLv4Inst78_io_z)
  );
  SnxnLv4Inst59 inst_SnxnLv4Inst79 ( // @[Snxn100k.scala 12929:34]
    .io_a(inst_SnxnLv4Inst79_io_a),
    .io_b(inst_SnxnLv4Inst79_io_b),
    .io_z(inst_SnxnLv4Inst79_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 12934:15]
  assign inst_SnxnLv4Inst76_io_a = io_a; // @[Snxn100k.scala 12918:27]
  assign inst_SnxnLv4Inst76_io_b = io_b; // @[Snxn100k.scala 12919:27]
  assign inst_SnxnLv4Inst77_io_a = io_a; // @[Snxn100k.scala 12922:27]
  assign inst_SnxnLv4Inst77_io_b = io_b; // @[Snxn100k.scala 12923:27]
  assign inst_SnxnLv4Inst78_io_a = io_a; // @[Snxn100k.scala 12926:27]
  assign inst_SnxnLv4Inst78_io_b = io_b; // @[Snxn100k.scala 12927:27]
  assign inst_SnxnLv4Inst79_io_a = io_a; // @[Snxn100k.scala 12930:27]
  assign inst_SnxnLv4Inst79_io_b = io_b; // @[Snxn100k.scala 12931:27]
endmodule
module SnxnLv2Inst4(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst16_io_a; // @[Snxn100k.scala 2694:34]
  wire  inst_SnxnLv3Inst16_io_b; // @[Snxn100k.scala 2694:34]
  wire  inst_SnxnLv3Inst16_io_z; // @[Snxn100k.scala 2694:34]
  wire  inst_SnxnLv3Inst17_io_a; // @[Snxn100k.scala 2698:34]
  wire  inst_SnxnLv3Inst17_io_b; // @[Snxn100k.scala 2698:34]
  wire  inst_SnxnLv3Inst17_io_z; // @[Snxn100k.scala 2698:34]
  wire  inst_SnxnLv3Inst18_io_a; // @[Snxn100k.scala 2702:34]
  wire  inst_SnxnLv3Inst18_io_b; // @[Snxn100k.scala 2702:34]
  wire  inst_SnxnLv3Inst18_io_z; // @[Snxn100k.scala 2702:34]
  wire  inst_SnxnLv3Inst19_io_a; // @[Snxn100k.scala 2706:34]
  wire  inst_SnxnLv3Inst19_io_b; // @[Snxn100k.scala 2706:34]
  wire  inst_SnxnLv3Inst19_io_z; // @[Snxn100k.scala 2706:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst16_io_z + inst_SnxnLv3Inst17_io_z; // @[Snxn100k.scala 2710:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst18_io_z; // @[Snxn100k.scala 2710:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst19_io_z; // @[Snxn100k.scala 2710:89]
  SnxnLv3Inst16 inst_SnxnLv3Inst16 ( // @[Snxn100k.scala 2694:34]
    .io_a(inst_SnxnLv3Inst16_io_a),
    .io_b(inst_SnxnLv3Inst16_io_b),
    .io_z(inst_SnxnLv3Inst16_io_z)
  );
  SnxnLv3Inst17 inst_SnxnLv3Inst17 ( // @[Snxn100k.scala 2698:34]
    .io_a(inst_SnxnLv3Inst17_io_a),
    .io_b(inst_SnxnLv3Inst17_io_b),
    .io_z(inst_SnxnLv3Inst17_io_z)
  );
  SnxnLv3Inst18 inst_SnxnLv3Inst18 ( // @[Snxn100k.scala 2702:34]
    .io_a(inst_SnxnLv3Inst18_io_a),
    .io_b(inst_SnxnLv3Inst18_io_b),
    .io_z(inst_SnxnLv3Inst18_io_z)
  );
  SnxnLv3Inst19 inst_SnxnLv3Inst19 ( // @[Snxn100k.scala 2706:34]
    .io_a(inst_SnxnLv3Inst19_io_a),
    .io_b(inst_SnxnLv3Inst19_io_b),
    .io_z(inst_SnxnLv3Inst19_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 2711:15]
  assign inst_SnxnLv3Inst16_io_a = io_a; // @[Snxn100k.scala 2695:27]
  assign inst_SnxnLv3Inst16_io_b = io_b; // @[Snxn100k.scala 2696:27]
  assign inst_SnxnLv3Inst17_io_a = io_a; // @[Snxn100k.scala 2699:27]
  assign inst_SnxnLv3Inst17_io_b = io_b; // @[Snxn100k.scala 2700:27]
  assign inst_SnxnLv3Inst18_io_a = io_a; // @[Snxn100k.scala 2703:27]
  assign inst_SnxnLv3Inst18_io_b = io_b; // @[Snxn100k.scala 2704:27]
  assign inst_SnxnLv3Inst19_io_a = io_a; // @[Snxn100k.scala 2707:27]
  assign inst_SnxnLv3Inst19_io_b = io_b; // @[Snxn100k.scala 2708:27]
endmodule
module SnxnLv3Inst20(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst80_io_a; // @[Snxn100k.scala 10739:34]
  wire  inst_SnxnLv4Inst80_io_b; // @[Snxn100k.scala 10739:34]
  wire  inst_SnxnLv4Inst80_io_z; // @[Snxn100k.scala 10739:34]
  wire  inst_SnxnLv4Inst81_io_a; // @[Snxn100k.scala 10743:34]
  wire  inst_SnxnLv4Inst81_io_b; // @[Snxn100k.scala 10743:34]
  wire  inst_SnxnLv4Inst81_io_z; // @[Snxn100k.scala 10743:34]
  wire  inst_SnxnLv4Inst82_io_a; // @[Snxn100k.scala 10747:34]
  wire  inst_SnxnLv4Inst82_io_b; // @[Snxn100k.scala 10747:34]
  wire  inst_SnxnLv4Inst82_io_z; // @[Snxn100k.scala 10747:34]
  wire  inst_SnxnLv4Inst83_io_a; // @[Snxn100k.scala 10751:34]
  wire  inst_SnxnLv4Inst83_io_b; // @[Snxn100k.scala 10751:34]
  wire  inst_SnxnLv4Inst83_io_z; // @[Snxn100k.scala 10751:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst80_io_z + inst_SnxnLv4Inst81_io_z; // @[Snxn100k.scala 10755:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst82_io_z; // @[Snxn100k.scala 10755:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst83_io_z; // @[Snxn100k.scala 10755:89]
  SnxnLv4Inst47 inst_SnxnLv4Inst80 ( // @[Snxn100k.scala 10739:34]
    .io_a(inst_SnxnLv4Inst80_io_a),
    .io_b(inst_SnxnLv4Inst80_io_b),
    .io_z(inst_SnxnLv4Inst80_io_z)
  );
  SnxnLv4Inst48 inst_SnxnLv4Inst81 ( // @[Snxn100k.scala 10743:34]
    .io_a(inst_SnxnLv4Inst81_io_a),
    .io_b(inst_SnxnLv4Inst81_io_b),
    .io_z(inst_SnxnLv4Inst81_io_z)
  );
  SnxnLv4Inst31 inst_SnxnLv4Inst82 ( // @[Snxn100k.scala 10747:34]
    .io_a(inst_SnxnLv4Inst82_io_a),
    .io_b(inst_SnxnLv4Inst82_io_b),
    .io_z(inst_SnxnLv4Inst82_io_z)
  );
  SnxnLv4Inst12 inst_SnxnLv4Inst83 ( // @[Snxn100k.scala 10751:34]
    .io_a(inst_SnxnLv4Inst83_io_a),
    .io_b(inst_SnxnLv4Inst83_io_b),
    .io_z(inst_SnxnLv4Inst83_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10756:15]
  assign inst_SnxnLv4Inst80_io_a = io_a; // @[Snxn100k.scala 10740:27]
  assign inst_SnxnLv4Inst80_io_b = io_b; // @[Snxn100k.scala 10741:27]
  assign inst_SnxnLv4Inst81_io_a = io_a; // @[Snxn100k.scala 10744:27]
  assign inst_SnxnLv4Inst81_io_b = io_b; // @[Snxn100k.scala 10745:27]
  assign inst_SnxnLv4Inst82_io_a = io_a; // @[Snxn100k.scala 10748:27]
  assign inst_SnxnLv4Inst82_io_b = io_b; // @[Snxn100k.scala 10749:27]
  assign inst_SnxnLv4Inst83_io_a = io_a; // @[Snxn100k.scala 10752:27]
  assign inst_SnxnLv4Inst83_io_b = io_b; // @[Snxn100k.scala 10753:27]
endmodule
module SnxnLv4Inst84(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 37027:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 37028:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 37029:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 37030:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 37031:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 37032:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 37033:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 37034:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 37035:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 37036:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 37037:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 37038:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 37039:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 37040:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 37041:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 37042:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 37043:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 37044:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 37045:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 37046:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 37047:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 37048:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 37049:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 37050:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 37051:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 37052:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 37053:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 37054:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 37055:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 37056:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 37057:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 37058:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 37059:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 37060:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 37061:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 37062:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 37063:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 37064:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 37065:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 37066:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 37067:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 37068:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 37069:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 37070:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 37071:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 37072:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 37073:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 37074:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 37075:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 37076:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 37077:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 37078:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 37079:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 37080:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 37081:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 37082:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 37083:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 37084:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 37085:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 37086:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 37087:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 37088:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 37089:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 37090:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 37091:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 37092:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 37093:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 37094:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 37095:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 37096:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 37097:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 37098:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 37099:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 37100:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 37101:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 37102:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 37103:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 37104:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 37105:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 37106:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 37107:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 37108:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 37109:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 37110:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 37111:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 37112:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 37113:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 37114:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 37115:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 37116:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 37117:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 37118:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 37119:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 37120:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 37121:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 37122:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 37123:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 37124:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 37125:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 37126:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 37127:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 37128:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 37129:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 37130:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 37131:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 37132:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 37133:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 37134:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 37135:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 37136:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 37137:20]
  assign io_z = ~x27; // @[Snxn100k.scala 37138:16]
endmodule
module SnxnLv4Inst86(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 37149:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 37150:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 37151:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 37152:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 37153:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 37154:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 37155:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 37156:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 37157:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 37158:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 37159:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 37160:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 37161:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 37162:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 37163:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 37164:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 37165:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 37166:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 37167:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 37168:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 37169:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 37170:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 37171:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 37172:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 37173:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 37174:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 37175:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 37176:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 37177:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 37178:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 37179:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 37180:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 37181:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 37182:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 37183:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 37184:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 37185:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 37186:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 37187:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 37188:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 37189:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 37190:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 37191:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 37192:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 37193:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 37194:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 37195:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 37196:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 37197:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 37198:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 37199:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 37200:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 37201:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 37202:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 37203:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 37204:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 37205:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 37206:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 37207:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 37208:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 37209:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 37210:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 37211:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 37212:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 37213:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 37214:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 37215:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 37216:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 37217:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 37218:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 37219:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 37220:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 37221:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 37222:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 37223:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 37224:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 37225:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 37226:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 37227:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 37228:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 37229:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 37230:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 37231:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 37232:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 37233:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 37234:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 37235:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 37236:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 37237:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 37238:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 37239:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 37240:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 37241:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 37242:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 37243:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 37244:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 37245:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 37246:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 37247:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 37248:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 37249:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 37250:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 37251:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 37252:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 37253:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 37254:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 37255:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 37256:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 37257:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 37258:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 37259:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 37260:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 37261:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 37262:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 37263:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 37264:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 37265:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 37266:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 37267:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 37268:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 37269:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 37270:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 37271:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 37272:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 37273:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 37274:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 37275:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 37276:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 37277:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 37278:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 37279:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 37280:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 37281:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 37282:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 37283:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 37284:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 37285:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 37286:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 37287:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 37288:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 37289:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 37290:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 37291:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 37292:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 37293:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 37294:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 37295:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 37296:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 37297:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 37298:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 37299:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 37300:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 37301:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 37302:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 37303:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 37304:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 37305:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 37306:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 37307:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 37308:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 37309:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 37310:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 37311:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 37312:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 37313:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 37314:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 37315:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 37316:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 37317:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 37318:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 37319:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 37320:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 37321:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 37322:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 37323:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 37324:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 37325:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 37326:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 37327:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 37328:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 37329:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 37330:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 37331:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 37332:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 37333:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 37334:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 37335:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 37336:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 37337:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 37338:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 37339:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 37340:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 37341:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 37342:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 37343:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 37344:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 37345:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 37346:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 37347:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 37348:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 37349:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 37350:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 37351:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 37352:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 37353:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 37354:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 37355:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 37356:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 37357:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 37358:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 37359:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 37360:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 37361:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 37362:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 37363:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 37364:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 37365:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 37366:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 37367:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 37368:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 37369:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 37370:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 37371:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 37372:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 37373:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 37374:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 37375:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 37376:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 37377:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 37378:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 37379:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 37380:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 37381:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 37382:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 37383:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 37384:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 37385:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 37386:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 37387:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 37388:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 37389:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 37390:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 37391:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 37392:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 37393:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 37394:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 37395:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 37396:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 37397:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 37398:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 37399:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 37400:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 37401:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 37402:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 37403:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 37404:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 37405:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 37406:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 37407:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 37408:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 37409:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 37410:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 37411:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 37412:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 37413:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 37414:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 37415:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 37416:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 37417:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 37418:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 37419:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 37420:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 37421:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 37422:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 37423:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 37424:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 37425:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 37426:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 37427:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 37428:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 37429:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 37430:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 37431:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 37432:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 37433:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 37434:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 37435:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 37436:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 37437:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 37438:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 37439:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 37440:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 37441:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 37442:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 37443:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 37444:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 37445:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 37446:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 37447:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 37448:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 37449:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 37450:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 37451:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 37452:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 37453:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 37454:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 37455:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 37456:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 37457:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 37458:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 37459:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 37460:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 37461:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 37462:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 37463:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 37464:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 37465:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 37466:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 37467:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 37468:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 37469:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 37470:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 37471:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 37472:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 37473:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 37474:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 37475:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 37476:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 37477:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 37478:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 37479:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 37480:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 37481:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 37482:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 37483:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 37484:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 37485:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 37486:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 37487:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 37488:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 37489:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 37490:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 37491:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 37492:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 37493:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 37494:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 37495:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 37496:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 37497:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 37498:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 37499:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 37500:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 37501:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 37502:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 37503:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 37504:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 37505:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 37506:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 37507:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 37508:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 37509:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 37510:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 37511:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 37512:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 37513:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 37514:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 37515:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 37516:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 37517:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 37518:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 37519:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 37520:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 37521:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 37522:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 37523:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 37524:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 37525:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 37526:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 37527:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 37528:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 37529:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 37530:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 37531:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 37532:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 37533:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 37534:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 37535:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 37536:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 37537:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 37538:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 37539:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 37540:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 37541:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 37542:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 37543:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 37544:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 37545:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 37546:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 37547:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 37548:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 37549:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 37550:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 37551:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 37552:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 37553:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 37554:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 37555:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 37556:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 37557:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 37558:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 37559:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 37560:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 37561:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 37562:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 37563:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 37564:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 37565:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 37566:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 37567:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 37568:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 37569:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 37570:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 37571:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 37572:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 37573:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 37574:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 37575:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 37576:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 37577:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 37578:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 37579:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 37580:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 37581:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 37582:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 37583:22]
  assign io_z = ~x108; // @[Snxn100k.scala 37584:17]
endmodule
module SnxnLv3Inst21(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst84_io_a; // @[Snxn100k.scala 11306:34]
  wire  inst_SnxnLv4Inst84_io_b; // @[Snxn100k.scala 11306:34]
  wire  inst_SnxnLv4Inst84_io_z; // @[Snxn100k.scala 11306:34]
  wire  inst_SnxnLv4Inst85_io_a; // @[Snxn100k.scala 11310:34]
  wire  inst_SnxnLv4Inst85_io_b; // @[Snxn100k.scala 11310:34]
  wire  inst_SnxnLv4Inst85_io_z; // @[Snxn100k.scala 11310:34]
  wire  inst_SnxnLv4Inst86_io_a; // @[Snxn100k.scala 11314:34]
  wire  inst_SnxnLv4Inst86_io_b; // @[Snxn100k.scala 11314:34]
  wire  inst_SnxnLv4Inst86_io_z; // @[Snxn100k.scala 11314:34]
  wire  inst_SnxnLv4Inst87_io_a; // @[Snxn100k.scala 11318:34]
  wire  inst_SnxnLv4Inst87_io_b; // @[Snxn100k.scala 11318:34]
  wire  inst_SnxnLv4Inst87_io_z; // @[Snxn100k.scala 11318:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst84_io_z + inst_SnxnLv4Inst85_io_z; // @[Snxn100k.scala 11322:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst86_io_z; // @[Snxn100k.scala 11322:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst87_io_z; // @[Snxn100k.scala 11322:89]
  SnxnLv4Inst84 inst_SnxnLv4Inst84 ( // @[Snxn100k.scala 11306:34]
    .io_a(inst_SnxnLv4Inst84_io_a),
    .io_b(inst_SnxnLv4Inst84_io_b),
    .io_z(inst_SnxnLv4Inst84_io_z)
  );
  SnxnLv4Inst56 inst_SnxnLv4Inst85 ( // @[Snxn100k.scala 11310:34]
    .io_a(inst_SnxnLv4Inst85_io_a),
    .io_b(inst_SnxnLv4Inst85_io_b),
    .io_z(inst_SnxnLv4Inst85_io_z)
  );
  SnxnLv4Inst86 inst_SnxnLv4Inst86 ( // @[Snxn100k.scala 11314:34]
    .io_a(inst_SnxnLv4Inst86_io_a),
    .io_b(inst_SnxnLv4Inst86_io_b),
    .io_z(inst_SnxnLv4Inst86_io_z)
  );
  SnxnLv4Inst36 inst_SnxnLv4Inst87 ( // @[Snxn100k.scala 11318:34]
    .io_a(inst_SnxnLv4Inst87_io_a),
    .io_b(inst_SnxnLv4Inst87_io_b),
    .io_z(inst_SnxnLv4Inst87_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11323:15]
  assign inst_SnxnLv4Inst84_io_a = io_a; // @[Snxn100k.scala 11307:27]
  assign inst_SnxnLv4Inst84_io_b = io_b; // @[Snxn100k.scala 11308:27]
  assign inst_SnxnLv4Inst85_io_a = io_a; // @[Snxn100k.scala 11311:27]
  assign inst_SnxnLv4Inst85_io_b = io_b; // @[Snxn100k.scala 11312:27]
  assign inst_SnxnLv4Inst86_io_a = io_a; // @[Snxn100k.scala 11315:27]
  assign inst_SnxnLv4Inst86_io_b = io_b; // @[Snxn100k.scala 11316:27]
  assign inst_SnxnLv4Inst87_io_a = io_a; // @[Snxn100k.scala 11319:27]
  assign inst_SnxnLv4Inst87_io_b = io_b; // @[Snxn100k.scala 11320:27]
endmodule
module SnxnLv4Inst90(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 35393:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 35394:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 35395:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 35396:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 35397:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 35398:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 35399:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 35400:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 35401:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 35402:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 35403:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 35404:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 35405:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 35406:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 35407:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 35408:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 35409:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 35410:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 35411:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 35412:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 35413:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 35414:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 35415:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 35416:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 35417:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 35418:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 35419:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 35420:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 35421:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 35422:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 35423:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 35424:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 35425:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 35426:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 35427:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 35428:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 35429:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 35430:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 35431:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 35432:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 35433:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 35434:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 35435:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 35436:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 35437:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 35438:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 35439:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 35440:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 35441:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 35442:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 35443:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 35444:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 35445:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 35446:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 35447:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 35448:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 35449:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 35450:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 35451:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 35452:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 35453:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 35454:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 35455:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 35456:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 35457:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 35458:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 35459:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 35460:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 35461:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 35462:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 35463:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 35464:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 35465:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 35466:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 35467:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 35468:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 35469:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 35470:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 35471:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 35472:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 35473:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 35474:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 35475:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 35476:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 35477:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 35478:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 35479:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 35480:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 35481:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 35482:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 35483:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 35484:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 35485:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 35486:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 35487:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 35488:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 35489:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 35490:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 35491:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 35492:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 35493:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 35494:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 35495:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 35496:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 35497:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 35498:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 35499:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 35500:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 35501:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 35502:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 35503:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 35504:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 35505:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 35506:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 35507:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 35508:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 35509:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 35510:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 35511:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 35512:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 35513:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 35514:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 35515:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 35516:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 35517:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 35518:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 35519:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 35520:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 35521:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 35522:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 35523:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 35524:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 35525:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 35526:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 35527:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 35528:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 35529:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 35530:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 35531:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 35532:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 35533:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 35534:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 35535:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 35536:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 35537:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 35538:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 35539:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 35540:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 35541:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 35542:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 35543:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 35544:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 35545:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 35546:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 35547:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 35548:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 35549:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 35550:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 35551:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 35552:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 35553:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 35554:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 35555:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 35556:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 35557:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 35558:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 35559:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 35560:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 35561:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 35562:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 35563:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 35564:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 35565:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 35566:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 35567:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 35568:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 35569:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 35570:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 35571:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 35572:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 35573:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 35574:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 35575:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 35576:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 35577:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 35578:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 35579:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 35580:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 35581:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 35582:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 35583:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 35584:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 35585:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 35586:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 35587:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 35588:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 35589:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 35590:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 35591:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 35592:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 35593:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 35594:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 35595:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 35596:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 35597:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 35598:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 35599:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 35600:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 35601:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 35602:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 35603:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 35604:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 35605:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 35606:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 35607:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 35608:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 35609:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 35610:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 35611:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 35612:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 35613:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 35614:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 35615:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 35616:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 35617:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 35618:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 35619:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 35620:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 35621:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 35622:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 35623:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 35624:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 35625:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 35626:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 35627:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 35628:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 35629:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 35630:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 35631:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 35632:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 35633:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 35634:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 35635:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 35636:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 35637:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 35638:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 35639:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 35640:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 35641:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 35642:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 35643:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 35644:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 35645:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 35646:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 35647:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 35648:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 35649:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 35650:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 35651:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 35652:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 35653:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 35654:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 35655:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 35656:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 35657:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 35658:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 35659:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 35660:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 35661:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 35662:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 35663:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 35664:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 35665:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 35666:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 35667:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 35668:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 35669:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 35670:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 35671:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 35672:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 35673:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 35674:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 35675:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 35676:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 35677:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 35678:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 35679:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 35680:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 35681:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 35682:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 35683:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 35684:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 35685:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 35686:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 35687:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 35688:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 35689:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 35690:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 35691:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 35692:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 35693:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 35694:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 35695:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 35696:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 35697:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 35698:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 35699:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 35700:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 35701:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 35702:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 35703:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 35704:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 35705:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 35706:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 35707:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 35708:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 35709:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 35710:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 35711:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 35712:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 35713:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 35714:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 35715:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 35716:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 35717:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 35718:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 35719:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 35720:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 35721:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 35722:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 35723:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 35724:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 35725:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 35726:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 35727:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 35728:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 35729:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 35730:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 35731:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 35732:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 35733:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 35734:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 35735:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 35736:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 35737:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 35738:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 35739:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 35740:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 35741:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 35742:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 35743:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 35744:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 35745:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 35746:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 35747:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 35748:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 35749:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 35750:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 35751:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 35752:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 35753:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 35754:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 35755:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 35756:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 35757:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 35758:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 35759:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 35760:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 35761:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 35762:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 35763:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 35764:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 35765:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 35766:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 35767:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 35768:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 35769:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 35770:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 35771:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 35772:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 35773:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 35774:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 35775:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 35776:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 35777:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 35778:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 35779:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 35780:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 35781:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 35782:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 35783:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 35784:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 35785:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 35786:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 35787:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 35788:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 35789:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 35790:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 35791:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 35792:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 35793:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 35794:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 35795:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 35796:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 35797:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 35798:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 35799:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 35800:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 35801:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 35802:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 35803:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 35804:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 35805:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 35806:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 35807:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 35808:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 35809:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 35810:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 35811:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 35812:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 35813:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 35814:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 35815:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 35816:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 35817:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 35818:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 35819:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 35820:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 35821:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 35822:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 35823:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 35824:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 35825:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 35826:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 35827:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 35828:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 35829:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 35830:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 35831:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 35832:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 35833:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 35834:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 35835:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 35836:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 35837:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 35838:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 35839:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 35840:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 35841:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 35842:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 35843:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 35844:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 35845:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 35846:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 35847:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 35848:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 35849:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 35850:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 35851:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 35852:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 35853:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 35854:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 35855:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 35856:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 35857:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 35858:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 35859:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 35860:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 35861:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 35862:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 35863:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 35864:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 35865:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 35866:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 35867:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 35868:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 35869:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 35870:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 35871:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 35872:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 35873:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 35874:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 35875:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 35876:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 35877:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 35878:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 35879:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 35880:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 35881:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 35882:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 35883:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 35884:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 35885:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 35886:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 35887:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 35888:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 35889:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 35890:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 35891:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 35892:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 35893:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 35894:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 35895:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 35896:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 35897:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 35898:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 35899:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 35900:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 35901:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 35902:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 35903:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 35904:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 35905:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 35906:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 35907:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 35908:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 35909:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 35910:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 35911:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 35912:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 35913:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 35914:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 35915:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 35916:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 35917:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 35918:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 35919:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 35920:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 35921:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 35922:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 35923:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 35924:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 35925:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 35926:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 35927:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 35928:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 35929:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 35930:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 35931:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 35932:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 35933:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 35934:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 35935:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 35936:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 35937:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 35938:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 35939:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 35940:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 35941:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 35942:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 35943:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 35944:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 35945:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 35946:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 35947:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 35948:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 35949:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 35950:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 35951:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 35952:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 35953:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 35954:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 35955:22]
  wire  invx140 = ~x140; // @[Snxn100k.scala 35956:17]
  wire  t141 = x140 + invx140; // @[Snxn100k.scala 35957:22]
  wire  inv141 = ~t141; // @[Snxn100k.scala 35958:17]
  wire  x141 = t141 ^ inv141; // @[Snxn100k.scala 35959:22]
  wire  invx141 = ~x141; // @[Snxn100k.scala 35960:17]
  wire  t142 = x141 + invx141; // @[Snxn100k.scala 35961:22]
  wire  inv142 = ~t142; // @[Snxn100k.scala 35962:17]
  wire  x142 = t142 ^ inv142; // @[Snxn100k.scala 35963:22]
  wire  invx142 = ~x142; // @[Snxn100k.scala 35964:17]
  wire  t143 = x142 + invx142; // @[Snxn100k.scala 35965:22]
  wire  inv143 = ~t143; // @[Snxn100k.scala 35966:17]
  wire  x143 = t143 ^ inv143; // @[Snxn100k.scala 35967:22]
  assign io_z = ~x143; // @[Snxn100k.scala 35968:17]
endmodule
module SnxnLv4Inst91(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 35979:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 35980:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 35981:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 35982:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 35983:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 35984:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 35985:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 35986:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 35987:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 35988:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 35989:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 35990:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 35991:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 35992:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 35993:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 35994:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 35995:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 35996:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 35997:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 35998:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 35999:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 36000:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 36001:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 36002:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 36003:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 36004:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 36005:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 36006:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 36007:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 36008:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 36009:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 36010:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 36011:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 36012:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 36013:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 36014:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 36015:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 36016:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 36017:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 36018:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 36019:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 36020:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 36021:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 36022:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 36023:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 36024:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 36025:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 36026:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 36027:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 36028:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 36029:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 36030:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 36031:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 36032:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 36033:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 36034:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 36035:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 36036:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 36037:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 36038:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 36039:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 36040:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 36041:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 36042:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 36043:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 36044:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 36045:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 36046:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 36047:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 36048:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 36049:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 36050:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 36051:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 36052:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 36053:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 36054:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 36055:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 36056:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 36057:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 36058:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 36059:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 36060:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 36061:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 36062:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 36063:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 36064:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 36065:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 36066:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 36067:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 36068:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 36069:20]
  assign io_z = ~x22; // @[Snxn100k.scala 36070:16]
endmodule
module SnxnLv3Inst22(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst88_io_a; // @[Snxn100k.scala 10312:34]
  wire  inst_SnxnLv4Inst88_io_b; // @[Snxn100k.scala 10312:34]
  wire  inst_SnxnLv4Inst88_io_z; // @[Snxn100k.scala 10312:34]
  wire  inst_SnxnLv4Inst89_io_a; // @[Snxn100k.scala 10316:34]
  wire  inst_SnxnLv4Inst89_io_b; // @[Snxn100k.scala 10316:34]
  wire  inst_SnxnLv4Inst89_io_z; // @[Snxn100k.scala 10316:34]
  wire  inst_SnxnLv4Inst90_io_a; // @[Snxn100k.scala 10320:34]
  wire  inst_SnxnLv4Inst90_io_b; // @[Snxn100k.scala 10320:34]
  wire  inst_SnxnLv4Inst90_io_z; // @[Snxn100k.scala 10320:34]
  wire  inst_SnxnLv4Inst91_io_a; // @[Snxn100k.scala 10324:34]
  wire  inst_SnxnLv4Inst91_io_b; // @[Snxn100k.scala 10324:34]
  wire  inst_SnxnLv4Inst91_io_z; // @[Snxn100k.scala 10324:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst88_io_z + inst_SnxnLv4Inst89_io_z; // @[Snxn100k.scala 10328:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst90_io_z; // @[Snxn100k.scala 10328:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst91_io_z; // @[Snxn100k.scala 10328:89]
  SnxnLv4Inst7 inst_SnxnLv4Inst88 ( // @[Snxn100k.scala 10312:34]
    .io_a(inst_SnxnLv4Inst88_io_a),
    .io_b(inst_SnxnLv4Inst88_io_b),
    .io_z(inst_SnxnLv4Inst88_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst89 ( // @[Snxn100k.scala 10316:34]
    .io_a(inst_SnxnLv4Inst89_io_a),
    .io_b(inst_SnxnLv4Inst89_io_b),
    .io_z(inst_SnxnLv4Inst89_io_z)
  );
  SnxnLv4Inst90 inst_SnxnLv4Inst90 ( // @[Snxn100k.scala 10320:34]
    .io_a(inst_SnxnLv4Inst90_io_a),
    .io_b(inst_SnxnLv4Inst90_io_b),
    .io_z(inst_SnxnLv4Inst90_io_z)
  );
  SnxnLv4Inst91 inst_SnxnLv4Inst91 ( // @[Snxn100k.scala 10324:34]
    .io_a(inst_SnxnLv4Inst91_io_a),
    .io_b(inst_SnxnLv4Inst91_io_b),
    .io_z(inst_SnxnLv4Inst91_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10329:15]
  assign inst_SnxnLv4Inst88_io_a = io_a; // @[Snxn100k.scala 10313:27]
  assign inst_SnxnLv4Inst88_io_b = io_b; // @[Snxn100k.scala 10314:27]
  assign inst_SnxnLv4Inst89_io_a = io_a; // @[Snxn100k.scala 10317:27]
  assign inst_SnxnLv4Inst89_io_b = io_b; // @[Snxn100k.scala 10318:27]
  assign inst_SnxnLv4Inst90_io_a = io_a; // @[Snxn100k.scala 10321:27]
  assign inst_SnxnLv4Inst90_io_b = io_b; // @[Snxn100k.scala 10322:27]
  assign inst_SnxnLv4Inst91_io_a = io_a; // @[Snxn100k.scala 10325:27]
  assign inst_SnxnLv4Inst91_io_b = io_b; // @[Snxn100k.scala 10326:27]
endmodule
module SnxnLv4Inst93(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 38643:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 38644:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 38645:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 38646:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 38647:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 38648:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 38649:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 38650:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 38651:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 38652:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 38653:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 38654:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 38655:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 38656:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 38657:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 38658:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 38659:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 38660:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 38661:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 38662:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 38663:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 38664:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 38665:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 38666:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 38667:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 38668:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 38669:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 38670:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 38671:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 38672:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 38673:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 38674:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 38675:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 38676:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 38677:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 38678:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 38679:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 38680:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 38681:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 38682:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 38683:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 38684:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 38685:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 38686:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 38687:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 38688:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 38689:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 38690:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 38691:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 38692:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 38693:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 38694:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 38695:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 38696:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 38697:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 38698:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 38699:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 38700:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 38701:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 38702:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 38703:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 38704:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 38705:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 38706:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 38707:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 38708:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 38709:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 38710:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 38711:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 38712:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 38713:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 38714:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 38715:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 38716:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 38717:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 38718:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 38719:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 38720:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 38721:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 38722:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 38723:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 38724:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 38725:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 38726:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 38727:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 38728:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 38729:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 38730:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 38731:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 38732:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 38733:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 38734:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 38735:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 38736:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 38737:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 38738:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 38739:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 38740:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 38741:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 38742:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 38743:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 38744:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 38745:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 38746:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 38747:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 38748:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 38749:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 38750:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 38751:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 38752:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 38753:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 38754:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 38755:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 38756:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 38757:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 38758:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 38759:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 38760:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 38761:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 38762:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 38763:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 38764:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 38765:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 38766:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 38767:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 38768:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 38769:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 38770:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 38771:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 38772:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 38773:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 38774:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 38775:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 38776:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 38777:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 38778:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 38779:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 38780:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 38781:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 38782:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 38783:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 38784:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 38785:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 38786:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 38787:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 38788:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 38789:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 38790:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 38791:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 38792:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 38793:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 38794:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 38795:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 38796:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 38797:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 38798:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 38799:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 38800:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 38801:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 38802:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 38803:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 38804:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 38805:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 38806:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 38807:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 38808:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 38809:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 38810:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 38811:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 38812:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 38813:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 38814:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 38815:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 38816:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 38817:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 38818:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 38819:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 38820:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 38821:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 38822:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 38823:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 38824:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 38825:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 38826:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 38827:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 38828:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 38829:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 38830:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 38831:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 38832:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 38833:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 38834:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 38835:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 38836:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 38837:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 38838:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 38839:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 38840:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 38841:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 38842:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 38843:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 38844:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 38845:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 38846:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 38847:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 38848:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 38849:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 38850:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 38851:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 38852:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 38853:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 38854:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 38855:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 38856:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 38857:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 38858:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 38859:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 38860:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 38861:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 38862:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 38863:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 38864:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 38865:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 38866:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 38867:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 38868:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 38869:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 38870:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 38871:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 38872:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 38873:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 38874:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 38875:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 38876:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 38877:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 38878:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 38879:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 38880:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 38881:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 38882:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 38883:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 38884:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 38885:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 38886:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 38887:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 38888:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 38889:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 38890:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 38891:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 38892:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 38893:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 38894:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 38895:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 38896:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 38897:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 38898:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 38899:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 38900:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 38901:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 38902:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 38903:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 38904:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 38905:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 38906:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 38907:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 38908:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 38909:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 38910:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 38911:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 38912:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 38913:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 38914:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 38915:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 38916:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 38917:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 38918:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 38919:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 38920:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 38921:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 38922:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 38923:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 38924:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 38925:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 38926:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 38927:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 38928:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 38929:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 38930:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 38931:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 38932:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 38933:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 38934:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 38935:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 38936:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 38937:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 38938:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 38939:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 38940:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 38941:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 38942:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 38943:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 38944:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 38945:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 38946:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 38947:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 38948:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 38949:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 38950:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 38951:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 38952:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 38953:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 38954:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 38955:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 38956:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 38957:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 38958:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 38959:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 38960:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 38961:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 38962:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 38963:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 38964:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 38965:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 38966:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 38967:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 38968:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 38969:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 38970:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 38971:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 38972:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 38973:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 38974:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 38975:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 38976:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 38977:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 38978:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 38979:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 38980:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 38981:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 38982:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 38983:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 38984:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 38985:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 38986:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 38987:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 38988:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 38989:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 38990:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 38991:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 38992:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 38993:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 38994:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 38995:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 38996:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 38997:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 38998:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 38999:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 39000:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 39001:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 39002:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 39003:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 39004:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 39005:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 39006:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 39007:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 39008:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 39009:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 39010:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 39011:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 39012:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 39013:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 39014:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 39015:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 39016:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 39017:20]
  assign io_z = ~x93; // @[Snxn100k.scala 39018:16]
endmodule
module SnxnLv4Inst94(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 38421:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 38422:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 38423:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 38424:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 38425:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 38426:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 38427:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 38428:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 38429:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 38430:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 38431:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 38432:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 38433:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 38434:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 38435:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 38436:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 38437:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 38438:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 38439:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 38440:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 38441:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 38442:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 38443:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 38444:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 38445:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 38446:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 38447:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 38448:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 38449:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 38450:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 38451:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 38452:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 38453:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 38454:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 38455:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 38456:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 38457:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 38458:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 38459:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 38460:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 38461:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 38462:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 38463:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 38464:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 38465:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 38466:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 38467:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 38468:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 38469:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 38470:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 38471:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 38472:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 38473:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 38474:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 38475:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 38476:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 38477:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 38478:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 38479:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 38480:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 38481:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 38482:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 38483:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 38484:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 38485:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 38486:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 38487:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 38488:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 38489:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 38490:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 38491:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 38492:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 38493:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 38494:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 38495:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 38496:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 38497:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 38498:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 38499:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 38500:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 38501:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 38502:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 38503:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 38504:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 38505:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 38506:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 38507:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 38508:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 38509:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 38510:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 38511:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 38512:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 38513:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 38514:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 38515:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 38516:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 38517:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 38518:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 38519:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 38520:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 38521:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 38522:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 38523:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 38524:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 38525:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 38526:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 38527:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 38528:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 38529:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 38530:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 38531:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 38532:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 38533:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 38534:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 38535:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 38536:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 38537:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 38538:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 38539:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 38540:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 38541:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 38542:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 38543:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 38544:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 38545:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 38546:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 38547:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 38548:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 38549:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 38550:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 38551:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 38552:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 38553:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 38554:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 38555:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 38556:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 38557:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 38558:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 38559:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 38560:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 38561:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 38562:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 38563:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 38564:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 38565:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 38566:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 38567:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 38568:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 38569:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 38570:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 38571:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 38572:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 38573:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 38574:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 38575:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 38576:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 38577:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 38578:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 38579:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 38580:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 38581:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 38582:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 38583:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 38584:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 38585:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 38586:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 38587:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 38588:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 38589:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 38590:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 38591:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 38592:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 38593:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 38594:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 38595:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 38596:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 38597:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 38598:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 38599:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 38600:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 38601:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 38602:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 38603:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 38604:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 38605:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 38606:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 38607:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 38608:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 38609:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 38610:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 38611:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 38612:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 38613:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 38614:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 38615:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 38616:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 38617:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 38618:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 38619:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 38620:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 38621:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 38622:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 38623:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 38624:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 38625:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 38626:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 38627:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 38628:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 38629:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 38630:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 38631:20]
  assign io_z = ~x52; // @[Snxn100k.scala 38632:16]
endmodule
module SnxnLv4Inst95(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 38263:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 38264:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 38265:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 38266:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 38267:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 38268:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 38269:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 38270:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 38271:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 38272:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 38273:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 38274:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 38275:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 38276:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 38277:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 38278:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 38279:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 38280:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 38281:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 38282:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 38283:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 38284:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 38285:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 38286:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 38287:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 38288:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 38289:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 38290:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 38291:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 38292:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 38293:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 38294:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 38295:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 38296:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 38297:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 38298:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 38299:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 38300:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 38301:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 38302:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 38303:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 38304:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 38305:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 38306:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 38307:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 38308:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 38309:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 38310:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 38311:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 38312:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 38313:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 38314:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 38315:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 38316:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 38317:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 38318:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 38319:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 38320:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 38321:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 38322:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 38323:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 38324:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 38325:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 38326:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 38327:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 38328:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 38329:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 38330:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 38331:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 38332:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 38333:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 38334:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 38335:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 38336:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 38337:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 38338:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 38339:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 38340:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 38341:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 38342:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 38343:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 38344:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 38345:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 38346:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 38347:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 38348:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 38349:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 38350:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 38351:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 38352:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 38353:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 38354:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 38355:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 38356:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 38357:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 38358:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 38359:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 38360:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 38361:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 38362:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 38363:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 38364:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 38365:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 38366:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 38367:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 38368:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 38369:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 38370:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 38371:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 38372:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 38373:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 38374:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 38375:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 38376:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 38377:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 38378:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 38379:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 38380:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 38381:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 38382:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 38383:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 38384:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 38385:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 38386:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 38387:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 38388:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 38389:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 38390:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 38391:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 38392:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 38393:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 38394:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 38395:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 38396:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 38397:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 38398:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 38399:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 38400:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 38401:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 38402:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 38403:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 38404:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 38405:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 38406:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 38407:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 38408:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 38409:20]
  assign io_z = ~x36; // @[Snxn100k.scala 38410:16]
endmodule
module SnxnLv3Inst23(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst92_io_a; // @[Snxn100k.scala 11409:34]
  wire  inst_SnxnLv4Inst92_io_b; // @[Snxn100k.scala 11409:34]
  wire  inst_SnxnLv4Inst92_io_z; // @[Snxn100k.scala 11409:34]
  wire  inst_SnxnLv4Inst93_io_a; // @[Snxn100k.scala 11413:34]
  wire  inst_SnxnLv4Inst93_io_b; // @[Snxn100k.scala 11413:34]
  wire  inst_SnxnLv4Inst93_io_z; // @[Snxn100k.scala 11413:34]
  wire  inst_SnxnLv4Inst94_io_a; // @[Snxn100k.scala 11417:34]
  wire  inst_SnxnLv4Inst94_io_b; // @[Snxn100k.scala 11417:34]
  wire  inst_SnxnLv4Inst94_io_z; // @[Snxn100k.scala 11417:34]
  wire  inst_SnxnLv4Inst95_io_a; // @[Snxn100k.scala 11421:34]
  wire  inst_SnxnLv4Inst95_io_b; // @[Snxn100k.scala 11421:34]
  wire  inst_SnxnLv4Inst95_io_z; // @[Snxn100k.scala 11421:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst92_io_z + inst_SnxnLv4Inst93_io_z; // @[Snxn100k.scala 11425:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst94_io_z; // @[Snxn100k.scala 11425:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst95_io_z; // @[Snxn100k.scala 11425:89]
  SnxnLv4Inst84 inst_SnxnLv4Inst92 ( // @[Snxn100k.scala 11409:34]
    .io_a(inst_SnxnLv4Inst92_io_a),
    .io_b(inst_SnxnLv4Inst92_io_b),
    .io_z(inst_SnxnLv4Inst92_io_z)
  );
  SnxnLv4Inst93 inst_SnxnLv4Inst93 ( // @[Snxn100k.scala 11413:34]
    .io_a(inst_SnxnLv4Inst93_io_a),
    .io_b(inst_SnxnLv4Inst93_io_b),
    .io_z(inst_SnxnLv4Inst93_io_z)
  );
  SnxnLv4Inst94 inst_SnxnLv4Inst94 ( // @[Snxn100k.scala 11417:34]
    .io_a(inst_SnxnLv4Inst94_io_a),
    .io_b(inst_SnxnLv4Inst94_io_b),
    .io_z(inst_SnxnLv4Inst94_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst95 ( // @[Snxn100k.scala 11421:34]
    .io_a(inst_SnxnLv4Inst95_io_a),
    .io_b(inst_SnxnLv4Inst95_io_b),
    .io_z(inst_SnxnLv4Inst95_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 11426:15]
  assign inst_SnxnLv4Inst92_io_a = io_a; // @[Snxn100k.scala 11410:27]
  assign inst_SnxnLv4Inst92_io_b = io_b; // @[Snxn100k.scala 11411:27]
  assign inst_SnxnLv4Inst93_io_a = io_a; // @[Snxn100k.scala 11414:27]
  assign inst_SnxnLv4Inst93_io_b = io_b; // @[Snxn100k.scala 11415:27]
  assign inst_SnxnLv4Inst94_io_a = io_a; // @[Snxn100k.scala 11418:27]
  assign inst_SnxnLv4Inst94_io_b = io_b; // @[Snxn100k.scala 11419:27]
  assign inst_SnxnLv4Inst95_io_a = io_a; // @[Snxn100k.scala 11422:27]
  assign inst_SnxnLv4Inst95_io_b = io_b; // @[Snxn100k.scala 11423:27]
endmodule
module SnxnLv2Inst5(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst20_io_a; // @[Snxn100k.scala 2211:34]
  wire  inst_SnxnLv3Inst20_io_b; // @[Snxn100k.scala 2211:34]
  wire  inst_SnxnLv3Inst20_io_z; // @[Snxn100k.scala 2211:34]
  wire  inst_SnxnLv3Inst21_io_a; // @[Snxn100k.scala 2215:34]
  wire  inst_SnxnLv3Inst21_io_b; // @[Snxn100k.scala 2215:34]
  wire  inst_SnxnLv3Inst21_io_z; // @[Snxn100k.scala 2215:34]
  wire  inst_SnxnLv3Inst22_io_a; // @[Snxn100k.scala 2219:34]
  wire  inst_SnxnLv3Inst22_io_b; // @[Snxn100k.scala 2219:34]
  wire  inst_SnxnLv3Inst22_io_z; // @[Snxn100k.scala 2219:34]
  wire  inst_SnxnLv3Inst23_io_a; // @[Snxn100k.scala 2223:34]
  wire  inst_SnxnLv3Inst23_io_b; // @[Snxn100k.scala 2223:34]
  wire  inst_SnxnLv3Inst23_io_z; // @[Snxn100k.scala 2223:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst20_io_z + inst_SnxnLv3Inst21_io_z; // @[Snxn100k.scala 2227:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst22_io_z; // @[Snxn100k.scala 2227:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst23_io_z; // @[Snxn100k.scala 2227:89]
  SnxnLv3Inst20 inst_SnxnLv3Inst20 ( // @[Snxn100k.scala 2211:34]
    .io_a(inst_SnxnLv3Inst20_io_a),
    .io_b(inst_SnxnLv3Inst20_io_b),
    .io_z(inst_SnxnLv3Inst20_io_z)
  );
  SnxnLv3Inst21 inst_SnxnLv3Inst21 ( // @[Snxn100k.scala 2215:34]
    .io_a(inst_SnxnLv3Inst21_io_a),
    .io_b(inst_SnxnLv3Inst21_io_b),
    .io_z(inst_SnxnLv3Inst21_io_z)
  );
  SnxnLv3Inst22 inst_SnxnLv3Inst22 ( // @[Snxn100k.scala 2219:34]
    .io_a(inst_SnxnLv3Inst22_io_a),
    .io_b(inst_SnxnLv3Inst22_io_b),
    .io_z(inst_SnxnLv3Inst22_io_z)
  );
  SnxnLv3Inst23 inst_SnxnLv3Inst23 ( // @[Snxn100k.scala 2223:34]
    .io_a(inst_SnxnLv3Inst23_io_a),
    .io_b(inst_SnxnLv3Inst23_io_b),
    .io_z(inst_SnxnLv3Inst23_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 2228:15]
  assign inst_SnxnLv3Inst20_io_a = io_a; // @[Snxn100k.scala 2212:27]
  assign inst_SnxnLv3Inst20_io_b = io_b; // @[Snxn100k.scala 2213:27]
  assign inst_SnxnLv3Inst21_io_a = io_a; // @[Snxn100k.scala 2216:27]
  assign inst_SnxnLv3Inst21_io_b = io_b; // @[Snxn100k.scala 2217:27]
  assign inst_SnxnLv3Inst22_io_a = io_a; // @[Snxn100k.scala 2220:27]
  assign inst_SnxnLv3Inst22_io_b = io_b; // @[Snxn100k.scala 2221:27]
  assign inst_SnxnLv3Inst23_io_a = io_a; // @[Snxn100k.scala 2224:27]
  assign inst_SnxnLv3Inst23_io_b = io_b; // @[Snxn100k.scala 2225:27]
endmodule
module SnxnLv4Inst97(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 44973:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 44974:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 44975:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 44976:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 44977:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 44978:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 44979:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 44980:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 44981:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 44982:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 44983:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 44984:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 44985:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 44986:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 44987:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 44988:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 44989:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 44990:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 44991:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 44992:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 44993:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 44994:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 44995:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 44996:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 44997:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 44998:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 44999:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 45000:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 45001:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 45002:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 45003:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 45004:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 45005:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 45006:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 45007:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 45008:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 45009:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 45010:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 45011:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 45012:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 45013:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 45014:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 45015:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 45016:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 45017:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 45018:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 45019:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 45020:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 45021:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 45022:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 45023:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 45024:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 45025:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 45026:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 45027:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 45028:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 45029:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 45030:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 45031:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 45032:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 45033:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 45034:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 45035:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 45036:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 45037:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 45038:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 45039:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 45040:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 45041:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 45042:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 45043:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 45044:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 45045:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 45046:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 45047:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 45048:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 45049:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 45050:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 45051:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 45052:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 45053:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 45054:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 45055:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 45056:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 45057:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 45058:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 45059:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 45060:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 45061:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 45062:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 45063:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 45064:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 45065:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 45066:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 45067:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 45068:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 45069:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 45070:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 45071:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 45072:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 45073:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 45074:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 45075:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 45076:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 45077:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 45078:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 45079:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 45080:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 45081:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 45082:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 45083:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 45084:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 45085:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 45086:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 45087:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 45088:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 45089:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 45090:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 45091:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 45092:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 45093:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 45094:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 45095:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 45096:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 45097:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 45098:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 45099:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 45100:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 45101:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 45102:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 45103:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 45104:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 45105:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 45106:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 45107:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 45108:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 45109:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 45110:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 45111:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 45112:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 45113:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 45114:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 45115:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 45116:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 45117:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 45118:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 45119:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 45120:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 45121:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 45122:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 45123:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 45124:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 45125:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 45126:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 45127:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 45128:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 45129:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 45130:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 45131:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 45132:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 45133:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 45134:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 45135:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 45136:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 45137:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 45138:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 45139:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 45140:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 45141:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 45142:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 45143:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 45144:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 45145:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 45146:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 45147:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 45148:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 45149:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 45150:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 45151:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 45152:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 45153:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 45154:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 45155:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 45156:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 45157:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 45158:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 45159:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 45160:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 45161:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 45162:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 45163:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 45164:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 45165:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 45166:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 45167:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 45168:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 45169:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 45170:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 45171:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 45172:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 45173:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 45174:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 45175:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 45176:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 45177:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 45178:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 45179:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 45180:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 45181:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 45182:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 45183:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 45184:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 45185:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 45186:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 45187:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 45188:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 45189:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 45190:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 45191:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 45192:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 45193:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 45194:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 45195:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 45196:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 45197:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 45198:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 45199:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 45200:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 45201:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 45202:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 45203:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 45204:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 45205:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 45206:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 45207:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 45208:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 45209:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 45210:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 45211:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 45212:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 45213:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 45214:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 45215:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 45216:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 45217:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 45218:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 45219:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 45220:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 45221:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 45222:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 45223:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 45224:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 45225:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 45226:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 45227:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 45228:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 45229:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 45230:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 45231:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 45232:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 45233:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 45234:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 45235:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 45236:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 45237:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 45238:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 45239:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 45240:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 45241:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 45242:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 45243:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 45244:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 45245:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 45246:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 45247:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 45248:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 45249:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 45250:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 45251:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 45252:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 45253:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 45254:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 45255:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 45256:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 45257:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 45258:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 45259:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 45260:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 45261:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 45262:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 45263:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 45264:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 45265:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 45266:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 45267:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 45268:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 45269:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 45270:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 45271:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 45272:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 45273:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 45274:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 45275:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 45276:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 45277:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 45278:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 45279:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 45280:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 45281:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 45282:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 45283:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 45284:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 45285:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 45286:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 45287:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 45288:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 45289:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 45290:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 45291:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 45292:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 45293:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 45294:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 45295:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 45296:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 45297:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 45298:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 45299:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 45300:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 45301:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 45302:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 45303:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 45304:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 45305:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 45306:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 45307:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 45308:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 45309:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 45310:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 45311:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 45312:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 45313:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 45314:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 45315:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 45316:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 45317:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 45318:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 45319:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 45320:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 45321:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 45322:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 45323:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 45324:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 45325:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 45326:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 45327:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 45328:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 45329:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 45330:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 45331:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 45332:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 45333:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 45334:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 45335:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 45336:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 45337:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 45338:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 45339:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 45340:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 45341:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 45342:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 45343:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 45344:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 45345:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 45346:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 45347:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 45348:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 45349:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 45350:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 45351:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 45352:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 45353:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 45354:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 45355:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 45356:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 45357:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 45358:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 45359:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 45360:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 45361:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 45362:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 45363:20]
  assign io_z = ~x97; // @[Snxn100k.scala 45364:16]
endmodule
module SnxnLv3Inst24(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst96_io_a; // @[Snxn100k.scala 13156:34]
  wire  inst_SnxnLv4Inst96_io_b; // @[Snxn100k.scala 13156:34]
  wire  inst_SnxnLv4Inst96_io_z; // @[Snxn100k.scala 13156:34]
  wire  inst_SnxnLv4Inst97_io_a; // @[Snxn100k.scala 13160:34]
  wire  inst_SnxnLv4Inst97_io_b; // @[Snxn100k.scala 13160:34]
  wire  inst_SnxnLv4Inst97_io_z; // @[Snxn100k.scala 13160:34]
  wire  inst_SnxnLv4Inst98_io_a; // @[Snxn100k.scala 13164:34]
  wire  inst_SnxnLv4Inst98_io_b; // @[Snxn100k.scala 13164:34]
  wire  inst_SnxnLv4Inst98_io_z; // @[Snxn100k.scala 13164:34]
  wire  inst_SnxnLv4Inst99_io_a; // @[Snxn100k.scala 13168:34]
  wire  inst_SnxnLv4Inst99_io_b; // @[Snxn100k.scala 13168:34]
  wire  inst_SnxnLv4Inst99_io_z; // @[Snxn100k.scala 13168:34]
  wire  _sum_T_1 = inst_SnxnLv4Inst96_io_z + inst_SnxnLv4Inst97_io_z; // @[Snxn100k.scala 13172:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst98_io_z; // @[Snxn100k.scala 13172:63]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst99_io_z; // @[Snxn100k.scala 13172:89]
  SnxnLv4Inst43 inst_SnxnLv4Inst96 ( // @[Snxn100k.scala 13156:34]
    .io_a(inst_SnxnLv4Inst96_io_a),
    .io_b(inst_SnxnLv4Inst96_io_b),
    .io_z(inst_SnxnLv4Inst96_io_z)
  );
  SnxnLv4Inst97 inst_SnxnLv4Inst97 ( // @[Snxn100k.scala 13160:34]
    .io_a(inst_SnxnLv4Inst97_io_a),
    .io_b(inst_SnxnLv4Inst97_io_b),
    .io_z(inst_SnxnLv4Inst97_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst98 ( // @[Snxn100k.scala 13164:34]
    .io_a(inst_SnxnLv4Inst98_io_a),
    .io_b(inst_SnxnLv4Inst98_io_b),
    .io_z(inst_SnxnLv4Inst98_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst99 ( // @[Snxn100k.scala 13168:34]
    .io_a(inst_SnxnLv4Inst99_io_a),
    .io_b(inst_SnxnLv4Inst99_io_b),
    .io_z(inst_SnxnLv4Inst99_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 13173:15]
  assign inst_SnxnLv4Inst96_io_a = io_a; // @[Snxn100k.scala 13157:27]
  assign inst_SnxnLv4Inst96_io_b = io_b; // @[Snxn100k.scala 13158:27]
  assign inst_SnxnLv4Inst97_io_a = io_a; // @[Snxn100k.scala 13161:27]
  assign inst_SnxnLv4Inst97_io_b = io_b; // @[Snxn100k.scala 13162:27]
  assign inst_SnxnLv4Inst98_io_a = io_a; // @[Snxn100k.scala 13165:27]
  assign inst_SnxnLv4Inst98_io_b = io_b; // @[Snxn100k.scala 13166:27]
  assign inst_SnxnLv4Inst99_io_a = io_a; // @[Snxn100k.scala 13169:27]
  assign inst_SnxnLv4Inst99_io_b = io_b; // @[Snxn100k.scala 13170:27]
endmodule
module SnxnLv4Inst101(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 46923:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 46924:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 46925:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 46926:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 46927:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 46928:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 46929:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 46930:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 46931:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 46932:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 46933:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 46934:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 46935:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 46936:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 46937:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 46938:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 46939:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 46940:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 46941:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 46942:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 46943:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 46944:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 46945:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 46946:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 46947:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 46948:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 46949:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 46950:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 46951:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 46952:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 46953:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 46954:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 46955:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 46956:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 46957:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 46958:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 46959:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 46960:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 46961:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 46962:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 46963:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 46964:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 46965:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 46966:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 46967:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 46968:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 46969:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 46970:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 46971:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 46972:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 46973:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 46974:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 46975:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 46976:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 46977:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 46978:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 46979:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 46980:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 46981:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 46982:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 46983:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 46984:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 46985:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 46986:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 46987:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 46988:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 46989:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 46990:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 46991:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 46992:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 46993:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 46994:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 46995:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 46996:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 46997:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 46998:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 46999:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 47000:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 47001:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 47002:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 47003:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 47004:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 47005:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 47006:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 47007:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 47008:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 47009:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 47010:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 47011:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 47012:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 47013:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 47014:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 47015:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 47016:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 47017:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 47018:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 47019:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 47020:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 47021:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 47022:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 47023:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 47024:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 47025:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 47026:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 47027:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 47028:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 47029:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 47030:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 47031:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 47032:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 47033:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 47034:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 47035:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 47036:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 47037:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 47038:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 47039:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 47040:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 47041:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 47042:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 47043:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 47044:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 47045:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 47046:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 47047:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 47048:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 47049:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 47050:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 47051:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 47052:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 47053:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 47054:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 47055:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 47056:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 47057:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 47058:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 47059:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 47060:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 47061:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 47062:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 47063:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 47064:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 47065:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 47066:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 47067:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 47068:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 47069:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 47070:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 47071:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 47072:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 47073:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 47074:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 47075:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 47076:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 47077:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 47078:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 47079:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 47080:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 47081:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 47082:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 47083:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 47084:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 47085:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 47086:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 47087:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 47088:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 47089:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 47090:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 47091:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 47092:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 47093:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 47094:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 47095:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 47096:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 47097:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 47098:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 47099:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 47100:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 47101:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 47102:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 47103:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 47104:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 47105:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 47106:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 47107:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 47108:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 47109:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 47110:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 47111:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 47112:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 47113:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 47114:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 47115:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 47116:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 47117:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 47118:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 47119:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 47120:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 47121:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 47122:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 47123:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 47124:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 47125:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 47126:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 47127:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 47128:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 47129:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 47130:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 47131:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 47132:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 47133:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 47134:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 47135:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 47136:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 47137:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 47138:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 47139:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 47140:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 47141:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 47142:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 47143:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 47144:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 47145:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 47146:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 47147:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 47148:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 47149:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 47150:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 47151:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 47152:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 47153:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 47154:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 47155:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 47156:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 47157:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 47158:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 47159:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 47160:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 47161:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 47162:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 47163:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 47164:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 47165:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 47166:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 47167:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 47168:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 47169:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 47170:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 47171:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 47172:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 47173:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 47174:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 47175:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 47176:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 47177:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 47178:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 47179:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 47180:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 47181:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 47182:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 47183:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 47184:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 47185:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 47186:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 47187:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 47188:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 47189:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 47190:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 47191:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 47192:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 47193:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 47194:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 47195:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 47196:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 47197:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 47198:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 47199:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 47200:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 47201:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 47202:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 47203:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 47204:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 47205:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 47206:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 47207:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 47208:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 47209:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 47210:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 47211:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 47212:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 47213:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 47214:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 47215:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 47216:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 47217:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 47218:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 47219:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 47220:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 47221:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 47222:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 47223:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 47224:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 47225:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 47226:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 47227:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 47228:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 47229:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 47230:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 47231:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 47232:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 47233:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 47234:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 47235:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 47236:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 47237:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 47238:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 47239:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 47240:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 47241:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 47242:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 47243:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 47244:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 47245:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 47246:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 47247:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 47248:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 47249:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 47250:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 47251:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 47252:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 47253:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 47254:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 47255:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 47256:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 47257:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 47258:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 47259:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 47260:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 47261:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 47262:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 47263:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 47264:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 47265:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 47266:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 47267:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 47268:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 47269:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 47270:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 47271:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 47272:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 47273:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 47274:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 47275:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 47276:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 47277:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 47278:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 47279:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 47280:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 47281:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 47282:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 47283:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 47284:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 47285:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 47286:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 47287:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 47288:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 47289:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 47290:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 47291:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 47292:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 47293:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 47294:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 47295:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 47296:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 47297:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 47298:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 47299:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 47300:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 47301:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 47302:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 47303:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 47304:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 47305:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 47306:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 47307:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 47308:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 47309:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 47310:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 47311:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 47312:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 47313:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 47314:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 47315:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 47316:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 47317:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 47318:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 47319:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 47320:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 47321:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 47322:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 47323:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 47324:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 47325:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 47326:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 47327:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 47328:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 47329:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 47330:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 47331:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 47332:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 47333:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 47334:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 47335:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 47336:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 47337:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 47338:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 47339:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 47340:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 47341:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 47342:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 47343:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 47344:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 47345:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 47346:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 47347:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 47348:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 47349:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 47350:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 47351:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 47352:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 47353:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 47354:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 47355:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 47356:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 47357:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 47358:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 47359:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 47360:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 47361:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 47362:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 47363:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 47364:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 47365:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 47366:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 47367:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 47368:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 47369:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 47370:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 47371:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 47372:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 47373:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 47374:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 47375:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 47376:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 47377:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 47378:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 47379:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 47380:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 47381:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 47382:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 47383:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 47384:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 47385:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 47386:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 47387:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 47388:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 47389:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 47390:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 47391:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 47392:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 47393:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 47394:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 47395:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 47396:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 47397:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 47398:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 47399:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 47400:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 47401:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 47402:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 47403:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 47404:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 47405:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 47406:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 47407:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 47408:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 47409:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 47410:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 47411:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 47412:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 47413:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 47414:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 47415:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 47416:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 47417:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 47418:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 47419:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 47420:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 47421:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 47422:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 47423:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 47424:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 47425:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 47426:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 47427:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 47428:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 47429:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 47430:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 47431:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 47432:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 47433:22]
  assign io_z = ~x127; // @[Snxn100k.scala 47434:17]
endmodule
module SnxnLv3Inst25(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst100_io_a; // @[Snxn100k.scala 13227:35]
  wire  inst_SnxnLv4Inst100_io_b; // @[Snxn100k.scala 13227:35]
  wire  inst_SnxnLv4Inst100_io_z; // @[Snxn100k.scala 13227:35]
  wire  inst_SnxnLv4Inst101_io_a; // @[Snxn100k.scala 13231:35]
  wire  inst_SnxnLv4Inst101_io_b; // @[Snxn100k.scala 13231:35]
  wire  inst_SnxnLv4Inst101_io_z; // @[Snxn100k.scala 13231:35]
  wire  inst_SnxnLv4Inst102_io_a; // @[Snxn100k.scala 13235:35]
  wire  inst_SnxnLv4Inst102_io_b; // @[Snxn100k.scala 13235:35]
  wire  inst_SnxnLv4Inst102_io_z; // @[Snxn100k.scala 13235:35]
  wire  inst_SnxnLv4Inst103_io_a; // @[Snxn100k.scala 13239:35]
  wire  inst_SnxnLv4Inst103_io_b; // @[Snxn100k.scala 13239:35]
  wire  inst_SnxnLv4Inst103_io_z; // @[Snxn100k.scala 13239:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst100_io_z + inst_SnxnLv4Inst101_io_z; // @[Snxn100k.scala 13243:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst102_io_z; // @[Snxn100k.scala 13243:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst103_io_z; // @[Snxn100k.scala 13243:92]
  SnxnLv4Inst69 inst_SnxnLv4Inst100 ( // @[Snxn100k.scala 13227:35]
    .io_a(inst_SnxnLv4Inst100_io_a),
    .io_b(inst_SnxnLv4Inst100_io_b),
    .io_z(inst_SnxnLv4Inst100_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst101 ( // @[Snxn100k.scala 13231:35]
    .io_a(inst_SnxnLv4Inst101_io_a),
    .io_b(inst_SnxnLv4Inst101_io_b),
    .io_z(inst_SnxnLv4Inst101_io_z)
  );
  SnxnLv4Inst97 inst_SnxnLv4Inst102 ( // @[Snxn100k.scala 13235:35]
    .io_a(inst_SnxnLv4Inst102_io_a),
    .io_b(inst_SnxnLv4Inst102_io_b),
    .io_z(inst_SnxnLv4Inst102_io_z)
  );
  SnxnLv4Inst94 inst_SnxnLv4Inst103 ( // @[Snxn100k.scala 13239:35]
    .io_a(inst_SnxnLv4Inst103_io_a),
    .io_b(inst_SnxnLv4Inst103_io_b),
    .io_z(inst_SnxnLv4Inst103_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 13244:15]
  assign inst_SnxnLv4Inst100_io_a = io_a; // @[Snxn100k.scala 13228:28]
  assign inst_SnxnLv4Inst100_io_b = io_b; // @[Snxn100k.scala 13229:28]
  assign inst_SnxnLv4Inst101_io_a = io_a; // @[Snxn100k.scala 13232:28]
  assign inst_SnxnLv4Inst101_io_b = io_b; // @[Snxn100k.scala 13233:28]
  assign inst_SnxnLv4Inst102_io_a = io_a; // @[Snxn100k.scala 13236:28]
  assign inst_SnxnLv4Inst102_io_b = io_b; // @[Snxn100k.scala 13237:28]
  assign inst_SnxnLv4Inst103_io_a = io_a; // @[Snxn100k.scala 13240:28]
  assign inst_SnxnLv4Inst103_io_b = io_b; // @[Snxn100k.scala 13241:28]
endmodule
module SnxnLv4Inst104(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 50107:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 50108:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 50109:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 50110:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 50111:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 50112:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 50113:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 50114:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 50115:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 50116:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 50117:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 50118:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 50119:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 50120:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 50121:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 50122:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 50123:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 50124:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 50125:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 50126:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 50127:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 50128:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 50129:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 50130:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 50131:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 50132:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 50133:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 50134:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 50135:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 50136:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 50137:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 50138:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 50139:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 50140:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 50141:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 50142:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 50143:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 50144:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 50145:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 50146:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 50147:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 50148:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 50149:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 50150:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 50151:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 50152:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 50153:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 50154:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 50155:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 50156:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 50157:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 50158:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 50159:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 50160:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 50161:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 50162:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 50163:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 50164:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 50165:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 50166:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 50167:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 50168:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 50169:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 50170:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 50171:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 50172:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 50173:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 50174:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 50175:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 50176:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 50177:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 50178:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 50179:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 50180:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 50181:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 50182:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 50183:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 50184:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 50185:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 50186:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 50187:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 50188:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 50189:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 50190:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 50191:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 50192:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 50193:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 50194:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 50195:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 50196:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 50197:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 50198:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 50199:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 50200:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 50201:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 50202:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 50203:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 50204:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 50205:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 50206:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 50207:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 50208:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 50209:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 50210:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 50211:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 50212:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 50213:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 50214:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 50215:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 50216:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 50217:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 50218:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 50219:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 50220:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 50221:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 50222:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 50223:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 50224:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 50225:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 50226:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 50227:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 50228:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 50229:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 50230:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 50231:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 50232:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 50233:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 50234:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 50235:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 50236:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 50237:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 50238:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 50239:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 50240:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 50241:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 50242:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 50243:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 50244:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 50245:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 50246:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 50247:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 50248:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 50249:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 50250:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 50251:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 50252:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 50253:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 50254:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 50255:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 50256:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 50257:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 50258:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 50259:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 50260:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 50261:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 50262:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 50263:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 50264:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 50265:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 50266:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 50267:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 50268:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 50269:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 50270:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 50271:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 50272:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 50273:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 50274:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 50275:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 50276:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 50277:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 50278:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 50279:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 50280:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 50281:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 50282:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 50283:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 50284:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 50285:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 50286:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 50287:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 50288:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 50289:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 50290:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 50291:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 50292:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 50293:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 50294:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 50295:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 50296:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 50297:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 50298:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 50299:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 50300:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 50301:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 50302:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 50303:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 50304:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 50305:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 50306:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 50307:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 50308:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 50309:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 50310:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 50311:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 50312:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 50313:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 50314:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 50315:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 50316:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 50317:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 50318:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 50319:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 50320:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 50321:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 50322:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 50323:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 50324:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 50325:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 50326:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 50327:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 50328:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 50329:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 50330:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 50331:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 50332:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 50333:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 50334:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 50335:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 50336:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 50337:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 50338:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 50339:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 50340:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 50341:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 50342:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 50343:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 50344:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 50345:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 50346:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 50347:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 50348:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 50349:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 50350:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 50351:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 50352:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 50353:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 50354:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 50355:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 50356:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 50357:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 50358:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 50359:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 50360:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 50361:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 50362:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 50363:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 50364:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 50365:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 50366:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 50367:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 50368:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 50369:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 50370:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 50371:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 50372:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 50373:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 50374:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 50375:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 50376:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 50377:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 50378:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 50379:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 50380:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 50381:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 50382:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 50383:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 50384:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 50385:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 50386:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 50387:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 50388:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 50389:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 50390:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 50391:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 50392:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 50393:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 50394:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 50395:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 50396:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 50397:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 50398:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 50399:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 50400:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 50401:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 50402:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 50403:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 50404:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 50405:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 50406:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 50407:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 50408:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 50409:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 50410:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 50411:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 50412:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 50413:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 50414:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 50415:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 50416:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 50417:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 50418:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 50419:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 50420:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 50421:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 50422:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 50423:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 50424:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 50425:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 50426:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 50427:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 50428:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 50429:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 50430:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 50431:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 50432:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 50433:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 50434:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 50435:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 50436:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 50437:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 50438:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 50439:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 50440:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 50441:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 50442:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 50443:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 50444:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 50445:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 50446:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 50447:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 50448:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 50449:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 50450:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 50451:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 50452:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 50453:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 50454:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 50455:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 50456:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 50457:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 50458:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 50459:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 50460:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 50461:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 50462:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 50463:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 50464:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 50465:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 50466:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 50467:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 50468:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 50469:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 50470:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 50471:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 50472:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 50473:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 50474:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 50475:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 50476:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 50477:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 50478:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 50479:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 50480:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 50481:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 50482:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 50483:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 50484:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 50485:20]
  assign io_z = ~x94; // @[Snxn100k.scala 50486:16]
endmodule
module SnxnLv4Inst107(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 49511:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 49512:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 49513:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 49514:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 49515:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 49516:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 49517:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 49518:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 49519:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 49520:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 49521:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 49522:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 49523:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 49524:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 49525:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 49526:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 49527:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 49528:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 49529:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 49530:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 49531:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 49532:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 49533:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 49534:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 49535:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 49536:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 49537:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 49538:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 49539:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 49540:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 49541:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 49542:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 49543:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 49544:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 49545:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 49546:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 49547:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 49548:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 49549:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 49550:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 49551:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 49552:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 49553:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 49554:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 49555:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 49556:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 49557:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 49558:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 49559:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 49560:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 49561:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 49562:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 49563:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 49564:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 49565:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 49566:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 49567:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 49568:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 49569:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 49570:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 49571:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 49572:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 49573:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 49574:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 49575:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 49576:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 49577:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 49578:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 49579:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 49580:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 49581:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 49582:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 49583:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 49584:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 49585:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 49586:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 49587:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 49588:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 49589:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 49590:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 49591:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 49592:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 49593:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 49594:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 49595:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 49596:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 49597:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 49598:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 49599:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 49600:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 49601:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 49602:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 49603:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 49604:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 49605:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 49606:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 49607:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 49608:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 49609:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 49610:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 49611:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 49612:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 49613:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 49614:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 49615:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 49616:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 49617:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 49618:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 49619:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 49620:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 49621:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 49622:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 49623:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 49624:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 49625:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 49626:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 49627:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 49628:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 49629:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 49630:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 49631:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 49632:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 49633:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 49634:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 49635:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 49636:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 49637:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 49638:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 49639:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 49640:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 49641:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 49642:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 49643:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 49644:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 49645:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 49646:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 49647:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 49648:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 49649:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 49650:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 49651:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 49652:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 49653:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 49654:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 49655:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 49656:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 49657:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 49658:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 49659:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 49660:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 49661:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 49662:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 49663:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 49664:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 49665:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 49666:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 49667:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 49668:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 49669:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 49670:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 49671:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 49672:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 49673:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 49674:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 49675:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 49676:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 49677:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 49678:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 49679:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 49680:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 49681:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 49682:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 49683:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 49684:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 49685:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 49686:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 49687:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 49688:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 49689:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 49690:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 49691:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 49692:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 49693:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 49694:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 49695:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 49696:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 49697:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 49698:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 49699:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 49700:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 49701:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 49702:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 49703:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 49704:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 49705:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 49706:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 49707:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 49708:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 49709:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 49710:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 49711:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 49712:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 49713:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 49714:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 49715:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 49716:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 49717:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 49718:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 49719:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 49720:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 49721:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 49722:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 49723:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 49724:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 49725:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 49726:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 49727:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 49728:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 49729:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 49730:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 49731:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 49732:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 49733:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 49734:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 49735:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 49736:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 49737:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 49738:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 49739:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 49740:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 49741:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 49742:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 49743:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 49744:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 49745:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 49746:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 49747:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 49748:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 49749:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 49750:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 49751:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 49752:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 49753:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 49754:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 49755:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 49756:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 49757:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 49758:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 49759:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 49760:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 49761:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 49762:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 49763:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 49764:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 49765:20]
  assign io_z = ~x63; // @[Snxn100k.scala 49766:16]
endmodule
module SnxnLv3Inst26(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst104_io_a; // @[Snxn100k.scala 14249:35]
  wire  inst_SnxnLv4Inst104_io_b; // @[Snxn100k.scala 14249:35]
  wire  inst_SnxnLv4Inst104_io_z; // @[Snxn100k.scala 14249:35]
  wire  inst_SnxnLv4Inst105_io_a; // @[Snxn100k.scala 14253:35]
  wire  inst_SnxnLv4Inst105_io_b; // @[Snxn100k.scala 14253:35]
  wire  inst_SnxnLv4Inst105_io_z; // @[Snxn100k.scala 14253:35]
  wire  inst_SnxnLv4Inst106_io_a; // @[Snxn100k.scala 14257:35]
  wire  inst_SnxnLv4Inst106_io_b; // @[Snxn100k.scala 14257:35]
  wire  inst_SnxnLv4Inst106_io_z; // @[Snxn100k.scala 14257:35]
  wire  inst_SnxnLv4Inst107_io_a; // @[Snxn100k.scala 14261:35]
  wire  inst_SnxnLv4Inst107_io_b; // @[Snxn100k.scala 14261:35]
  wire  inst_SnxnLv4Inst107_io_z; // @[Snxn100k.scala 14261:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst104_io_z + inst_SnxnLv4Inst105_io_z; // @[Snxn100k.scala 14265:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst106_io_z; // @[Snxn100k.scala 14265:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst107_io_z; // @[Snxn100k.scala 14265:92]
  SnxnLv4Inst104 inst_SnxnLv4Inst104 ( // @[Snxn100k.scala 14249:35]
    .io_a(inst_SnxnLv4Inst104_io_a),
    .io_b(inst_SnxnLv4Inst104_io_b),
    .io_z(inst_SnxnLv4Inst104_io_z)
  );
  SnxnLv4Inst41 inst_SnxnLv4Inst105 ( // @[Snxn100k.scala 14253:35]
    .io_a(inst_SnxnLv4Inst105_io_a),
    .io_b(inst_SnxnLv4Inst105_io_b),
    .io_z(inst_SnxnLv4Inst105_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst106 ( // @[Snxn100k.scala 14257:35]
    .io_a(inst_SnxnLv4Inst106_io_a),
    .io_b(inst_SnxnLv4Inst106_io_b),
    .io_z(inst_SnxnLv4Inst106_io_z)
  );
  SnxnLv4Inst107 inst_SnxnLv4Inst107 ( // @[Snxn100k.scala 14261:35]
    .io_a(inst_SnxnLv4Inst107_io_a),
    .io_b(inst_SnxnLv4Inst107_io_b),
    .io_z(inst_SnxnLv4Inst107_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14266:15]
  assign inst_SnxnLv4Inst104_io_a = io_a; // @[Snxn100k.scala 14250:28]
  assign inst_SnxnLv4Inst104_io_b = io_b; // @[Snxn100k.scala 14251:28]
  assign inst_SnxnLv4Inst105_io_a = io_a; // @[Snxn100k.scala 14254:28]
  assign inst_SnxnLv4Inst105_io_b = io_b; // @[Snxn100k.scala 14255:28]
  assign inst_SnxnLv4Inst106_io_a = io_a; // @[Snxn100k.scala 14258:28]
  assign inst_SnxnLv4Inst106_io_b = io_b; // @[Snxn100k.scala 14259:28]
  assign inst_SnxnLv4Inst107_io_a = io_a; // @[Snxn100k.scala 14262:28]
  assign inst_SnxnLv4Inst107_io_b = io_b; // @[Snxn100k.scala 14263:28]
endmodule
module SnxnLv4Inst108(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 47815:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 47816:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 47817:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 47818:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 47819:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 47820:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 47821:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 47822:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 47823:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 47824:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 47825:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 47826:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 47827:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 47828:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 47829:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 47830:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 47831:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 47832:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 47833:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 47834:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 47835:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 47836:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 47837:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 47838:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 47839:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 47840:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 47841:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 47842:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 47843:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 47844:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 47845:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 47846:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 47847:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 47848:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 47849:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 47850:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 47851:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 47852:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 47853:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 47854:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 47855:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 47856:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 47857:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 47858:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 47859:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 47860:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 47861:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 47862:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 47863:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 47864:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 47865:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 47866:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 47867:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 47868:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 47869:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 47870:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 47871:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 47872:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 47873:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 47874:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 47875:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 47876:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 47877:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 47878:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 47879:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 47880:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 47881:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 47882:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 47883:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 47884:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 47885:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 47886:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 47887:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 47888:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 47889:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 47890:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 47891:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 47892:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 47893:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 47894:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 47895:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 47896:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 47897:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 47898:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 47899:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 47900:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 47901:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 47902:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 47903:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 47904:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 47905:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 47906:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 47907:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 47908:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 47909:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 47910:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 47911:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 47912:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 47913:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 47914:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 47915:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 47916:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 47917:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 47918:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 47919:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 47920:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 47921:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 47922:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 47923:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 47924:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 47925:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 47926:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 47927:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 47928:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 47929:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 47930:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 47931:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 47932:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 47933:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 47934:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 47935:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 47936:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 47937:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 47938:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 47939:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 47940:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 47941:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 47942:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 47943:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 47944:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 47945:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 47946:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 47947:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 47948:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 47949:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 47950:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 47951:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 47952:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 47953:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 47954:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 47955:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 47956:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 47957:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 47958:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 47959:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 47960:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 47961:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 47962:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 47963:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 47964:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 47965:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 47966:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 47967:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 47968:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 47969:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 47970:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 47971:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 47972:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 47973:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 47974:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 47975:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 47976:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 47977:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 47978:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 47979:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 47980:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 47981:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 47982:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 47983:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 47984:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 47985:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 47986:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 47987:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 47988:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 47989:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 47990:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 47991:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 47992:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 47993:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 47994:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 47995:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 47996:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 47997:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 47998:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 47999:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 48000:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 48001:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 48002:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 48003:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 48004:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 48005:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 48006:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 48007:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 48008:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 48009:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 48010:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 48011:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 48012:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 48013:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 48014:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 48015:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 48016:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 48017:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 48018:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 48019:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 48020:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 48021:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 48022:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 48023:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 48024:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 48025:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 48026:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 48027:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 48028:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 48029:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 48030:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 48031:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 48032:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 48033:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 48034:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 48035:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 48036:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 48037:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 48038:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 48039:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 48040:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 48041:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 48042:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 48043:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 48044:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 48045:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 48046:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 48047:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 48048:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 48049:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 48050:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 48051:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 48052:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 48053:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 48054:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 48055:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 48056:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 48057:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 48058:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 48059:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 48060:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 48061:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 48062:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 48063:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 48064:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 48065:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 48066:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 48067:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 48068:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 48069:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 48070:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 48071:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 48072:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 48073:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 48074:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 48075:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 48076:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 48077:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 48078:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 48079:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 48080:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 48081:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 48082:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 48083:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 48084:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 48085:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 48086:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 48087:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 48088:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 48089:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 48090:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 48091:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 48092:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 48093:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 48094:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 48095:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 48096:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 48097:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 48098:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 48099:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 48100:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 48101:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 48102:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 48103:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 48104:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 48105:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 48106:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 48107:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 48108:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 48109:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 48110:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 48111:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 48112:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 48113:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 48114:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 48115:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 48116:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 48117:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 48118:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 48119:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 48120:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 48121:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 48122:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 48123:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 48124:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 48125:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 48126:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 48127:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 48128:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 48129:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 48130:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 48131:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 48132:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 48133:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 48134:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 48135:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 48136:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 48137:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 48138:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 48139:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 48140:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 48141:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 48142:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 48143:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 48144:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 48145:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 48146:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 48147:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 48148:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 48149:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 48150:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 48151:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 48152:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 48153:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 48154:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 48155:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 48156:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 48157:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 48158:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 48159:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 48160:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 48161:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 48162:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 48163:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 48164:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 48165:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 48166:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 48167:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 48168:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 48169:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 48170:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 48171:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 48172:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 48173:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 48174:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 48175:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 48176:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 48177:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 48178:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 48179:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 48180:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 48181:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 48182:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 48183:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 48184:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 48185:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 48186:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 48187:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 48188:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 48189:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 48190:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 48191:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 48192:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 48193:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 48194:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 48195:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 48196:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 48197:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 48198:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 48199:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 48200:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 48201:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 48202:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 48203:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 48204:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 48205:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 48206:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 48207:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 48208:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 48209:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 48210:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 48211:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 48212:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 48213:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 48214:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 48215:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 48216:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 48217:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 48218:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 48219:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 48220:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 48221:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 48222:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 48223:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 48224:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 48225:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 48226:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 48227:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 48228:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 48229:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 48230:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 48231:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 48232:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 48233:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 48234:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 48235:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 48236:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 48237:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 48238:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 48239:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 48240:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 48241:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 48242:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 48243:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 48244:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 48245:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 48246:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 48247:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 48248:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 48249:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 48250:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 48251:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 48252:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 48253:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 48254:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 48255:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 48256:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 48257:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 48258:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 48259:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 48260:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 48261:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 48262:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 48263:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 48264:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 48265:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 48266:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 48267:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 48268:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 48269:22]
  assign io_z = ~x113; // @[Snxn100k.scala 48270:17]
endmodule
module SnxnLv3Inst27(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst108_io_a; // @[Snxn100k.scala 13690:35]
  wire  inst_SnxnLv4Inst108_io_b; // @[Snxn100k.scala 13690:35]
  wire  inst_SnxnLv4Inst108_io_z; // @[Snxn100k.scala 13690:35]
  wire  inst_SnxnLv4Inst109_io_a; // @[Snxn100k.scala 13694:35]
  wire  inst_SnxnLv4Inst109_io_b; // @[Snxn100k.scala 13694:35]
  wire  inst_SnxnLv4Inst109_io_z; // @[Snxn100k.scala 13694:35]
  wire  inst_SnxnLv4Inst110_io_a; // @[Snxn100k.scala 13698:35]
  wire  inst_SnxnLv4Inst110_io_b; // @[Snxn100k.scala 13698:35]
  wire  inst_SnxnLv4Inst110_io_z; // @[Snxn100k.scala 13698:35]
  wire  inst_SnxnLv4Inst111_io_a; // @[Snxn100k.scala 13702:35]
  wire  inst_SnxnLv4Inst111_io_b; // @[Snxn100k.scala 13702:35]
  wire  inst_SnxnLv4Inst111_io_z; // @[Snxn100k.scala 13702:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst108_io_z + inst_SnxnLv4Inst109_io_z; // @[Snxn100k.scala 13706:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst110_io_z; // @[Snxn100k.scala 13706:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst111_io_z; // @[Snxn100k.scala 13706:92]
  SnxnLv4Inst108 inst_SnxnLv4Inst108 ( // @[Snxn100k.scala 13690:35]
    .io_a(inst_SnxnLv4Inst108_io_a),
    .io_b(inst_SnxnLv4Inst108_io_b),
    .io_z(inst_SnxnLv4Inst108_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst109 ( // @[Snxn100k.scala 13694:35]
    .io_a(inst_SnxnLv4Inst109_io_a),
    .io_b(inst_SnxnLv4Inst109_io_b),
    .io_z(inst_SnxnLv4Inst109_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst110 ( // @[Snxn100k.scala 13698:35]
    .io_a(inst_SnxnLv4Inst110_io_a),
    .io_b(inst_SnxnLv4Inst110_io_b),
    .io_z(inst_SnxnLv4Inst110_io_z)
  );
  SnxnLv4Inst12 inst_SnxnLv4Inst111 ( // @[Snxn100k.scala 13702:35]
    .io_a(inst_SnxnLv4Inst111_io_a),
    .io_b(inst_SnxnLv4Inst111_io_b),
    .io_z(inst_SnxnLv4Inst111_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 13707:15]
  assign inst_SnxnLv4Inst108_io_a = io_a; // @[Snxn100k.scala 13691:28]
  assign inst_SnxnLv4Inst108_io_b = io_b; // @[Snxn100k.scala 13692:28]
  assign inst_SnxnLv4Inst109_io_a = io_a; // @[Snxn100k.scala 13695:28]
  assign inst_SnxnLv4Inst109_io_b = io_b; // @[Snxn100k.scala 13696:28]
  assign inst_SnxnLv4Inst110_io_a = io_a; // @[Snxn100k.scala 13699:28]
  assign inst_SnxnLv4Inst110_io_b = io_b; // @[Snxn100k.scala 13700:28]
  assign inst_SnxnLv4Inst111_io_a = io_a; // @[Snxn100k.scala 13703:28]
  assign inst_SnxnLv4Inst111_io_b = io_b; // @[Snxn100k.scala 13704:28]
endmodule
module SnxnLv2Inst6(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst24_io_a; // @[Snxn100k.scala 3253:34]
  wire  inst_SnxnLv3Inst24_io_b; // @[Snxn100k.scala 3253:34]
  wire  inst_SnxnLv3Inst24_io_z; // @[Snxn100k.scala 3253:34]
  wire  inst_SnxnLv3Inst25_io_a; // @[Snxn100k.scala 3257:34]
  wire  inst_SnxnLv3Inst25_io_b; // @[Snxn100k.scala 3257:34]
  wire  inst_SnxnLv3Inst25_io_z; // @[Snxn100k.scala 3257:34]
  wire  inst_SnxnLv3Inst26_io_a; // @[Snxn100k.scala 3261:34]
  wire  inst_SnxnLv3Inst26_io_b; // @[Snxn100k.scala 3261:34]
  wire  inst_SnxnLv3Inst26_io_z; // @[Snxn100k.scala 3261:34]
  wire  inst_SnxnLv3Inst27_io_a; // @[Snxn100k.scala 3265:34]
  wire  inst_SnxnLv3Inst27_io_b; // @[Snxn100k.scala 3265:34]
  wire  inst_SnxnLv3Inst27_io_z; // @[Snxn100k.scala 3265:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst24_io_z + inst_SnxnLv3Inst25_io_z; // @[Snxn100k.scala 3269:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst26_io_z; // @[Snxn100k.scala 3269:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst27_io_z; // @[Snxn100k.scala 3269:89]
  SnxnLv3Inst24 inst_SnxnLv3Inst24 ( // @[Snxn100k.scala 3253:34]
    .io_a(inst_SnxnLv3Inst24_io_a),
    .io_b(inst_SnxnLv3Inst24_io_b),
    .io_z(inst_SnxnLv3Inst24_io_z)
  );
  SnxnLv3Inst25 inst_SnxnLv3Inst25 ( // @[Snxn100k.scala 3257:34]
    .io_a(inst_SnxnLv3Inst25_io_a),
    .io_b(inst_SnxnLv3Inst25_io_b),
    .io_z(inst_SnxnLv3Inst25_io_z)
  );
  SnxnLv3Inst26 inst_SnxnLv3Inst26 ( // @[Snxn100k.scala 3261:34]
    .io_a(inst_SnxnLv3Inst26_io_a),
    .io_b(inst_SnxnLv3Inst26_io_b),
    .io_z(inst_SnxnLv3Inst26_io_z)
  );
  SnxnLv3Inst27 inst_SnxnLv3Inst27 ( // @[Snxn100k.scala 3265:34]
    .io_a(inst_SnxnLv3Inst27_io_a),
    .io_b(inst_SnxnLv3Inst27_io_b),
    .io_z(inst_SnxnLv3Inst27_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 3270:15]
  assign inst_SnxnLv3Inst24_io_a = io_a; // @[Snxn100k.scala 3254:27]
  assign inst_SnxnLv3Inst24_io_b = io_b; // @[Snxn100k.scala 3255:27]
  assign inst_SnxnLv3Inst25_io_a = io_a; // @[Snxn100k.scala 3258:27]
  assign inst_SnxnLv3Inst25_io_b = io_b; // @[Snxn100k.scala 3259:27]
  assign inst_SnxnLv3Inst26_io_a = io_a; // @[Snxn100k.scala 3262:27]
  assign inst_SnxnLv3Inst26_io_b = io_b; // @[Snxn100k.scala 3263:27]
  assign inst_SnxnLv3Inst27_io_a = io_a; // @[Snxn100k.scala 3266:27]
  assign inst_SnxnLv3Inst27_io_b = io_b; // @[Snxn100k.scala 3267:27]
endmodule
module SnxnLv4Inst113(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 32397:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 32398:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 32399:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 32400:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 32401:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 32402:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 32403:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 32404:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 32405:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 32406:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 32407:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 32408:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 32409:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 32410:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 32411:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 32412:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 32413:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 32414:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 32415:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 32416:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 32417:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 32418:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 32419:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 32420:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 32421:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 32422:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 32423:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 32424:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 32425:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 32426:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 32427:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 32428:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 32429:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 32430:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 32431:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 32432:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 32433:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 32434:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 32435:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 32436:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 32437:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 32438:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 32439:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 32440:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 32441:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 32442:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 32443:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 32444:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 32445:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 32446:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 32447:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 32448:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 32449:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 32450:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 32451:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 32452:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 32453:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 32454:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 32455:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 32456:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 32457:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 32458:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 32459:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 32460:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 32461:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 32462:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 32463:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 32464:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 32465:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 32466:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 32467:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 32468:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 32469:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 32470:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 32471:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 32472:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 32473:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 32474:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 32475:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 32476:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 32477:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 32478:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 32479:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 32480:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 32481:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 32482:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 32483:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 32484:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 32485:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 32486:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 32487:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 32488:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 32489:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 32490:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 32491:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 32492:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 32493:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 32494:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 32495:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 32496:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 32497:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 32498:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 32499:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 32500:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 32501:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 32502:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 32503:20]
  assign io_z = ~x26; // @[Snxn100k.scala 32504:16]
endmodule
module SnxnLv4Inst114(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 32859:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 32860:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 32861:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 32862:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 32863:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 32864:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 32865:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 32866:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 32867:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 32868:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 32869:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 32870:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 32871:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 32872:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 32873:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 32874:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 32875:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 32876:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 32877:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 32878:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 32879:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 32880:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 32881:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 32882:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 32883:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 32884:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 32885:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 32886:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 32887:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 32888:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 32889:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 32890:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 32891:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 32892:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 32893:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 32894:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 32895:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 32896:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 32897:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 32898:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 32899:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 32900:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 32901:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 32902:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 32903:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 32904:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 32905:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 32906:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 32907:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 32908:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 32909:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 32910:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 32911:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 32912:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 32913:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 32914:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 32915:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 32916:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 32917:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 32918:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 32919:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 32920:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 32921:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 32922:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 32923:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 32924:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 32925:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 32926:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 32927:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 32928:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 32929:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 32930:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 32931:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 32932:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 32933:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 32934:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 32935:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 32936:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 32937:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 32938:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 32939:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 32940:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 32941:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 32942:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 32943:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 32944:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 32945:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 32946:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 32947:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 32948:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 32949:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 32950:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 32951:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 32952:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 32953:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 32954:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 32955:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 32956:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 32957:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 32958:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 32959:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 32960:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 32961:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 32962:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 32963:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 32964:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 32965:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 32966:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 32967:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 32968:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 32969:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 32970:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 32971:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 32972:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 32973:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 32974:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 32975:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 32976:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 32977:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 32978:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 32979:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 32980:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 32981:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 32982:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 32983:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 32984:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 32985:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 32986:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 32987:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 32988:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 32989:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 32990:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 32991:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 32992:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 32993:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 32994:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 32995:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 32996:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 32997:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 32998:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 32999:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 33000:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 33001:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 33002:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 33003:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 33004:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 33005:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 33006:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 33007:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 33008:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 33009:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 33010:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 33011:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 33012:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 33013:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 33014:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 33015:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 33016:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 33017:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 33018:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 33019:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 33020:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 33021:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 33022:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 33023:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 33024:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 33025:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 33026:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 33027:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 33028:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 33029:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 33030:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 33031:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 33032:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 33033:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 33034:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 33035:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 33036:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 33037:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 33038:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 33039:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 33040:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 33041:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 33042:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 33043:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 33044:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 33045:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 33046:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 33047:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 33048:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 33049:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 33050:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 33051:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 33052:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 33053:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 33054:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 33055:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 33056:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 33057:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 33058:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 33059:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 33060:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 33061:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 33062:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 33063:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 33064:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 33065:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 33066:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 33067:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 33068:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 33069:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 33070:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 33071:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 33072:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 33073:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 33074:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 33075:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 33076:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 33077:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 33078:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 33079:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 33080:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 33081:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 33082:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 33083:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 33084:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 33085:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 33086:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 33087:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 33088:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 33089:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 33090:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 33091:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 33092:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 33093:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 33094:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 33095:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 33096:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 33097:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 33098:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 33099:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 33100:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 33101:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 33102:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 33103:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 33104:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 33105:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 33106:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 33107:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 33108:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 33109:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 33110:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 33111:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 33112:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 33113:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 33114:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 33115:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 33116:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 33117:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 33118:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 33119:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 33120:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 33121:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 33122:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 33123:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 33124:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 33125:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 33126:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 33127:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 33128:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 33129:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 33130:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 33131:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 33132:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 33133:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 33134:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 33135:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 33136:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 33137:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 33138:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 33139:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 33140:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 33141:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 33142:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 33143:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 33144:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 33145:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 33146:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 33147:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 33148:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 33149:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 33150:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 33151:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 33152:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 33153:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 33154:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 33155:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 33156:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 33157:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 33158:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 33159:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 33160:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 33161:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 33162:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 33163:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 33164:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 33165:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 33166:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 33167:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 33168:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 33169:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 33170:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 33171:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 33172:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 33173:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 33174:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 33175:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 33176:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 33177:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 33178:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 33179:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 33180:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 33181:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 33182:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 33183:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 33184:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 33185:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 33186:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 33187:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 33188:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 33189:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 33190:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 33191:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 33192:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 33193:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 33194:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 33195:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 33196:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 33197:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 33198:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 33199:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 33200:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 33201:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 33202:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 33203:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 33204:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 33205:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 33206:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 33207:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 33208:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 33209:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 33210:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 33211:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 33212:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 33213:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 33214:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 33215:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 33216:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 33217:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 33218:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 33219:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 33220:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 33221:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 33222:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 33223:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 33224:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 33225:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 33226:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 33227:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 33228:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 33229:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 33230:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 33231:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 33232:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 33233:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 33234:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 33235:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 33236:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 33237:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 33238:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 33239:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 33240:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 33241:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 33242:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 33243:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 33244:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 33245:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 33246:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 33247:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 33248:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 33249:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 33250:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 33251:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 33252:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 33253:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 33254:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 33255:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 33256:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 33257:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 33258:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 33259:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 33260:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 33261:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 33262:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 33263:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 33264:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 33265:22]
  assign io_z = ~x101; // @[Snxn100k.scala 33266:17]
endmodule
module SnxnLv3Inst28(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst112_io_a; // @[Snxn100k.scala 9758:35]
  wire  inst_SnxnLv4Inst112_io_b; // @[Snxn100k.scala 9758:35]
  wire  inst_SnxnLv4Inst112_io_z; // @[Snxn100k.scala 9758:35]
  wire  inst_SnxnLv4Inst113_io_a; // @[Snxn100k.scala 9762:35]
  wire  inst_SnxnLv4Inst113_io_b; // @[Snxn100k.scala 9762:35]
  wire  inst_SnxnLv4Inst113_io_z; // @[Snxn100k.scala 9762:35]
  wire  inst_SnxnLv4Inst114_io_a; // @[Snxn100k.scala 9766:35]
  wire  inst_SnxnLv4Inst114_io_b; // @[Snxn100k.scala 9766:35]
  wire  inst_SnxnLv4Inst114_io_z; // @[Snxn100k.scala 9766:35]
  wire  inst_SnxnLv4Inst115_io_a; // @[Snxn100k.scala 9770:35]
  wire  inst_SnxnLv4Inst115_io_b; // @[Snxn100k.scala 9770:35]
  wire  inst_SnxnLv4Inst115_io_z; // @[Snxn100k.scala 9770:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst112_io_z + inst_SnxnLv4Inst113_io_z; // @[Snxn100k.scala 9774:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst114_io_z; // @[Snxn100k.scala 9774:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst115_io_z; // @[Snxn100k.scala 9774:92]
  SnxnLv4Inst31 inst_SnxnLv4Inst112 ( // @[Snxn100k.scala 9758:35]
    .io_a(inst_SnxnLv4Inst112_io_a),
    .io_b(inst_SnxnLv4Inst112_io_b),
    .io_z(inst_SnxnLv4Inst112_io_z)
  );
  SnxnLv4Inst113 inst_SnxnLv4Inst113 ( // @[Snxn100k.scala 9762:35]
    .io_a(inst_SnxnLv4Inst113_io_a),
    .io_b(inst_SnxnLv4Inst113_io_b),
    .io_z(inst_SnxnLv4Inst113_io_z)
  );
  SnxnLv4Inst114 inst_SnxnLv4Inst114 ( // @[Snxn100k.scala 9766:35]
    .io_a(inst_SnxnLv4Inst114_io_a),
    .io_b(inst_SnxnLv4Inst114_io_b),
    .io_z(inst_SnxnLv4Inst114_io_z)
  );
  SnxnLv4Inst113 inst_SnxnLv4Inst115 ( // @[Snxn100k.scala 9770:35]
    .io_a(inst_SnxnLv4Inst115_io_a),
    .io_b(inst_SnxnLv4Inst115_io_b),
    .io_z(inst_SnxnLv4Inst115_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 9775:15]
  assign inst_SnxnLv4Inst112_io_a = io_a; // @[Snxn100k.scala 9759:28]
  assign inst_SnxnLv4Inst112_io_b = io_b; // @[Snxn100k.scala 9760:28]
  assign inst_SnxnLv4Inst113_io_a = io_a; // @[Snxn100k.scala 9763:28]
  assign inst_SnxnLv4Inst113_io_b = io_b; // @[Snxn100k.scala 9764:28]
  assign inst_SnxnLv4Inst114_io_a = io_a; // @[Snxn100k.scala 9767:28]
  assign inst_SnxnLv4Inst114_io_b = io_b; // @[Snxn100k.scala 9768:28]
  assign inst_SnxnLv4Inst115_io_a = io_a; // @[Snxn100k.scala 9771:28]
  assign inst_SnxnLv4Inst115_io_b = io_b; // @[Snxn100k.scala 9772:28]
endmodule
module SnxnLv4Inst119(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 30945:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 30946:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 30947:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 30948:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 30949:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 30950:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 30951:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 30952:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 30953:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 30954:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 30955:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 30956:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 30957:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 30958:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 30959:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 30960:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 30961:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 30962:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 30963:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 30964:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 30965:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 30966:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 30967:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 30968:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 30969:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 30970:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 30971:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 30972:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 30973:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 30974:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 30975:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 30976:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 30977:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 30978:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 30979:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 30980:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 30981:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 30982:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 30983:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 30984:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 30985:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 30986:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 30987:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 30988:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 30989:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 30990:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 30991:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 30992:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 30993:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 30994:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 30995:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 30996:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 30997:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 30998:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 30999:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 31000:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 31001:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 31002:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 31003:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 31004:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 31005:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 31006:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 31007:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 31008:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 31009:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 31010:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 31011:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 31012:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 31013:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 31014:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 31015:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 31016:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 31017:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 31018:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 31019:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 31020:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 31021:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 31022:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 31023:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 31024:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 31025:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 31026:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 31027:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 31028:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 31029:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 31030:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 31031:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 31032:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 31033:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 31034:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 31035:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 31036:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 31037:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 31038:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 31039:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 31040:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 31041:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 31042:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 31043:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 31044:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 31045:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 31046:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 31047:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 31048:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 31049:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 31050:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 31051:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 31052:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 31053:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 31054:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 31055:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 31056:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 31057:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 31058:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 31059:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 31060:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 31061:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 31062:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 31063:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 31064:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 31065:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 31066:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 31067:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 31068:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 31069:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 31070:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 31071:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 31072:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 31073:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 31074:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 31075:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 31076:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 31077:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 31078:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 31079:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 31080:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 31081:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 31082:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 31083:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 31084:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 31085:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 31086:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 31087:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 31088:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 31089:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 31090:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 31091:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 31092:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 31093:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 31094:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 31095:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 31096:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 31097:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 31098:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 31099:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 31100:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 31101:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 31102:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 31103:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 31104:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 31105:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 31106:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 31107:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 31108:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 31109:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 31110:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 31111:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 31112:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 31113:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 31114:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 31115:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 31116:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 31117:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 31118:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 31119:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 31120:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 31121:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 31122:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 31123:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 31124:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 31125:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 31126:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 31127:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 31128:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 31129:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 31130:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 31131:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 31132:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 31133:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 31134:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 31135:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 31136:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 31137:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 31138:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 31139:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 31140:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 31141:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 31142:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 31143:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 31144:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 31145:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 31146:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 31147:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 31148:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 31149:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 31150:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 31151:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 31152:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 31153:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 31154:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 31155:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 31156:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 31157:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 31158:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 31159:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 31160:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 31161:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 31162:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 31163:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 31164:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 31165:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 31166:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 31167:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 31168:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 31169:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 31170:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 31171:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 31172:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 31173:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 31174:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 31175:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 31176:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 31177:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 31178:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 31179:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 31180:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 31181:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 31182:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 31183:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 31184:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 31185:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 31186:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 31187:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 31188:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 31189:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 31190:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 31191:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 31192:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 31193:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 31194:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 31195:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 31196:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 31197:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 31198:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 31199:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 31200:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 31201:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 31202:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 31203:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 31204:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 31205:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 31206:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 31207:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 31208:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 31209:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 31210:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 31211:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 31212:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 31213:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 31214:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 31215:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 31216:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 31217:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 31218:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 31219:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 31220:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 31221:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 31222:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 31223:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 31224:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 31225:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 31226:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 31227:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 31228:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 31229:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 31230:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 31231:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 31232:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 31233:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 31234:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 31235:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 31236:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 31237:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 31238:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 31239:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 31240:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 31241:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 31242:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 31243:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 31244:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 31245:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 31246:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 31247:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 31248:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 31249:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 31250:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 31251:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 31252:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 31253:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 31254:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 31255:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 31256:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 31257:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 31258:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 31259:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 31260:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 31261:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 31262:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 31263:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 31264:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 31265:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 31266:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 31267:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 31268:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 31269:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 31270:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 31271:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 31272:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 31273:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 31274:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 31275:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 31276:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 31277:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 31278:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 31279:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 31280:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 31281:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 31282:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 31283:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 31284:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 31285:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 31286:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 31287:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 31288:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 31289:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 31290:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 31291:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 31292:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 31293:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 31294:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 31295:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 31296:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 31297:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 31298:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 31299:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 31300:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 31301:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 31302:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 31303:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 31304:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 31305:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 31306:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 31307:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 31308:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 31309:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 31310:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 31311:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 31312:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 31313:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 31314:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 31315:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 31316:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 31317:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 31318:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 31319:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 31320:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 31321:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 31322:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 31323:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 31324:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 31325:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 31326:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 31327:20]
  assign io_z = ~x95; // @[Snxn100k.scala 31328:16]
endmodule
module SnxnLv3Inst29(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst116_io_a; // @[Snxn100k.scala 9024:35]
  wire  inst_SnxnLv4Inst116_io_b; // @[Snxn100k.scala 9024:35]
  wire  inst_SnxnLv4Inst116_io_z; // @[Snxn100k.scala 9024:35]
  wire  inst_SnxnLv4Inst117_io_a; // @[Snxn100k.scala 9028:35]
  wire  inst_SnxnLv4Inst117_io_b; // @[Snxn100k.scala 9028:35]
  wire  inst_SnxnLv4Inst117_io_z; // @[Snxn100k.scala 9028:35]
  wire  inst_SnxnLv4Inst118_io_a; // @[Snxn100k.scala 9032:35]
  wire  inst_SnxnLv4Inst118_io_b; // @[Snxn100k.scala 9032:35]
  wire  inst_SnxnLv4Inst118_io_z; // @[Snxn100k.scala 9032:35]
  wire  inst_SnxnLv4Inst119_io_a; // @[Snxn100k.scala 9036:35]
  wire  inst_SnxnLv4Inst119_io_b; // @[Snxn100k.scala 9036:35]
  wire  inst_SnxnLv4Inst119_io_z; // @[Snxn100k.scala 9036:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst116_io_z + inst_SnxnLv4Inst117_io_z; // @[Snxn100k.scala 9040:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst118_io_z; // @[Snxn100k.scala 9040:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst119_io_z; // @[Snxn100k.scala 9040:92]
  SnxnLv4Inst104 inst_SnxnLv4Inst116 ( // @[Snxn100k.scala 9024:35]
    .io_a(inst_SnxnLv4Inst116_io_a),
    .io_b(inst_SnxnLv4Inst116_io_b),
    .io_z(inst_SnxnLv4Inst116_io_z)
  );
  SnxnLv4Inst27 inst_SnxnLv4Inst117 ( // @[Snxn100k.scala 9028:35]
    .io_a(inst_SnxnLv4Inst117_io_a),
    .io_b(inst_SnxnLv4Inst117_io_b),
    .io_z(inst_SnxnLv4Inst117_io_z)
  );
  SnxnLv4Inst40 inst_SnxnLv4Inst118 ( // @[Snxn100k.scala 9032:35]
    .io_a(inst_SnxnLv4Inst118_io_a),
    .io_b(inst_SnxnLv4Inst118_io_b),
    .io_z(inst_SnxnLv4Inst118_io_z)
  );
  SnxnLv4Inst119 inst_SnxnLv4Inst119 ( // @[Snxn100k.scala 9036:35]
    .io_a(inst_SnxnLv4Inst119_io_a),
    .io_b(inst_SnxnLv4Inst119_io_b),
    .io_z(inst_SnxnLv4Inst119_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 9041:15]
  assign inst_SnxnLv4Inst116_io_a = io_a; // @[Snxn100k.scala 9025:28]
  assign inst_SnxnLv4Inst116_io_b = io_b; // @[Snxn100k.scala 9026:28]
  assign inst_SnxnLv4Inst117_io_a = io_a; // @[Snxn100k.scala 9029:28]
  assign inst_SnxnLv4Inst117_io_b = io_b; // @[Snxn100k.scala 9030:28]
  assign inst_SnxnLv4Inst118_io_a = io_a; // @[Snxn100k.scala 9033:28]
  assign inst_SnxnLv4Inst118_io_b = io_b; // @[Snxn100k.scala 9034:28]
  assign inst_SnxnLv4Inst119_io_a = io_a; // @[Snxn100k.scala 9037:28]
  assign inst_SnxnLv4Inst119_io_b = io_b; // @[Snxn100k.scala 9038:28]
endmodule
module SnxnLv4Inst120(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 31389:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 31390:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 31391:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 31392:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 31393:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 31394:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 31395:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 31396:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 31397:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 31398:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 31399:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 31400:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 31401:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 31402:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 31403:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 31404:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 31405:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 31406:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 31407:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 31408:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 31409:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 31410:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 31411:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 31412:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 31413:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 31414:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 31415:18]
  assign io_z = ~x6; // @[Snxn100k.scala 31416:15]
endmodule
module SnxnLv4Inst122(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 32319:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 32320:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 32321:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 32322:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 32323:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 32324:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 32325:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 32326:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 32327:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 32328:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 32329:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 32330:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 32331:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 32332:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 32333:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 32334:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 32335:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 32336:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 32337:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 32338:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 32339:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 32340:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 32341:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 32342:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 32343:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 32344:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 32345:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 32346:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 32347:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 32348:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 32349:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 32350:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 32351:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 32352:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 32353:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 32354:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 32355:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 32356:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 32357:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 32358:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 32359:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 32360:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 32361:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 32362:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 32363:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 32364:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 32365:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 32366:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 32367:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 32368:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 32369:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 32370:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 32371:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 32372:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 32373:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 32374:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 32375:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 32376:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 32377:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 32378:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 32379:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 32380:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 32381:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 32382:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 32383:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 32384:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 32385:20]
  assign io_z = ~x16; // @[Snxn100k.scala 32386:16]
endmodule
module SnxnLv3Inst30(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst120_io_a; // @[Snxn100k.scala 9391:35]
  wire  inst_SnxnLv4Inst120_io_b; // @[Snxn100k.scala 9391:35]
  wire  inst_SnxnLv4Inst120_io_z; // @[Snxn100k.scala 9391:35]
  wire  inst_SnxnLv4Inst121_io_a; // @[Snxn100k.scala 9395:35]
  wire  inst_SnxnLv4Inst121_io_b; // @[Snxn100k.scala 9395:35]
  wire  inst_SnxnLv4Inst121_io_z; // @[Snxn100k.scala 9395:35]
  wire  inst_SnxnLv4Inst122_io_a; // @[Snxn100k.scala 9399:35]
  wire  inst_SnxnLv4Inst122_io_b; // @[Snxn100k.scala 9399:35]
  wire  inst_SnxnLv4Inst122_io_z; // @[Snxn100k.scala 9399:35]
  wire  inst_SnxnLv4Inst123_io_a; // @[Snxn100k.scala 9403:35]
  wire  inst_SnxnLv4Inst123_io_b; // @[Snxn100k.scala 9403:35]
  wire  inst_SnxnLv4Inst123_io_z; // @[Snxn100k.scala 9403:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst120_io_z + inst_SnxnLv4Inst121_io_z; // @[Snxn100k.scala 9407:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst122_io_z; // @[Snxn100k.scala 9407:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst123_io_z; // @[Snxn100k.scala 9407:92]
  SnxnLv4Inst120 inst_SnxnLv4Inst120 ( // @[Snxn100k.scala 9391:35]
    .io_a(inst_SnxnLv4Inst120_io_a),
    .io_b(inst_SnxnLv4Inst120_io_b),
    .io_z(inst_SnxnLv4Inst120_io_z)
  );
  SnxnLv4Inst52 inst_SnxnLv4Inst121 ( // @[Snxn100k.scala 9395:35]
    .io_a(inst_SnxnLv4Inst121_io_a),
    .io_b(inst_SnxnLv4Inst121_io_b),
    .io_z(inst_SnxnLv4Inst121_io_z)
  );
  SnxnLv4Inst122 inst_SnxnLv4Inst122 ( // @[Snxn100k.scala 9399:35]
    .io_a(inst_SnxnLv4Inst122_io_a),
    .io_b(inst_SnxnLv4Inst122_io_b),
    .io_z(inst_SnxnLv4Inst122_io_z)
  );
  SnxnLv4Inst32 inst_SnxnLv4Inst123 ( // @[Snxn100k.scala 9403:35]
    .io_a(inst_SnxnLv4Inst123_io_a),
    .io_b(inst_SnxnLv4Inst123_io_b),
    .io_z(inst_SnxnLv4Inst123_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 9408:15]
  assign inst_SnxnLv4Inst120_io_a = io_a; // @[Snxn100k.scala 9392:28]
  assign inst_SnxnLv4Inst120_io_b = io_b; // @[Snxn100k.scala 9393:28]
  assign inst_SnxnLv4Inst121_io_a = io_a; // @[Snxn100k.scala 9396:28]
  assign inst_SnxnLv4Inst121_io_b = io_b; // @[Snxn100k.scala 9397:28]
  assign inst_SnxnLv4Inst122_io_a = io_a; // @[Snxn100k.scala 9400:28]
  assign inst_SnxnLv4Inst122_io_b = io_b; // @[Snxn100k.scala 9401:28]
  assign inst_SnxnLv4Inst123_io_a = io_a; // @[Snxn100k.scala 9404:28]
  assign inst_SnxnLv4Inst123_io_b = io_b; // @[Snxn100k.scala 9405:28]
endmodule
module SnxnLv4Inst124(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 33277:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 33278:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 33279:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 33280:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 33281:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 33282:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 33283:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 33284:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 33285:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 33286:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 33287:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 33288:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 33289:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 33290:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 33291:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 33292:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 33293:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 33294:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 33295:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 33296:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 33297:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 33298:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 33299:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 33300:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 33301:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 33302:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 33303:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 33304:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 33305:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 33306:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 33307:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 33308:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 33309:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 33310:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 33311:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 33312:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 33313:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 33314:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 33315:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 33316:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 33317:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 33318:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 33319:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 33320:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 33321:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 33322:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 33323:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 33324:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 33325:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 33326:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 33327:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 33328:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 33329:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 33330:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 33331:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 33332:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 33333:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 33334:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 33335:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 33336:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 33337:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 33338:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 33339:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 33340:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 33341:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 33342:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 33343:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 33344:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 33345:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 33346:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 33347:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 33348:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 33349:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 33350:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 33351:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 33352:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 33353:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 33354:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 33355:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 33356:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 33357:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 33358:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 33359:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 33360:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 33361:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 33362:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 33363:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 33364:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 33365:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 33366:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 33367:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 33368:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 33369:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 33370:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 33371:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 33372:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 33373:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 33374:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 33375:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 33376:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 33377:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 33378:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 33379:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 33380:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 33381:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 33382:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 33383:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 33384:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 33385:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 33386:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 33387:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 33388:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 33389:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 33390:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 33391:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 33392:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 33393:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 33394:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 33395:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 33396:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 33397:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 33398:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 33399:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 33400:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 33401:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 33402:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 33403:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 33404:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 33405:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 33406:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 33407:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 33408:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 33409:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 33410:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 33411:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 33412:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 33413:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 33414:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 33415:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 33416:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 33417:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 33418:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 33419:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 33420:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 33421:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 33422:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 33423:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 33424:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 33425:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 33426:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 33427:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 33428:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 33429:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 33430:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 33431:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 33432:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 33433:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 33434:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 33435:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 33436:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 33437:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 33438:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 33439:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 33440:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 33441:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 33442:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 33443:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 33444:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 33445:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 33446:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 33447:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 33448:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 33449:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 33450:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 33451:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 33452:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 33453:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 33454:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 33455:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 33456:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 33457:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 33458:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 33459:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 33460:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 33461:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 33462:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 33463:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 33464:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 33465:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 33466:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 33467:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 33468:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 33469:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 33470:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 33471:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 33472:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 33473:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 33474:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 33475:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 33476:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 33477:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 33478:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 33479:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 33480:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 33481:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 33482:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 33483:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 33484:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 33485:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 33486:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 33487:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 33488:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 33489:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 33490:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 33491:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 33492:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 33493:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 33494:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 33495:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 33496:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 33497:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 33498:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 33499:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 33500:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 33501:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 33502:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 33503:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 33504:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 33505:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 33506:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 33507:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 33508:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 33509:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 33510:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 33511:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 33512:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 33513:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 33514:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 33515:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 33516:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 33517:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 33518:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 33519:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 33520:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 33521:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 33522:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 33523:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 33524:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 33525:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 33526:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 33527:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 33528:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 33529:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 33530:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 33531:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 33532:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 33533:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 33534:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 33535:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 33536:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 33537:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 33538:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 33539:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 33540:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 33541:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 33542:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 33543:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 33544:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 33545:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 33546:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 33547:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 33548:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 33549:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 33550:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 33551:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 33552:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 33553:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 33554:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 33555:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 33556:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 33557:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 33558:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 33559:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 33560:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 33561:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 33562:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 33563:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 33564:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 33565:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 33566:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 33567:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 33568:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 33569:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 33570:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 33571:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 33572:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 33573:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 33574:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 33575:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 33576:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 33577:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 33578:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 33579:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 33580:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 33581:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 33582:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 33583:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 33584:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 33585:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 33586:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 33587:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 33588:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 33589:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 33590:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 33591:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 33592:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 33593:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 33594:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 33595:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 33596:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 33597:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 33598:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 33599:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 33600:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 33601:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 33602:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 33603:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 33604:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 33605:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 33606:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 33607:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 33608:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 33609:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 33610:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 33611:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 33612:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 33613:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 33614:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 33615:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 33616:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 33617:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 33618:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 33619:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 33620:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 33621:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 33622:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 33623:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 33624:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 33625:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 33626:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 33627:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 33628:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 33629:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 33630:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 33631:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 33632:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 33633:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 33634:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 33635:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 33636:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 33637:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 33638:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 33639:20]
  assign io_z = ~x90; // @[Snxn100k.scala 33640:16]
endmodule
module SnxnLv4Inst127(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 34751:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 34752:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 34753:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 34754:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 34755:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 34756:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 34757:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 34758:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 34759:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 34760:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 34761:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 34762:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 34763:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 34764:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 34765:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 34766:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 34767:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 34768:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 34769:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 34770:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 34771:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 34772:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 34773:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 34774:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 34775:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 34776:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 34777:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 34778:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 34779:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 34780:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 34781:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 34782:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 34783:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 34784:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 34785:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 34786:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 34787:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 34788:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 34789:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 34790:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 34791:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 34792:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 34793:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 34794:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 34795:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 34796:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 34797:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 34798:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 34799:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 34800:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 34801:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 34802:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 34803:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 34804:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 34805:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 34806:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 34807:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 34808:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 34809:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 34810:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 34811:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 34812:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 34813:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 34814:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 34815:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 34816:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 34817:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 34818:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 34819:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 34820:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 34821:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 34822:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 34823:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 34824:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 34825:20]
  assign io_z = ~x18; // @[Snxn100k.scala 34826:16]
endmodule
module SnxnLv3Inst31(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst124_io_a; // @[Snxn100k.scala 10157:35]
  wire  inst_SnxnLv4Inst124_io_b; // @[Snxn100k.scala 10157:35]
  wire  inst_SnxnLv4Inst124_io_z; // @[Snxn100k.scala 10157:35]
  wire  inst_SnxnLv4Inst125_io_a; // @[Snxn100k.scala 10161:35]
  wire  inst_SnxnLv4Inst125_io_b; // @[Snxn100k.scala 10161:35]
  wire  inst_SnxnLv4Inst125_io_z; // @[Snxn100k.scala 10161:35]
  wire  inst_SnxnLv4Inst126_io_a; // @[Snxn100k.scala 10165:35]
  wire  inst_SnxnLv4Inst126_io_b; // @[Snxn100k.scala 10165:35]
  wire  inst_SnxnLv4Inst126_io_z; // @[Snxn100k.scala 10165:35]
  wire  inst_SnxnLv4Inst127_io_a; // @[Snxn100k.scala 10169:35]
  wire  inst_SnxnLv4Inst127_io_b; // @[Snxn100k.scala 10169:35]
  wire  inst_SnxnLv4Inst127_io_z; // @[Snxn100k.scala 10169:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst124_io_z + inst_SnxnLv4Inst125_io_z; // @[Snxn100k.scala 10173:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst126_io_z; // @[Snxn100k.scala 10173:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst127_io_z; // @[Snxn100k.scala 10173:92]
  SnxnLv4Inst124 inst_SnxnLv4Inst124 ( // @[Snxn100k.scala 10157:35]
    .io_a(inst_SnxnLv4Inst124_io_a),
    .io_b(inst_SnxnLv4Inst124_io_b),
    .io_z(inst_SnxnLv4Inst124_io_z)
  );
  SnxnLv4Inst24 inst_SnxnLv4Inst125 ( // @[Snxn100k.scala 10161:35]
    .io_a(inst_SnxnLv4Inst125_io_a),
    .io_b(inst_SnxnLv4Inst125_io_b),
    .io_z(inst_SnxnLv4Inst125_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst126 ( // @[Snxn100k.scala 10165:35]
    .io_a(inst_SnxnLv4Inst126_io_a),
    .io_b(inst_SnxnLv4Inst126_io_b),
    .io_z(inst_SnxnLv4Inst126_io_z)
  );
  SnxnLv4Inst127 inst_SnxnLv4Inst127 ( // @[Snxn100k.scala 10169:35]
    .io_a(inst_SnxnLv4Inst127_io_a),
    .io_b(inst_SnxnLv4Inst127_io_b),
    .io_z(inst_SnxnLv4Inst127_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 10174:15]
  assign inst_SnxnLv4Inst124_io_a = io_a; // @[Snxn100k.scala 10158:28]
  assign inst_SnxnLv4Inst124_io_b = io_b; // @[Snxn100k.scala 10159:28]
  assign inst_SnxnLv4Inst125_io_a = io_a; // @[Snxn100k.scala 10162:28]
  assign inst_SnxnLv4Inst125_io_b = io_b; // @[Snxn100k.scala 10163:28]
  assign inst_SnxnLv4Inst126_io_a = io_a; // @[Snxn100k.scala 10166:28]
  assign inst_SnxnLv4Inst126_io_b = io_b; // @[Snxn100k.scala 10167:28]
  assign inst_SnxnLv4Inst127_io_a = io_a; // @[Snxn100k.scala 10170:28]
  assign inst_SnxnLv4Inst127_io_b = io_b; // @[Snxn100k.scala 10171:28]
endmodule
module SnxnLv2Inst7(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst28_io_a; // @[Snxn100k.scala 1852:34]
  wire  inst_SnxnLv3Inst28_io_b; // @[Snxn100k.scala 1852:34]
  wire  inst_SnxnLv3Inst28_io_z; // @[Snxn100k.scala 1852:34]
  wire  inst_SnxnLv3Inst29_io_a; // @[Snxn100k.scala 1856:34]
  wire  inst_SnxnLv3Inst29_io_b; // @[Snxn100k.scala 1856:34]
  wire  inst_SnxnLv3Inst29_io_z; // @[Snxn100k.scala 1856:34]
  wire  inst_SnxnLv3Inst30_io_a; // @[Snxn100k.scala 1860:34]
  wire  inst_SnxnLv3Inst30_io_b; // @[Snxn100k.scala 1860:34]
  wire  inst_SnxnLv3Inst30_io_z; // @[Snxn100k.scala 1860:34]
  wire  inst_SnxnLv3Inst31_io_a; // @[Snxn100k.scala 1864:34]
  wire  inst_SnxnLv3Inst31_io_b; // @[Snxn100k.scala 1864:34]
  wire  inst_SnxnLv3Inst31_io_z; // @[Snxn100k.scala 1864:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst28_io_z + inst_SnxnLv3Inst29_io_z; // @[Snxn100k.scala 1868:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst30_io_z; // @[Snxn100k.scala 1868:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst31_io_z; // @[Snxn100k.scala 1868:89]
  SnxnLv3Inst28 inst_SnxnLv3Inst28 ( // @[Snxn100k.scala 1852:34]
    .io_a(inst_SnxnLv3Inst28_io_a),
    .io_b(inst_SnxnLv3Inst28_io_b),
    .io_z(inst_SnxnLv3Inst28_io_z)
  );
  SnxnLv3Inst29 inst_SnxnLv3Inst29 ( // @[Snxn100k.scala 1856:34]
    .io_a(inst_SnxnLv3Inst29_io_a),
    .io_b(inst_SnxnLv3Inst29_io_b),
    .io_z(inst_SnxnLv3Inst29_io_z)
  );
  SnxnLv3Inst30 inst_SnxnLv3Inst30 ( // @[Snxn100k.scala 1860:34]
    .io_a(inst_SnxnLv3Inst30_io_a),
    .io_b(inst_SnxnLv3Inst30_io_b),
    .io_z(inst_SnxnLv3Inst30_io_z)
  );
  SnxnLv3Inst31 inst_SnxnLv3Inst31 ( // @[Snxn100k.scala 1864:34]
    .io_a(inst_SnxnLv3Inst31_io_a),
    .io_b(inst_SnxnLv3Inst31_io_b),
    .io_z(inst_SnxnLv3Inst31_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1869:15]
  assign inst_SnxnLv3Inst28_io_a = io_a; // @[Snxn100k.scala 1853:27]
  assign inst_SnxnLv3Inst28_io_b = io_b; // @[Snxn100k.scala 1854:27]
  assign inst_SnxnLv3Inst29_io_a = io_a; // @[Snxn100k.scala 1857:27]
  assign inst_SnxnLv3Inst29_io_b = io_b; // @[Snxn100k.scala 1858:27]
  assign inst_SnxnLv3Inst30_io_a = io_a; // @[Snxn100k.scala 1861:27]
  assign inst_SnxnLv3Inst30_io_b = io_b; // @[Snxn100k.scala 1862:27]
  assign inst_SnxnLv3Inst31_io_a = io_a; // @[Snxn100k.scala 1865:27]
  assign inst_SnxnLv3Inst31_io_b = io_b; // @[Snxn100k.scala 1866:27]
endmodule
module SnxnLv1Inst1(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst4_io_a; // @[Snxn100k.scala 616:33]
  wire  inst_SnxnLv2Inst4_io_b; // @[Snxn100k.scala 616:33]
  wire  inst_SnxnLv2Inst4_io_z; // @[Snxn100k.scala 616:33]
  wire  inst_SnxnLv2Inst5_io_a; // @[Snxn100k.scala 620:33]
  wire  inst_SnxnLv2Inst5_io_b; // @[Snxn100k.scala 620:33]
  wire  inst_SnxnLv2Inst5_io_z; // @[Snxn100k.scala 620:33]
  wire  inst_SnxnLv2Inst6_io_a; // @[Snxn100k.scala 624:33]
  wire  inst_SnxnLv2Inst6_io_b; // @[Snxn100k.scala 624:33]
  wire  inst_SnxnLv2Inst6_io_z; // @[Snxn100k.scala 624:33]
  wire  inst_SnxnLv2Inst7_io_a; // @[Snxn100k.scala 628:33]
  wire  inst_SnxnLv2Inst7_io_b; // @[Snxn100k.scala 628:33]
  wire  inst_SnxnLv2Inst7_io_z; // @[Snxn100k.scala 628:33]
  wire  _sum_T_1 = inst_SnxnLv2Inst4_io_z + inst_SnxnLv2Inst5_io_z; // @[Snxn100k.scala 632:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst6_io_z; // @[Snxn100k.scala 632:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst7_io_z; // @[Snxn100k.scala 632:86]
  SnxnLv2Inst4 inst_SnxnLv2Inst4 ( // @[Snxn100k.scala 616:33]
    .io_a(inst_SnxnLv2Inst4_io_a),
    .io_b(inst_SnxnLv2Inst4_io_b),
    .io_z(inst_SnxnLv2Inst4_io_z)
  );
  SnxnLv2Inst5 inst_SnxnLv2Inst5 ( // @[Snxn100k.scala 620:33]
    .io_a(inst_SnxnLv2Inst5_io_a),
    .io_b(inst_SnxnLv2Inst5_io_b),
    .io_z(inst_SnxnLv2Inst5_io_z)
  );
  SnxnLv2Inst6 inst_SnxnLv2Inst6 ( // @[Snxn100k.scala 624:33]
    .io_a(inst_SnxnLv2Inst6_io_a),
    .io_b(inst_SnxnLv2Inst6_io_b),
    .io_z(inst_SnxnLv2Inst6_io_z)
  );
  SnxnLv2Inst7 inst_SnxnLv2Inst7 ( // @[Snxn100k.scala 628:33]
    .io_a(inst_SnxnLv2Inst7_io_a),
    .io_b(inst_SnxnLv2Inst7_io_b),
    .io_z(inst_SnxnLv2Inst7_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 633:15]
  assign inst_SnxnLv2Inst4_io_a = io_a; // @[Snxn100k.scala 617:26]
  assign inst_SnxnLv2Inst4_io_b = io_b; // @[Snxn100k.scala 618:26]
  assign inst_SnxnLv2Inst5_io_a = io_a; // @[Snxn100k.scala 621:26]
  assign inst_SnxnLv2Inst5_io_b = io_b; // @[Snxn100k.scala 622:26]
  assign inst_SnxnLv2Inst6_io_a = io_a; // @[Snxn100k.scala 625:26]
  assign inst_SnxnLv2Inst6_io_b = io_b; // @[Snxn100k.scala 626:26]
  assign inst_SnxnLv2Inst7_io_a = io_a; // @[Snxn100k.scala 629:26]
  assign inst_SnxnLv2Inst7_io_b = io_b; // @[Snxn100k.scala 630:26]
endmodule
module SnxnLv4Inst129(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 101905:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 101906:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 101907:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 101908:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 101909:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 101910:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 101911:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 101912:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 101913:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 101914:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 101915:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 101916:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 101917:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 101918:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 101919:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 101920:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 101921:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 101922:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 101923:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 101924:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 101925:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 101926:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 101927:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 101928:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 101929:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 101930:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 101931:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 101932:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 101933:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 101934:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 101935:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 101936:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 101937:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 101938:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 101939:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 101940:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 101941:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 101942:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 101943:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 101944:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 101945:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 101946:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 101947:20]
  assign io_z = ~x10; // @[Snxn100k.scala 101948:16]
endmodule
module SnxnLv4Inst130(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 102405:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 102406:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 102407:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 102408:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 102409:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 102410:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 102411:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 102412:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 102413:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 102414:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 102415:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 102416:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 102417:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 102418:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 102419:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 102420:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 102421:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 102422:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 102423:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 102424:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 102425:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 102426:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 102427:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 102428:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 102429:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 102430:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 102431:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 102432:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 102433:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 102434:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 102435:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 102436:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 102437:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 102438:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 102439:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 102440:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 102441:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 102442:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 102443:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 102444:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 102445:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 102446:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 102447:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 102448:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 102449:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 102450:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 102451:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 102452:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 102453:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 102454:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 102455:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 102456:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 102457:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 102458:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 102459:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 102460:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 102461:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 102462:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 102463:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 102464:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 102465:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 102466:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 102467:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 102468:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 102469:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 102470:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 102471:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 102472:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 102473:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 102474:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 102475:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 102476:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 102477:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 102478:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 102479:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 102480:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 102481:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 102482:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 102483:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 102484:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 102485:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 102486:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 102487:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 102488:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 102489:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 102490:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 102491:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 102492:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 102493:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 102494:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 102495:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 102496:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 102497:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 102498:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 102499:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 102500:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 102501:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 102502:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 102503:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 102504:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 102505:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 102506:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 102507:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 102508:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 102509:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 102510:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 102511:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 102512:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 102513:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 102514:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 102515:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 102516:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 102517:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 102518:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 102519:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 102520:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 102521:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 102522:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 102523:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 102524:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 102525:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 102526:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 102527:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 102528:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 102529:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 102530:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 102531:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 102532:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 102533:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 102534:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 102535:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 102536:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 102537:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 102538:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 102539:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 102540:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 102541:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 102542:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 102543:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 102544:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 102545:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 102546:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 102547:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 102548:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 102549:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 102550:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 102551:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 102552:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 102553:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 102554:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 102555:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 102556:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 102557:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 102558:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 102559:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 102560:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 102561:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 102562:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 102563:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 102564:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 102565:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 102566:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 102567:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 102568:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 102569:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 102570:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 102571:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 102572:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 102573:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 102574:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 102575:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 102576:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 102577:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 102578:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 102579:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 102580:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 102581:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 102582:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 102583:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 102584:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 102585:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 102586:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 102587:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 102588:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 102589:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 102590:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 102591:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 102592:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 102593:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 102594:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 102595:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 102596:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 102597:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 102598:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 102599:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 102600:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 102601:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 102602:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 102603:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 102604:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 102605:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 102606:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 102607:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 102608:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 102609:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 102610:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 102611:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 102612:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 102613:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 102614:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 102615:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 102616:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 102617:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 102618:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 102619:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 102620:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 102621:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 102622:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 102623:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 102624:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 102625:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 102626:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 102627:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 102628:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 102629:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 102630:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 102631:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 102632:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 102633:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 102634:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 102635:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 102636:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 102637:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 102638:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 102639:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 102640:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 102641:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 102642:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 102643:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 102644:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 102645:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 102646:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 102647:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 102648:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 102649:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 102650:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 102651:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 102652:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 102653:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 102654:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 102655:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 102656:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 102657:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 102658:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 102659:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 102660:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 102661:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 102662:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 102663:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 102664:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 102665:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 102666:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 102667:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 102668:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 102669:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 102670:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 102671:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 102672:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 102673:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 102674:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 102675:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 102676:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 102677:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 102678:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 102679:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 102680:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 102681:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 102682:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 102683:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 102684:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 102685:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 102686:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 102687:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 102688:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 102689:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 102690:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 102691:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 102692:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 102693:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 102694:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 102695:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 102696:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 102697:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 102698:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 102699:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 102700:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 102701:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 102702:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 102703:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 102704:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 102705:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 102706:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 102707:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 102708:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 102709:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 102710:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 102711:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 102712:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 102713:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 102714:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 102715:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 102716:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 102717:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 102718:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 102719:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 102720:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 102721:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 102722:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 102723:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 102724:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 102725:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 102726:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 102727:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 102728:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 102729:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 102730:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 102731:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 102732:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 102733:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 102734:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 102735:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 102736:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 102737:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 102738:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 102739:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 102740:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 102741:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 102742:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 102743:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 102744:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 102745:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 102746:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 102747:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 102748:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 102749:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 102750:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 102751:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 102752:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 102753:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 102754:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 102755:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 102756:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 102757:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 102758:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 102759:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 102760:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 102761:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 102762:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 102763:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 102764:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 102765:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 102766:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 102767:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 102768:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 102769:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 102770:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 102771:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 102772:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 102773:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 102774:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 102775:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 102776:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 102777:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 102778:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 102779:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 102780:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 102781:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 102782:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 102783:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 102784:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 102785:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 102786:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 102787:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 102788:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 102789:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 102790:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 102791:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 102792:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 102793:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 102794:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 102795:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 102796:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 102797:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 102798:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 102799:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 102800:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 102801:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 102802:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 102803:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 102804:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 102805:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 102806:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 102807:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 102808:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 102809:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 102810:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 102811:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 102812:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 102813:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 102814:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 102815:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 102816:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 102817:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 102818:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 102819:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 102820:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 102821:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 102822:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 102823:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 102824:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 102825:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 102826:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 102827:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 102828:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 102829:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 102830:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 102831:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 102832:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 102833:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 102834:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 102835:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 102836:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 102837:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 102838:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 102839:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 102840:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 102841:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 102842:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 102843:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 102844:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 102845:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 102846:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 102847:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 102848:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 102849:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 102850:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 102851:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 102852:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 102853:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 102854:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 102855:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 102856:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 102857:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 102858:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 102859:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 102860:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 102861:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 102862:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 102863:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 102864:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 102865:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 102866:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 102867:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 102868:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 102869:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 102870:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 102871:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 102872:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 102873:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 102874:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 102875:22]
  assign io_z = ~x117; // @[Snxn100k.scala 102876:17]
endmodule
module SnxnLv3Inst32(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst128_io_a; // @[Snxn100k.scala 29149:35]
  wire  inst_SnxnLv4Inst128_io_b; // @[Snxn100k.scala 29149:35]
  wire  inst_SnxnLv4Inst128_io_z; // @[Snxn100k.scala 29149:35]
  wire  inst_SnxnLv4Inst129_io_a; // @[Snxn100k.scala 29153:35]
  wire  inst_SnxnLv4Inst129_io_b; // @[Snxn100k.scala 29153:35]
  wire  inst_SnxnLv4Inst129_io_z; // @[Snxn100k.scala 29153:35]
  wire  inst_SnxnLv4Inst130_io_a; // @[Snxn100k.scala 29157:35]
  wire  inst_SnxnLv4Inst130_io_b; // @[Snxn100k.scala 29157:35]
  wire  inst_SnxnLv4Inst130_io_z; // @[Snxn100k.scala 29157:35]
  wire  inst_SnxnLv4Inst131_io_a; // @[Snxn100k.scala 29161:35]
  wire  inst_SnxnLv4Inst131_io_b; // @[Snxn100k.scala 29161:35]
  wire  inst_SnxnLv4Inst131_io_z; // @[Snxn100k.scala 29161:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst128_io_z + inst_SnxnLv4Inst129_io_z; // @[Snxn100k.scala 29165:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst130_io_z; // @[Snxn100k.scala 29165:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst131_io_z; // @[Snxn100k.scala 29165:92]
  SnxnLv4Inst38 inst_SnxnLv4Inst128 ( // @[Snxn100k.scala 29149:35]
    .io_a(inst_SnxnLv4Inst128_io_a),
    .io_b(inst_SnxnLv4Inst128_io_b),
    .io_z(inst_SnxnLv4Inst128_io_z)
  );
  SnxnLv4Inst129 inst_SnxnLv4Inst129 ( // @[Snxn100k.scala 29153:35]
    .io_a(inst_SnxnLv4Inst129_io_a),
    .io_b(inst_SnxnLv4Inst129_io_b),
    .io_z(inst_SnxnLv4Inst129_io_z)
  );
  SnxnLv4Inst130 inst_SnxnLv4Inst130 ( // @[Snxn100k.scala 29157:35]
    .io_a(inst_SnxnLv4Inst130_io_a),
    .io_b(inst_SnxnLv4Inst130_io_b),
    .io_z(inst_SnxnLv4Inst130_io_z)
  );
  SnxnLv4Inst86 inst_SnxnLv4Inst131 ( // @[Snxn100k.scala 29161:35]
    .io_a(inst_SnxnLv4Inst131_io_a),
    .io_b(inst_SnxnLv4Inst131_io_b),
    .io_z(inst_SnxnLv4Inst131_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 29166:15]
  assign inst_SnxnLv4Inst128_io_a = io_a; // @[Snxn100k.scala 29150:28]
  assign inst_SnxnLv4Inst128_io_b = io_b; // @[Snxn100k.scala 29151:28]
  assign inst_SnxnLv4Inst129_io_a = io_a; // @[Snxn100k.scala 29154:28]
  assign inst_SnxnLv4Inst129_io_b = io_b; // @[Snxn100k.scala 29155:28]
  assign inst_SnxnLv4Inst130_io_a = io_a; // @[Snxn100k.scala 29158:28]
  assign inst_SnxnLv4Inst130_io_b = io_b; // @[Snxn100k.scala 29159:28]
  assign inst_SnxnLv4Inst131_io_a = io_a; // @[Snxn100k.scala 29162:28]
  assign inst_SnxnLv4Inst131_io_b = io_b; // @[Snxn100k.scala 29163:28]
endmodule
module SnxnLv4Inst134(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 99839:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 99840:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 99841:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 99842:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 99843:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 99844:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 99845:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 99846:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 99847:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 99848:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 99849:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 99850:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 99851:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 99852:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 99853:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 99854:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 99855:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 99856:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 99857:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 99858:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 99859:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 99860:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 99861:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 99862:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 99863:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 99864:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 99865:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 99866:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 99867:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 99868:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 99869:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 99870:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 99871:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 99872:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 99873:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 99874:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 99875:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 99876:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 99877:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 99878:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 99879:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 99880:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 99881:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 99882:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 99883:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 99884:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 99885:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 99886:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 99887:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 99888:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 99889:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 99890:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 99891:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 99892:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 99893:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 99894:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 99895:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 99896:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 99897:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 99898:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 99899:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 99900:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 99901:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 99902:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 99903:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 99904:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 99905:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 99906:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 99907:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 99908:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 99909:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 99910:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 99911:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 99912:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 99913:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 99914:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 99915:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 99916:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 99917:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 99918:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 99919:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 99920:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 99921:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 99922:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 99923:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 99924:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 99925:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 99926:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 99927:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 99928:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 99929:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 99930:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 99931:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 99932:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 99933:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 99934:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 99935:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 99936:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 99937:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 99938:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 99939:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 99940:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 99941:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 99942:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 99943:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 99944:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 99945:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 99946:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 99947:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 99948:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 99949:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 99950:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 99951:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 99952:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 99953:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 99954:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 99955:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 99956:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 99957:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 99958:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 99959:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 99960:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 99961:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 99962:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 99963:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 99964:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 99965:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 99966:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 99967:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 99968:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 99969:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 99970:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 99971:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 99972:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 99973:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 99974:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 99975:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 99976:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 99977:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 99978:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 99979:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 99980:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 99981:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 99982:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 99983:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 99984:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 99985:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 99986:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 99987:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 99988:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 99989:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 99990:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 99991:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 99992:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 99993:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 99994:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 99995:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 99996:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 99997:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 99998:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 99999:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 100000:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 100001:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 100002:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 100003:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 100004:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 100005:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 100006:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 100007:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 100008:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 100009:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 100010:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 100011:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 100012:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 100013:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 100014:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 100015:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 100016:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 100017:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 100018:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 100019:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 100020:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 100021:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 100022:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 100023:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 100024:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 100025:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 100026:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 100027:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 100028:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 100029:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 100030:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 100031:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 100032:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 100033:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 100034:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 100035:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 100036:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 100037:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 100038:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 100039:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 100040:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 100041:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 100042:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 100043:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 100044:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 100045:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 100046:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 100047:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 100048:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 100049:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 100050:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 100051:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 100052:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 100053:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 100054:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 100055:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 100056:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 100057:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 100058:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 100059:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 100060:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 100061:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 100062:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 100063:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 100064:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 100065:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 100066:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 100067:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 100068:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 100069:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 100070:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 100071:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 100072:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 100073:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 100074:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 100075:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 100076:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 100077:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 100078:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 100079:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 100080:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 100081:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 100082:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 100083:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 100084:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 100085:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 100086:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 100087:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 100088:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 100089:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 100090:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 100091:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 100092:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 100093:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 100094:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 100095:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 100096:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 100097:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 100098:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 100099:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 100100:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 100101:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 100102:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 100103:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 100104:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 100105:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 100106:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 100107:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 100108:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 100109:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 100110:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 100111:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 100112:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 100113:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 100114:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 100115:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 100116:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 100117:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 100118:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 100119:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 100120:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 100121:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 100122:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 100123:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 100124:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 100125:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 100126:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 100127:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 100128:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 100129:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 100130:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 100131:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 100132:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 100133:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 100134:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 100135:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 100136:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 100137:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 100138:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 100139:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 100140:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 100141:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 100142:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 100143:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 100144:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 100145:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 100146:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 100147:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 100148:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 100149:20]
  assign io_z = ~x77; // @[Snxn100k.scala 100150:16]
endmodule
module SnxnLv3Inst33(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst132_io_a; // @[Snxn100k.scala 28626:35]
  wire  inst_SnxnLv4Inst132_io_b; // @[Snxn100k.scala 28626:35]
  wire  inst_SnxnLv4Inst132_io_z; // @[Snxn100k.scala 28626:35]
  wire  inst_SnxnLv4Inst133_io_a; // @[Snxn100k.scala 28630:35]
  wire  inst_SnxnLv4Inst133_io_b; // @[Snxn100k.scala 28630:35]
  wire  inst_SnxnLv4Inst133_io_z; // @[Snxn100k.scala 28630:35]
  wire  inst_SnxnLv4Inst134_io_a; // @[Snxn100k.scala 28634:35]
  wire  inst_SnxnLv4Inst134_io_b; // @[Snxn100k.scala 28634:35]
  wire  inst_SnxnLv4Inst134_io_z; // @[Snxn100k.scala 28634:35]
  wire  inst_SnxnLv4Inst135_io_a; // @[Snxn100k.scala 28638:35]
  wire  inst_SnxnLv4Inst135_io_b; // @[Snxn100k.scala 28638:35]
  wire  inst_SnxnLv4Inst135_io_z; // @[Snxn100k.scala 28638:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst132_io_z + inst_SnxnLv4Inst133_io_z; // @[Snxn100k.scala 28642:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst134_io_z; // @[Snxn100k.scala 28642:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst135_io_z; // @[Snxn100k.scala 28642:92]
  SnxnLv4Inst33 inst_SnxnLv4Inst132 ( // @[Snxn100k.scala 28626:35]
    .io_a(inst_SnxnLv4Inst132_io_a),
    .io_b(inst_SnxnLv4Inst132_io_b),
    .io_z(inst_SnxnLv4Inst132_io_z)
  );
  SnxnLv4Inst51 inst_SnxnLv4Inst133 ( // @[Snxn100k.scala 28630:35]
    .io_a(inst_SnxnLv4Inst133_io_a),
    .io_b(inst_SnxnLv4Inst133_io_b),
    .io_z(inst_SnxnLv4Inst133_io_z)
  );
  SnxnLv4Inst134 inst_SnxnLv4Inst134 ( // @[Snxn100k.scala 28634:35]
    .io_a(inst_SnxnLv4Inst134_io_a),
    .io_b(inst_SnxnLv4Inst134_io_b),
    .io_z(inst_SnxnLv4Inst134_io_z)
  );
  SnxnLv4Inst18 inst_SnxnLv4Inst135 ( // @[Snxn100k.scala 28638:35]
    .io_a(inst_SnxnLv4Inst135_io_a),
    .io_b(inst_SnxnLv4Inst135_io_b),
    .io_z(inst_SnxnLv4Inst135_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 28643:15]
  assign inst_SnxnLv4Inst132_io_a = io_a; // @[Snxn100k.scala 28627:28]
  assign inst_SnxnLv4Inst132_io_b = io_b; // @[Snxn100k.scala 28628:28]
  assign inst_SnxnLv4Inst133_io_a = io_a; // @[Snxn100k.scala 28631:28]
  assign inst_SnxnLv4Inst133_io_b = io_b; // @[Snxn100k.scala 28632:28]
  assign inst_SnxnLv4Inst134_io_a = io_a; // @[Snxn100k.scala 28635:28]
  assign inst_SnxnLv4Inst134_io_b = io_b; // @[Snxn100k.scala 28636:28]
  assign inst_SnxnLv4Inst135_io_a = io_a; // @[Snxn100k.scala 28639:28]
  assign inst_SnxnLv4Inst135_io_b = io_b; // @[Snxn100k.scala 28640:28]
endmodule
module SnxnLv3Inst34(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst136_io_a; // @[Snxn100k.scala 30343:35]
  wire  inst_SnxnLv4Inst136_io_b; // @[Snxn100k.scala 30343:35]
  wire  inst_SnxnLv4Inst136_io_z; // @[Snxn100k.scala 30343:35]
  wire  inst_SnxnLv4Inst137_io_a; // @[Snxn100k.scala 30347:35]
  wire  inst_SnxnLv4Inst137_io_b; // @[Snxn100k.scala 30347:35]
  wire  inst_SnxnLv4Inst137_io_z; // @[Snxn100k.scala 30347:35]
  wire  inst_SnxnLv4Inst138_io_a; // @[Snxn100k.scala 30351:35]
  wire  inst_SnxnLv4Inst138_io_b; // @[Snxn100k.scala 30351:35]
  wire  inst_SnxnLv4Inst138_io_z; // @[Snxn100k.scala 30351:35]
  wire  inst_SnxnLv4Inst139_io_a; // @[Snxn100k.scala 30355:35]
  wire  inst_SnxnLv4Inst139_io_b; // @[Snxn100k.scala 30355:35]
  wire  inst_SnxnLv4Inst139_io_z; // @[Snxn100k.scala 30355:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst136_io_z + inst_SnxnLv4Inst137_io_z; // @[Snxn100k.scala 30359:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst138_io_z; // @[Snxn100k.scala 30359:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst139_io_z; // @[Snxn100k.scala 30359:92]
  SnxnLv4Inst47 inst_SnxnLv4Inst136 ( // @[Snxn100k.scala 30343:35]
    .io_a(inst_SnxnLv4Inst136_io_a),
    .io_b(inst_SnxnLv4Inst136_io_b),
    .io_z(inst_SnxnLv4Inst136_io_z)
  );
  SnxnLv4Inst24 inst_SnxnLv4Inst137 ( // @[Snxn100k.scala 30347:35]
    .io_a(inst_SnxnLv4Inst137_io_a),
    .io_b(inst_SnxnLv4Inst137_io_b),
    .io_z(inst_SnxnLv4Inst137_io_z)
  );
  SnxnLv4Inst114 inst_SnxnLv4Inst138 ( // @[Snxn100k.scala 30351:35]
    .io_a(inst_SnxnLv4Inst138_io_a),
    .io_b(inst_SnxnLv4Inst138_io_b),
    .io_z(inst_SnxnLv4Inst138_io_z)
  );
  SnxnLv4Inst56 inst_SnxnLv4Inst139 ( // @[Snxn100k.scala 30355:35]
    .io_a(inst_SnxnLv4Inst139_io_a),
    .io_b(inst_SnxnLv4Inst139_io_b),
    .io_z(inst_SnxnLv4Inst139_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 30360:15]
  assign inst_SnxnLv4Inst136_io_a = io_a; // @[Snxn100k.scala 30344:28]
  assign inst_SnxnLv4Inst136_io_b = io_b; // @[Snxn100k.scala 30345:28]
  assign inst_SnxnLv4Inst137_io_a = io_a; // @[Snxn100k.scala 30348:28]
  assign inst_SnxnLv4Inst137_io_b = io_b; // @[Snxn100k.scala 30349:28]
  assign inst_SnxnLv4Inst138_io_a = io_a; // @[Snxn100k.scala 30352:28]
  assign inst_SnxnLv4Inst138_io_b = io_b; // @[Snxn100k.scala 30353:28]
  assign inst_SnxnLv4Inst139_io_a = io_a; // @[Snxn100k.scala 30356:28]
  assign inst_SnxnLv4Inst139_io_b = io_b; // @[Snxn100k.scala 30357:28]
endmodule
module SnxnLv4Inst140(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 103215:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 103216:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 103217:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 103218:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 103219:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 103220:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 103221:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 103222:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 103223:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 103224:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 103225:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 103226:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 103227:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 103228:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 103229:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 103230:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 103231:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 103232:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 103233:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 103234:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 103235:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 103236:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 103237:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 103238:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 103239:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 103240:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 103241:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 103242:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 103243:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 103244:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 103245:18]
  assign io_z = ~x7; // @[Snxn100k.scala 103246:15]
endmodule
module SnxnLv4Inst142(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 102917:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 102918:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 102919:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 102920:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 102921:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 102922:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 102923:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 102924:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 102925:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 102926:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 102927:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 102928:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 102929:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 102930:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 102931:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 102932:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 102933:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 102934:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 102935:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 102936:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 102937:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 102938:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 102939:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 102940:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 102941:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 102942:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 102943:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 102944:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 102945:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 102946:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 102947:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 102948:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 102949:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 102950:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 102951:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 102952:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 102953:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 102954:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 102955:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 102956:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 102957:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 102958:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 102959:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 102960:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 102961:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 102962:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 102963:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 102964:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 102965:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 102966:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 102967:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 102968:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 102969:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 102970:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 102971:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 102972:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 102973:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 102974:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 102975:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 102976:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 102977:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 102978:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 102979:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 102980:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 102981:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 102982:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 102983:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 102984:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 102985:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 102986:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 102987:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 102988:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 102989:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 102990:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 102991:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 102992:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 102993:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 102994:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 102995:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 102996:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 102997:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 102998:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 102999:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 103000:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 103001:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 103002:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 103003:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 103004:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 103005:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 103006:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 103007:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 103008:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 103009:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 103010:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 103011:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 103012:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 103013:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 103014:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 103015:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 103016:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 103017:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 103018:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 103019:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 103020:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 103021:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 103022:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 103023:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 103024:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 103025:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 103026:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 103027:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 103028:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 103029:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 103030:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 103031:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 103032:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 103033:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 103034:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 103035:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 103036:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 103037:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 103038:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 103039:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 103040:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 103041:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 103042:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 103043:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 103044:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 103045:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 103046:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 103047:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 103048:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 103049:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 103050:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 103051:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 103052:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 103053:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 103054:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 103055:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 103056:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 103057:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 103058:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 103059:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 103060:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 103061:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 103062:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 103063:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 103064:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 103065:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 103066:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 103067:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 103068:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 103069:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 103070:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 103071:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 103072:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 103073:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 103074:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 103075:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 103076:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 103077:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 103078:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 103079:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 103080:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 103081:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 103082:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 103083:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 103084:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 103085:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 103086:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 103087:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 103088:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 103089:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 103090:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 103091:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 103092:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 103093:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 103094:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 103095:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 103096:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 103097:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 103098:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 103099:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 103100:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 103101:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 103102:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 103103:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 103104:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 103105:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 103106:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 103107:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 103108:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 103109:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 103110:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 103111:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 103112:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 103113:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 103114:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 103115:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 103116:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 103117:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 103118:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 103119:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 103120:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 103121:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 103122:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 103123:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 103124:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 103125:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 103126:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 103127:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 103128:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 103129:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 103130:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 103131:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 103132:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 103133:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 103134:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 103135:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 103136:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 103137:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 103138:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 103139:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 103140:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 103141:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 103142:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 103143:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 103144:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 103145:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 103146:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 103147:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 103148:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 103149:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 103150:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 103151:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 103152:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 103153:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 103154:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 103155:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 103156:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 103157:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 103158:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 103159:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 103160:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 103161:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 103162:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 103163:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 103164:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 103165:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 103166:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 103167:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 103168:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 103169:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 103170:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 103171:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 103172:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 103173:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 103174:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 103175:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 103176:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 103177:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 103178:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 103179:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 103180:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 103181:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 103182:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 103183:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 103184:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 103185:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 103186:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 103187:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 103188:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 103189:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 103190:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 103191:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 103192:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 103193:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 103194:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 103195:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 103196:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 103197:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 103198:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 103199:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 103200:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 103201:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 103202:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 103203:20]
  assign io_z = ~x71; // @[Snxn100k.scala 103204:16]
endmodule
module SnxnLv3Inst35(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst140_io_a; // @[Snxn100k.scala 29744:35]
  wire  inst_SnxnLv4Inst140_io_b; // @[Snxn100k.scala 29744:35]
  wire  inst_SnxnLv4Inst140_io_z; // @[Snxn100k.scala 29744:35]
  wire  inst_SnxnLv4Inst141_io_a; // @[Snxn100k.scala 29748:35]
  wire  inst_SnxnLv4Inst141_io_b; // @[Snxn100k.scala 29748:35]
  wire  inst_SnxnLv4Inst141_io_z; // @[Snxn100k.scala 29748:35]
  wire  inst_SnxnLv4Inst142_io_a; // @[Snxn100k.scala 29752:35]
  wire  inst_SnxnLv4Inst142_io_b; // @[Snxn100k.scala 29752:35]
  wire  inst_SnxnLv4Inst142_io_z; // @[Snxn100k.scala 29752:35]
  wire  inst_SnxnLv4Inst143_io_a; // @[Snxn100k.scala 29756:35]
  wire  inst_SnxnLv4Inst143_io_b; // @[Snxn100k.scala 29756:35]
  wire  inst_SnxnLv4Inst143_io_z; // @[Snxn100k.scala 29756:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst140_io_z + inst_SnxnLv4Inst141_io_z; // @[Snxn100k.scala 29760:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst142_io_z; // @[Snxn100k.scala 29760:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst143_io_z; // @[Snxn100k.scala 29760:92]
  SnxnLv4Inst140 inst_SnxnLv4Inst140 ( // @[Snxn100k.scala 29744:35]
    .io_a(inst_SnxnLv4Inst140_io_a),
    .io_b(inst_SnxnLv4Inst140_io_b),
    .io_z(inst_SnxnLv4Inst140_io_z)
  );
  SnxnLv4Inst49 inst_SnxnLv4Inst141 ( // @[Snxn100k.scala 29748:35]
    .io_a(inst_SnxnLv4Inst141_io_a),
    .io_b(inst_SnxnLv4Inst141_io_b),
    .io_z(inst_SnxnLv4Inst141_io_z)
  );
  SnxnLv4Inst142 inst_SnxnLv4Inst142 ( // @[Snxn100k.scala 29752:35]
    .io_a(inst_SnxnLv4Inst142_io_a),
    .io_b(inst_SnxnLv4Inst142_io_b),
    .io_z(inst_SnxnLv4Inst142_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst143 ( // @[Snxn100k.scala 29756:35]
    .io_a(inst_SnxnLv4Inst143_io_a),
    .io_b(inst_SnxnLv4Inst143_io_b),
    .io_z(inst_SnxnLv4Inst143_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 29761:15]
  assign inst_SnxnLv4Inst140_io_a = io_a; // @[Snxn100k.scala 29745:28]
  assign inst_SnxnLv4Inst140_io_b = io_b; // @[Snxn100k.scala 29746:28]
  assign inst_SnxnLv4Inst141_io_a = io_a; // @[Snxn100k.scala 29749:28]
  assign inst_SnxnLv4Inst141_io_b = io_b; // @[Snxn100k.scala 29750:28]
  assign inst_SnxnLv4Inst142_io_a = io_a; // @[Snxn100k.scala 29753:28]
  assign inst_SnxnLv4Inst142_io_b = io_b; // @[Snxn100k.scala 29754:28]
  assign inst_SnxnLv4Inst143_io_a = io_a; // @[Snxn100k.scala 29757:28]
  assign inst_SnxnLv4Inst143_io_b = io_b; // @[Snxn100k.scala 29758:28]
endmodule
module SnxnLv2Inst8(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst32_io_a; // @[Snxn100k.scala 8781:34]
  wire  inst_SnxnLv3Inst32_io_b; // @[Snxn100k.scala 8781:34]
  wire  inst_SnxnLv3Inst32_io_z; // @[Snxn100k.scala 8781:34]
  wire  inst_SnxnLv3Inst33_io_a; // @[Snxn100k.scala 8785:34]
  wire  inst_SnxnLv3Inst33_io_b; // @[Snxn100k.scala 8785:34]
  wire  inst_SnxnLv3Inst33_io_z; // @[Snxn100k.scala 8785:34]
  wire  inst_SnxnLv3Inst34_io_a; // @[Snxn100k.scala 8789:34]
  wire  inst_SnxnLv3Inst34_io_b; // @[Snxn100k.scala 8789:34]
  wire  inst_SnxnLv3Inst34_io_z; // @[Snxn100k.scala 8789:34]
  wire  inst_SnxnLv3Inst35_io_a; // @[Snxn100k.scala 8793:34]
  wire  inst_SnxnLv3Inst35_io_b; // @[Snxn100k.scala 8793:34]
  wire  inst_SnxnLv3Inst35_io_z; // @[Snxn100k.scala 8793:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst32_io_z + inst_SnxnLv3Inst33_io_z; // @[Snxn100k.scala 8797:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst34_io_z; // @[Snxn100k.scala 8797:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst35_io_z; // @[Snxn100k.scala 8797:89]
  SnxnLv3Inst32 inst_SnxnLv3Inst32 ( // @[Snxn100k.scala 8781:34]
    .io_a(inst_SnxnLv3Inst32_io_a),
    .io_b(inst_SnxnLv3Inst32_io_b),
    .io_z(inst_SnxnLv3Inst32_io_z)
  );
  SnxnLv3Inst33 inst_SnxnLv3Inst33 ( // @[Snxn100k.scala 8785:34]
    .io_a(inst_SnxnLv3Inst33_io_a),
    .io_b(inst_SnxnLv3Inst33_io_b),
    .io_z(inst_SnxnLv3Inst33_io_z)
  );
  SnxnLv3Inst34 inst_SnxnLv3Inst34 ( // @[Snxn100k.scala 8789:34]
    .io_a(inst_SnxnLv3Inst34_io_a),
    .io_b(inst_SnxnLv3Inst34_io_b),
    .io_z(inst_SnxnLv3Inst34_io_z)
  );
  SnxnLv3Inst35 inst_SnxnLv3Inst35 ( // @[Snxn100k.scala 8793:34]
    .io_a(inst_SnxnLv3Inst35_io_a),
    .io_b(inst_SnxnLv3Inst35_io_b),
    .io_z(inst_SnxnLv3Inst35_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 8798:15]
  assign inst_SnxnLv3Inst32_io_a = io_a; // @[Snxn100k.scala 8782:27]
  assign inst_SnxnLv3Inst32_io_b = io_b; // @[Snxn100k.scala 8783:27]
  assign inst_SnxnLv3Inst33_io_a = io_a; // @[Snxn100k.scala 8786:27]
  assign inst_SnxnLv3Inst33_io_b = io_b; // @[Snxn100k.scala 8787:27]
  assign inst_SnxnLv3Inst34_io_a = io_a; // @[Snxn100k.scala 8790:27]
  assign inst_SnxnLv3Inst34_io_b = io_b; // @[Snxn100k.scala 8791:27]
  assign inst_SnxnLv3Inst35_io_a = io_a; // @[Snxn100k.scala 8794:27]
  assign inst_SnxnLv3Inst35_io_b = io_b; // @[Snxn100k.scala 8795:27]
endmodule
module SnxnLv4Inst146(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 83309:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 83310:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 83311:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 83312:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 83313:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 83314:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 83315:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 83316:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 83317:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 83318:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 83319:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 83320:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 83321:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 83322:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 83323:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 83324:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 83325:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 83326:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 83327:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 83328:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 83329:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 83330:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 83331:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 83332:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 83333:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 83334:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 83335:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 83336:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 83337:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 83338:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 83339:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 83340:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 83341:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 83342:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 83343:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 83344:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 83345:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 83346:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 83347:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 83348:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 83349:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 83350:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 83351:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 83352:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 83353:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 83354:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 83355:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 83356:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 83357:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 83358:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 83359:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 83360:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 83361:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 83362:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 83363:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 83364:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 83365:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 83366:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 83367:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 83368:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 83369:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 83370:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 83371:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 83372:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 83373:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 83374:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 83375:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 83376:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 83377:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 83378:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 83379:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 83380:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 83381:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 83382:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 83383:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 83384:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 83385:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 83386:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 83387:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 83388:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 83389:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 83390:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 83391:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 83392:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 83393:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 83394:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 83395:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 83396:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 83397:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 83398:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 83399:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 83400:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 83401:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 83402:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 83403:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 83404:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 83405:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 83406:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 83407:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 83408:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 83409:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 83410:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 83411:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 83412:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 83413:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 83414:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 83415:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 83416:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 83417:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 83418:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 83419:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 83420:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 83421:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 83422:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 83423:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 83424:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 83425:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 83426:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 83427:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 83428:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 83429:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 83430:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 83431:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 83432:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 83433:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 83434:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 83435:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 83436:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 83437:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 83438:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 83439:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 83440:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 83441:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 83442:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 83443:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 83444:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 83445:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 83446:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 83447:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 83448:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 83449:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 83450:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 83451:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 83452:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 83453:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 83454:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 83455:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 83456:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 83457:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 83458:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 83459:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 83460:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 83461:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 83462:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 83463:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 83464:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 83465:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 83466:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 83467:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 83468:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 83469:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 83470:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 83471:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 83472:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 83473:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 83474:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 83475:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 83476:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 83477:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 83478:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 83479:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 83480:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 83481:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 83482:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 83483:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 83484:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 83485:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 83486:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 83487:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 83488:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 83489:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 83490:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 83491:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 83492:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 83493:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 83494:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 83495:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 83496:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 83497:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 83498:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 83499:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 83500:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 83501:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 83502:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 83503:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 83504:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 83505:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 83506:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 83507:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 83508:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 83509:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 83510:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 83511:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 83512:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 83513:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 83514:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 83515:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 83516:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 83517:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 83518:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 83519:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 83520:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 83521:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 83522:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 83523:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 83524:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 83525:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 83526:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 83527:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 83528:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 83529:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 83530:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 83531:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 83532:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 83533:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 83534:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 83535:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 83536:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 83537:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 83538:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 83539:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 83540:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 83541:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 83542:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 83543:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 83544:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 83545:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 83546:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 83547:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 83548:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 83549:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 83550:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 83551:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 83552:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 83553:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 83554:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 83555:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 83556:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 83557:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 83558:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 83559:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 83560:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 83561:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 83562:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 83563:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 83564:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 83565:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 83566:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 83567:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 83568:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 83569:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 83570:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 83571:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 83572:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 83573:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 83574:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 83575:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 83576:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 83577:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 83578:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 83579:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 83580:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 83581:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 83582:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 83583:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 83584:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 83585:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 83586:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 83587:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 83588:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 83589:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 83590:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 83591:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 83592:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 83593:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 83594:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 83595:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 83596:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 83597:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 83598:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 83599:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 83600:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 83601:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 83602:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 83603:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 83604:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 83605:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 83606:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 83607:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 83608:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 83609:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 83610:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 83611:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 83612:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 83613:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 83614:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 83615:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 83616:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 83617:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 83618:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 83619:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 83620:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 83621:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 83622:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 83623:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 83624:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 83625:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 83626:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 83627:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 83628:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 83629:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 83630:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 83631:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 83632:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 83633:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 83634:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 83635:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 83636:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 83637:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 83638:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 83639:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 83640:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 83641:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 83642:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 83643:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 83644:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 83645:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 83646:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 83647:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 83648:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 83649:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 83650:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 83651:20]
  assign io_z = ~x85; // @[Snxn100k.scala 83652:16]
endmodule
module SnxnLv4Inst147(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 83663:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 83664:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 83665:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 83666:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 83667:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 83668:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 83669:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 83670:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 83671:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 83672:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 83673:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 83674:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 83675:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 83676:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 83677:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 83678:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 83679:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 83680:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 83681:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 83682:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 83683:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 83684:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 83685:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 83686:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 83687:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 83688:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 83689:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 83690:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 83691:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 83692:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 83693:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 83694:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 83695:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 83696:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 83697:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 83698:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 83699:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 83700:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 83701:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 83702:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 83703:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 83704:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 83705:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 83706:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 83707:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 83708:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 83709:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 83710:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 83711:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 83712:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 83713:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 83714:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 83715:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 83716:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 83717:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 83718:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 83719:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 83720:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 83721:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 83722:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 83723:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 83724:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 83725:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 83726:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 83727:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 83728:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 83729:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 83730:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 83731:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 83732:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 83733:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 83734:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 83735:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 83736:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 83737:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 83738:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 83739:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 83740:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 83741:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 83742:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 83743:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 83744:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 83745:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 83746:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 83747:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 83748:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 83749:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 83750:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 83751:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 83752:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 83753:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 83754:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 83755:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 83756:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 83757:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 83758:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 83759:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 83760:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 83761:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 83762:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 83763:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 83764:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 83765:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 83766:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 83767:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 83768:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 83769:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 83770:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 83771:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 83772:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 83773:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 83774:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 83775:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 83776:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 83777:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 83778:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 83779:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 83780:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 83781:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 83782:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 83783:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 83784:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 83785:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 83786:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 83787:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 83788:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 83789:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 83790:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 83791:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 83792:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 83793:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 83794:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 83795:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 83796:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 83797:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 83798:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 83799:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 83800:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 83801:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 83802:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 83803:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 83804:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 83805:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 83806:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 83807:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 83808:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 83809:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 83810:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 83811:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 83812:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 83813:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 83814:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 83815:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 83816:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 83817:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 83818:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 83819:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 83820:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 83821:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 83822:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 83823:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 83824:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 83825:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 83826:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 83827:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 83828:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 83829:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 83830:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 83831:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 83832:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 83833:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 83834:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 83835:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 83836:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 83837:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 83838:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 83839:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 83840:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 83841:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 83842:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 83843:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 83844:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 83845:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 83846:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 83847:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 83848:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 83849:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 83850:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 83851:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 83852:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 83853:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 83854:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 83855:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 83856:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 83857:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 83858:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 83859:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 83860:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 83861:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 83862:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 83863:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 83864:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 83865:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 83866:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 83867:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 83868:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 83869:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 83870:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 83871:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 83872:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 83873:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 83874:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 83875:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 83876:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 83877:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 83878:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 83879:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 83880:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 83881:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 83882:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 83883:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 83884:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 83885:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 83886:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 83887:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 83888:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 83889:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 83890:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 83891:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 83892:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 83893:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 83894:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 83895:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 83896:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 83897:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 83898:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 83899:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 83900:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 83901:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 83902:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 83903:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 83904:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 83905:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 83906:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 83907:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 83908:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 83909:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 83910:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 83911:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 83912:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 83913:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 83914:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 83915:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 83916:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 83917:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 83918:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 83919:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 83920:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 83921:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 83922:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 83923:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 83924:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 83925:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 83926:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 83927:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 83928:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 83929:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 83930:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 83931:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 83932:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 83933:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 83934:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 83935:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 83936:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 83937:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 83938:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 83939:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 83940:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 83941:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 83942:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 83943:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 83944:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 83945:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 83946:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 83947:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 83948:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 83949:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 83950:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 83951:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 83952:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 83953:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 83954:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 83955:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 83956:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 83957:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 83958:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 83959:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 83960:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 83961:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 83962:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 83963:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 83964:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 83965:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 83966:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 83967:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 83968:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 83969:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 83970:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 83971:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 83972:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 83973:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 83974:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 83975:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 83976:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 83977:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 83978:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 83979:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 83980:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 83981:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 83982:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 83983:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 83984:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 83985:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 83986:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 83987:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 83988:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 83989:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 83990:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 83991:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 83992:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 83993:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 83994:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 83995:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 83996:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 83997:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 83998:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 83999:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 84000:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 84001:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 84002:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 84003:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 84004:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 84005:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 84006:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 84007:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 84008:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 84009:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 84010:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 84011:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 84012:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 84013:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 84014:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 84015:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 84016:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 84017:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 84018:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 84019:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 84020:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 84021:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 84022:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 84023:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 84024:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 84025:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 84026:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 84027:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 84028:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 84029:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 84030:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 84031:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 84032:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 84033:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 84034:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 84035:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 84036:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 84037:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 84038:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 84039:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 84040:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 84041:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 84042:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 84043:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 84044:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 84045:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 84046:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 84047:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 84048:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 84049:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 84050:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 84051:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 84052:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 84053:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 84054:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 84055:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 84056:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 84057:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 84058:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 84059:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 84060:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 84061:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 84062:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 84063:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 84064:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 84065:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 84066:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 84067:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 84068:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 84069:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 84070:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 84071:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 84072:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 84073:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 84074:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 84075:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 84076:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 84077:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 84078:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 84079:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 84080:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 84081:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 84082:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 84083:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 84084:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 84085:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 84086:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 84087:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 84088:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 84089:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 84090:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 84091:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 84092:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 84093:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 84094:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 84095:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 84096:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 84097:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 84098:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 84099:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 84100:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 84101:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 84102:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 84103:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 84104:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 84105:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 84106:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 84107:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 84108:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 84109:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 84110:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 84111:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 84112:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 84113:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 84114:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 84115:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 84116:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 84117:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 84118:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 84119:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 84120:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 84121:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 84122:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 84123:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 84124:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 84125:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 84126:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 84127:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 84128:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 84129:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 84130:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 84131:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 84132:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 84133:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 84134:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 84135:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 84136:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 84137:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 84138:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 84139:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 84140:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 84141:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 84142:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 84143:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 84144:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 84145:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 84146:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 84147:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 84148:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 84149:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 84150:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 84151:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 84152:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 84153:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 84154:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 84155:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 84156:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 84157:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 84158:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 84159:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 84160:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 84161:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 84162:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 84163:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 84164:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 84165:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 84166:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 84167:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 84168:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 84169:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 84170:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 84171:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 84172:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 84173:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 84174:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 84175:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 84176:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 84177:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 84178:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 84179:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 84180:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 84181:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 84182:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 84183:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 84184:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 84185:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 84186:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 84187:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 84188:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 84189:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 84190:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 84191:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 84192:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 84193:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 84194:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 84195:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 84196:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 84197:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 84198:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 84199:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 84200:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 84201:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 84202:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 84203:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 84204:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 84205:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 84206:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 84207:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 84208:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 84209:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 84210:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 84211:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 84212:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 84213:22]
  wire  invx137 = ~x137; // @[Snxn100k.scala 84214:17]
  wire  t138 = x137 + invx137; // @[Snxn100k.scala 84215:22]
  wire  inv138 = ~t138; // @[Snxn100k.scala 84216:17]
  wire  x138 = t138 ^ inv138; // @[Snxn100k.scala 84217:22]
  wire  invx138 = ~x138; // @[Snxn100k.scala 84218:17]
  wire  t139 = x138 + invx138; // @[Snxn100k.scala 84219:22]
  wire  inv139 = ~t139; // @[Snxn100k.scala 84220:17]
  wire  x139 = t139 ^ inv139; // @[Snxn100k.scala 84221:22]
  wire  invx139 = ~x139; // @[Snxn100k.scala 84222:17]
  wire  t140 = x139 + invx139; // @[Snxn100k.scala 84223:22]
  wire  inv140 = ~t140; // @[Snxn100k.scala 84224:17]
  wire  x140 = t140 ^ inv140; // @[Snxn100k.scala 84225:22]
  assign io_z = ~x140; // @[Snxn100k.scala 84226:17]
endmodule
module SnxnLv3Inst36(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst144_io_a; // @[Snxn100k.scala 25150:35]
  wire  inst_SnxnLv4Inst144_io_b; // @[Snxn100k.scala 25150:35]
  wire  inst_SnxnLv4Inst144_io_z; // @[Snxn100k.scala 25150:35]
  wire  inst_SnxnLv4Inst145_io_a; // @[Snxn100k.scala 25154:35]
  wire  inst_SnxnLv4Inst145_io_b; // @[Snxn100k.scala 25154:35]
  wire  inst_SnxnLv4Inst145_io_z; // @[Snxn100k.scala 25154:35]
  wire  inst_SnxnLv4Inst146_io_a; // @[Snxn100k.scala 25158:35]
  wire  inst_SnxnLv4Inst146_io_b; // @[Snxn100k.scala 25158:35]
  wire  inst_SnxnLv4Inst146_io_z; // @[Snxn100k.scala 25158:35]
  wire  inst_SnxnLv4Inst147_io_a; // @[Snxn100k.scala 25162:35]
  wire  inst_SnxnLv4Inst147_io_b; // @[Snxn100k.scala 25162:35]
  wire  inst_SnxnLv4Inst147_io_z; // @[Snxn100k.scala 25162:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst144_io_z + inst_SnxnLv4Inst145_io_z; // @[Snxn100k.scala 25166:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst146_io_z; // @[Snxn100k.scala 25166:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst147_io_z; // @[Snxn100k.scala 25166:92]
  SnxnLv4Inst5 inst_SnxnLv4Inst144 ( // @[Snxn100k.scala 25150:35]
    .io_a(inst_SnxnLv4Inst144_io_a),
    .io_b(inst_SnxnLv4Inst144_io_b),
    .io_z(inst_SnxnLv4Inst144_io_z)
  );
  SnxnLv4Inst90 inst_SnxnLv4Inst145 ( // @[Snxn100k.scala 25154:35]
    .io_a(inst_SnxnLv4Inst145_io_a),
    .io_b(inst_SnxnLv4Inst145_io_b),
    .io_z(inst_SnxnLv4Inst145_io_z)
  );
  SnxnLv4Inst146 inst_SnxnLv4Inst146 ( // @[Snxn100k.scala 25158:35]
    .io_a(inst_SnxnLv4Inst146_io_a),
    .io_b(inst_SnxnLv4Inst146_io_b),
    .io_z(inst_SnxnLv4Inst146_io_z)
  );
  SnxnLv4Inst147 inst_SnxnLv4Inst147 ( // @[Snxn100k.scala 25162:35]
    .io_a(inst_SnxnLv4Inst147_io_a),
    .io_b(inst_SnxnLv4Inst147_io_b),
    .io_z(inst_SnxnLv4Inst147_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25167:15]
  assign inst_SnxnLv4Inst144_io_a = io_a; // @[Snxn100k.scala 25151:28]
  assign inst_SnxnLv4Inst144_io_b = io_b; // @[Snxn100k.scala 25152:28]
  assign inst_SnxnLv4Inst145_io_a = io_a; // @[Snxn100k.scala 25155:28]
  assign inst_SnxnLv4Inst145_io_b = io_b; // @[Snxn100k.scala 25156:28]
  assign inst_SnxnLv4Inst146_io_a = io_a; // @[Snxn100k.scala 25159:28]
  assign inst_SnxnLv4Inst146_io_b = io_b; // @[Snxn100k.scala 25160:28]
  assign inst_SnxnLv4Inst147_io_a = io_a; // @[Snxn100k.scala 25163:28]
  assign inst_SnxnLv4Inst147_io_b = io_b; // @[Snxn100k.scala 25164:28]
endmodule
module SnxnLv4Inst151(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 86257:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 86258:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 86259:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 86260:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 86261:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 86262:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 86263:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 86264:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 86265:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 86266:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 86267:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 86268:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 86269:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 86270:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 86271:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 86272:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 86273:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 86274:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 86275:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 86276:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 86277:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 86278:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 86279:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 86280:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 86281:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 86282:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 86283:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 86284:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 86285:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 86286:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 86287:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 86288:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 86289:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 86290:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 86291:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 86292:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 86293:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 86294:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 86295:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 86296:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 86297:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 86298:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 86299:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 86300:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 86301:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 86302:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 86303:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 86304:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 86305:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 86306:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 86307:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 86308:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 86309:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 86310:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 86311:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 86312:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 86313:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 86314:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 86315:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 86316:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 86317:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 86318:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 86319:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 86320:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 86321:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 86322:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 86323:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 86324:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 86325:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 86326:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 86327:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 86328:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 86329:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 86330:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 86331:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 86332:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 86333:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 86334:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 86335:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 86336:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 86337:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 86338:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 86339:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 86340:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 86341:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 86342:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 86343:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 86344:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 86345:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 86346:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 86347:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 86348:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 86349:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 86350:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 86351:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 86352:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 86353:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 86354:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 86355:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 86356:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 86357:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 86358:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 86359:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 86360:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 86361:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 86362:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 86363:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 86364:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 86365:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 86366:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 86367:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 86368:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 86369:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 86370:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 86371:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 86372:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 86373:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 86374:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 86375:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 86376:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 86377:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 86378:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 86379:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 86380:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 86381:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 86382:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 86383:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 86384:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 86385:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 86386:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 86387:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 86388:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 86389:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 86390:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 86391:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 86392:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 86393:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 86394:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 86395:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 86396:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 86397:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 86398:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 86399:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 86400:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 86401:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 86402:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 86403:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 86404:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 86405:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 86406:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 86407:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 86408:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 86409:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 86410:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 86411:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 86412:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 86413:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 86414:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 86415:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 86416:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 86417:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 86418:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 86419:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 86420:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 86421:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 86422:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 86423:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 86424:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 86425:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 86426:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 86427:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 86428:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 86429:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 86430:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 86431:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 86432:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 86433:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 86434:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 86435:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 86436:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 86437:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 86438:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 86439:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 86440:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 86441:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 86442:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 86443:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 86444:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 86445:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 86446:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 86447:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 86448:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 86449:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 86450:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 86451:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 86452:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 86453:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 86454:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 86455:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 86456:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 86457:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 86458:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 86459:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 86460:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 86461:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 86462:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 86463:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 86464:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 86465:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 86466:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 86467:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 86468:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 86469:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 86470:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 86471:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 86472:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 86473:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 86474:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 86475:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 86476:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 86477:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 86478:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 86479:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 86480:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 86481:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 86482:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 86483:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 86484:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 86485:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 86486:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 86487:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 86488:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 86489:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 86490:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 86491:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 86492:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 86493:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 86494:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 86495:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 86496:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 86497:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 86498:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 86499:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 86500:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 86501:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 86502:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 86503:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 86504:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 86505:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 86506:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 86507:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 86508:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 86509:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 86510:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 86511:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 86512:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 86513:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 86514:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 86515:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 86516:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 86517:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 86518:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 86519:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 86520:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 86521:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 86522:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 86523:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 86524:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 86525:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 86526:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 86527:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 86528:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 86529:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 86530:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 86531:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 86532:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 86533:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 86534:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 86535:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 86536:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 86537:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 86538:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 86539:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 86540:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 86541:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 86542:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 86543:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 86544:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 86545:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 86546:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 86547:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 86548:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 86549:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 86550:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 86551:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 86552:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 86553:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 86554:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 86555:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 86556:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 86557:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 86558:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 86559:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 86560:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 86561:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 86562:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 86563:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 86564:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 86565:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 86566:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 86567:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 86568:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 86569:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 86570:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 86571:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 86572:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 86573:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 86574:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 86575:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 86576:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 86577:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 86578:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 86579:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 86580:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 86581:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 86582:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 86583:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 86584:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 86585:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 86586:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 86587:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 86588:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 86589:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 86590:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 86591:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 86592:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 86593:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 86594:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 86595:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 86596:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 86597:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 86598:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 86599:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 86600:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 86601:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 86602:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 86603:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 86604:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 86605:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 86606:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 86607:20]
  assign io_z = ~x87; // @[Snxn100k.scala 86608:16]
endmodule
module SnxnLv3Inst37(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst148_io_a; // @[Snxn100k.scala 25964:35]
  wire  inst_SnxnLv4Inst148_io_b; // @[Snxn100k.scala 25964:35]
  wire  inst_SnxnLv4Inst148_io_z; // @[Snxn100k.scala 25964:35]
  wire  inst_SnxnLv4Inst149_io_a; // @[Snxn100k.scala 25968:35]
  wire  inst_SnxnLv4Inst149_io_b; // @[Snxn100k.scala 25968:35]
  wire  inst_SnxnLv4Inst149_io_z; // @[Snxn100k.scala 25968:35]
  wire  inst_SnxnLv4Inst150_io_a; // @[Snxn100k.scala 25972:35]
  wire  inst_SnxnLv4Inst150_io_b; // @[Snxn100k.scala 25972:35]
  wire  inst_SnxnLv4Inst150_io_z; // @[Snxn100k.scala 25972:35]
  wire  inst_SnxnLv4Inst151_io_a; // @[Snxn100k.scala 25976:35]
  wire  inst_SnxnLv4Inst151_io_b; // @[Snxn100k.scala 25976:35]
  wire  inst_SnxnLv4Inst151_io_z; // @[Snxn100k.scala 25976:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst148_io_z + inst_SnxnLv4Inst149_io_z; // @[Snxn100k.scala 25980:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst150_io_z; // @[Snxn100k.scala 25980:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst151_io_z; // @[Snxn100k.scala 25980:92]
  SnxnLv4Inst49 inst_SnxnLv4Inst148 ( // @[Snxn100k.scala 25964:35]
    .io_a(inst_SnxnLv4Inst148_io_a),
    .io_b(inst_SnxnLv4Inst148_io_b),
    .io_z(inst_SnxnLv4Inst148_io_z)
  );
  SnxnLv4Inst2 inst_SnxnLv4Inst149 ( // @[Snxn100k.scala 25968:35]
    .io_a(inst_SnxnLv4Inst149_io_a),
    .io_b(inst_SnxnLv4Inst149_io_b),
    .io_z(inst_SnxnLv4Inst149_io_z)
  );
  SnxnLv4Inst41 inst_SnxnLv4Inst150 ( // @[Snxn100k.scala 25972:35]
    .io_a(inst_SnxnLv4Inst150_io_a),
    .io_b(inst_SnxnLv4Inst150_io_b),
    .io_z(inst_SnxnLv4Inst150_io_z)
  );
  SnxnLv4Inst151 inst_SnxnLv4Inst151 ( // @[Snxn100k.scala 25976:35]
    .io_a(inst_SnxnLv4Inst151_io_a),
    .io_b(inst_SnxnLv4Inst151_io_b),
    .io_z(inst_SnxnLv4Inst151_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25981:15]
  assign inst_SnxnLv4Inst148_io_a = io_a; // @[Snxn100k.scala 25965:28]
  assign inst_SnxnLv4Inst148_io_b = io_b; // @[Snxn100k.scala 25966:28]
  assign inst_SnxnLv4Inst149_io_a = io_a; // @[Snxn100k.scala 25969:28]
  assign inst_SnxnLv4Inst149_io_b = io_b; // @[Snxn100k.scala 25970:28]
  assign inst_SnxnLv4Inst150_io_a = io_a; // @[Snxn100k.scala 25973:28]
  assign inst_SnxnLv4Inst150_io_b = io_b; // @[Snxn100k.scala 25974:28]
  assign inst_SnxnLv4Inst151_io_a = io_a; // @[Snxn100k.scala 25977:28]
  assign inst_SnxnLv4Inst151_io_b = io_b; // @[Snxn100k.scala 25978:28]
endmodule
module SnxnLv4Inst152(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 87841:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 87842:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 87843:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 87844:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 87845:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 87846:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 87847:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 87848:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 87849:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 87850:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 87851:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 87852:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 87853:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 87854:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 87855:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 87856:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 87857:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 87858:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 87859:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 87860:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 87861:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 87862:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 87863:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 87864:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 87865:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 87866:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 87867:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 87868:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 87869:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 87870:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 87871:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 87872:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 87873:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 87874:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 87875:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 87876:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 87877:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 87878:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 87879:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 87880:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 87881:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 87882:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 87883:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 87884:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 87885:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 87886:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 87887:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 87888:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 87889:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 87890:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 87891:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 87892:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 87893:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 87894:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 87895:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 87896:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 87897:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 87898:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 87899:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 87900:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 87901:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 87902:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 87903:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 87904:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 87905:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 87906:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 87907:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 87908:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 87909:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 87910:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 87911:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 87912:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 87913:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 87914:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 87915:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 87916:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 87917:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 87918:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 87919:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 87920:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 87921:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 87922:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 87923:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 87924:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 87925:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 87926:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 87927:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 87928:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 87929:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 87930:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 87931:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 87932:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 87933:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 87934:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 87935:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 87936:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 87937:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 87938:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 87939:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 87940:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 87941:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 87942:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 87943:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 87944:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 87945:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 87946:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 87947:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 87948:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 87949:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 87950:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 87951:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 87952:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 87953:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 87954:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 87955:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 87956:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 87957:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 87958:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 87959:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 87960:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 87961:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 87962:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 87963:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 87964:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 87965:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 87966:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 87967:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 87968:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 87969:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 87970:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 87971:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 87972:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 87973:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 87974:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 87975:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 87976:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 87977:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 87978:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 87979:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 87980:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 87981:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 87982:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 87983:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 87984:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 87985:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 87986:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 87987:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 87988:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 87989:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 87990:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 87991:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 87992:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 87993:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 87994:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 87995:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 87996:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 87997:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 87998:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 87999:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 88000:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 88001:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 88002:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 88003:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 88004:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 88005:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 88006:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 88007:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 88008:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 88009:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 88010:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 88011:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 88012:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 88013:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 88014:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 88015:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 88016:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 88017:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 88018:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 88019:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 88020:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 88021:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 88022:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 88023:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 88024:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 88025:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 88026:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 88027:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 88028:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 88029:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 88030:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 88031:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 88032:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 88033:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 88034:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 88035:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 88036:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 88037:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 88038:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 88039:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 88040:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 88041:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 88042:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 88043:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 88044:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 88045:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 88046:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 88047:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 88048:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 88049:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 88050:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 88051:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 88052:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 88053:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 88054:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 88055:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 88056:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 88057:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 88058:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 88059:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 88060:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 88061:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 88062:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 88063:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 88064:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 88065:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 88066:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 88067:20]
  assign io_z = ~x56; // @[Snxn100k.scala 88068:16]
endmodule
module SnxnLv4Inst154(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 88141:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 88142:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 88143:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 88144:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 88145:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 88146:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 88147:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 88148:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 88149:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 88150:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 88151:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 88152:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 88153:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 88154:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 88155:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 88156:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 88157:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 88158:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 88159:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 88160:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 88161:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 88162:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 88163:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 88164:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 88165:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 88166:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 88167:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 88168:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 88169:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 88170:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 88171:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 88172:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 88173:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 88174:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 88175:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 88176:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 88177:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 88178:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 88179:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 88180:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 88181:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 88182:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 88183:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 88184:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 88185:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 88186:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 88187:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 88188:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 88189:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 88190:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 88191:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 88192:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 88193:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 88194:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 88195:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 88196:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 88197:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 88198:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 88199:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 88200:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 88201:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 88202:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 88203:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 88204:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 88205:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 88206:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 88207:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 88208:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 88209:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 88210:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 88211:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 88212:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 88213:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 88214:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 88215:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 88216:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 88217:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 88218:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 88219:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 88220:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 88221:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 88222:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 88223:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 88224:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 88225:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 88226:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 88227:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 88228:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 88229:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 88230:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 88231:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 88232:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 88233:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 88234:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 88235:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 88236:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 88237:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 88238:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 88239:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 88240:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 88241:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 88242:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 88243:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 88244:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 88245:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 88246:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 88247:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 88248:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 88249:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 88250:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 88251:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 88252:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 88253:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 88254:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 88255:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 88256:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 88257:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 88258:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 88259:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 88260:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 88261:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 88262:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 88263:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 88264:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 88265:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 88266:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 88267:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 88268:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 88269:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 88270:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 88271:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 88272:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 88273:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 88274:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 88275:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 88276:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 88277:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 88278:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 88279:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 88280:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 88281:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 88282:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 88283:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 88284:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 88285:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 88286:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 88287:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 88288:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 88289:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 88290:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 88291:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 88292:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 88293:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 88294:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 88295:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 88296:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 88297:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 88298:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 88299:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 88300:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 88301:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 88302:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 88303:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 88304:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 88305:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 88306:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 88307:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 88308:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 88309:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 88310:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 88311:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 88312:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 88313:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 88314:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 88315:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 88316:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 88317:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 88318:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 88319:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 88320:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 88321:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 88322:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 88323:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 88324:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 88325:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 88326:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 88327:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 88328:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 88329:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 88330:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 88331:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 88332:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 88333:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 88334:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 88335:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 88336:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 88337:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 88338:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 88339:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 88340:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 88341:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 88342:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 88343:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 88344:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 88345:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 88346:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 88347:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 88348:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 88349:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 88350:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 88351:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 88352:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 88353:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 88354:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 88355:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 88356:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 88357:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 88358:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 88359:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 88360:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 88361:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 88362:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 88363:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 88364:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 88365:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 88366:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 88367:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 88368:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 88369:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 88370:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 88371:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 88372:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 88373:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 88374:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 88375:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 88376:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 88377:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 88378:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 88379:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 88380:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 88381:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 88382:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 88383:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 88384:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 88385:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 88386:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 88387:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 88388:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 88389:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 88390:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 88391:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 88392:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 88393:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 88394:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 88395:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 88396:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 88397:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 88398:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 88399:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 88400:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 88401:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 88402:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 88403:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 88404:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 88405:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 88406:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 88407:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 88408:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 88409:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 88410:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 88411:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 88412:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 88413:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 88414:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 88415:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 88416:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 88417:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 88418:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 88419:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 88420:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 88421:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 88422:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 88423:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 88424:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 88425:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 88426:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 88427:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 88428:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 88429:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 88430:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 88431:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 88432:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 88433:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 88434:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 88435:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 88436:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 88437:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 88438:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 88439:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 88440:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 88441:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 88442:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 88443:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 88444:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 88445:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 88446:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 88447:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 88448:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 88449:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 88450:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 88451:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 88452:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 88453:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 88454:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 88455:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 88456:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 88457:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 88458:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 88459:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 88460:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 88461:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 88462:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 88463:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 88464:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 88465:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 88466:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 88467:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 88468:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 88469:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 88470:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 88471:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 88472:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 88473:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 88474:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 88475:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 88476:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 88477:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 88478:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 88479:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 88480:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 88481:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 88482:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 88483:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 88484:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 88485:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 88486:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 88487:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 88488:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 88489:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 88490:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 88491:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 88492:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 88493:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 88494:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 88495:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 88496:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 88497:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 88498:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 88499:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 88500:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 88501:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 88502:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 88503:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 88504:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 88505:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 88506:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 88507:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 88508:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 88509:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 88510:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 88511:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 88512:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 88513:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 88514:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 88515:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 88516:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 88517:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 88518:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 88519:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 88520:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 88521:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 88522:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 88523:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 88524:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 88525:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 88526:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 88527:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 88528:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 88529:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 88530:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 88531:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 88532:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 88533:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 88534:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 88535:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 88536:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 88537:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 88538:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 88539:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 88540:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 88541:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 88542:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 88543:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 88544:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 88545:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 88546:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 88547:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 88548:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 88549:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 88550:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 88551:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 88552:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 88553:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 88554:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 88555:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 88556:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 88557:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 88558:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 88559:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 88560:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 88561:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 88562:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 88563:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 88564:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 88565:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 88566:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 88567:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 88568:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 88569:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 88570:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 88571:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 88572:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 88573:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 88574:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 88575:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 88576:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 88577:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 88578:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 88579:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 88580:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 88581:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 88582:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 88583:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 88584:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 88585:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 88586:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 88587:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 88588:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 88589:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 88590:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 88591:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 88592:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 88593:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 88594:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 88595:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 88596:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 88597:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 88598:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 88599:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 88600:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 88601:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 88602:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 88603:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 88604:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 88605:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 88606:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 88607:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 88608:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 88609:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 88610:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 88611:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 88612:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 88613:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 88614:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 88615:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 88616:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 88617:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 88618:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 88619:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 88620:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 88621:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 88622:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 88623:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 88624:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 88625:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 88626:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 88627:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 88628:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 88629:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 88630:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 88631:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 88632:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 88633:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 88634:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 88635:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 88636:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 88637:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 88638:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 88639:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 88640:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 88641:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 88642:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 88643:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 88644:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 88645:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 88646:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 88647:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 88648:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 88649:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 88650:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 88651:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 88652:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 88653:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 88654:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 88655:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 88656:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 88657:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 88658:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 88659:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 88660:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 88661:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 88662:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 88663:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 88664:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 88665:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 88666:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 88667:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 88668:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 88669:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 88670:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 88671:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 88672:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 88673:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 88674:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 88675:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 88676:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 88677:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 88678:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 88679:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 88680:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 88681:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 88682:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 88683:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 88684:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 88685:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 88686:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 88687:22]
  wire  invx136 = ~x136; // @[Snxn100k.scala 88688:17]
  wire  t137 = x136 + invx136; // @[Snxn100k.scala 88689:22]
  wire  inv137 = ~t137; // @[Snxn100k.scala 88690:17]
  wire  x137 = t137 ^ inv137; // @[Snxn100k.scala 88691:22]
  assign io_z = ~x137; // @[Snxn100k.scala 88692:17]
endmodule
module SnxnLv3Inst38(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst152_io_a; // @[Snxn100k.scala 26071:35]
  wire  inst_SnxnLv4Inst152_io_b; // @[Snxn100k.scala 26071:35]
  wire  inst_SnxnLv4Inst152_io_z; // @[Snxn100k.scala 26071:35]
  wire  inst_SnxnLv4Inst153_io_a; // @[Snxn100k.scala 26075:35]
  wire  inst_SnxnLv4Inst153_io_b; // @[Snxn100k.scala 26075:35]
  wire  inst_SnxnLv4Inst153_io_z; // @[Snxn100k.scala 26075:35]
  wire  inst_SnxnLv4Inst154_io_a; // @[Snxn100k.scala 26079:35]
  wire  inst_SnxnLv4Inst154_io_b; // @[Snxn100k.scala 26079:35]
  wire  inst_SnxnLv4Inst154_io_z; // @[Snxn100k.scala 26079:35]
  wire  inst_SnxnLv4Inst155_io_a; // @[Snxn100k.scala 26083:35]
  wire  inst_SnxnLv4Inst155_io_b; // @[Snxn100k.scala 26083:35]
  wire  inst_SnxnLv4Inst155_io_z; // @[Snxn100k.scala 26083:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst152_io_z + inst_SnxnLv4Inst153_io_z; // @[Snxn100k.scala 26087:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst154_io_z; // @[Snxn100k.scala 26087:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst155_io_z; // @[Snxn100k.scala 26087:92]
  SnxnLv4Inst152 inst_SnxnLv4Inst152 ( // @[Snxn100k.scala 26071:35]
    .io_a(inst_SnxnLv4Inst152_io_a),
    .io_b(inst_SnxnLv4Inst152_io_b),
    .io_z(inst_SnxnLv4Inst152_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst153 ( // @[Snxn100k.scala 26075:35]
    .io_a(inst_SnxnLv4Inst153_io_a),
    .io_b(inst_SnxnLv4Inst153_io_b),
    .io_z(inst_SnxnLv4Inst153_io_z)
  );
  SnxnLv4Inst154 inst_SnxnLv4Inst154 ( // @[Snxn100k.scala 26079:35]
    .io_a(inst_SnxnLv4Inst154_io_a),
    .io_b(inst_SnxnLv4Inst154_io_b),
    .io_z(inst_SnxnLv4Inst154_io_z)
  );
  SnxnLv4Inst42 inst_SnxnLv4Inst155 ( // @[Snxn100k.scala 26083:35]
    .io_a(inst_SnxnLv4Inst155_io_a),
    .io_b(inst_SnxnLv4Inst155_io_b),
    .io_z(inst_SnxnLv4Inst155_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26088:15]
  assign inst_SnxnLv4Inst152_io_a = io_a; // @[Snxn100k.scala 26072:28]
  assign inst_SnxnLv4Inst152_io_b = io_b; // @[Snxn100k.scala 26073:28]
  assign inst_SnxnLv4Inst153_io_a = io_a; // @[Snxn100k.scala 26076:28]
  assign inst_SnxnLv4Inst153_io_b = io_b; // @[Snxn100k.scala 26077:28]
  assign inst_SnxnLv4Inst154_io_a = io_a; // @[Snxn100k.scala 26080:28]
  assign inst_SnxnLv4Inst154_io_b = io_b; // @[Snxn100k.scala 26081:28]
  assign inst_SnxnLv4Inst155_io_a = io_a; // @[Snxn100k.scala 26084:28]
  assign inst_SnxnLv4Inst155_io_b = io_b; // @[Snxn100k.scala 26085:28]
endmodule
module SnxnLv4Inst156(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 85497:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 85498:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 85499:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 85500:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 85501:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 85502:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 85503:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 85504:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 85505:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 85506:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 85507:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 85508:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 85509:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 85510:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 85511:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 85512:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 85513:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 85514:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 85515:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 85516:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 85517:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 85518:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 85519:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 85520:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 85521:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 85522:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 85523:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 85524:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 85525:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 85526:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 85527:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 85528:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 85529:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 85530:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 85531:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 85532:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 85533:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 85534:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 85535:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 85536:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 85537:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 85538:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 85539:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 85540:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 85541:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 85542:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 85543:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 85544:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 85545:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 85546:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 85547:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 85548:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 85549:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 85550:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 85551:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 85552:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 85553:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 85554:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 85555:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 85556:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 85557:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 85558:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 85559:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 85560:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 85561:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 85562:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 85563:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 85564:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 85565:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 85566:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 85567:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 85568:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 85569:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 85570:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 85571:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 85572:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 85573:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 85574:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 85575:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 85576:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 85577:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 85578:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 85579:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 85580:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 85581:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 85582:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 85583:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 85584:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 85585:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 85586:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 85587:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 85588:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 85589:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 85590:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 85591:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 85592:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 85593:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 85594:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 85595:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 85596:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 85597:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 85598:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 85599:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 85600:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 85601:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 85602:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 85603:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 85604:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 85605:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 85606:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 85607:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 85608:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 85609:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 85610:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 85611:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 85612:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 85613:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 85614:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 85615:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 85616:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 85617:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 85618:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 85619:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 85620:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 85621:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 85622:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 85623:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 85624:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 85625:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 85626:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 85627:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 85628:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 85629:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 85630:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 85631:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 85632:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 85633:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 85634:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 85635:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 85636:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 85637:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 85638:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 85639:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 85640:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 85641:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 85642:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 85643:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 85644:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 85645:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 85646:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 85647:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 85648:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 85649:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 85650:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 85651:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 85652:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 85653:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 85654:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 85655:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 85656:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 85657:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 85658:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 85659:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 85660:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 85661:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 85662:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 85663:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 85664:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 85665:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 85666:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 85667:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 85668:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 85669:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 85670:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 85671:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 85672:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 85673:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 85674:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 85675:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 85676:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 85677:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 85678:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 85679:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 85680:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 85681:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 85682:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 85683:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 85684:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 85685:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 85686:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 85687:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 85688:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 85689:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 85690:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 85691:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 85692:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 85693:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 85694:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 85695:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 85696:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 85697:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 85698:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 85699:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 85700:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 85701:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 85702:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 85703:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 85704:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 85705:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 85706:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 85707:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 85708:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 85709:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 85710:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 85711:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 85712:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 85713:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 85714:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 85715:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 85716:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 85717:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 85718:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 85719:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 85720:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 85721:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 85722:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 85723:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 85724:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 85725:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 85726:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 85727:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 85728:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 85729:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 85730:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 85731:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 85732:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 85733:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 85734:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 85735:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 85736:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 85737:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 85738:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 85739:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 85740:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 85741:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 85742:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 85743:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 85744:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 85745:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 85746:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 85747:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 85748:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 85749:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 85750:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 85751:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 85752:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 85753:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 85754:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 85755:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 85756:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 85757:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 85758:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 85759:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 85760:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 85761:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 85762:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 85763:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 85764:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 85765:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 85766:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 85767:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 85768:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 85769:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 85770:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 85771:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 85772:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 85773:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 85774:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 85775:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 85776:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 85777:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 85778:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 85779:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 85780:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 85781:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 85782:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 85783:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 85784:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 85785:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 85786:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 85787:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 85788:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 85789:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 85790:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 85791:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 85792:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 85793:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 85794:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 85795:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 85796:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 85797:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 85798:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 85799:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 85800:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 85801:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 85802:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 85803:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 85804:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 85805:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 85806:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 85807:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 85808:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 85809:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 85810:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 85811:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 85812:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 85813:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 85814:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 85815:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 85816:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 85817:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 85818:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 85819:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 85820:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 85821:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 85822:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 85823:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 85824:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 85825:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 85826:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 85827:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 85828:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 85829:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 85830:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 85831:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 85832:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 85833:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 85834:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 85835:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 85836:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 85837:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 85838:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 85839:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 85840:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 85841:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 85842:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 85843:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 85844:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 85845:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 85846:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 85847:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 85848:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 85849:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 85850:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 85851:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 85852:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 85853:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 85854:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 85855:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 85856:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 85857:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 85858:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 85859:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 85860:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 85861:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 85862:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 85863:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 85864:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 85865:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 85866:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 85867:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 85868:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 85869:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 85870:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 85871:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 85872:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 85873:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 85874:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 85875:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 85876:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 85877:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 85878:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 85879:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 85880:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 85881:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 85882:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 85883:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 85884:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 85885:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 85886:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 85887:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 85888:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 85889:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 85890:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 85891:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 85892:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 85893:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 85894:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 85895:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 85896:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 85897:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 85898:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 85899:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 85900:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 85901:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 85902:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 85903:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 85904:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 85905:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 85906:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 85907:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 85908:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 85909:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 85910:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 85911:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 85912:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 85913:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 85914:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 85915:22]
  assign io_z = ~x104; // @[Snxn100k.scala 85916:17]
endmodule
module SnxnLv4Inst158(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 84823:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 84824:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 84825:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 84826:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 84827:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 84828:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 84829:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 84830:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 84831:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 84832:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 84833:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 84834:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 84835:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 84836:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 84837:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 84838:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 84839:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 84840:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 84841:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 84842:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 84843:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 84844:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 84845:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 84846:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 84847:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 84848:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 84849:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 84850:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 84851:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 84852:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 84853:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 84854:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 84855:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 84856:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 84857:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 84858:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 84859:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 84860:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 84861:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 84862:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 84863:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 84864:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 84865:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 84866:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 84867:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 84868:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 84869:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 84870:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 84871:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 84872:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 84873:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 84874:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 84875:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 84876:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 84877:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 84878:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 84879:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 84880:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 84881:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 84882:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 84883:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 84884:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 84885:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 84886:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 84887:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 84888:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 84889:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 84890:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 84891:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 84892:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 84893:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 84894:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 84895:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 84896:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 84897:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 84898:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 84899:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 84900:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 84901:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 84902:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 84903:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 84904:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 84905:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 84906:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 84907:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 84908:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 84909:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 84910:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 84911:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 84912:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 84913:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 84914:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 84915:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 84916:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 84917:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 84918:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 84919:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 84920:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 84921:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 84922:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 84923:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 84924:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 84925:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 84926:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 84927:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 84928:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 84929:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 84930:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 84931:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 84932:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 84933:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 84934:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 84935:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 84936:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 84937:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 84938:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 84939:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 84940:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 84941:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 84942:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 84943:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 84944:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 84945:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 84946:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 84947:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 84948:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 84949:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 84950:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 84951:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 84952:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 84953:20]
  assign io_z = ~x32; // @[Snxn100k.scala 84954:16]
endmodule
module SnxnLv4Inst159(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 84965:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 84966:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 84967:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 84968:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 84969:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 84970:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 84971:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 84972:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 84973:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 84974:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 84975:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 84976:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 84977:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 84978:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 84979:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 84980:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 84981:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 84982:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 84983:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 84984:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 84985:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 84986:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 84987:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 84988:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 84989:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 84990:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 84991:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 84992:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 84993:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 84994:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 84995:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 84996:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 84997:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 84998:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 84999:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 85000:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 85001:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 85002:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 85003:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 85004:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 85005:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 85006:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 85007:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 85008:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 85009:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 85010:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 85011:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 85012:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 85013:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 85014:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 85015:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 85016:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 85017:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 85018:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 85019:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 85020:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 85021:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 85022:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 85023:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 85024:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 85025:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 85026:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 85027:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 85028:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 85029:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 85030:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 85031:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 85032:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 85033:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 85034:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 85035:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 85036:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 85037:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 85038:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 85039:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 85040:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 85041:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 85042:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 85043:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 85044:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 85045:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 85046:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 85047:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 85048:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 85049:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 85050:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 85051:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 85052:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 85053:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 85054:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 85055:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 85056:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 85057:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 85058:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 85059:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 85060:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 85061:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 85062:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 85063:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 85064:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 85065:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 85066:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 85067:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 85068:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 85069:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 85070:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 85071:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 85072:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 85073:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 85074:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 85075:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 85076:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 85077:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 85078:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 85079:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 85080:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 85081:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 85082:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 85083:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 85084:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 85085:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 85086:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 85087:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 85088:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 85089:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 85090:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 85091:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 85092:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 85093:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 85094:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 85095:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 85096:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 85097:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 85098:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 85099:20]
  assign io_z = ~x33; // @[Snxn100k.scala 85100:16]
endmodule
module SnxnLv3Inst39(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst156_io_a; // @[Snxn100k.scala 25481:35]
  wire  inst_SnxnLv4Inst156_io_b; // @[Snxn100k.scala 25481:35]
  wire  inst_SnxnLv4Inst156_io_z; // @[Snxn100k.scala 25481:35]
  wire  inst_SnxnLv4Inst157_io_a; // @[Snxn100k.scala 25485:35]
  wire  inst_SnxnLv4Inst157_io_b; // @[Snxn100k.scala 25485:35]
  wire  inst_SnxnLv4Inst157_io_z; // @[Snxn100k.scala 25485:35]
  wire  inst_SnxnLv4Inst158_io_a; // @[Snxn100k.scala 25489:35]
  wire  inst_SnxnLv4Inst158_io_b; // @[Snxn100k.scala 25489:35]
  wire  inst_SnxnLv4Inst158_io_z; // @[Snxn100k.scala 25489:35]
  wire  inst_SnxnLv4Inst159_io_a; // @[Snxn100k.scala 25493:35]
  wire  inst_SnxnLv4Inst159_io_b; // @[Snxn100k.scala 25493:35]
  wire  inst_SnxnLv4Inst159_io_z; // @[Snxn100k.scala 25493:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst156_io_z + inst_SnxnLv4Inst157_io_z; // @[Snxn100k.scala 25497:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst158_io_z; // @[Snxn100k.scala 25497:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst159_io_z; // @[Snxn100k.scala 25497:92]
  SnxnLv4Inst156 inst_SnxnLv4Inst156 ( // @[Snxn100k.scala 25481:35]
    .io_a(inst_SnxnLv4Inst156_io_a),
    .io_b(inst_SnxnLv4Inst156_io_b),
    .io_z(inst_SnxnLv4Inst156_io_z)
  );
  SnxnLv4Inst93 inst_SnxnLv4Inst157 ( // @[Snxn100k.scala 25485:35]
    .io_a(inst_SnxnLv4Inst157_io_a),
    .io_b(inst_SnxnLv4Inst157_io_b),
    .io_z(inst_SnxnLv4Inst157_io_z)
  );
  SnxnLv4Inst158 inst_SnxnLv4Inst158 ( // @[Snxn100k.scala 25489:35]
    .io_a(inst_SnxnLv4Inst158_io_a),
    .io_b(inst_SnxnLv4Inst158_io_b),
    .io_z(inst_SnxnLv4Inst158_io_z)
  );
  SnxnLv4Inst159 inst_SnxnLv4Inst159 ( // @[Snxn100k.scala 25493:35]
    .io_a(inst_SnxnLv4Inst159_io_a),
    .io_b(inst_SnxnLv4Inst159_io_b),
    .io_z(inst_SnxnLv4Inst159_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 25498:15]
  assign inst_SnxnLv4Inst156_io_a = io_a; // @[Snxn100k.scala 25482:28]
  assign inst_SnxnLv4Inst156_io_b = io_b; // @[Snxn100k.scala 25483:28]
  assign inst_SnxnLv4Inst157_io_a = io_a; // @[Snxn100k.scala 25486:28]
  assign inst_SnxnLv4Inst157_io_b = io_b; // @[Snxn100k.scala 25487:28]
  assign inst_SnxnLv4Inst158_io_a = io_a; // @[Snxn100k.scala 25490:28]
  assign inst_SnxnLv4Inst158_io_b = io_b; // @[Snxn100k.scala 25491:28]
  assign inst_SnxnLv4Inst159_io_a = io_a; // @[Snxn100k.scala 25494:28]
  assign inst_SnxnLv4Inst159_io_b = io_b; // @[Snxn100k.scala 25495:28]
endmodule
module SnxnLv2Inst9(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst36_io_a; // @[Snxn100k.scala 7452:34]
  wire  inst_SnxnLv3Inst36_io_b; // @[Snxn100k.scala 7452:34]
  wire  inst_SnxnLv3Inst36_io_z; // @[Snxn100k.scala 7452:34]
  wire  inst_SnxnLv3Inst37_io_a; // @[Snxn100k.scala 7456:34]
  wire  inst_SnxnLv3Inst37_io_b; // @[Snxn100k.scala 7456:34]
  wire  inst_SnxnLv3Inst37_io_z; // @[Snxn100k.scala 7456:34]
  wire  inst_SnxnLv3Inst38_io_a; // @[Snxn100k.scala 7460:34]
  wire  inst_SnxnLv3Inst38_io_b; // @[Snxn100k.scala 7460:34]
  wire  inst_SnxnLv3Inst38_io_z; // @[Snxn100k.scala 7460:34]
  wire  inst_SnxnLv3Inst39_io_a; // @[Snxn100k.scala 7464:34]
  wire  inst_SnxnLv3Inst39_io_b; // @[Snxn100k.scala 7464:34]
  wire  inst_SnxnLv3Inst39_io_z; // @[Snxn100k.scala 7464:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst36_io_z + inst_SnxnLv3Inst37_io_z; // @[Snxn100k.scala 7468:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst38_io_z; // @[Snxn100k.scala 7468:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst39_io_z; // @[Snxn100k.scala 7468:89]
  SnxnLv3Inst36 inst_SnxnLv3Inst36 ( // @[Snxn100k.scala 7452:34]
    .io_a(inst_SnxnLv3Inst36_io_a),
    .io_b(inst_SnxnLv3Inst36_io_b),
    .io_z(inst_SnxnLv3Inst36_io_z)
  );
  SnxnLv3Inst37 inst_SnxnLv3Inst37 ( // @[Snxn100k.scala 7456:34]
    .io_a(inst_SnxnLv3Inst37_io_a),
    .io_b(inst_SnxnLv3Inst37_io_b),
    .io_z(inst_SnxnLv3Inst37_io_z)
  );
  SnxnLv3Inst38 inst_SnxnLv3Inst38 ( // @[Snxn100k.scala 7460:34]
    .io_a(inst_SnxnLv3Inst38_io_a),
    .io_b(inst_SnxnLv3Inst38_io_b),
    .io_z(inst_SnxnLv3Inst38_io_z)
  );
  SnxnLv3Inst39 inst_SnxnLv3Inst39 ( // @[Snxn100k.scala 7464:34]
    .io_a(inst_SnxnLv3Inst39_io_a),
    .io_b(inst_SnxnLv3Inst39_io_b),
    .io_z(inst_SnxnLv3Inst39_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7469:15]
  assign inst_SnxnLv3Inst36_io_a = io_a; // @[Snxn100k.scala 7453:27]
  assign inst_SnxnLv3Inst36_io_b = io_b; // @[Snxn100k.scala 7454:27]
  assign inst_SnxnLv3Inst37_io_a = io_a; // @[Snxn100k.scala 7457:27]
  assign inst_SnxnLv3Inst37_io_b = io_b; // @[Snxn100k.scala 7458:27]
  assign inst_SnxnLv3Inst38_io_a = io_a; // @[Snxn100k.scala 7461:27]
  assign inst_SnxnLv3Inst38_io_b = io_b; // @[Snxn100k.scala 7462:27]
  assign inst_SnxnLv3Inst39_io_a = io_a; // @[Snxn100k.scala 7465:27]
  assign inst_SnxnLv3Inst39_io_b = io_b; // @[Snxn100k.scala 7466:27]
endmodule
module SnxnLv4Inst162(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 90951:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 90952:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 90953:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 90954:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 90955:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 90956:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 90957:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 90958:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 90959:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 90960:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 90961:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 90962:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 90963:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 90964:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 90965:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 90966:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 90967:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 90968:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 90969:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 90970:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 90971:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 90972:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 90973:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 90974:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 90975:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 90976:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 90977:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 90978:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 90979:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 90980:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 90981:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 90982:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 90983:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 90984:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 90985:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 90986:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 90987:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 90988:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 90989:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 90990:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 90991:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 90992:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 90993:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 90994:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 90995:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 90996:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 90997:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 90998:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 90999:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 91000:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 91001:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 91002:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 91003:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 91004:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 91005:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 91006:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 91007:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 91008:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 91009:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 91010:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 91011:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 91012:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 91013:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 91014:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 91015:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 91016:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 91017:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 91018:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 91019:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 91020:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 91021:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 91022:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 91023:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 91024:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 91025:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 91026:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 91027:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 91028:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 91029:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 91030:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 91031:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 91032:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 91033:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 91034:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 91035:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 91036:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 91037:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 91038:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 91039:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 91040:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 91041:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 91042:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 91043:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 91044:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 91045:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 91046:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 91047:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 91048:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 91049:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 91050:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 91051:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 91052:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 91053:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 91054:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 91055:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 91056:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 91057:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 91058:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 91059:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 91060:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 91061:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 91062:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 91063:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 91064:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 91065:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 91066:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 91067:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 91068:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 91069:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 91070:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 91071:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 91072:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 91073:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 91074:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 91075:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 91076:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 91077:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 91078:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 91079:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 91080:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 91081:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 91082:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 91083:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 91084:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 91085:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 91086:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 91087:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 91088:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 91089:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 91090:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 91091:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 91092:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 91093:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 91094:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 91095:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 91096:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 91097:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 91098:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 91099:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 91100:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 91101:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 91102:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 91103:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 91104:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 91105:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 91106:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 91107:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 91108:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 91109:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 91110:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 91111:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 91112:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 91113:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 91114:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 91115:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 91116:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 91117:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 91118:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 91119:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 91120:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 91121:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 91122:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 91123:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 91124:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 91125:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 91126:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 91127:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 91128:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 91129:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 91130:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 91131:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 91132:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 91133:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 91134:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 91135:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 91136:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 91137:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 91138:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 91139:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 91140:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 91141:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 91142:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 91143:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 91144:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 91145:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 91146:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 91147:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 91148:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 91149:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 91150:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 91151:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 91152:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 91153:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 91154:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 91155:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 91156:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 91157:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 91158:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 91159:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 91160:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 91161:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 91162:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 91163:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 91164:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 91165:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 91166:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 91167:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 91168:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 91169:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 91170:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 91171:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 91172:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 91173:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 91174:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 91175:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 91176:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 91177:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 91178:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 91179:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 91180:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 91181:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 91182:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 91183:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 91184:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 91185:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 91186:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 91187:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 91188:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 91189:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 91190:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 91191:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 91192:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 91193:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 91194:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 91195:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 91196:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 91197:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 91198:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 91199:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 91200:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 91201:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 91202:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 91203:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 91204:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 91205:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 91206:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 91207:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 91208:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 91209:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 91210:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 91211:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 91212:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 91213:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 91214:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 91215:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 91216:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 91217:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 91218:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 91219:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 91220:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 91221:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 91222:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 91223:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 91224:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 91225:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 91226:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 91227:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 91228:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 91229:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 91230:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 91231:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 91232:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 91233:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 91234:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 91235:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 91236:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 91237:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 91238:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 91239:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 91240:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 91241:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 91242:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 91243:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 91244:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 91245:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 91246:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 91247:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 91248:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 91249:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 91250:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 91251:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 91252:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 91253:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 91254:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 91255:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 91256:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 91257:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 91258:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 91259:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 91260:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 91261:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 91262:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 91263:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 91264:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 91265:20]
  assign io_z = ~x78; // @[Snxn100k.scala 91266:16]
endmodule
module SnxnLv3Inst40(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst160_io_a; // @[Snxn100k.scala 26996:35]
  wire  inst_SnxnLv4Inst160_io_b; // @[Snxn100k.scala 26996:35]
  wire  inst_SnxnLv4Inst160_io_z; // @[Snxn100k.scala 26996:35]
  wire  inst_SnxnLv4Inst161_io_a; // @[Snxn100k.scala 27000:35]
  wire  inst_SnxnLv4Inst161_io_b; // @[Snxn100k.scala 27000:35]
  wire  inst_SnxnLv4Inst161_io_z; // @[Snxn100k.scala 27000:35]
  wire  inst_SnxnLv4Inst162_io_a; // @[Snxn100k.scala 27004:35]
  wire  inst_SnxnLv4Inst162_io_b; // @[Snxn100k.scala 27004:35]
  wire  inst_SnxnLv4Inst162_io_z; // @[Snxn100k.scala 27004:35]
  wire  inst_SnxnLv4Inst163_io_a; // @[Snxn100k.scala 27008:35]
  wire  inst_SnxnLv4Inst163_io_b; // @[Snxn100k.scala 27008:35]
  wire  inst_SnxnLv4Inst163_io_z; // @[Snxn100k.scala 27008:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst160_io_z + inst_SnxnLv4Inst161_io_z; // @[Snxn100k.scala 27012:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst162_io_z; // @[Snxn100k.scala 27012:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst163_io_z; // @[Snxn100k.scala 27012:92]
  SnxnLv4Inst86 inst_SnxnLv4Inst160 ( // @[Snxn100k.scala 26996:35]
    .io_a(inst_SnxnLv4Inst160_io_a),
    .io_b(inst_SnxnLv4Inst160_io_b),
    .io_z(inst_SnxnLv4Inst160_io_z)
  );
  SnxnLv4Inst69 inst_SnxnLv4Inst161 ( // @[Snxn100k.scala 27000:35]
    .io_a(inst_SnxnLv4Inst161_io_a),
    .io_b(inst_SnxnLv4Inst161_io_b),
    .io_z(inst_SnxnLv4Inst161_io_z)
  );
  SnxnLv4Inst162 inst_SnxnLv4Inst162 ( // @[Snxn100k.scala 27004:35]
    .io_a(inst_SnxnLv4Inst162_io_a),
    .io_b(inst_SnxnLv4Inst162_io_b),
    .io_z(inst_SnxnLv4Inst162_io_z)
  );
  SnxnLv4Inst12 inst_SnxnLv4Inst163 ( // @[Snxn100k.scala 27008:35]
    .io_a(inst_SnxnLv4Inst163_io_a),
    .io_b(inst_SnxnLv4Inst163_io_b),
    .io_z(inst_SnxnLv4Inst163_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27013:15]
  assign inst_SnxnLv4Inst160_io_a = io_a; // @[Snxn100k.scala 26997:28]
  assign inst_SnxnLv4Inst160_io_b = io_b; // @[Snxn100k.scala 26998:28]
  assign inst_SnxnLv4Inst161_io_a = io_a; // @[Snxn100k.scala 27001:28]
  assign inst_SnxnLv4Inst161_io_b = io_b; // @[Snxn100k.scala 27002:28]
  assign inst_SnxnLv4Inst162_io_a = io_a; // @[Snxn100k.scala 27005:28]
  assign inst_SnxnLv4Inst162_io_b = io_b; // @[Snxn100k.scala 27006:28]
  assign inst_SnxnLv4Inst163_io_a = io_a; // @[Snxn100k.scala 27009:28]
  assign inst_SnxnLv4Inst163_io_b = io_b; // @[Snxn100k.scala 27010:28]
endmodule
module SnxnLv4Inst164(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 89293:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 89294:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 89295:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 89296:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 89297:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 89298:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 89299:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 89300:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 89301:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 89302:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 89303:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 89304:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 89305:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 89306:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 89307:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 89308:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 89309:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 89310:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 89311:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 89312:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 89313:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 89314:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 89315:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 89316:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 89317:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 89318:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 89319:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 89320:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 89321:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 89322:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 89323:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 89324:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 89325:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 89326:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 89327:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 89328:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 89329:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 89330:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 89331:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 89332:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 89333:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 89334:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 89335:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 89336:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 89337:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 89338:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 89339:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 89340:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 89341:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 89342:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 89343:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 89344:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 89345:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 89346:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 89347:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 89348:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 89349:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 89350:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 89351:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 89352:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 89353:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 89354:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 89355:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 89356:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 89357:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 89358:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 89359:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 89360:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 89361:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 89362:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 89363:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 89364:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 89365:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 89366:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 89367:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 89368:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 89369:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 89370:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 89371:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 89372:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 89373:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 89374:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 89375:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 89376:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 89377:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 89378:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 89379:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 89380:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 89381:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 89382:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 89383:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 89384:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 89385:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 89386:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 89387:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 89388:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 89389:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 89390:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 89391:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 89392:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 89393:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 89394:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 89395:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 89396:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 89397:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 89398:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 89399:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 89400:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 89401:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 89402:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 89403:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 89404:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 89405:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 89406:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 89407:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 89408:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 89409:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 89410:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 89411:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 89412:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 89413:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 89414:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 89415:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 89416:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 89417:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 89418:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 89419:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 89420:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 89421:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 89422:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 89423:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 89424:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 89425:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 89426:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 89427:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 89428:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 89429:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 89430:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 89431:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 89432:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 89433:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 89434:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 89435:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 89436:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 89437:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 89438:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 89439:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 89440:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 89441:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 89442:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 89443:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 89444:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 89445:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 89446:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 89447:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 89448:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 89449:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 89450:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 89451:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 89452:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 89453:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 89454:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 89455:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 89456:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 89457:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 89458:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 89459:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 89460:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 89461:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 89462:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 89463:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 89464:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 89465:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 89466:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 89467:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 89468:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 89469:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 89470:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 89471:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 89472:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 89473:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 89474:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 89475:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 89476:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 89477:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 89478:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 89479:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 89480:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 89481:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 89482:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 89483:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 89484:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 89485:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 89486:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 89487:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 89488:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 89489:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 89490:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 89491:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 89492:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 89493:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 89494:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 89495:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 89496:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 89497:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 89498:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 89499:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 89500:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 89501:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 89502:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 89503:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 89504:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 89505:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 89506:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 89507:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 89508:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 89509:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 89510:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 89511:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 89512:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 89513:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 89514:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 89515:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 89516:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 89517:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 89518:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 89519:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 89520:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 89521:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 89522:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 89523:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 89524:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 89525:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 89526:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 89527:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 89528:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 89529:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 89530:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 89531:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 89532:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 89533:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 89534:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 89535:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 89536:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 89537:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 89538:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 89539:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 89540:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 89541:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 89542:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 89543:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 89544:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 89545:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 89546:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 89547:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 89548:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 89549:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 89550:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 89551:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 89552:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 89553:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 89554:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 89555:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 89556:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 89557:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 89558:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 89559:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 89560:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 89561:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 89562:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 89563:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 89564:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 89565:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 89566:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 89567:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 89568:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 89569:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 89570:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 89571:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 89572:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 89573:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 89574:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 89575:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 89576:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 89577:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 89578:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 89579:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 89580:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 89581:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 89582:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 89583:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 89584:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 89585:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 89586:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 89587:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 89588:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 89589:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 89590:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 89591:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 89592:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 89593:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 89594:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 89595:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 89596:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 89597:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 89598:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 89599:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 89600:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 89601:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 89602:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 89603:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 89604:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 89605:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 89606:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 89607:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 89608:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 89609:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 89610:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 89611:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 89612:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 89613:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 89614:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 89615:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 89616:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 89617:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 89618:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 89619:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 89620:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 89621:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 89622:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 89623:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 89624:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 89625:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 89626:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 89627:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 89628:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 89629:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 89630:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 89631:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 89632:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 89633:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 89634:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 89635:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 89636:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 89637:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 89638:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 89639:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 89640:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 89641:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 89642:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 89643:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 89644:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 89645:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 89646:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 89647:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 89648:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 89649:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 89650:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 89651:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 89652:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 89653:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 89654:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 89655:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 89656:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 89657:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 89658:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 89659:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 89660:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 89661:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 89662:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 89663:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 89664:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 89665:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 89666:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 89667:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 89668:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 89669:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 89670:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 89671:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 89672:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 89673:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 89674:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 89675:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 89676:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 89677:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 89678:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 89679:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 89680:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 89681:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 89682:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 89683:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 89684:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 89685:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 89686:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 89687:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 89688:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 89689:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 89690:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 89691:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 89692:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 89693:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 89694:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 89695:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 89696:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 89697:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 89698:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 89699:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 89700:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 89701:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 89702:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 89703:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 89704:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 89705:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 89706:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 89707:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 89708:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 89709:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 89710:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 89711:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 89712:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 89713:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 89714:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 89715:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 89716:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 89717:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 89718:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 89719:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 89720:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 89721:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 89722:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 89723:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 89724:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 89725:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 89726:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 89727:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 89728:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 89729:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 89730:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 89731:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 89732:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 89733:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 89734:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 89735:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 89736:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 89737:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 89738:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 89739:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 89740:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 89741:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 89742:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 89743:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 89744:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 89745:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 89746:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 89747:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 89748:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 89749:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 89750:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 89751:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 89752:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 89753:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 89754:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 89755:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 89756:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 89757:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 89758:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 89759:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 89760:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 89761:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 89762:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 89763:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 89764:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 89765:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 89766:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 89767:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 89768:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 89769:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 89770:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 89771:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 89772:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 89773:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 89774:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 89775:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 89776:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 89777:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 89778:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 89779:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 89780:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 89781:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 89782:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 89783:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 89784:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 89785:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 89786:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 89787:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 89788:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 89789:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 89790:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 89791:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 89792:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 89793:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 89794:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 89795:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 89796:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 89797:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 89798:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 89799:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 89800:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 89801:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 89802:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 89803:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 89804:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 89805:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 89806:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 89807:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 89808:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 89809:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 89810:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 89811:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 89812:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 89813:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 89814:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 89815:22]
  wire  invx130 = ~x130; // @[Snxn100k.scala 89816:17]
  wire  t131 = x130 + invx130; // @[Snxn100k.scala 89817:22]
  wire  inv131 = ~t131; // @[Snxn100k.scala 89818:17]
  wire  x131 = t131 ^ inv131; // @[Snxn100k.scala 89819:22]
  wire  invx131 = ~x131; // @[Snxn100k.scala 89820:17]
  wire  t132 = x131 + invx131; // @[Snxn100k.scala 89821:22]
  wire  inv132 = ~t132; // @[Snxn100k.scala 89822:17]
  wire  x132 = t132 ^ inv132; // @[Snxn100k.scala 89823:22]
  wire  invx132 = ~x132; // @[Snxn100k.scala 89824:17]
  wire  t133 = x132 + invx132; // @[Snxn100k.scala 89825:22]
  wire  inv133 = ~t133; // @[Snxn100k.scala 89826:17]
  wire  x133 = t133 ^ inv133; // @[Snxn100k.scala 89827:22]
  wire  invx133 = ~x133; // @[Snxn100k.scala 89828:17]
  wire  t134 = x133 + invx133; // @[Snxn100k.scala 89829:22]
  wire  inv134 = ~t134; // @[Snxn100k.scala 89830:17]
  wire  x134 = t134 ^ inv134; // @[Snxn100k.scala 89831:22]
  wire  invx134 = ~x134; // @[Snxn100k.scala 89832:17]
  wire  t135 = x134 + invx134; // @[Snxn100k.scala 89833:22]
  wire  inv135 = ~t135; // @[Snxn100k.scala 89834:17]
  wire  x135 = t135 ^ inv135; // @[Snxn100k.scala 89835:22]
  wire  invx135 = ~x135; // @[Snxn100k.scala 89836:17]
  wire  t136 = x135 + invx135; // @[Snxn100k.scala 89837:22]
  wire  inv136 = ~t136; // @[Snxn100k.scala 89838:17]
  wire  x136 = t136 ^ inv136; // @[Snxn100k.scala 89839:22]
  assign io_z = ~x136; // @[Snxn100k.scala 89840:17]
endmodule
module SnxnLv3Inst41(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst164_io_a; // @[Snxn100k.scala 26290:35]
  wire  inst_SnxnLv4Inst164_io_b; // @[Snxn100k.scala 26290:35]
  wire  inst_SnxnLv4Inst164_io_z; // @[Snxn100k.scala 26290:35]
  wire  inst_SnxnLv4Inst165_io_a; // @[Snxn100k.scala 26294:35]
  wire  inst_SnxnLv4Inst165_io_b; // @[Snxn100k.scala 26294:35]
  wire  inst_SnxnLv4Inst165_io_z; // @[Snxn100k.scala 26294:35]
  wire  inst_SnxnLv4Inst166_io_a; // @[Snxn100k.scala 26298:35]
  wire  inst_SnxnLv4Inst166_io_b; // @[Snxn100k.scala 26298:35]
  wire  inst_SnxnLv4Inst166_io_z; // @[Snxn100k.scala 26298:35]
  wire  inst_SnxnLv4Inst167_io_a; // @[Snxn100k.scala 26302:35]
  wire  inst_SnxnLv4Inst167_io_b; // @[Snxn100k.scala 26302:35]
  wire  inst_SnxnLv4Inst167_io_z; // @[Snxn100k.scala 26302:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst164_io_z + inst_SnxnLv4Inst165_io_z; // @[Snxn100k.scala 26306:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst166_io_z; // @[Snxn100k.scala 26306:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst167_io_z; // @[Snxn100k.scala 26306:92]
  SnxnLv4Inst164 inst_SnxnLv4Inst164 ( // @[Snxn100k.scala 26290:35]
    .io_a(inst_SnxnLv4Inst164_io_a),
    .io_b(inst_SnxnLv4Inst164_io_b),
    .io_z(inst_SnxnLv4Inst164_io_z)
  );
  SnxnLv4Inst15 inst_SnxnLv4Inst165 ( // @[Snxn100k.scala 26294:35]
    .io_a(inst_SnxnLv4Inst165_io_a),
    .io_b(inst_SnxnLv4Inst165_io_b),
    .io_z(inst_SnxnLv4Inst165_io_z)
  );
  SnxnLv4Inst42 inst_SnxnLv4Inst166 ( // @[Snxn100k.scala 26298:35]
    .io_a(inst_SnxnLv4Inst166_io_a),
    .io_b(inst_SnxnLv4Inst166_io_b),
    .io_z(inst_SnxnLv4Inst166_io_z)
  );
  SnxnLv4Inst8 inst_SnxnLv4Inst167 ( // @[Snxn100k.scala 26302:35]
    .io_a(inst_SnxnLv4Inst167_io_a),
    .io_b(inst_SnxnLv4Inst167_io_b),
    .io_z(inst_SnxnLv4Inst167_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26307:15]
  assign inst_SnxnLv4Inst164_io_a = io_a; // @[Snxn100k.scala 26291:28]
  assign inst_SnxnLv4Inst164_io_b = io_b; // @[Snxn100k.scala 26292:28]
  assign inst_SnxnLv4Inst165_io_a = io_a; // @[Snxn100k.scala 26295:28]
  assign inst_SnxnLv4Inst165_io_b = io_b; // @[Snxn100k.scala 26296:28]
  assign inst_SnxnLv4Inst166_io_a = io_a; // @[Snxn100k.scala 26299:28]
  assign inst_SnxnLv4Inst166_io_b = io_b; // @[Snxn100k.scala 26300:28]
  assign inst_SnxnLv4Inst167_io_a = io_a; // @[Snxn100k.scala 26303:28]
  assign inst_SnxnLv4Inst167_io_b = io_b; // @[Snxn100k.scala 26304:28]
endmodule
module SnxnLv4Inst168(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 89851:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 89852:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 89853:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 89854:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 89855:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 89856:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 89857:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 89858:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 89859:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 89860:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 89861:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 89862:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 89863:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 89864:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 89865:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 89866:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 89867:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 89868:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 89869:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 89870:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 89871:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 89872:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 89873:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 89874:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 89875:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 89876:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 89877:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 89878:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 89879:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 89880:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 89881:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 89882:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 89883:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 89884:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 89885:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 89886:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 89887:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 89888:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 89889:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 89890:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 89891:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 89892:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 89893:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 89894:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 89895:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 89896:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 89897:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 89898:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 89899:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 89900:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 89901:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 89902:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 89903:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 89904:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 89905:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 89906:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 89907:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 89908:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 89909:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 89910:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 89911:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 89912:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 89913:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 89914:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 89915:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 89916:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 89917:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 89918:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 89919:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 89920:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 89921:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 89922:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 89923:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 89924:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 89925:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 89926:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 89927:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 89928:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 89929:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 89930:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 89931:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 89932:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 89933:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 89934:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 89935:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 89936:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 89937:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 89938:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 89939:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 89940:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 89941:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 89942:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 89943:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 89944:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 89945:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 89946:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 89947:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 89948:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 89949:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 89950:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 89951:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 89952:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 89953:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 89954:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 89955:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 89956:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 89957:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 89958:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 89959:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 89960:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 89961:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 89962:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 89963:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 89964:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 89965:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 89966:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 89967:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 89968:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 89969:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 89970:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 89971:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 89972:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 89973:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 89974:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 89975:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 89976:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 89977:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 89978:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 89979:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 89980:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 89981:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 89982:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 89983:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 89984:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 89985:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 89986:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 89987:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 89988:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 89989:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 89990:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 89991:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 89992:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 89993:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 89994:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 89995:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 89996:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 89997:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 89998:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 89999:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 90000:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 90001:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 90002:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 90003:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 90004:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 90005:20]
  assign io_z = ~x38; // @[Snxn100k.scala 90006:16]
endmodule
module SnxnLv4Inst171(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 90017:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 90018:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 90019:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 90020:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 90021:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 90022:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 90023:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 90024:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 90025:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 90026:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 90027:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 90028:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 90029:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 90030:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 90031:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 90032:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 90033:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 90034:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 90035:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 90036:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 90037:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 90038:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 90039:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 90040:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 90041:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 90042:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 90043:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 90044:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 90045:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 90046:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 90047:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 90048:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 90049:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 90050:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 90051:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 90052:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 90053:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 90054:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 90055:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 90056:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 90057:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 90058:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 90059:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 90060:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 90061:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 90062:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 90063:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 90064:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 90065:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 90066:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 90067:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 90068:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 90069:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 90070:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 90071:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 90072:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 90073:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 90074:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 90075:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 90076:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 90077:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 90078:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 90079:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 90080:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 90081:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 90082:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 90083:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 90084:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 90085:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 90086:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 90087:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 90088:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 90089:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 90090:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 90091:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 90092:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 90093:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 90094:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 90095:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 90096:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 90097:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 90098:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 90099:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 90100:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 90101:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 90102:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 90103:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 90104:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 90105:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 90106:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 90107:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 90108:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 90109:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 90110:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 90111:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 90112:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 90113:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 90114:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 90115:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 90116:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 90117:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 90118:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 90119:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 90120:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 90121:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 90122:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 90123:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 90124:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 90125:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 90126:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 90127:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 90128:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 90129:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 90130:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 90131:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 90132:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 90133:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 90134:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 90135:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 90136:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 90137:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 90138:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 90139:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 90140:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 90141:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 90142:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 90143:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 90144:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 90145:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 90146:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 90147:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 90148:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 90149:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 90150:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 90151:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 90152:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 90153:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 90154:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 90155:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 90156:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 90157:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 90158:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 90159:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 90160:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 90161:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 90162:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 90163:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 90164:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 90165:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 90166:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 90167:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 90168:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 90169:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 90170:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 90171:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 90172:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 90173:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 90174:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 90175:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 90176:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 90177:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 90178:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 90179:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 90180:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 90181:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 90182:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 90183:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 90184:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 90185:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 90186:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 90187:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 90188:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 90189:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 90190:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 90191:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 90192:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 90193:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 90194:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 90195:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 90196:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 90197:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 90198:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 90199:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 90200:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 90201:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 90202:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 90203:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 90204:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 90205:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 90206:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 90207:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 90208:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 90209:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 90210:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 90211:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 90212:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 90213:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 90214:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 90215:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 90216:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 90217:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 90218:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 90219:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 90220:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 90221:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 90222:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 90223:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 90224:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 90225:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 90226:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 90227:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 90228:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 90229:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 90230:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 90231:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 90232:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 90233:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 90234:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 90235:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 90236:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 90237:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 90238:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 90239:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 90240:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 90241:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 90242:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 90243:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 90244:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 90245:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 90246:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 90247:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 90248:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 90249:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 90250:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 90251:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 90252:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 90253:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 90254:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 90255:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 90256:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 90257:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 90258:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 90259:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 90260:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 90261:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 90262:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 90263:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 90264:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 90265:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 90266:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 90267:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 90268:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 90269:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 90270:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 90271:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 90272:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 90273:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 90274:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 90275:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 90276:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 90277:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 90278:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 90279:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 90280:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 90281:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 90282:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 90283:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 90284:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 90285:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 90286:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 90287:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 90288:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 90289:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 90290:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 90291:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 90292:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 90293:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 90294:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 90295:20]
  assign io_z = ~x69; // @[Snxn100k.scala 90296:16]
endmodule
module SnxnLv3Inst42(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst168_io_a; // @[Snxn100k.scala 26601:35]
  wire  inst_SnxnLv4Inst168_io_b; // @[Snxn100k.scala 26601:35]
  wire  inst_SnxnLv4Inst168_io_z; // @[Snxn100k.scala 26601:35]
  wire  inst_SnxnLv4Inst169_io_a; // @[Snxn100k.scala 26605:35]
  wire  inst_SnxnLv4Inst169_io_b; // @[Snxn100k.scala 26605:35]
  wire  inst_SnxnLv4Inst169_io_z; // @[Snxn100k.scala 26605:35]
  wire  inst_SnxnLv4Inst170_io_a; // @[Snxn100k.scala 26609:35]
  wire  inst_SnxnLv4Inst170_io_b; // @[Snxn100k.scala 26609:35]
  wire  inst_SnxnLv4Inst170_io_z; // @[Snxn100k.scala 26609:35]
  wire  inst_SnxnLv4Inst171_io_a; // @[Snxn100k.scala 26613:35]
  wire  inst_SnxnLv4Inst171_io_b; // @[Snxn100k.scala 26613:35]
  wire  inst_SnxnLv4Inst171_io_z; // @[Snxn100k.scala 26613:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst168_io_z + inst_SnxnLv4Inst169_io_z; // @[Snxn100k.scala 26617:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst170_io_z; // @[Snxn100k.scala 26617:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst171_io_z; // @[Snxn100k.scala 26617:92]
  SnxnLv4Inst168 inst_SnxnLv4Inst168 ( // @[Snxn100k.scala 26601:35]
    .io_a(inst_SnxnLv4Inst168_io_a),
    .io_b(inst_SnxnLv4Inst168_io_b),
    .io_z(inst_SnxnLv4Inst168_io_z)
  );
  SnxnLv4Inst36 inst_SnxnLv4Inst169 ( // @[Snxn100k.scala 26605:35]
    .io_a(inst_SnxnLv4Inst169_io_a),
    .io_b(inst_SnxnLv4Inst169_io_b),
    .io_z(inst_SnxnLv4Inst169_io_z)
  );
  SnxnLv4Inst48 inst_SnxnLv4Inst170 ( // @[Snxn100k.scala 26609:35]
    .io_a(inst_SnxnLv4Inst170_io_a),
    .io_b(inst_SnxnLv4Inst170_io_b),
    .io_z(inst_SnxnLv4Inst170_io_z)
  );
  SnxnLv4Inst171 inst_SnxnLv4Inst171 ( // @[Snxn100k.scala 26613:35]
    .io_a(inst_SnxnLv4Inst171_io_a),
    .io_b(inst_SnxnLv4Inst171_io_b),
    .io_z(inst_SnxnLv4Inst171_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 26618:15]
  assign inst_SnxnLv4Inst168_io_a = io_a; // @[Snxn100k.scala 26602:28]
  assign inst_SnxnLv4Inst168_io_b = io_b; // @[Snxn100k.scala 26603:28]
  assign inst_SnxnLv4Inst169_io_a = io_a; // @[Snxn100k.scala 26606:28]
  assign inst_SnxnLv4Inst169_io_b = io_b; // @[Snxn100k.scala 26607:28]
  assign inst_SnxnLv4Inst170_io_a = io_a; // @[Snxn100k.scala 26610:28]
  assign inst_SnxnLv4Inst170_io_b = io_b; // @[Snxn100k.scala 26611:28]
  assign inst_SnxnLv4Inst171_io_a = io_a; // @[Snxn100k.scala 26614:28]
  assign inst_SnxnLv4Inst171_io_b = io_b; // @[Snxn100k.scala 26615:28]
endmodule
module SnxnLv4Inst174(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 92499:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 92500:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 92501:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 92502:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 92503:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 92504:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 92505:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 92506:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 92507:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 92508:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 92509:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 92510:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 92511:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 92512:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 92513:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 92514:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 92515:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 92516:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 92517:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 92518:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 92519:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 92520:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 92521:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 92522:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 92523:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 92524:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 92525:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 92526:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 92527:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 92528:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 92529:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 92530:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 92531:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 92532:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 92533:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 92534:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 92535:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 92536:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 92537:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 92538:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 92539:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 92540:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 92541:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 92542:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 92543:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 92544:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 92545:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 92546:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 92547:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 92548:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 92549:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 92550:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 92551:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 92552:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 92553:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 92554:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 92555:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 92556:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 92557:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 92558:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 92559:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 92560:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 92561:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 92562:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 92563:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 92564:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 92565:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 92566:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 92567:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 92568:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 92569:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 92570:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 92571:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 92572:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 92573:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 92574:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 92575:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 92576:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 92577:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 92578:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 92579:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 92580:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 92581:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 92582:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 92583:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 92584:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 92585:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 92586:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 92587:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 92588:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 92589:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 92590:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 92591:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 92592:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 92593:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 92594:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 92595:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 92596:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 92597:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 92598:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 92599:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 92600:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 92601:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 92602:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 92603:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 92604:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 92605:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 92606:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 92607:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 92608:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 92609:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 92610:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 92611:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 92612:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 92613:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 92614:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 92615:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 92616:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 92617:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 92618:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 92619:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 92620:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 92621:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 92622:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 92623:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 92624:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 92625:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 92626:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 92627:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 92628:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 92629:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 92630:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 92631:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 92632:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 92633:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 92634:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 92635:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 92636:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 92637:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 92638:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 92639:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 92640:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 92641:20]
  assign io_z = ~x35; // @[Snxn100k.scala 92642:16]
endmodule
module SnxnLv4Inst175(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 93023:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 93024:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 93025:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 93026:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 93027:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 93028:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 93029:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 93030:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 93031:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 93032:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 93033:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 93034:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 93035:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 93036:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 93037:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 93038:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 93039:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 93040:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 93041:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 93042:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 93043:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 93044:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 93045:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 93046:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 93047:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 93048:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 93049:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 93050:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 93051:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 93052:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 93053:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 93054:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 93055:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 93056:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 93057:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 93058:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 93059:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 93060:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 93061:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 93062:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 93063:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 93064:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 93065:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 93066:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 93067:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 93068:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 93069:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 93070:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 93071:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 93072:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 93073:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 93074:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 93075:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 93076:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 93077:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 93078:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 93079:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 93080:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 93081:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 93082:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 93083:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 93084:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 93085:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 93086:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 93087:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 93088:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 93089:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 93090:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 93091:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 93092:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 93093:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 93094:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 93095:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 93096:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 93097:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 93098:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 93099:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 93100:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 93101:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 93102:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 93103:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 93104:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 93105:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 93106:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 93107:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 93108:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 93109:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 93110:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 93111:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 93112:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 93113:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 93114:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 93115:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 93116:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 93117:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 93118:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 93119:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 93120:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 93121:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 93122:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 93123:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 93124:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 93125:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 93126:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 93127:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 93128:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 93129:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 93130:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 93131:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 93132:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 93133:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 93134:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 93135:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 93136:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 93137:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 93138:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 93139:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 93140:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 93141:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 93142:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 93143:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 93144:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 93145:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 93146:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 93147:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 93148:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 93149:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 93150:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 93151:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 93152:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 93153:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 93154:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 93155:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 93156:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 93157:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 93158:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 93159:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 93160:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 93161:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 93162:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 93163:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 93164:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 93165:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 93166:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 93167:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 93168:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 93169:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 93170:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 93171:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 93172:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 93173:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 93174:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 93175:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 93176:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 93177:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 93178:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 93179:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 93180:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 93181:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 93182:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 93183:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 93184:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 93185:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 93186:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 93187:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 93188:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 93189:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 93190:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 93191:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 93192:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 93193:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 93194:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 93195:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 93196:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 93197:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 93198:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 93199:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 93200:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 93201:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 93202:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 93203:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 93204:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 93205:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 93206:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 93207:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 93208:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 93209:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 93210:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 93211:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 93212:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 93213:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 93214:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 93215:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 93216:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 93217:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 93218:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 93219:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 93220:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 93221:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 93222:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 93223:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 93224:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 93225:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 93226:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 93227:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 93228:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 93229:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 93230:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 93231:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 93232:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 93233:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 93234:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 93235:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 93236:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 93237:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 93238:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 93239:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 93240:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 93241:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 93242:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 93243:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 93244:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 93245:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 93246:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 93247:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 93248:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 93249:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 93250:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 93251:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 93252:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 93253:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 93254:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 93255:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 93256:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 93257:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 93258:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 93259:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 93260:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 93261:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 93262:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 93263:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 93264:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 93265:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 93266:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 93267:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 93268:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 93269:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 93270:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 93271:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 93272:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 93273:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 93274:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 93275:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 93276:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 93277:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 93278:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 93279:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 93280:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 93281:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 93282:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 93283:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 93284:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 93285:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 93286:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 93287:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 93288:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 93289:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 93290:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 93291:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 93292:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 93293:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 93294:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 93295:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 93296:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 93297:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 93298:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 93299:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 93300:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 93301:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 93302:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 93303:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 93304:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 93305:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 93306:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 93307:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 93308:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 93309:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 93310:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 93311:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 93312:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 93313:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 93314:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 93315:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 93316:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 93317:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 93318:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 93319:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 93320:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 93321:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 93322:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 93323:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 93324:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 93325:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 93326:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 93327:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 93328:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 93329:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 93330:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 93331:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 93332:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 93333:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 93334:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 93335:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 93336:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 93337:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 93338:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 93339:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 93340:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 93341:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 93342:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 93343:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 93344:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 93345:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 93346:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 93347:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 93348:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 93349:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 93350:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 93351:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 93352:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 93353:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 93354:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 93355:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 93356:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 93357:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 93358:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 93359:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 93360:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 93361:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 93362:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 93363:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 93364:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 93365:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 93366:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 93367:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 93368:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 93369:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 93370:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 93371:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 93372:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 93373:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 93374:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 93375:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 93376:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 93377:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 93378:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 93379:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 93380:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 93381:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 93382:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 93383:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 93384:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 93385:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 93386:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 93387:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 93388:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 93389:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 93390:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 93391:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 93392:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 93393:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 93394:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 93395:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 93396:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 93397:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 93398:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 93399:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 93400:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 93401:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 93402:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 93403:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 93404:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 93405:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 93406:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 93407:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 93408:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 93409:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 93410:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 93411:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 93412:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 93413:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 93414:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 93415:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 93416:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 93417:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 93418:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 93419:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 93420:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 93421:20]
  assign io_z = ~x99; // @[Snxn100k.scala 93422:16]
endmodule
module SnxnLv3Inst43(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst172_io_a; // @[Snxn100k.scala 27075:35]
  wire  inst_SnxnLv4Inst172_io_b; // @[Snxn100k.scala 27075:35]
  wire  inst_SnxnLv4Inst172_io_z; // @[Snxn100k.scala 27075:35]
  wire  inst_SnxnLv4Inst173_io_a; // @[Snxn100k.scala 27079:35]
  wire  inst_SnxnLv4Inst173_io_b; // @[Snxn100k.scala 27079:35]
  wire  inst_SnxnLv4Inst173_io_z; // @[Snxn100k.scala 27079:35]
  wire  inst_SnxnLv4Inst174_io_a; // @[Snxn100k.scala 27083:35]
  wire  inst_SnxnLv4Inst174_io_b; // @[Snxn100k.scala 27083:35]
  wire  inst_SnxnLv4Inst174_io_z; // @[Snxn100k.scala 27083:35]
  wire  inst_SnxnLv4Inst175_io_a; // @[Snxn100k.scala 27087:35]
  wire  inst_SnxnLv4Inst175_io_b; // @[Snxn100k.scala 27087:35]
  wire  inst_SnxnLv4Inst175_io_z; // @[Snxn100k.scala 27087:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst172_io_z + inst_SnxnLv4Inst173_io_z; // @[Snxn100k.scala 27091:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst174_io_z; // @[Snxn100k.scala 27091:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst175_io_z; // @[Snxn100k.scala 27091:92]
  SnxnLv4Inst101 inst_SnxnLv4Inst172 ( // @[Snxn100k.scala 27075:35]
    .io_a(inst_SnxnLv4Inst172_io_a),
    .io_b(inst_SnxnLv4Inst172_io_b),
    .io_z(inst_SnxnLv4Inst172_io_z)
  );
  SnxnLv4Inst12 inst_SnxnLv4Inst173 ( // @[Snxn100k.scala 27079:35]
    .io_a(inst_SnxnLv4Inst173_io_a),
    .io_b(inst_SnxnLv4Inst173_io_b),
    .io_z(inst_SnxnLv4Inst173_io_z)
  );
  SnxnLv4Inst174 inst_SnxnLv4Inst174 ( // @[Snxn100k.scala 27083:35]
    .io_a(inst_SnxnLv4Inst174_io_a),
    .io_b(inst_SnxnLv4Inst174_io_b),
    .io_z(inst_SnxnLv4Inst174_io_z)
  );
  SnxnLv4Inst175 inst_SnxnLv4Inst175 ( // @[Snxn100k.scala 27087:35]
    .io_a(inst_SnxnLv4Inst175_io_a),
    .io_b(inst_SnxnLv4Inst175_io_b),
    .io_z(inst_SnxnLv4Inst175_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27092:15]
  assign inst_SnxnLv4Inst172_io_a = io_a; // @[Snxn100k.scala 27076:28]
  assign inst_SnxnLv4Inst172_io_b = io_b; // @[Snxn100k.scala 27077:28]
  assign inst_SnxnLv4Inst173_io_a = io_a; // @[Snxn100k.scala 27080:28]
  assign inst_SnxnLv4Inst173_io_b = io_b; // @[Snxn100k.scala 27081:28]
  assign inst_SnxnLv4Inst174_io_a = io_a; // @[Snxn100k.scala 27084:28]
  assign inst_SnxnLv4Inst174_io_b = io_b; // @[Snxn100k.scala 27085:28]
  assign inst_SnxnLv4Inst175_io_a = io_a; // @[Snxn100k.scala 27088:28]
  assign inst_SnxnLv4Inst175_io_b = io_b; // @[Snxn100k.scala 27089:28]
endmodule
module SnxnLv2Inst10(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst40_io_a; // @[Snxn100k.scala 7875:34]
  wire  inst_SnxnLv3Inst40_io_b; // @[Snxn100k.scala 7875:34]
  wire  inst_SnxnLv3Inst40_io_z; // @[Snxn100k.scala 7875:34]
  wire  inst_SnxnLv3Inst41_io_a; // @[Snxn100k.scala 7879:34]
  wire  inst_SnxnLv3Inst41_io_b; // @[Snxn100k.scala 7879:34]
  wire  inst_SnxnLv3Inst41_io_z; // @[Snxn100k.scala 7879:34]
  wire  inst_SnxnLv3Inst42_io_a; // @[Snxn100k.scala 7883:34]
  wire  inst_SnxnLv3Inst42_io_b; // @[Snxn100k.scala 7883:34]
  wire  inst_SnxnLv3Inst42_io_z; // @[Snxn100k.scala 7883:34]
  wire  inst_SnxnLv3Inst43_io_a; // @[Snxn100k.scala 7887:34]
  wire  inst_SnxnLv3Inst43_io_b; // @[Snxn100k.scala 7887:34]
  wire  inst_SnxnLv3Inst43_io_z; // @[Snxn100k.scala 7887:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst40_io_z + inst_SnxnLv3Inst41_io_z; // @[Snxn100k.scala 7891:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst42_io_z; // @[Snxn100k.scala 7891:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst43_io_z; // @[Snxn100k.scala 7891:89]
  SnxnLv3Inst40 inst_SnxnLv3Inst40 ( // @[Snxn100k.scala 7875:34]
    .io_a(inst_SnxnLv3Inst40_io_a),
    .io_b(inst_SnxnLv3Inst40_io_b),
    .io_z(inst_SnxnLv3Inst40_io_z)
  );
  SnxnLv3Inst41 inst_SnxnLv3Inst41 ( // @[Snxn100k.scala 7879:34]
    .io_a(inst_SnxnLv3Inst41_io_a),
    .io_b(inst_SnxnLv3Inst41_io_b),
    .io_z(inst_SnxnLv3Inst41_io_z)
  );
  SnxnLv3Inst42 inst_SnxnLv3Inst42 ( // @[Snxn100k.scala 7883:34]
    .io_a(inst_SnxnLv3Inst42_io_a),
    .io_b(inst_SnxnLv3Inst42_io_b),
    .io_z(inst_SnxnLv3Inst42_io_z)
  );
  SnxnLv3Inst43 inst_SnxnLv3Inst43 ( // @[Snxn100k.scala 7887:34]
    .io_a(inst_SnxnLv3Inst43_io_a),
    .io_b(inst_SnxnLv3Inst43_io_b),
    .io_z(inst_SnxnLv3Inst43_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 7892:15]
  assign inst_SnxnLv3Inst40_io_a = io_a; // @[Snxn100k.scala 7876:27]
  assign inst_SnxnLv3Inst40_io_b = io_b; // @[Snxn100k.scala 7877:27]
  assign inst_SnxnLv3Inst41_io_a = io_a; // @[Snxn100k.scala 7880:27]
  assign inst_SnxnLv3Inst41_io_b = io_b; // @[Snxn100k.scala 7881:27]
  assign inst_SnxnLv3Inst42_io_a = io_a; // @[Snxn100k.scala 7884:27]
  assign inst_SnxnLv3Inst42_io_b = io_b; // @[Snxn100k.scala 7885:27]
  assign inst_SnxnLv3Inst43_io_a = io_a; // @[Snxn100k.scala 7888:27]
  assign inst_SnxnLv3Inst43_io_b = io_b; // @[Snxn100k.scala 7889:27]
endmodule
module SnxnLv3Inst44(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst176_io_a; // @[Snxn100k.scala 27457:35]
  wire  inst_SnxnLv4Inst176_io_b; // @[Snxn100k.scala 27457:35]
  wire  inst_SnxnLv4Inst176_io_z; // @[Snxn100k.scala 27457:35]
  wire  inst_SnxnLv4Inst177_io_a; // @[Snxn100k.scala 27461:35]
  wire  inst_SnxnLv4Inst177_io_b; // @[Snxn100k.scala 27461:35]
  wire  inst_SnxnLv4Inst177_io_z; // @[Snxn100k.scala 27461:35]
  wire  inst_SnxnLv4Inst178_io_a; // @[Snxn100k.scala 27465:35]
  wire  inst_SnxnLv4Inst178_io_b; // @[Snxn100k.scala 27465:35]
  wire  inst_SnxnLv4Inst178_io_z; // @[Snxn100k.scala 27465:35]
  wire  inst_SnxnLv4Inst179_io_a; // @[Snxn100k.scala 27469:35]
  wire  inst_SnxnLv4Inst179_io_b; // @[Snxn100k.scala 27469:35]
  wire  inst_SnxnLv4Inst179_io_z; // @[Snxn100k.scala 27469:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst176_io_z + inst_SnxnLv4Inst177_io_z; // @[Snxn100k.scala 27473:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst178_io_z; // @[Snxn100k.scala 27473:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst179_io_z; // @[Snxn100k.scala 27473:92]
  SnxnLv4Inst90 inst_SnxnLv4Inst176 ( // @[Snxn100k.scala 27457:35]
    .io_a(inst_SnxnLv4Inst176_io_a),
    .io_b(inst_SnxnLv4Inst176_io_b),
    .io_z(inst_SnxnLv4Inst176_io_z)
  );
  SnxnLv4Inst54 inst_SnxnLv4Inst177 ( // @[Snxn100k.scala 27461:35]
    .io_a(inst_SnxnLv4Inst177_io_a),
    .io_b(inst_SnxnLv4Inst177_io_b),
    .io_z(inst_SnxnLv4Inst177_io_z)
  );
  SnxnLv4Inst67 inst_SnxnLv4Inst178 ( // @[Snxn100k.scala 27465:35]
    .io_a(inst_SnxnLv4Inst178_io_a),
    .io_b(inst_SnxnLv4Inst178_io_b),
    .io_z(inst_SnxnLv4Inst178_io_z)
  );
  SnxnLv4Inst9 inst_SnxnLv4Inst179 ( // @[Snxn100k.scala 27469:35]
    .io_a(inst_SnxnLv4Inst179_io_a),
    .io_b(inst_SnxnLv4Inst179_io_b),
    .io_z(inst_SnxnLv4Inst179_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27474:15]
  assign inst_SnxnLv4Inst176_io_a = io_a; // @[Snxn100k.scala 27458:28]
  assign inst_SnxnLv4Inst176_io_b = io_b; // @[Snxn100k.scala 27459:28]
  assign inst_SnxnLv4Inst177_io_a = io_a; // @[Snxn100k.scala 27462:28]
  assign inst_SnxnLv4Inst177_io_b = io_b; // @[Snxn100k.scala 27463:28]
  assign inst_SnxnLv4Inst178_io_a = io_a; // @[Snxn100k.scala 27466:28]
  assign inst_SnxnLv4Inst178_io_b = io_b; // @[Snxn100k.scala 27467:28]
  assign inst_SnxnLv4Inst179_io_a = io_a; // @[Snxn100k.scala 27470:28]
  assign inst_SnxnLv4Inst179_io_b = io_b; // @[Snxn100k.scala 27471:28]
endmodule
module SnxnLv4Inst181(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 98017:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 98018:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 98019:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 98020:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 98021:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 98022:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 98023:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 98024:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 98025:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 98026:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 98027:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 98028:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 98029:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 98030:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 98031:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 98032:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 98033:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 98034:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 98035:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 98036:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 98037:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 98038:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 98039:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 98040:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 98041:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 98042:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 98043:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 98044:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 98045:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 98046:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 98047:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 98048:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 98049:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 98050:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 98051:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 98052:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 98053:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 98054:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 98055:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 98056:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 98057:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 98058:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 98059:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 98060:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 98061:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 98062:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 98063:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 98064:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 98065:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 98066:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 98067:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 98068:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 98069:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 98070:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 98071:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 98072:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 98073:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 98074:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 98075:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 98076:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 98077:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 98078:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 98079:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 98080:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 98081:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 98082:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 98083:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 98084:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 98085:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 98086:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 98087:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 98088:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 98089:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 98090:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 98091:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 98092:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 98093:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 98094:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 98095:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 98096:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 98097:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 98098:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 98099:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 98100:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 98101:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 98102:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 98103:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 98104:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 98105:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 98106:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 98107:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 98108:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 98109:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 98110:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 98111:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 98112:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 98113:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 98114:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 98115:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 98116:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 98117:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 98118:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 98119:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 98120:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 98121:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 98122:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 98123:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 98124:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 98125:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 98126:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 98127:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 98128:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 98129:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 98130:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 98131:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 98132:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 98133:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 98134:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 98135:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 98136:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 98137:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 98138:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 98139:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 98140:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 98141:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 98142:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 98143:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 98144:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 98145:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 98146:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 98147:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 98148:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 98149:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 98150:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 98151:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 98152:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 98153:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 98154:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 98155:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 98156:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 98157:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 98158:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 98159:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 98160:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 98161:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 98162:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 98163:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 98164:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 98165:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 98166:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 98167:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 98168:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 98169:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 98170:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 98171:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 98172:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 98173:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 98174:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 98175:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 98176:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 98177:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 98178:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 98179:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 98180:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 98181:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 98182:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 98183:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 98184:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 98185:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 98186:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 98187:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 98188:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 98189:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 98190:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 98191:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 98192:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 98193:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 98194:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 98195:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 98196:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 98197:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 98198:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 98199:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 98200:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 98201:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 98202:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 98203:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 98204:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 98205:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 98206:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 98207:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 98208:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 98209:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 98210:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 98211:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 98212:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 98213:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 98214:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 98215:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 98216:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 98217:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 98218:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 98219:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 98220:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 98221:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 98222:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 98223:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 98224:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 98225:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 98226:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 98227:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 98228:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 98229:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 98230:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 98231:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 98232:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 98233:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 98234:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 98235:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 98236:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 98237:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 98238:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 98239:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 98240:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 98241:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 98242:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 98243:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 98244:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 98245:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 98246:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 98247:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 98248:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 98249:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 98250:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 98251:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 98252:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 98253:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 98254:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 98255:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 98256:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 98257:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 98258:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 98259:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 98260:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 98261:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 98262:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 98263:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 98264:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 98265:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 98266:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 98267:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 98268:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 98269:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 98270:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 98271:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 98272:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 98273:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 98274:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 98275:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 98276:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 98277:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 98278:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 98279:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 98280:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 98281:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 98282:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 98283:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 98284:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 98285:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 98286:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 98287:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 98288:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 98289:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 98290:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 98291:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 98292:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 98293:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 98294:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 98295:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 98296:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 98297:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 98298:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 98299:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 98300:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 98301:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 98302:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 98303:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 98304:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 98305:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 98306:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 98307:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 98308:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 98309:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 98310:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 98311:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 98312:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 98313:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 98314:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 98315:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 98316:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 98317:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 98318:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 98319:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 98320:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 98321:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 98322:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 98323:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 98324:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 98325:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 98326:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 98327:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 98328:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 98329:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 98330:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 98331:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 98332:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 98333:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 98334:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 98335:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 98336:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 98337:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 98338:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 98339:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 98340:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 98341:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 98342:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 98343:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 98344:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 98345:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 98346:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 98347:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 98348:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 98349:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 98350:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 98351:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 98352:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 98353:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 98354:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 98355:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 98356:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 98357:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 98358:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 98359:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 98360:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 98361:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 98362:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 98363:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 98364:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 98365:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 98366:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 98367:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 98368:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 98369:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 98370:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 98371:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 98372:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 98373:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 98374:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 98375:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 98376:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 98377:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 98378:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 98379:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 98380:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 98381:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 98382:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 98383:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 98384:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 98385:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 98386:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 98387:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 98388:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 98389:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 98390:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 98391:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 98392:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 98393:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 98394:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 98395:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 98396:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 98397:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 98398:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 98399:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 98400:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 98401:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 98402:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 98403:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 98404:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 98405:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 98406:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 98407:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 98408:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 98409:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 98410:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 98411:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 98412:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 98413:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 98414:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 98415:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 98416:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 98417:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 98418:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 98419:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 98420:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 98421:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 98422:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 98423:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 98424:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 98425:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 98426:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 98427:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 98428:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 98429:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 98430:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 98431:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 98432:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 98433:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 98434:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 98435:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 98436:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 98437:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 98438:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 98439:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 98440:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 98441:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 98442:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 98443:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 98444:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 98445:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 98446:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 98447:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 98448:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 98449:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 98450:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 98451:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 98452:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 98453:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 98454:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 98455:22]
  assign io_z = ~x109; // @[Snxn100k.scala 98456:17]
endmodule
module SnxnLv3Inst45(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst180_io_a; // @[Snxn100k.scala 27728:35]
  wire  inst_SnxnLv4Inst180_io_b; // @[Snxn100k.scala 27728:35]
  wire  inst_SnxnLv4Inst180_io_z; // @[Snxn100k.scala 27728:35]
  wire  inst_SnxnLv4Inst181_io_a; // @[Snxn100k.scala 27732:35]
  wire  inst_SnxnLv4Inst181_io_b; // @[Snxn100k.scala 27732:35]
  wire  inst_SnxnLv4Inst181_io_z; // @[Snxn100k.scala 27732:35]
  wire  inst_SnxnLv4Inst182_io_a; // @[Snxn100k.scala 27736:35]
  wire  inst_SnxnLv4Inst182_io_b; // @[Snxn100k.scala 27736:35]
  wire  inst_SnxnLv4Inst182_io_z; // @[Snxn100k.scala 27736:35]
  wire  inst_SnxnLv4Inst183_io_a; // @[Snxn100k.scala 27740:35]
  wire  inst_SnxnLv4Inst183_io_b; // @[Snxn100k.scala 27740:35]
  wire  inst_SnxnLv4Inst183_io_z; // @[Snxn100k.scala 27740:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst180_io_z + inst_SnxnLv4Inst181_io_z; // @[Snxn100k.scala 27744:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst182_io_z; // @[Snxn100k.scala 27744:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst183_io_z; // @[Snxn100k.scala 27744:92]
  SnxnLv4Inst31 inst_SnxnLv4Inst180 ( // @[Snxn100k.scala 27728:35]
    .io_a(inst_SnxnLv4Inst180_io_a),
    .io_b(inst_SnxnLv4Inst180_io_b),
    .io_z(inst_SnxnLv4Inst180_io_z)
  );
  SnxnLv4Inst181 inst_SnxnLv4Inst181 ( // @[Snxn100k.scala 27732:35]
    .io_a(inst_SnxnLv4Inst181_io_a),
    .io_b(inst_SnxnLv4Inst181_io_b),
    .io_z(inst_SnxnLv4Inst181_io_z)
  );
  SnxnLv4Inst26 inst_SnxnLv4Inst182 ( // @[Snxn100k.scala 27736:35]
    .io_a(inst_SnxnLv4Inst182_io_a),
    .io_b(inst_SnxnLv4Inst182_io_b),
    .io_z(inst_SnxnLv4Inst182_io_z)
  );
  SnxnLv4Inst162 inst_SnxnLv4Inst183 ( // @[Snxn100k.scala 27740:35]
    .io_a(inst_SnxnLv4Inst183_io_a),
    .io_b(inst_SnxnLv4Inst183_io_b),
    .io_z(inst_SnxnLv4Inst183_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27745:15]
  assign inst_SnxnLv4Inst180_io_a = io_a; // @[Snxn100k.scala 27729:28]
  assign inst_SnxnLv4Inst180_io_b = io_b; // @[Snxn100k.scala 27730:28]
  assign inst_SnxnLv4Inst181_io_a = io_a; // @[Snxn100k.scala 27733:28]
  assign inst_SnxnLv4Inst181_io_b = io_b; // @[Snxn100k.scala 27734:28]
  assign inst_SnxnLv4Inst182_io_a = io_a; // @[Snxn100k.scala 27737:28]
  assign inst_SnxnLv4Inst182_io_b = io_b; // @[Snxn100k.scala 27738:28]
  assign inst_SnxnLv4Inst183_io_a = io_a; // @[Snxn100k.scala 27741:28]
  assign inst_SnxnLv4Inst183_io_b = io_b; // @[Snxn100k.scala 27742:28]
endmodule
module SnxnLv4Inst184(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 98887:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 98888:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 98889:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 98890:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 98891:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 98892:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 98893:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 98894:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 98895:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 98896:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 98897:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 98898:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 98899:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 98900:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 98901:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 98902:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 98903:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 98904:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 98905:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 98906:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 98907:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 98908:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 98909:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 98910:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 98911:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 98912:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 98913:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 98914:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 98915:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 98916:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 98917:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 98918:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 98919:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 98920:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 98921:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 98922:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 98923:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 98924:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 98925:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 98926:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 98927:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 98928:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 98929:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 98930:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 98931:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 98932:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 98933:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 98934:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 98935:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 98936:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 98937:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 98938:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 98939:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 98940:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 98941:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 98942:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 98943:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 98944:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 98945:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 98946:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 98947:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 98948:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 98949:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 98950:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 98951:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 98952:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 98953:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 98954:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 98955:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 98956:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 98957:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 98958:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 98959:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 98960:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 98961:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 98962:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 98963:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 98964:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 98965:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 98966:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 98967:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 98968:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 98969:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 98970:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 98971:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 98972:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 98973:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 98974:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 98975:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 98976:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 98977:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 98978:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 98979:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 98980:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 98981:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 98982:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 98983:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 98984:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 98985:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 98986:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 98987:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 98988:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 98989:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 98990:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 98991:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 98992:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 98993:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 98994:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 98995:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 98996:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 98997:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 98998:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 98999:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 99000:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 99001:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 99002:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 99003:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 99004:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 99005:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 99006:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 99007:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 99008:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 99009:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 99010:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 99011:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 99012:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 99013:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 99014:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 99015:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 99016:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 99017:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 99018:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 99019:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 99020:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 99021:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 99022:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 99023:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 99024:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 99025:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 99026:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 99027:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 99028:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 99029:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 99030:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 99031:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 99032:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 99033:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 99034:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 99035:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 99036:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 99037:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 99038:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 99039:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 99040:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 99041:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 99042:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 99043:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 99044:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 99045:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 99046:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 99047:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 99048:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 99049:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 99050:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 99051:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 99052:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 99053:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 99054:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 99055:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 99056:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 99057:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 99058:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 99059:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 99060:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 99061:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 99062:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 99063:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 99064:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 99065:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 99066:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 99067:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 99068:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 99069:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 99070:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 99071:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 99072:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 99073:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 99074:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 99075:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 99076:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 99077:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 99078:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 99079:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 99080:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 99081:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 99082:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 99083:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 99084:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 99085:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 99086:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 99087:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 99088:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 99089:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 99090:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 99091:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 99092:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 99093:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 99094:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 99095:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 99096:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 99097:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 99098:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 99099:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 99100:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 99101:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 99102:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 99103:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 99104:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 99105:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 99106:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 99107:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 99108:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 99109:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 99110:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 99111:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 99112:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 99113:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 99114:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 99115:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 99116:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 99117:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 99118:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 99119:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 99120:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 99121:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 99122:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 99123:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 99124:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 99125:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 99126:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 99127:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 99128:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 99129:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 99130:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 99131:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 99132:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 99133:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 99134:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 99135:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 99136:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 99137:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 99138:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 99139:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 99140:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 99141:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 99142:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 99143:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 99144:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 99145:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 99146:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 99147:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 99148:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 99149:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 99150:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 99151:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 99152:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 99153:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 99154:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 99155:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 99156:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 99157:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 99158:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 99159:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 99160:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 99161:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 99162:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 99163:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 99164:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 99165:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 99166:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 99167:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 99168:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 99169:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 99170:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 99171:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 99172:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 99173:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 99174:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 99175:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 99176:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 99177:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 99178:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 99179:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 99180:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 99181:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 99182:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 99183:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 99184:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 99185:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 99186:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 99187:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 99188:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 99189:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 99190:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 99191:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 99192:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 99193:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 99194:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 99195:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 99196:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 99197:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 99198:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 99199:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 99200:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 99201:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 99202:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 99203:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 99204:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 99205:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 99206:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 99207:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 99208:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 99209:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 99210:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 99211:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 99212:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 99213:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 99214:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 99215:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 99216:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 99217:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 99218:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 99219:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 99220:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 99221:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 99222:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 99223:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 99224:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 99225:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 99226:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 99227:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 99228:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 99229:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 99230:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 99231:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 99232:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 99233:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 99234:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 99235:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 99236:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 99237:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 99238:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 99239:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 99240:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 99241:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 99242:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 99243:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 99244:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 99245:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 99246:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 99247:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 99248:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 99249:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 99250:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 99251:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 99252:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 99253:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 99254:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 99255:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 99256:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 99257:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 99258:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 99259:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 99260:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 99261:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 99262:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 99263:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 99264:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 99265:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 99266:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 99267:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 99268:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 99269:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 99270:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 99271:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 99272:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 99273:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 99274:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 99275:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 99276:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 99277:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 99278:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 99279:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 99280:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 99281:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 99282:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 99283:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 99284:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 99285:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 99286:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 99287:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 99288:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 99289:22]
  assign io_z = ~x100; // @[Snxn100k.scala 99290:17]
endmodule
module SnxnLv3Inst46(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst184_io_a; // @[Snxn100k.scala 28167:35]
  wire  inst_SnxnLv4Inst184_io_b; // @[Snxn100k.scala 28167:35]
  wire  inst_SnxnLv4Inst184_io_z; // @[Snxn100k.scala 28167:35]
  wire  inst_SnxnLv4Inst185_io_a; // @[Snxn100k.scala 28171:35]
  wire  inst_SnxnLv4Inst185_io_b; // @[Snxn100k.scala 28171:35]
  wire  inst_SnxnLv4Inst185_io_z; // @[Snxn100k.scala 28171:35]
  wire  inst_SnxnLv4Inst186_io_a; // @[Snxn100k.scala 28175:35]
  wire  inst_SnxnLv4Inst186_io_b; // @[Snxn100k.scala 28175:35]
  wire  inst_SnxnLv4Inst186_io_z; // @[Snxn100k.scala 28175:35]
  wire  inst_SnxnLv4Inst187_io_a; // @[Snxn100k.scala 28179:35]
  wire  inst_SnxnLv4Inst187_io_b; // @[Snxn100k.scala 28179:35]
  wire  inst_SnxnLv4Inst187_io_z; // @[Snxn100k.scala 28179:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst184_io_z + inst_SnxnLv4Inst185_io_z; // @[Snxn100k.scala 28183:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst186_io_z; // @[Snxn100k.scala 28183:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst187_io_z; // @[Snxn100k.scala 28183:92]
  SnxnLv4Inst184 inst_SnxnLv4Inst184 ( // @[Snxn100k.scala 28167:35]
    .io_a(inst_SnxnLv4Inst184_io_a),
    .io_b(inst_SnxnLv4Inst184_io_b),
    .io_z(inst_SnxnLv4Inst184_io_z)
  );
  SnxnLv4Inst58 inst_SnxnLv4Inst185 ( // @[Snxn100k.scala 28171:35]
    .io_a(inst_SnxnLv4Inst185_io_a),
    .io_b(inst_SnxnLv4Inst185_io_b),
    .io_z(inst_SnxnLv4Inst185_io_z)
  );
  SnxnLv4Inst76 inst_SnxnLv4Inst186 ( // @[Snxn100k.scala 28175:35]
    .io_a(inst_SnxnLv4Inst186_io_a),
    .io_b(inst_SnxnLv4Inst186_io_b),
    .io_z(inst_SnxnLv4Inst186_io_z)
  );
  SnxnLv4Inst74 inst_SnxnLv4Inst187 ( // @[Snxn100k.scala 28179:35]
    .io_a(inst_SnxnLv4Inst187_io_a),
    .io_b(inst_SnxnLv4Inst187_io_b),
    .io_z(inst_SnxnLv4Inst187_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 28184:15]
  assign inst_SnxnLv4Inst184_io_a = io_a; // @[Snxn100k.scala 28168:28]
  assign inst_SnxnLv4Inst184_io_b = io_b; // @[Snxn100k.scala 28169:28]
  assign inst_SnxnLv4Inst185_io_a = io_a; // @[Snxn100k.scala 28172:28]
  assign inst_SnxnLv4Inst185_io_b = io_b; // @[Snxn100k.scala 28173:28]
  assign inst_SnxnLv4Inst186_io_a = io_a; // @[Snxn100k.scala 28176:28]
  assign inst_SnxnLv4Inst186_io_b = io_b; // @[Snxn100k.scala 28177:28]
  assign inst_SnxnLv4Inst187_io_a = io_a; // @[Snxn100k.scala 28180:28]
  assign inst_SnxnLv4Inst187_io_b = io_b; // @[Snxn100k.scala 28181:28]
endmodule
module SnxnLv4Inst189(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 94193:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 94194:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 94195:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 94196:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 94197:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 94198:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 94199:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 94200:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 94201:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 94202:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 94203:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 94204:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 94205:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 94206:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 94207:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 94208:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 94209:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 94210:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 94211:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 94212:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 94213:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 94214:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 94215:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 94216:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 94217:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 94218:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 94219:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 94220:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 94221:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 94222:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 94223:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 94224:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 94225:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 94226:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 94227:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 94228:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 94229:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 94230:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 94231:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 94232:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 94233:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 94234:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 94235:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 94236:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 94237:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 94238:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 94239:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 94240:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 94241:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 94242:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 94243:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 94244:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 94245:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 94246:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 94247:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 94248:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 94249:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 94250:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 94251:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 94252:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 94253:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 94254:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 94255:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 94256:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 94257:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 94258:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 94259:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 94260:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 94261:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 94262:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 94263:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 94264:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 94265:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 94266:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 94267:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 94268:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 94269:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 94270:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 94271:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 94272:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 94273:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 94274:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 94275:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 94276:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 94277:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 94278:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 94279:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 94280:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 94281:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 94282:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 94283:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 94284:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 94285:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 94286:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 94287:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 94288:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 94289:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 94290:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 94291:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 94292:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 94293:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 94294:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 94295:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 94296:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 94297:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 94298:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 94299:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 94300:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 94301:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 94302:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 94303:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 94304:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 94305:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 94306:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 94307:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 94308:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 94309:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 94310:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 94311:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 94312:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 94313:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 94314:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 94315:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 94316:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 94317:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 94318:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 94319:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 94320:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 94321:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 94322:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 94323:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 94324:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 94325:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 94326:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 94327:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 94328:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 94329:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 94330:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 94331:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 94332:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 94333:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 94334:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 94335:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 94336:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 94337:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 94338:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 94339:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 94340:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 94341:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 94342:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 94343:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 94344:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 94345:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 94346:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 94347:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 94348:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 94349:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 94350:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 94351:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 94352:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 94353:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 94354:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 94355:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 94356:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 94357:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 94358:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 94359:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 94360:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 94361:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 94362:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 94363:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 94364:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 94365:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 94366:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 94367:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 94368:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 94369:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 94370:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 94371:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 94372:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 94373:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 94374:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 94375:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 94376:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 94377:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 94378:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 94379:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 94380:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 94381:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 94382:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 94383:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 94384:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 94385:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 94386:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 94387:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 94388:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 94389:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 94390:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 94391:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 94392:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 94393:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 94394:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 94395:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 94396:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 94397:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 94398:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 94399:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 94400:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 94401:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 94402:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 94403:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 94404:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 94405:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 94406:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 94407:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 94408:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 94409:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 94410:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 94411:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 94412:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 94413:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 94414:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 94415:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 94416:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 94417:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 94418:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 94419:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 94420:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 94421:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 94422:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 94423:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 94424:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 94425:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 94426:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 94427:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 94428:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 94429:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 94430:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 94431:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 94432:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 94433:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 94434:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 94435:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 94436:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 94437:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 94438:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 94439:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 94440:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 94441:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 94442:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 94443:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 94444:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 94445:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 94446:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 94447:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 94448:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 94449:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 94450:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 94451:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 94452:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 94453:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 94454:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 94455:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 94456:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 94457:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 94458:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 94459:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 94460:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 94461:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 94462:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 94463:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 94464:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 94465:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 94466:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 94467:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 94468:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 94469:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 94470:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 94471:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 94472:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 94473:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 94474:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 94475:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 94476:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 94477:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 94478:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 94479:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 94480:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 94481:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 94482:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 94483:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 94484:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 94485:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 94486:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 94487:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 94488:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 94489:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 94490:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 94491:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 94492:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 94493:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 94494:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 94495:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 94496:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 94497:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 94498:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 94499:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 94500:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 94501:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 94502:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 94503:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 94504:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 94505:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 94506:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 94507:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 94508:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 94509:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 94510:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 94511:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 94512:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 94513:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 94514:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 94515:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 94516:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 94517:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 94518:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 94519:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 94520:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 94521:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 94522:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 94523:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 94524:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 94525:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 94526:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 94527:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 94528:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 94529:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 94530:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 94531:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 94532:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 94533:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 94534:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 94535:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 94536:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 94537:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 94538:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 94539:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 94540:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 94541:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 94542:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 94543:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 94544:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 94545:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 94546:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 94547:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 94548:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 94549:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 94550:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 94551:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 94552:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 94553:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 94554:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 94555:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 94556:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 94557:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 94558:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 94559:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 94560:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 94561:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 94562:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 94563:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 94564:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 94565:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 94566:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 94567:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 94568:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 94569:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 94570:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 94571:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 94572:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 94573:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 94574:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 94575:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 94576:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 94577:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 94578:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 94579:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 94580:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 94581:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 94582:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 94583:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 94584:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 94585:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 94586:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 94587:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 94588:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 94589:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 94590:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 94591:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 94592:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 94593:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 94594:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 94595:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 94596:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 94597:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 94598:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 94599:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 94600:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 94601:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 94602:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 94603:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 94604:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 94605:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 94606:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 94607:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 94608:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 94609:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 94610:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 94611:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 94612:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 94613:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 94614:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 94615:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 94616:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 94617:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 94618:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 94619:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 94620:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 94621:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 94622:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 94623:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 94624:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 94625:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 94626:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 94627:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 94628:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 94629:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 94630:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 94631:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 94632:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 94633:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 94634:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 94635:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 94636:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 94637:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 94638:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 94639:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 94640:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 94641:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 94642:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 94643:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 94644:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 94645:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 94646:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 94647:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 94648:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 94649:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 94650:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 94651:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 94652:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 94653:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 94654:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 94655:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 94656:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 94657:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 94658:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 94659:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 94660:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 94661:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 94662:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 94663:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 94664:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 94665:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 94666:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 94667:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 94668:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 94669:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 94670:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 94671:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 94672:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 94673:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 94674:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 94675:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 94676:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 94677:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 94678:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 94679:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 94680:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 94681:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 94682:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 94683:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 94684:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 94685:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 94686:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 94687:22]
  assign io_z = ~x123; // @[Snxn100k.scala 94688:17]
endmodule
module SnxnLv3Inst47(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst188_io_a; // @[Snxn100k.scala 27258:35]
  wire  inst_SnxnLv4Inst188_io_b; // @[Snxn100k.scala 27258:35]
  wire  inst_SnxnLv4Inst188_io_z; // @[Snxn100k.scala 27258:35]
  wire  inst_SnxnLv4Inst189_io_a; // @[Snxn100k.scala 27262:35]
  wire  inst_SnxnLv4Inst189_io_b; // @[Snxn100k.scala 27262:35]
  wire  inst_SnxnLv4Inst189_io_z; // @[Snxn100k.scala 27262:35]
  wire  inst_SnxnLv4Inst190_io_a; // @[Snxn100k.scala 27266:35]
  wire  inst_SnxnLv4Inst190_io_b; // @[Snxn100k.scala 27266:35]
  wire  inst_SnxnLv4Inst190_io_z; // @[Snxn100k.scala 27266:35]
  wire  inst_SnxnLv4Inst191_io_a; // @[Snxn100k.scala 27270:35]
  wire  inst_SnxnLv4Inst191_io_b; // @[Snxn100k.scala 27270:35]
  wire  inst_SnxnLv4Inst191_io_z; // @[Snxn100k.scala 27270:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst188_io_z + inst_SnxnLv4Inst189_io_z; // @[Snxn100k.scala 27274:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst190_io_z; // @[Snxn100k.scala 27274:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst191_io_z; // @[Snxn100k.scala 27274:92]
  SnxnLv4Inst0 inst_SnxnLv4Inst188 ( // @[Snxn100k.scala 27258:35]
    .io_a(inst_SnxnLv4Inst188_io_a),
    .io_b(inst_SnxnLv4Inst188_io_b),
    .io_z(inst_SnxnLv4Inst188_io_z)
  );
  SnxnLv4Inst189 inst_SnxnLv4Inst189 ( // @[Snxn100k.scala 27262:35]
    .io_a(inst_SnxnLv4Inst189_io_a),
    .io_b(inst_SnxnLv4Inst189_io_b),
    .io_z(inst_SnxnLv4Inst189_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst190 ( // @[Snxn100k.scala 27266:35]
    .io_a(inst_SnxnLv4Inst190_io_a),
    .io_b(inst_SnxnLv4Inst190_io_b),
    .io_z(inst_SnxnLv4Inst190_io_z)
  );
  SnxnLv4Inst152 inst_SnxnLv4Inst191 ( // @[Snxn100k.scala 27270:35]
    .io_a(inst_SnxnLv4Inst191_io_a),
    .io_b(inst_SnxnLv4Inst191_io_b),
    .io_z(inst_SnxnLv4Inst191_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 27275:15]
  assign inst_SnxnLv4Inst188_io_a = io_a; // @[Snxn100k.scala 27259:28]
  assign inst_SnxnLv4Inst188_io_b = io_b; // @[Snxn100k.scala 27260:28]
  assign inst_SnxnLv4Inst189_io_a = io_a; // @[Snxn100k.scala 27263:28]
  assign inst_SnxnLv4Inst189_io_b = io_b; // @[Snxn100k.scala 27264:28]
  assign inst_SnxnLv4Inst190_io_a = io_a; // @[Snxn100k.scala 27267:28]
  assign inst_SnxnLv4Inst190_io_b = io_b; // @[Snxn100k.scala 27268:28]
  assign inst_SnxnLv4Inst191_io_a = io_a; // @[Snxn100k.scala 27271:28]
  assign inst_SnxnLv4Inst191_io_b = io_b; // @[Snxn100k.scala 27272:28]
endmodule
module SnxnLv2Inst11(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst44_io_a; // @[Snxn100k.scala 8306:34]
  wire  inst_SnxnLv3Inst44_io_b; // @[Snxn100k.scala 8306:34]
  wire  inst_SnxnLv3Inst44_io_z; // @[Snxn100k.scala 8306:34]
  wire  inst_SnxnLv3Inst45_io_a; // @[Snxn100k.scala 8310:34]
  wire  inst_SnxnLv3Inst45_io_b; // @[Snxn100k.scala 8310:34]
  wire  inst_SnxnLv3Inst45_io_z; // @[Snxn100k.scala 8310:34]
  wire  inst_SnxnLv3Inst46_io_a; // @[Snxn100k.scala 8314:34]
  wire  inst_SnxnLv3Inst46_io_b; // @[Snxn100k.scala 8314:34]
  wire  inst_SnxnLv3Inst46_io_z; // @[Snxn100k.scala 8314:34]
  wire  inst_SnxnLv3Inst47_io_a; // @[Snxn100k.scala 8318:34]
  wire  inst_SnxnLv3Inst47_io_b; // @[Snxn100k.scala 8318:34]
  wire  inst_SnxnLv3Inst47_io_z; // @[Snxn100k.scala 8318:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst44_io_z + inst_SnxnLv3Inst45_io_z; // @[Snxn100k.scala 8322:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst46_io_z; // @[Snxn100k.scala 8322:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst47_io_z; // @[Snxn100k.scala 8322:89]
  SnxnLv3Inst44 inst_SnxnLv3Inst44 ( // @[Snxn100k.scala 8306:34]
    .io_a(inst_SnxnLv3Inst44_io_a),
    .io_b(inst_SnxnLv3Inst44_io_b),
    .io_z(inst_SnxnLv3Inst44_io_z)
  );
  SnxnLv3Inst45 inst_SnxnLv3Inst45 ( // @[Snxn100k.scala 8310:34]
    .io_a(inst_SnxnLv3Inst45_io_a),
    .io_b(inst_SnxnLv3Inst45_io_b),
    .io_z(inst_SnxnLv3Inst45_io_z)
  );
  SnxnLv3Inst46 inst_SnxnLv3Inst46 ( // @[Snxn100k.scala 8314:34]
    .io_a(inst_SnxnLv3Inst46_io_a),
    .io_b(inst_SnxnLv3Inst46_io_b),
    .io_z(inst_SnxnLv3Inst46_io_z)
  );
  SnxnLv3Inst47 inst_SnxnLv3Inst47 ( // @[Snxn100k.scala 8318:34]
    .io_a(inst_SnxnLv3Inst47_io_a),
    .io_b(inst_SnxnLv3Inst47_io_b),
    .io_z(inst_SnxnLv3Inst47_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 8323:15]
  assign inst_SnxnLv3Inst44_io_a = io_a; // @[Snxn100k.scala 8307:27]
  assign inst_SnxnLv3Inst44_io_b = io_b; // @[Snxn100k.scala 8308:27]
  assign inst_SnxnLv3Inst45_io_a = io_a; // @[Snxn100k.scala 8311:27]
  assign inst_SnxnLv3Inst45_io_b = io_b; // @[Snxn100k.scala 8312:27]
  assign inst_SnxnLv3Inst46_io_a = io_a; // @[Snxn100k.scala 8315:27]
  assign inst_SnxnLv3Inst46_io_b = io_b; // @[Snxn100k.scala 8316:27]
  assign inst_SnxnLv3Inst47_io_a = io_a; // @[Snxn100k.scala 8319:27]
  assign inst_SnxnLv3Inst47_io_b = io_b; // @[Snxn100k.scala 8320:27]
endmodule
module SnxnLv1Inst2(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst8_io_a; // @[Snxn100k.scala 1585:33]
  wire  inst_SnxnLv2Inst8_io_b; // @[Snxn100k.scala 1585:33]
  wire  inst_SnxnLv2Inst8_io_z; // @[Snxn100k.scala 1585:33]
  wire  inst_SnxnLv2Inst9_io_a; // @[Snxn100k.scala 1589:33]
  wire  inst_SnxnLv2Inst9_io_b; // @[Snxn100k.scala 1589:33]
  wire  inst_SnxnLv2Inst9_io_z; // @[Snxn100k.scala 1589:33]
  wire  inst_SnxnLv2Inst10_io_a; // @[Snxn100k.scala 1593:34]
  wire  inst_SnxnLv2Inst10_io_b; // @[Snxn100k.scala 1593:34]
  wire  inst_SnxnLv2Inst10_io_z; // @[Snxn100k.scala 1593:34]
  wire  inst_SnxnLv2Inst11_io_a; // @[Snxn100k.scala 1597:34]
  wire  inst_SnxnLv2Inst11_io_b; // @[Snxn100k.scala 1597:34]
  wire  inst_SnxnLv2Inst11_io_z; // @[Snxn100k.scala 1597:34]
  wire  _sum_T_1 = inst_SnxnLv2Inst8_io_z + inst_SnxnLv2Inst9_io_z; // @[Snxn100k.scala 1601:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst10_io_z; // @[Snxn100k.scala 1601:61]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst11_io_z; // @[Snxn100k.scala 1601:87]
  SnxnLv2Inst8 inst_SnxnLv2Inst8 ( // @[Snxn100k.scala 1585:33]
    .io_a(inst_SnxnLv2Inst8_io_a),
    .io_b(inst_SnxnLv2Inst8_io_b),
    .io_z(inst_SnxnLv2Inst8_io_z)
  );
  SnxnLv2Inst9 inst_SnxnLv2Inst9 ( // @[Snxn100k.scala 1589:33]
    .io_a(inst_SnxnLv2Inst9_io_a),
    .io_b(inst_SnxnLv2Inst9_io_b),
    .io_z(inst_SnxnLv2Inst9_io_z)
  );
  SnxnLv2Inst10 inst_SnxnLv2Inst10 ( // @[Snxn100k.scala 1593:34]
    .io_a(inst_SnxnLv2Inst10_io_a),
    .io_b(inst_SnxnLv2Inst10_io_b),
    .io_z(inst_SnxnLv2Inst10_io_z)
  );
  SnxnLv2Inst11 inst_SnxnLv2Inst11 ( // @[Snxn100k.scala 1597:34]
    .io_a(inst_SnxnLv2Inst11_io_a),
    .io_b(inst_SnxnLv2Inst11_io_b),
    .io_z(inst_SnxnLv2Inst11_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 1602:15]
  assign inst_SnxnLv2Inst8_io_a = io_a; // @[Snxn100k.scala 1586:26]
  assign inst_SnxnLv2Inst8_io_b = io_b; // @[Snxn100k.scala 1587:26]
  assign inst_SnxnLv2Inst9_io_a = io_a; // @[Snxn100k.scala 1590:26]
  assign inst_SnxnLv2Inst9_io_b = io_b; // @[Snxn100k.scala 1591:26]
  assign inst_SnxnLv2Inst10_io_a = io_a; // @[Snxn100k.scala 1594:27]
  assign inst_SnxnLv2Inst10_io_b = io_b; // @[Snxn100k.scala 1595:27]
  assign inst_SnxnLv2Inst11_io_a = io_a; // @[Snxn100k.scala 1598:27]
  assign inst_SnxnLv2Inst11_io_b = io_b; // @[Snxn100k.scala 1599:27]
endmodule
module SnxnLv3Inst48(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst192_io_a; // @[Snxn100k.scala 17621:35]
  wire  inst_SnxnLv4Inst192_io_b; // @[Snxn100k.scala 17621:35]
  wire  inst_SnxnLv4Inst192_io_z; // @[Snxn100k.scala 17621:35]
  wire  inst_SnxnLv4Inst193_io_a; // @[Snxn100k.scala 17625:35]
  wire  inst_SnxnLv4Inst193_io_b; // @[Snxn100k.scala 17625:35]
  wire  inst_SnxnLv4Inst193_io_z; // @[Snxn100k.scala 17625:35]
  wire  inst_SnxnLv4Inst194_io_a; // @[Snxn100k.scala 17629:35]
  wire  inst_SnxnLv4Inst194_io_b; // @[Snxn100k.scala 17629:35]
  wire  inst_SnxnLv4Inst194_io_z; // @[Snxn100k.scala 17629:35]
  wire  inst_SnxnLv4Inst195_io_a; // @[Snxn100k.scala 17633:35]
  wire  inst_SnxnLv4Inst195_io_b; // @[Snxn100k.scala 17633:35]
  wire  inst_SnxnLv4Inst195_io_z; // @[Snxn100k.scala 17633:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst192_io_z + inst_SnxnLv4Inst193_io_z; // @[Snxn100k.scala 17637:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst194_io_z; // @[Snxn100k.scala 17637:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst195_io_z; // @[Snxn100k.scala 17637:92]
  SnxnLv4Inst0 inst_SnxnLv4Inst192 ( // @[Snxn100k.scala 17621:35]
    .io_a(inst_SnxnLv4Inst192_io_a),
    .io_b(inst_SnxnLv4Inst192_io_b),
    .io_z(inst_SnxnLv4Inst192_io_z)
  );
  SnxnLv4Inst17 inst_SnxnLv4Inst193 ( // @[Snxn100k.scala 17625:35]
    .io_a(inst_SnxnLv4Inst193_io_a),
    .io_b(inst_SnxnLv4Inst193_io_b),
    .io_z(inst_SnxnLv4Inst193_io_z)
  );
  SnxnLv4Inst32 inst_SnxnLv4Inst194 ( // @[Snxn100k.scala 17629:35]
    .io_a(inst_SnxnLv4Inst194_io_a),
    .io_b(inst_SnxnLv4Inst194_io_b),
    .io_z(inst_SnxnLv4Inst194_io_z)
  );
  SnxnLv4Inst32 inst_SnxnLv4Inst195 ( // @[Snxn100k.scala 17633:35]
    .io_a(inst_SnxnLv4Inst195_io_a),
    .io_b(inst_SnxnLv4Inst195_io_b),
    .io_z(inst_SnxnLv4Inst195_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17638:15]
  assign inst_SnxnLv4Inst192_io_a = io_a; // @[Snxn100k.scala 17622:28]
  assign inst_SnxnLv4Inst192_io_b = io_b; // @[Snxn100k.scala 17623:28]
  assign inst_SnxnLv4Inst193_io_a = io_a; // @[Snxn100k.scala 17626:28]
  assign inst_SnxnLv4Inst193_io_b = io_b; // @[Snxn100k.scala 17627:28]
  assign inst_SnxnLv4Inst194_io_a = io_a; // @[Snxn100k.scala 17630:28]
  assign inst_SnxnLv4Inst194_io_b = io_b; // @[Snxn100k.scala 17631:28]
  assign inst_SnxnLv4Inst195_io_a = io_a; // @[Snxn100k.scala 17634:28]
  assign inst_SnxnLv4Inst195_io_b = io_b; // @[Snxn100k.scala 17635:28]
endmodule
module SnxnLv4Inst197(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 58245:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 58246:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 58247:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 58248:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 58249:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 58250:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 58251:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 58252:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 58253:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 58254:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 58255:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 58256:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 58257:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 58258:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 58259:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 58260:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 58261:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 58262:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 58263:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 58264:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 58265:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 58266:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 58267:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 58268:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 58269:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 58270:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 58271:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 58272:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 58273:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 58274:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 58275:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 58276:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 58277:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 58278:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 58279:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 58280:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 58281:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 58282:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 58283:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 58284:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 58285:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 58286:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 58287:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 58288:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 58289:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 58290:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 58291:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 58292:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 58293:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 58294:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 58295:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 58296:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 58297:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 58298:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 58299:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 58300:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 58301:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 58302:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 58303:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 58304:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 58305:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 58306:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 58307:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 58308:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 58309:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 58310:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 58311:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 58312:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 58313:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 58314:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 58315:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 58316:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 58317:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 58318:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 58319:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 58320:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 58321:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 58322:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 58323:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 58324:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 58325:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 58326:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 58327:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 58328:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 58329:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 58330:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 58331:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 58332:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 58333:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 58334:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 58335:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 58336:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 58337:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 58338:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 58339:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 58340:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 58341:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 58342:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 58343:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 58344:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 58345:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 58346:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 58347:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 58348:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 58349:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 58350:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 58351:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 58352:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 58353:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 58354:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 58355:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 58356:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 58357:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 58358:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 58359:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 58360:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 58361:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 58362:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 58363:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 58364:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 58365:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 58366:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 58367:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 58368:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 58369:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 58370:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 58371:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 58372:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 58373:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 58374:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 58375:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 58376:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 58377:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 58378:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 58379:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 58380:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 58381:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 58382:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 58383:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 58384:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 58385:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 58386:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 58387:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 58388:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 58389:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 58390:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 58391:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 58392:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 58393:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 58394:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 58395:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 58396:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 58397:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 58398:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 58399:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 58400:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 58401:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 58402:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 58403:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 58404:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 58405:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 58406:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 58407:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 58408:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 58409:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 58410:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 58411:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 58412:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 58413:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 58414:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 58415:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 58416:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 58417:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 58418:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 58419:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 58420:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 58421:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 58422:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 58423:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 58424:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 58425:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 58426:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 58427:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 58428:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 58429:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 58430:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 58431:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 58432:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 58433:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 58434:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 58435:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 58436:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 58437:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 58438:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 58439:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 58440:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 58441:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 58442:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 58443:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 58444:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 58445:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 58446:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 58447:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 58448:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 58449:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 58450:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 58451:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 58452:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 58453:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 58454:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 58455:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 58456:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 58457:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 58458:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 58459:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 58460:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 58461:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 58462:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 58463:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 58464:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 58465:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 58466:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 58467:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 58468:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 58469:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 58470:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 58471:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 58472:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 58473:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 58474:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 58475:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 58476:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 58477:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 58478:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 58479:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 58480:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 58481:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 58482:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 58483:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 58484:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 58485:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 58486:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 58487:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 58488:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 58489:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 58490:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 58491:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 58492:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 58493:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 58494:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 58495:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 58496:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 58497:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 58498:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 58499:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 58500:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 58501:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 58502:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 58503:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 58504:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 58505:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 58506:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 58507:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 58508:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 58509:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 58510:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 58511:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 58512:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 58513:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 58514:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 58515:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 58516:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 58517:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 58518:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 58519:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 58520:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 58521:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 58522:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 58523:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 58524:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 58525:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 58526:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 58527:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 58528:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 58529:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 58530:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 58531:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 58532:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 58533:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 58534:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 58535:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 58536:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 58537:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 58538:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 58539:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 58540:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 58541:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 58542:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 58543:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 58544:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 58545:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 58546:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 58547:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 58548:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 58549:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 58550:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 58551:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 58552:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 58553:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 58554:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 58555:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 58556:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 58557:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 58558:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 58559:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 58560:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 58561:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 58562:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 58563:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 58564:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 58565:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 58566:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 58567:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 58568:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 58569:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 58570:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 58571:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 58572:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 58573:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 58574:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 58575:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 58576:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 58577:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 58578:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 58579:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 58580:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 58581:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 58582:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 58583:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 58584:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 58585:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 58586:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 58587:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 58588:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 58589:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 58590:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 58591:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 58592:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 58593:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 58594:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 58595:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 58596:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 58597:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 58598:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 58599:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 58600:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 58601:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 58602:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 58603:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 58604:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 58605:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 58606:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 58607:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 58608:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 58609:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 58610:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 58611:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 58612:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 58613:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 58614:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 58615:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 58616:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 58617:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 58618:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 58619:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 58620:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 58621:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 58622:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 58623:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 58624:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 58625:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 58626:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 58627:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 58628:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 58629:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 58630:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 58631:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 58632:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 58633:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 58634:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 58635:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 58636:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 58637:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 58638:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 58639:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 58640:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 58641:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 58642:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 58643:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 58644:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 58645:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 58646:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 58647:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 58648:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 58649:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 58650:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 58651:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 58652:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 58653:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 58654:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 58655:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 58656:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 58657:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 58658:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 58659:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 58660:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 58661:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 58662:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 58663:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 58664:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 58665:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 58666:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 58667:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 58668:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 58669:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 58670:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 58671:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 58672:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 58673:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 58674:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 58675:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 58676:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 58677:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 58678:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 58679:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 58680:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 58681:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 58682:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 58683:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 58684:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 58685:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 58686:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 58687:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 58688:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 58689:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 58690:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 58691:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 58692:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 58693:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 58694:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 58695:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 58696:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 58697:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 58698:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 58699:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 58700:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 58701:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 58702:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 58703:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 58704:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 58705:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 58706:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 58707:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 58708:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 58709:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 58710:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 58711:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 58712:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 58713:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 58714:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 58715:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 58716:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 58717:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 58718:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 58719:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 58720:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 58721:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 58722:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 58723:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 58724:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 58725:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 58726:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 58727:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 58728:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 58729:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 58730:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 58731:22]
  wire  invx121 = ~x121; // @[Snxn100k.scala 58732:17]
  wire  t122 = x121 + invx121; // @[Snxn100k.scala 58733:22]
  wire  inv122 = ~t122; // @[Snxn100k.scala 58734:17]
  wire  x122 = t122 ^ inv122; // @[Snxn100k.scala 58735:22]
  wire  invx122 = ~x122; // @[Snxn100k.scala 58736:17]
  wire  t123 = x122 + invx122; // @[Snxn100k.scala 58737:22]
  wire  inv123 = ~t123; // @[Snxn100k.scala 58738:17]
  wire  x123 = t123 ^ inv123; // @[Snxn100k.scala 58739:22]
  wire  invx123 = ~x123; // @[Snxn100k.scala 58740:17]
  wire  t124 = x123 + invx123; // @[Snxn100k.scala 58741:22]
  wire  inv124 = ~t124; // @[Snxn100k.scala 58742:17]
  wire  x124 = t124 ^ inv124; // @[Snxn100k.scala 58743:22]
  wire  invx124 = ~x124; // @[Snxn100k.scala 58744:17]
  wire  t125 = x124 + invx124; // @[Snxn100k.scala 58745:22]
  wire  inv125 = ~t125; // @[Snxn100k.scala 58746:17]
  wire  x125 = t125 ^ inv125; // @[Snxn100k.scala 58747:22]
  wire  invx125 = ~x125; // @[Snxn100k.scala 58748:17]
  wire  t126 = x125 + invx125; // @[Snxn100k.scala 58749:22]
  wire  inv126 = ~t126; // @[Snxn100k.scala 58750:17]
  wire  x126 = t126 ^ inv126; // @[Snxn100k.scala 58751:22]
  wire  invx126 = ~x126; // @[Snxn100k.scala 58752:17]
  wire  t127 = x126 + invx126; // @[Snxn100k.scala 58753:22]
  wire  inv127 = ~t127; // @[Snxn100k.scala 58754:17]
  wire  x127 = t127 ^ inv127; // @[Snxn100k.scala 58755:22]
  wire  invx127 = ~x127; // @[Snxn100k.scala 58756:17]
  wire  t128 = x127 + invx127; // @[Snxn100k.scala 58757:22]
  wire  inv128 = ~t128; // @[Snxn100k.scala 58758:17]
  wire  x128 = t128 ^ inv128; // @[Snxn100k.scala 58759:22]
  wire  invx128 = ~x128; // @[Snxn100k.scala 58760:17]
  wire  t129 = x128 + invx128; // @[Snxn100k.scala 58761:22]
  wire  inv129 = ~t129; // @[Snxn100k.scala 58762:17]
  wire  x129 = t129 ^ inv129; // @[Snxn100k.scala 58763:22]
  wire  invx129 = ~x129; // @[Snxn100k.scala 58764:17]
  wire  t130 = x129 + invx129; // @[Snxn100k.scala 58765:22]
  wire  inv130 = ~t130; // @[Snxn100k.scala 58766:17]
  wire  x130 = t130 ^ inv130; // @[Snxn100k.scala 58767:22]
  assign io_z = ~x130; // @[Snxn100k.scala 58768:17]
endmodule
module SnxnLv3Inst49(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst196_io_a; // @[Snxn100k.scala 17090:35]
  wire  inst_SnxnLv4Inst196_io_b; // @[Snxn100k.scala 17090:35]
  wire  inst_SnxnLv4Inst196_io_z; // @[Snxn100k.scala 17090:35]
  wire  inst_SnxnLv4Inst197_io_a; // @[Snxn100k.scala 17094:35]
  wire  inst_SnxnLv4Inst197_io_b; // @[Snxn100k.scala 17094:35]
  wire  inst_SnxnLv4Inst197_io_z; // @[Snxn100k.scala 17094:35]
  wire  inst_SnxnLv4Inst198_io_a; // @[Snxn100k.scala 17098:35]
  wire  inst_SnxnLv4Inst198_io_b; // @[Snxn100k.scala 17098:35]
  wire  inst_SnxnLv4Inst198_io_z; // @[Snxn100k.scala 17098:35]
  wire  inst_SnxnLv4Inst199_io_a; // @[Snxn100k.scala 17102:35]
  wire  inst_SnxnLv4Inst199_io_b; // @[Snxn100k.scala 17102:35]
  wire  inst_SnxnLv4Inst199_io_z; // @[Snxn100k.scala 17102:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst196_io_z + inst_SnxnLv4Inst197_io_z; // @[Snxn100k.scala 17106:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst198_io_z; // @[Snxn100k.scala 17106:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst199_io_z; // @[Snxn100k.scala 17106:92]
  SnxnLv4Inst36 inst_SnxnLv4Inst196 ( // @[Snxn100k.scala 17090:35]
    .io_a(inst_SnxnLv4Inst196_io_a),
    .io_b(inst_SnxnLv4Inst196_io_b),
    .io_z(inst_SnxnLv4Inst196_io_z)
  );
  SnxnLv4Inst197 inst_SnxnLv4Inst197 ( // @[Snxn100k.scala 17094:35]
    .io_a(inst_SnxnLv4Inst197_io_a),
    .io_b(inst_SnxnLv4Inst197_io_b),
    .io_z(inst_SnxnLv4Inst197_io_z)
  );
  SnxnLv4Inst1 inst_SnxnLv4Inst198 ( // @[Snxn100k.scala 17098:35]
    .io_a(inst_SnxnLv4Inst198_io_a),
    .io_b(inst_SnxnLv4Inst198_io_b),
    .io_z(inst_SnxnLv4Inst198_io_z)
  );
  SnxnLv4Inst56 inst_SnxnLv4Inst199 ( // @[Snxn100k.scala 17102:35]
    .io_a(inst_SnxnLv4Inst199_io_a),
    .io_b(inst_SnxnLv4Inst199_io_b),
    .io_z(inst_SnxnLv4Inst199_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17107:15]
  assign inst_SnxnLv4Inst196_io_a = io_a; // @[Snxn100k.scala 17091:28]
  assign inst_SnxnLv4Inst196_io_b = io_b; // @[Snxn100k.scala 17092:28]
  assign inst_SnxnLv4Inst197_io_a = io_a; // @[Snxn100k.scala 17095:28]
  assign inst_SnxnLv4Inst197_io_b = io_b; // @[Snxn100k.scala 17096:28]
  assign inst_SnxnLv4Inst198_io_a = io_a; // @[Snxn100k.scala 17099:28]
  assign inst_SnxnLv4Inst198_io_b = io_b; // @[Snxn100k.scala 17100:28]
  assign inst_SnxnLv4Inst199_io_a = io_a; // @[Snxn100k.scala 17103:28]
  assign inst_SnxnLv4Inst199_io_b = io_b; // @[Snxn100k.scala 17104:28]
endmodule
module SnxnLv4Inst200(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 56281:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 56282:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 56283:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 56284:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 56285:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 56286:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 56287:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 56288:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 56289:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 56290:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 56291:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 56292:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 56293:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 56294:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 56295:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 56296:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 56297:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 56298:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 56299:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 56300:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 56301:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 56302:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 56303:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 56304:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 56305:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 56306:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 56307:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 56308:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 56309:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 56310:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 56311:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 56312:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 56313:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 56314:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 56315:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 56316:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 56317:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 56318:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 56319:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 56320:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 56321:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 56322:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 56323:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 56324:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 56325:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 56326:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 56327:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 56328:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 56329:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 56330:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 56331:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 56332:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 56333:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 56334:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 56335:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 56336:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 56337:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 56338:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 56339:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 56340:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 56341:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 56342:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 56343:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 56344:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 56345:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 56346:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 56347:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 56348:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 56349:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 56350:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 56351:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 56352:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 56353:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 56354:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 56355:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 56356:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 56357:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 56358:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 56359:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 56360:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 56361:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 56362:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 56363:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 56364:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 56365:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 56366:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 56367:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 56368:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 56369:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 56370:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 56371:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 56372:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 56373:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 56374:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 56375:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 56376:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 56377:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 56378:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 56379:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 56380:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 56381:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 56382:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 56383:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 56384:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 56385:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 56386:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 56387:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 56388:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 56389:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 56390:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 56391:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 56392:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 56393:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 56394:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 56395:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 56396:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 56397:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 56398:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 56399:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 56400:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 56401:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 56402:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 56403:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 56404:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 56405:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 56406:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 56407:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 56408:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 56409:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 56410:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 56411:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 56412:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 56413:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 56414:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 56415:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 56416:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 56417:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 56418:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 56419:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 56420:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 56421:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 56422:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 56423:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 56424:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 56425:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 56426:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 56427:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 56428:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 56429:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 56430:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 56431:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 56432:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 56433:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 56434:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 56435:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 56436:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 56437:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 56438:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 56439:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 56440:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 56441:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 56442:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 56443:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 56444:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 56445:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 56446:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 56447:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 56448:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 56449:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 56450:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 56451:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 56452:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 56453:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 56454:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 56455:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 56456:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 56457:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 56458:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 56459:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 56460:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 56461:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 56462:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 56463:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 56464:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 56465:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 56466:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 56467:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 56468:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 56469:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 56470:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 56471:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 56472:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 56473:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 56474:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 56475:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 56476:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 56477:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 56478:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 56479:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 56480:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 56481:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 56482:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 56483:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 56484:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 56485:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 56486:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 56487:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 56488:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 56489:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 56490:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 56491:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 56492:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 56493:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 56494:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 56495:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 56496:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 56497:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 56498:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 56499:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 56500:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 56501:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 56502:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 56503:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 56504:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 56505:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 56506:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 56507:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 56508:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 56509:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 56510:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 56511:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 56512:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 56513:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 56514:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 56515:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 56516:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 56517:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 56518:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 56519:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 56520:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 56521:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 56522:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 56523:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 56524:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 56525:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 56526:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 56527:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 56528:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 56529:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 56530:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 56531:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 56532:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 56533:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 56534:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 56535:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 56536:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 56537:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 56538:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 56539:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 56540:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 56541:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 56542:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 56543:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 56544:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 56545:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 56546:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 56547:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 56548:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 56549:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 56550:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 56551:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 56552:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 56553:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 56554:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 56555:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 56556:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 56557:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 56558:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 56559:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 56560:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 56561:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 56562:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 56563:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 56564:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 56565:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 56566:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 56567:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 56568:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 56569:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 56570:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 56571:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 56572:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 56573:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 56574:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 56575:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 56576:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 56577:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 56578:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 56579:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 56580:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 56581:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 56582:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 56583:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 56584:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 56585:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 56586:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 56587:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 56588:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 56589:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 56590:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 56591:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 56592:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 56593:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 56594:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 56595:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 56596:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 56597:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 56598:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 56599:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 56600:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 56601:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 56602:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 56603:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 56604:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 56605:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 56606:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 56607:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 56608:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 56609:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 56610:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 56611:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 56612:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 56613:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 56614:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 56615:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 56616:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 56617:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 56618:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 56619:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 56620:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 56621:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 56622:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 56623:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 56624:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 56625:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 56626:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 56627:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 56628:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 56629:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 56630:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 56631:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 56632:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 56633:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 56634:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 56635:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 56636:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 56637:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 56638:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 56639:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 56640:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 56641:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 56642:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 56643:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 56644:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 56645:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 56646:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 56647:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 56648:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 56649:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 56650:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 56651:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 56652:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 56653:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 56654:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 56655:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 56656:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 56657:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 56658:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 56659:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 56660:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 56661:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 56662:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 56663:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 56664:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 56665:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 56666:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 56667:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 56668:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 56669:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 56670:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 56671:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 56672:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 56673:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 56674:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 56675:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 56676:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 56677:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 56678:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 56679:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 56680:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 56681:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 56682:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 56683:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 56684:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 56685:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 56686:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 56687:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 56688:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 56689:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 56690:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 56691:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 56692:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 56693:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 56694:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 56695:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 56696:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 56697:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 56698:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 56699:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 56700:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 56701:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 56702:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 56703:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 56704:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 56705:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 56706:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 56707:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 56708:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 56709:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 56710:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 56711:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 56712:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 56713:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 56714:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 56715:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 56716:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 56717:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 56718:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 56719:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 56720:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 56721:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 56722:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 56723:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 56724:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 56725:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 56726:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 56727:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 56728:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 56729:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 56730:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 56731:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 56732:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 56733:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 56734:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 56735:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 56736:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 56737:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 56738:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 56739:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 56740:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 56741:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 56742:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 56743:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 56744:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 56745:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 56746:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 56747:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 56748:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 56749:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 56750:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 56751:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 56752:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 56753:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 56754:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 56755:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 56756:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 56757:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 56758:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 56759:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 56760:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 56761:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 56762:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 56763:22]
  assign io_z = ~x120; // @[Snxn100k.scala 56764:17]
endmodule
module SnxnLv3Inst50(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst200_io_a; // @[Snxn100k.scala 16096:35]
  wire  inst_SnxnLv4Inst200_io_b; // @[Snxn100k.scala 16096:35]
  wire  inst_SnxnLv4Inst200_io_z; // @[Snxn100k.scala 16096:35]
  wire  inst_SnxnLv4Inst201_io_a; // @[Snxn100k.scala 16100:35]
  wire  inst_SnxnLv4Inst201_io_b; // @[Snxn100k.scala 16100:35]
  wire  inst_SnxnLv4Inst201_io_z; // @[Snxn100k.scala 16100:35]
  wire  inst_SnxnLv4Inst202_io_a; // @[Snxn100k.scala 16104:35]
  wire  inst_SnxnLv4Inst202_io_b; // @[Snxn100k.scala 16104:35]
  wire  inst_SnxnLv4Inst202_io_z; // @[Snxn100k.scala 16104:35]
  wire  inst_SnxnLv4Inst203_io_a; // @[Snxn100k.scala 16108:35]
  wire  inst_SnxnLv4Inst203_io_b; // @[Snxn100k.scala 16108:35]
  wire  inst_SnxnLv4Inst203_io_z; // @[Snxn100k.scala 16108:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst200_io_z + inst_SnxnLv4Inst201_io_z; // @[Snxn100k.scala 16112:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst202_io_z; // @[Snxn100k.scala 16112:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst203_io_z; // @[Snxn100k.scala 16112:92]
  SnxnLv4Inst200 inst_SnxnLv4Inst200 ( // @[Snxn100k.scala 16096:35]
    .io_a(inst_SnxnLv4Inst200_io_a),
    .io_b(inst_SnxnLv4Inst200_io_b),
    .io_z(inst_SnxnLv4Inst200_io_z)
  );
  SnxnLv4Inst77 inst_SnxnLv4Inst201 ( // @[Snxn100k.scala 16100:35]
    .io_a(inst_SnxnLv4Inst201_io_a),
    .io_b(inst_SnxnLv4Inst201_io_b),
    .io_z(inst_SnxnLv4Inst201_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst202 ( // @[Snxn100k.scala 16104:35]
    .io_a(inst_SnxnLv4Inst202_io_a),
    .io_b(inst_SnxnLv4Inst202_io_b),
    .io_z(inst_SnxnLv4Inst202_io_z)
  );
  SnxnLv4Inst171 inst_SnxnLv4Inst203 ( // @[Snxn100k.scala 16108:35]
    .io_a(inst_SnxnLv4Inst203_io_a),
    .io_b(inst_SnxnLv4Inst203_io_b),
    .io_z(inst_SnxnLv4Inst203_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 16113:15]
  assign inst_SnxnLv4Inst200_io_a = io_a; // @[Snxn100k.scala 16097:28]
  assign inst_SnxnLv4Inst200_io_b = io_b; // @[Snxn100k.scala 16098:28]
  assign inst_SnxnLv4Inst201_io_a = io_a; // @[Snxn100k.scala 16101:28]
  assign inst_SnxnLv4Inst201_io_b = io_b; // @[Snxn100k.scala 16102:28]
  assign inst_SnxnLv4Inst202_io_a = io_a; // @[Snxn100k.scala 16105:28]
  assign inst_SnxnLv4Inst202_io_b = io_b; // @[Snxn100k.scala 16106:28]
  assign inst_SnxnLv4Inst203_io_a = io_a; // @[Snxn100k.scala 16109:28]
  assign inst_SnxnLv4Inst203_io_b = io_b; // @[Snxn100k.scala 16110:28]
endmodule
module SnxnLv4Inst204(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 57795:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 57796:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 57797:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 57798:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 57799:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 57800:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 57801:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 57802:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 57803:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 57804:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 57805:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 57806:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 57807:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 57808:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 57809:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 57810:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 57811:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 57812:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 57813:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 57814:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 57815:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 57816:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 57817:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 57818:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 57819:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 57820:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 57821:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 57822:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 57823:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 57824:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 57825:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 57826:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 57827:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 57828:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 57829:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 57830:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 57831:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 57832:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 57833:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 57834:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 57835:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 57836:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 57837:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 57838:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 57839:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 57840:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 57841:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 57842:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 57843:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 57844:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 57845:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 57846:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 57847:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 57848:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 57849:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 57850:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 57851:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 57852:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 57853:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 57854:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 57855:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 57856:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 57857:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 57858:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 57859:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 57860:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 57861:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 57862:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 57863:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 57864:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 57865:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 57866:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 57867:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 57868:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 57869:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 57870:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 57871:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 57872:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 57873:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 57874:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 57875:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 57876:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 57877:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 57878:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 57879:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 57880:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 57881:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 57882:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 57883:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 57884:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 57885:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 57886:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 57887:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 57888:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 57889:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 57890:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 57891:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 57892:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 57893:20]
  assign io_z = ~x24; // @[Snxn100k.scala 57894:16]
endmodule
module SnxnLv4Inst207(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 57335:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 57336:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 57337:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 57338:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 57339:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 57340:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 57341:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 57342:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 57343:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 57344:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 57345:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 57346:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 57347:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 57348:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 57349:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 57350:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 57351:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 57352:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 57353:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 57354:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 57355:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 57356:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 57357:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 57358:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 57359:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 57360:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 57361:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 57362:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 57363:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 57364:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 57365:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 57366:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 57367:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 57368:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 57369:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 57370:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 57371:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 57372:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 57373:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 57374:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 57375:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 57376:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 57377:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 57378:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 57379:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 57380:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 57381:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 57382:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 57383:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 57384:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 57385:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 57386:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 57387:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 57388:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 57389:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 57390:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 57391:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 57392:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 57393:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 57394:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 57395:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 57396:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 57397:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 57398:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 57399:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 57400:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 57401:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 57402:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 57403:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 57404:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 57405:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 57406:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 57407:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 57408:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 57409:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 57410:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 57411:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 57412:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 57413:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 57414:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 57415:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 57416:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 57417:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 57418:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 57419:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 57420:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 57421:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 57422:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 57423:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 57424:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 57425:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 57426:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 57427:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 57428:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 57429:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 57430:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 57431:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 57432:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 57433:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 57434:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 57435:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 57436:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 57437:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 57438:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 57439:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 57440:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 57441:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 57442:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 57443:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 57444:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 57445:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 57446:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 57447:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 57448:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 57449:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 57450:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 57451:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 57452:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 57453:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 57454:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 57455:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 57456:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 57457:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 57458:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 57459:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 57460:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 57461:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 57462:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 57463:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 57464:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 57465:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 57466:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 57467:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 57468:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 57469:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 57470:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 57471:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 57472:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 57473:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 57474:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 57475:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 57476:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 57477:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 57478:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 57479:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 57480:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 57481:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 57482:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 57483:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 57484:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 57485:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 57486:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 57487:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 57488:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 57489:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 57490:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 57491:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 57492:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 57493:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 57494:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 57495:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 57496:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 57497:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 57498:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 57499:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 57500:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 57501:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 57502:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 57503:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 57504:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 57505:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 57506:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 57507:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 57508:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 57509:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 57510:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 57511:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 57512:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 57513:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 57514:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 57515:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 57516:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 57517:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 57518:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 57519:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 57520:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 57521:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 57522:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 57523:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 57524:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 57525:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 57526:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 57527:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 57528:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 57529:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 57530:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 57531:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 57532:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 57533:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 57534:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 57535:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 57536:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 57537:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 57538:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 57539:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 57540:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 57541:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 57542:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 57543:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 57544:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 57545:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 57546:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 57547:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 57548:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 57549:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 57550:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 57551:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 57552:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 57553:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 57554:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 57555:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 57556:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 57557:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 57558:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 57559:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 57560:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 57561:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 57562:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 57563:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 57564:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 57565:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 57566:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 57567:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 57568:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 57569:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 57570:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 57571:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 57572:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 57573:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 57574:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 57575:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 57576:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 57577:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 57578:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 57579:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 57580:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 57581:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 57582:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 57583:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 57584:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 57585:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 57586:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 57587:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 57588:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 57589:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 57590:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 57591:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 57592:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 57593:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 57594:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 57595:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 57596:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 57597:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 57598:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 57599:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 57600:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 57601:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 57602:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 57603:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 57604:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 57605:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 57606:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 57607:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 57608:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 57609:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 57610:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 57611:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 57612:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 57613:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 57614:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 57615:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 57616:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 57617:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 57618:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 57619:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 57620:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 57621:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 57622:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 57623:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 57624:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 57625:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 57626:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 57627:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 57628:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 57629:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 57630:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 57631:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 57632:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 57633:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 57634:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 57635:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 57636:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 57637:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 57638:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 57639:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 57640:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 57641:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 57642:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 57643:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 57644:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 57645:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 57646:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 57647:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 57648:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 57649:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 57650:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 57651:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 57652:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 57653:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 57654:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 57655:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 57656:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 57657:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 57658:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 57659:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 57660:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 57661:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 57662:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 57663:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 57664:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 57665:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 57666:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 57667:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 57668:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 57669:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 57670:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 57671:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 57672:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 57673:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 57674:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 57675:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 57676:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 57677:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 57678:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 57679:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 57680:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 57681:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 57682:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 57683:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 57684:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 57685:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 57686:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 57687:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 57688:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 57689:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 57690:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 57691:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 57692:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 57693:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 57694:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 57695:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 57696:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 57697:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 57698:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 57699:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 57700:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 57701:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 57702:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 57703:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 57704:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 57705:20]
  assign io_z = ~x92; // @[Snxn100k.scala 57706:16]
endmodule
module SnxnLv3Inst51(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst204_io_a; // @[Snxn100k.scala 16575:35]
  wire  inst_SnxnLv4Inst204_io_b; // @[Snxn100k.scala 16575:35]
  wire  inst_SnxnLv4Inst204_io_z; // @[Snxn100k.scala 16575:35]
  wire  inst_SnxnLv4Inst205_io_a; // @[Snxn100k.scala 16579:35]
  wire  inst_SnxnLv4Inst205_io_b; // @[Snxn100k.scala 16579:35]
  wire  inst_SnxnLv4Inst205_io_z; // @[Snxn100k.scala 16579:35]
  wire  inst_SnxnLv4Inst206_io_a; // @[Snxn100k.scala 16583:35]
  wire  inst_SnxnLv4Inst206_io_b; // @[Snxn100k.scala 16583:35]
  wire  inst_SnxnLv4Inst206_io_z; // @[Snxn100k.scala 16583:35]
  wire  inst_SnxnLv4Inst207_io_a; // @[Snxn100k.scala 16587:35]
  wire  inst_SnxnLv4Inst207_io_b; // @[Snxn100k.scala 16587:35]
  wire  inst_SnxnLv4Inst207_io_z; // @[Snxn100k.scala 16587:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst204_io_z + inst_SnxnLv4Inst205_io_z; // @[Snxn100k.scala 16591:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst206_io_z; // @[Snxn100k.scala 16591:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst207_io_z; // @[Snxn100k.scala 16591:92]
  SnxnLv4Inst204 inst_SnxnLv4Inst204 ( // @[Snxn100k.scala 16575:35]
    .io_a(inst_SnxnLv4Inst204_io_a),
    .io_b(inst_SnxnLv4Inst204_io_b),
    .io_z(inst_SnxnLv4Inst204_io_z)
  );
  SnxnLv4Inst122 inst_SnxnLv4Inst205 ( // @[Snxn100k.scala 16579:35]
    .io_a(inst_SnxnLv4Inst205_io_a),
    .io_b(inst_SnxnLv4Inst205_io_b),
    .io_z(inst_SnxnLv4Inst205_io_z)
  );
  SnxnLv4Inst120 inst_SnxnLv4Inst206 ( // @[Snxn100k.scala 16583:35]
    .io_a(inst_SnxnLv4Inst206_io_a),
    .io_b(inst_SnxnLv4Inst206_io_b),
    .io_z(inst_SnxnLv4Inst206_io_z)
  );
  SnxnLv4Inst207 inst_SnxnLv4Inst207 ( // @[Snxn100k.scala 16587:35]
    .io_a(inst_SnxnLv4Inst207_io_a),
    .io_b(inst_SnxnLv4Inst207_io_b),
    .io_z(inst_SnxnLv4Inst207_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 16592:15]
  assign inst_SnxnLv4Inst204_io_a = io_a; // @[Snxn100k.scala 16576:28]
  assign inst_SnxnLv4Inst204_io_b = io_b; // @[Snxn100k.scala 16577:28]
  assign inst_SnxnLv4Inst205_io_a = io_a; // @[Snxn100k.scala 16580:28]
  assign inst_SnxnLv4Inst205_io_b = io_b; // @[Snxn100k.scala 16581:28]
  assign inst_SnxnLv4Inst206_io_a = io_a; // @[Snxn100k.scala 16584:28]
  assign inst_SnxnLv4Inst206_io_b = io_b; // @[Snxn100k.scala 16585:28]
  assign inst_SnxnLv4Inst207_io_a = io_a; // @[Snxn100k.scala 16588:28]
  assign inst_SnxnLv4Inst207_io_b = io_b; // @[Snxn100k.scala 16589:28]
endmodule
module SnxnLv2Inst12(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst48_io_a; // @[Snxn100k.scala 4271:34]
  wire  inst_SnxnLv3Inst48_io_b; // @[Snxn100k.scala 4271:34]
  wire  inst_SnxnLv3Inst48_io_z; // @[Snxn100k.scala 4271:34]
  wire  inst_SnxnLv3Inst49_io_a; // @[Snxn100k.scala 4275:34]
  wire  inst_SnxnLv3Inst49_io_b; // @[Snxn100k.scala 4275:34]
  wire  inst_SnxnLv3Inst49_io_z; // @[Snxn100k.scala 4275:34]
  wire  inst_SnxnLv3Inst50_io_a; // @[Snxn100k.scala 4279:34]
  wire  inst_SnxnLv3Inst50_io_b; // @[Snxn100k.scala 4279:34]
  wire  inst_SnxnLv3Inst50_io_z; // @[Snxn100k.scala 4279:34]
  wire  inst_SnxnLv3Inst51_io_a; // @[Snxn100k.scala 4283:34]
  wire  inst_SnxnLv3Inst51_io_b; // @[Snxn100k.scala 4283:34]
  wire  inst_SnxnLv3Inst51_io_z; // @[Snxn100k.scala 4283:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst48_io_z + inst_SnxnLv3Inst49_io_z; // @[Snxn100k.scala 4287:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst50_io_z; // @[Snxn100k.scala 4287:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst51_io_z; // @[Snxn100k.scala 4287:89]
  SnxnLv3Inst48 inst_SnxnLv3Inst48 ( // @[Snxn100k.scala 4271:34]
    .io_a(inst_SnxnLv3Inst48_io_a),
    .io_b(inst_SnxnLv3Inst48_io_b),
    .io_z(inst_SnxnLv3Inst48_io_z)
  );
  SnxnLv3Inst49 inst_SnxnLv3Inst49 ( // @[Snxn100k.scala 4275:34]
    .io_a(inst_SnxnLv3Inst49_io_a),
    .io_b(inst_SnxnLv3Inst49_io_b),
    .io_z(inst_SnxnLv3Inst49_io_z)
  );
  SnxnLv3Inst50 inst_SnxnLv3Inst50 ( // @[Snxn100k.scala 4279:34]
    .io_a(inst_SnxnLv3Inst50_io_a),
    .io_b(inst_SnxnLv3Inst50_io_b),
    .io_z(inst_SnxnLv3Inst50_io_z)
  );
  SnxnLv3Inst51 inst_SnxnLv3Inst51 ( // @[Snxn100k.scala 4283:34]
    .io_a(inst_SnxnLv3Inst51_io_a),
    .io_b(inst_SnxnLv3Inst51_io_b),
    .io_z(inst_SnxnLv3Inst51_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 4288:15]
  assign inst_SnxnLv3Inst48_io_a = io_a; // @[Snxn100k.scala 4272:27]
  assign inst_SnxnLv3Inst48_io_b = io_b; // @[Snxn100k.scala 4273:27]
  assign inst_SnxnLv3Inst49_io_a = io_a; // @[Snxn100k.scala 4276:27]
  assign inst_SnxnLv3Inst49_io_b = io_b; // @[Snxn100k.scala 4277:27]
  assign inst_SnxnLv3Inst50_io_a = io_a; // @[Snxn100k.scala 4280:27]
  assign inst_SnxnLv3Inst50_io_b = io_b; // @[Snxn100k.scala 4281:27]
  assign inst_SnxnLv3Inst51_io_a = io_a; // @[Snxn100k.scala 4284:27]
  assign inst_SnxnLv3Inst51_io_b = io_b; // @[Snxn100k.scala 4285:27]
endmodule
module SnxnLv4Inst210(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 50727:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 50728:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 50729:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 50730:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 50731:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 50732:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 50733:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 50734:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 50735:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 50736:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 50737:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 50738:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 50739:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 50740:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 50741:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 50742:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 50743:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 50744:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 50745:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 50746:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 50747:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 50748:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 50749:18]
  assign io_z = ~x5; // @[Snxn100k.scala 50750:15]
endmodule
module SnxnLv4Inst211(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 50761:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 50762:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 50763:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 50764:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 50765:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 50766:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 50767:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 50768:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 50769:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 50770:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 50771:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 50772:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 50773:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 50774:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 50775:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 50776:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 50777:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 50778:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 50779:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 50780:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 50781:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 50782:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 50783:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 50784:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 50785:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 50786:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 50787:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 50788:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 50789:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 50790:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 50791:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 50792:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 50793:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 50794:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 50795:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 50796:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 50797:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 50798:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 50799:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 50800:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 50801:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 50802:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 50803:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 50804:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 50805:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 50806:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 50807:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 50808:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 50809:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 50810:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 50811:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 50812:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 50813:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 50814:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 50815:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 50816:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 50817:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 50818:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 50819:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 50820:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 50821:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 50822:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 50823:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 50824:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 50825:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 50826:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 50827:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 50828:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 50829:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 50830:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 50831:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 50832:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 50833:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 50834:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 50835:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 50836:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 50837:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 50838:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 50839:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 50840:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 50841:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 50842:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 50843:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 50844:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 50845:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 50846:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 50847:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 50848:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 50849:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 50850:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 50851:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 50852:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 50853:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 50854:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 50855:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 50856:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 50857:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 50858:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 50859:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 50860:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 50861:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 50862:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 50863:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 50864:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 50865:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 50866:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 50867:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 50868:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 50869:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 50870:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 50871:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 50872:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 50873:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 50874:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 50875:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 50876:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 50877:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 50878:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 50879:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 50880:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 50881:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 50882:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 50883:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 50884:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 50885:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 50886:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 50887:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 50888:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 50889:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 50890:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 50891:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 50892:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 50893:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 50894:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 50895:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 50896:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 50897:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 50898:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 50899:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 50900:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 50901:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 50902:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 50903:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 50904:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 50905:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 50906:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 50907:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 50908:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 50909:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 50910:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 50911:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 50912:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 50913:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 50914:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 50915:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 50916:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 50917:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 50918:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 50919:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 50920:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 50921:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 50922:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 50923:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 50924:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 50925:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 50926:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 50927:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 50928:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 50929:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 50930:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 50931:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 50932:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 50933:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 50934:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 50935:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 50936:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 50937:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 50938:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 50939:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 50940:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 50941:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 50942:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 50943:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 50944:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 50945:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 50946:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 50947:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 50948:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 50949:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 50950:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 50951:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 50952:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 50953:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 50954:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 50955:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 50956:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 50957:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 50958:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 50959:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 50960:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 50961:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 50962:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 50963:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 50964:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 50965:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 50966:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 50967:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 50968:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 50969:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 50970:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 50971:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 50972:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 50973:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 50974:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 50975:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 50976:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 50977:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 50978:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 50979:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 50980:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 50981:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 50982:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 50983:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 50984:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 50985:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 50986:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 50987:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 50988:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 50989:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 50990:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 50991:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 50992:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 50993:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 50994:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 50995:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 50996:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 50997:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 50998:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 50999:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 51000:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 51001:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 51002:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 51003:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 51004:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 51005:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 51006:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 51007:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 51008:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 51009:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 51010:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 51011:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 51012:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 51013:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 51014:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 51015:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 51016:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 51017:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 51018:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 51019:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 51020:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 51021:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 51022:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 51023:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 51024:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 51025:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 51026:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 51027:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 51028:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 51029:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 51030:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 51031:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 51032:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 51033:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 51034:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 51035:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 51036:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 51037:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 51038:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 51039:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 51040:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 51041:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 51042:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 51043:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 51044:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 51045:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 51046:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 51047:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 51048:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 51049:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 51050:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 51051:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 51052:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 51053:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 51054:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 51055:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 51056:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 51057:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 51058:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 51059:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 51060:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 51061:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 51062:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 51063:20]
  assign io_z = ~x75; // @[Snxn100k.scala 51064:16]
endmodule
module SnxnLv3Inst52(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst208_io_a; // @[Snxn100k.scala 14464:35]
  wire  inst_SnxnLv4Inst208_io_b; // @[Snxn100k.scala 14464:35]
  wire  inst_SnxnLv4Inst208_io_z; // @[Snxn100k.scala 14464:35]
  wire  inst_SnxnLv4Inst209_io_a; // @[Snxn100k.scala 14468:35]
  wire  inst_SnxnLv4Inst209_io_b; // @[Snxn100k.scala 14468:35]
  wire  inst_SnxnLv4Inst209_io_z; // @[Snxn100k.scala 14468:35]
  wire  inst_SnxnLv4Inst210_io_a; // @[Snxn100k.scala 14472:35]
  wire  inst_SnxnLv4Inst210_io_b; // @[Snxn100k.scala 14472:35]
  wire  inst_SnxnLv4Inst210_io_z; // @[Snxn100k.scala 14472:35]
  wire  inst_SnxnLv4Inst211_io_a; // @[Snxn100k.scala 14476:35]
  wire  inst_SnxnLv4Inst211_io_b; // @[Snxn100k.scala 14476:35]
  wire  inst_SnxnLv4Inst211_io_z; // @[Snxn100k.scala 14476:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst208_io_z + inst_SnxnLv4Inst209_io_z; // @[Snxn100k.scala 14480:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst210_io_z; // @[Snxn100k.scala 14480:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst211_io_z; // @[Snxn100k.scala 14480:92]
  SnxnLv4Inst33 inst_SnxnLv4Inst208 ( // @[Snxn100k.scala 14464:35]
    .io_a(inst_SnxnLv4Inst208_io_a),
    .io_b(inst_SnxnLv4Inst208_io_b),
    .io_z(inst_SnxnLv4Inst208_io_z)
  );
  SnxnLv4Inst47 inst_SnxnLv4Inst209 ( // @[Snxn100k.scala 14468:35]
    .io_a(inst_SnxnLv4Inst209_io_a),
    .io_b(inst_SnxnLv4Inst209_io_b),
    .io_z(inst_SnxnLv4Inst209_io_z)
  );
  SnxnLv4Inst210 inst_SnxnLv4Inst210 ( // @[Snxn100k.scala 14472:35]
    .io_a(inst_SnxnLv4Inst210_io_a),
    .io_b(inst_SnxnLv4Inst210_io_b),
    .io_z(inst_SnxnLv4Inst210_io_z)
  );
  SnxnLv4Inst211 inst_SnxnLv4Inst211 ( // @[Snxn100k.scala 14476:35]
    .io_a(inst_SnxnLv4Inst211_io_a),
    .io_b(inst_SnxnLv4Inst211_io_b),
    .io_z(inst_SnxnLv4Inst211_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14481:15]
  assign inst_SnxnLv4Inst208_io_a = io_a; // @[Snxn100k.scala 14465:28]
  assign inst_SnxnLv4Inst208_io_b = io_b; // @[Snxn100k.scala 14466:28]
  assign inst_SnxnLv4Inst209_io_a = io_a; // @[Snxn100k.scala 14469:28]
  assign inst_SnxnLv4Inst209_io_b = io_b; // @[Snxn100k.scala 14470:28]
  assign inst_SnxnLv4Inst210_io_a = io_a; // @[Snxn100k.scala 14473:28]
  assign inst_SnxnLv4Inst210_io_b = io_b; // @[Snxn100k.scala 14474:28]
  assign inst_SnxnLv4Inst211_io_a = io_a; // @[Snxn100k.scala 14477:28]
  assign inst_SnxnLv4Inst211_io_b = io_b; // @[Snxn100k.scala 14478:28]
endmodule
module SnxnLv3Inst53(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst212_io_a; // @[Snxn100k.scala 14827:35]
  wire  inst_SnxnLv4Inst212_io_b; // @[Snxn100k.scala 14827:35]
  wire  inst_SnxnLv4Inst212_io_z; // @[Snxn100k.scala 14827:35]
  wire  inst_SnxnLv4Inst213_io_a; // @[Snxn100k.scala 14831:35]
  wire  inst_SnxnLv4Inst213_io_b; // @[Snxn100k.scala 14831:35]
  wire  inst_SnxnLv4Inst213_io_z; // @[Snxn100k.scala 14831:35]
  wire  inst_SnxnLv4Inst214_io_a; // @[Snxn100k.scala 14835:35]
  wire  inst_SnxnLv4Inst214_io_b; // @[Snxn100k.scala 14835:35]
  wire  inst_SnxnLv4Inst214_io_z; // @[Snxn100k.scala 14835:35]
  wire  inst_SnxnLv4Inst215_io_a; // @[Snxn100k.scala 14839:35]
  wire  inst_SnxnLv4Inst215_io_b; // @[Snxn100k.scala 14839:35]
  wire  inst_SnxnLv4Inst215_io_z; // @[Snxn100k.scala 14839:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst212_io_z + inst_SnxnLv4Inst213_io_z; // @[Snxn100k.scala 14843:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst214_io_z; // @[Snxn100k.scala 14843:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst215_io_z; // @[Snxn100k.scala 14843:92]
  SnxnLv4Inst93 inst_SnxnLv4Inst212 ( // @[Snxn100k.scala 14827:35]
    .io_a(inst_SnxnLv4Inst212_io_a),
    .io_b(inst_SnxnLv4Inst212_io_b),
    .io_z(inst_SnxnLv4Inst212_io_z)
  );
  SnxnLv4Inst6 inst_SnxnLv4Inst213 ( // @[Snxn100k.scala 14831:35]
    .io_a(inst_SnxnLv4Inst213_io_a),
    .io_b(inst_SnxnLv4Inst213_io_b),
    .io_z(inst_SnxnLv4Inst213_io_z)
  );
  SnxnLv4Inst119 inst_SnxnLv4Inst214 ( // @[Snxn100k.scala 14835:35]
    .io_a(inst_SnxnLv4Inst214_io_a),
    .io_b(inst_SnxnLv4Inst214_io_b),
    .io_z(inst_SnxnLv4Inst214_io_z)
  );
  SnxnLv4Inst16 inst_SnxnLv4Inst215 ( // @[Snxn100k.scala 14839:35]
    .io_a(inst_SnxnLv4Inst215_io_a),
    .io_b(inst_SnxnLv4Inst215_io_b),
    .io_z(inst_SnxnLv4Inst215_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 14844:15]
  assign inst_SnxnLv4Inst212_io_a = io_a; // @[Snxn100k.scala 14828:28]
  assign inst_SnxnLv4Inst212_io_b = io_b; // @[Snxn100k.scala 14829:28]
  assign inst_SnxnLv4Inst213_io_a = io_a; // @[Snxn100k.scala 14832:28]
  assign inst_SnxnLv4Inst213_io_b = io_b; // @[Snxn100k.scala 14833:28]
  assign inst_SnxnLv4Inst214_io_a = io_a; // @[Snxn100k.scala 14836:28]
  assign inst_SnxnLv4Inst214_io_b = io_b; // @[Snxn100k.scala 14837:28]
  assign inst_SnxnLv4Inst215_io_a = io_a; // @[Snxn100k.scala 14840:28]
  assign inst_SnxnLv4Inst215_io_b = io_b; // @[Snxn100k.scala 14841:28]
endmodule
module SnxnLv4Inst218(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 54417:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 54418:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 54419:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 54420:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 54421:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 54422:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 54423:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 54424:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 54425:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 54426:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 54427:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 54428:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 54429:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 54430:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 54431:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 54432:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 54433:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 54434:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 54435:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 54436:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 54437:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 54438:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 54439:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 54440:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 54441:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 54442:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 54443:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 54444:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 54445:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 54446:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 54447:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 54448:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 54449:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 54450:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 54451:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 54452:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 54453:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 54454:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 54455:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 54456:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 54457:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 54458:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 54459:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 54460:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 54461:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 54462:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 54463:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 54464:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 54465:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 54466:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 54467:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 54468:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 54469:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 54470:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 54471:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 54472:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 54473:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 54474:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 54475:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 54476:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 54477:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 54478:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 54479:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 54480:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 54481:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 54482:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 54483:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 54484:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 54485:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 54486:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 54487:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 54488:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 54489:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 54490:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 54491:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 54492:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 54493:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 54494:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 54495:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 54496:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 54497:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 54498:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 54499:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 54500:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 54501:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 54502:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 54503:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 54504:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 54505:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 54506:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 54507:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 54508:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 54509:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 54510:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 54511:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 54512:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 54513:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 54514:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 54515:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 54516:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 54517:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 54518:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 54519:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 54520:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 54521:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 54522:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 54523:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 54524:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 54525:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 54526:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 54527:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 54528:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 54529:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 54530:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 54531:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 54532:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 54533:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 54534:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 54535:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 54536:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 54537:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 54538:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 54539:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 54540:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 54541:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 54542:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 54543:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 54544:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 54545:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 54546:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 54547:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 54548:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 54549:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 54550:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 54551:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 54552:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 54553:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 54554:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 54555:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 54556:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 54557:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 54558:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 54559:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 54560:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 54561:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 54562:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 54563:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 54564:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 54565:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 54566:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 54567:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 54568:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 54569:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 54570:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 54571:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 54572:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 54573:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 54574:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 54575:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 54576:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 54577:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 54578:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 54579:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 54580:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 54581:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 54582:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 54583:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 54584:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 54585:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 54586:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 54587:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 54588:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 54589:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 54590:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 54591:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 54592:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 54593:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 54594:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 54595:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 54596:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 54597:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 54598:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 54599:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 54600:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 54601:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 54602:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 54603:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 54604:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 54605:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 54606:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 54607:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 54608:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 54609:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 54610:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 54611:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 54612:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 54613:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 54614:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 54615:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 54616:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 54617:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 54618:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 54619:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 54620:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 54621:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 54622:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 54623:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 54624:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 54625:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 54626:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 54627:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 54628:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 54629:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 54630:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 54631:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 54632:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 54633:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 54634:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 54635:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 54636:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 54637:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 54638:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 54639:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 54640:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 54641:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 54642:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 54643:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 54644:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 54645:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 54646:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 54647:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 54648:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 54649:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 54650:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 54651:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 54652:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 54653:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 54654:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 54655:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 54656:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 54657:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 54658:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 54659:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 54660:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 54661:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 54662:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 54663:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 54664:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 54665:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 54666:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 54667:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 54668:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 54669:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 54670:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 54671:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 54672:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 54673:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 54674:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 54675:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 54676:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 54677:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 54678:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 54679:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 54680:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 54681:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 54682:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 54683:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 54684:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 54685:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 54686:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 54687:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 54688:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 54689:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 54690:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 54691:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 54692:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 54693:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 54694:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 54695:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 54696:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 54697:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 54698:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 54699:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 54700:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 54701:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 54702:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 54703:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 54704:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 54705:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 54706:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 54707:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 54708:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 54709:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 54710:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 54711:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 54712:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 54713:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 54714:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 54715:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 54716:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 54717:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 54718:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 54719:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 54720:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 54721:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 54722:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 54723:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 54724:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 54725:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 54726:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 54727:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 54728:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 54729:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 54730:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 54731:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 54732:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 54733:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 54734:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 54735:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 54736:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 54737:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 54738:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 54739:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 54740:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 54741:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 54742:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 54743:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 54744:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 54745:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 54746:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 54747:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 54748:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 54749:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 54750:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 54751:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 54752:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 54753:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 54754:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 54755:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 54756:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 54757:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 54758:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 54759:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 54760:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 54761:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 54762:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 54763:20]
  assign io_z = ~x86; // @[Snxn100k.scala 54764:16]
endmodule
module SnxnLv4Inst219(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 54775:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 54776:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 54777:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 54778:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 54779:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 54780:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 54781:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 54782:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 54783:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 54784:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 54785:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 54786:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 54787:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 54788:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 54789:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 54790:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 54791:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 54792:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 54793:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 54794:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 54795:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 54796:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 54797:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 54798:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 54799:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 54800:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 54801:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 54802:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 54803:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 54804:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 54805:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 54806:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 54807:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 54808:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 54809:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 54810:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 54811:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 54812:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 54813:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 54814:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 54815:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 54816:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 54817:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 54818:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 54819:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 54820:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 54821:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 54822:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 54823:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 54824:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 54825:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 54826:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 54827:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 54828:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 54829:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 54830:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 54831:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 54832:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 54833:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 54834:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 54835:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 54836:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 54837:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 54838:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 54839:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 54840:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 54841:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 54842:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 54843:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 54844:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 54845:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 54846:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 54847:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 54848:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 54849:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 54850:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 54851:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 54852:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 54853:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 54854:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 54855:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 54856:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 54857:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 54858:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 54859:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 54860:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 54861:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 54862:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 54863:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 54864:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 54865:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 54866:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 54867:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 54868:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 54869:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 54870:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 54871:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 54872:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 54873:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 54874:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 54875:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 54876:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 54877:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 54878:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 54879:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 54880:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 54881:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 54882:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 54883:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 54884:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 54885:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 54886:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 54887:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 54888:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 54889:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 54890:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 54891:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 54892:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 54893:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 54894:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 54895:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 54896:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 54897:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 54898:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 54899:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 54900:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 54901:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 54902:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 54903:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 54904:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 54905:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 54906:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 54907:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 54908:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 54909:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 54910:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 54911:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 54912:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 54913:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 54914:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 54915:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 54916:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 54917:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 54918:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 54919:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 54920:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 54921:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 54922:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 54923:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 54924:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 54925:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 54926:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 54927:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 54928:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 54929:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 54930:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 54931:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 54932:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 54933:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 54934:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 54935:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 54936:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 54937:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 54938:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 54939:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 54940:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 54941:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 54942:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 54943:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 54944:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 54945:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 54946:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 54947:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 54948:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 54949:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 54950:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 54951:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 54952:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 54953:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 54954:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 54955:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 54956:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 54957:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 54958:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 54959:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 54960:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 54961:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 54962:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 54963:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 54964:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 54965:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 54966:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 54967:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 54968:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 54969:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 54970:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 54971:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 54972:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 54973:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 54974:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 54975:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 54976:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 54977:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 54978:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 54979:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 54980:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 54981:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 54982:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 54983:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 54984:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 54985:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 54986:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 54987:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 54988:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 54989:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 54990:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 54991:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 54992:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 54993:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 54994:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 54995:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 54996:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 54997:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 54998:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 54999:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 55000:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 55001:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 55002:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 55003:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 55004:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 55005:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 55006:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 55007:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 55008:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 55009:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 55010:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 55011:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 55012:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 55013:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 55014:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 55015:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 55016:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 55017:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 55018:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 55019:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 55020:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 55021:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 55022:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 55023:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 55024:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 55025:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 55026:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 55027:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 55028:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 55029:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 55030:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 55031:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 55032:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 55033:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 55034:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 55035:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 55036:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 55037:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 55038:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 55039:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 55040:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 55041:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 55042:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 55043:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 55044:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 55045:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 55046:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 55047:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 55048:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 55049:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 55050:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 55051:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 55052:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 55053:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 55054:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 55055:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 55056:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 55057:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 55058:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 55059:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 55060:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 55061:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 55062:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 55063:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 55064:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 55065:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 55066:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 55067:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 55068:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 55069:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 55070:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 55071:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 55072:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 55073:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 55074:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 55075:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 55076:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 55077:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 55078:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 55079:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 55080:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 55081:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 55082:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 55083:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 55084:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 55085:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 55086:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 55087:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 55088:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 55089:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 55090:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 55091:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 55092:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 55093:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 55094:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 55095:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 55096:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 55097:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 55098:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 55099:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 55100:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 55101:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 55102:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 55103:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 55104:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 55105:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 55106:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 55107:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 55108:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 55109:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 55110:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 55111:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 55112:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 55113:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 55114:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 55115:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 55116:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 55117:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 55118:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 55119:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 55120:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 55121:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 55122:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 55123:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 55124:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 55125:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 55126:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 55127:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 55128:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 55129:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 55130:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 55131:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 55132:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 55133:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 55134:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 55135:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 55136:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 55137:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 55138:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 55139:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 55140:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 55141:20]
  assign io_z = ~x91; // @[Snxn100k.scala 55142:16]
endmodule
module SnxnLv3Inst54(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst216_io_a; // @[Snxn100k.scala 15753:35]
  wire  inst_SnxnLv4Inst216_io_b; // @[Snxn100k.scala 15753:35]
  wire  inst_SnxnLv4Inst216_io_z; // @[Snxn100k.scala 15753:35]
  wire  inst_SnxnLv4Inst217_io_a; // @[Snxn100k.scala 15757:35]
  wire  inst_SnxnLv4Inst217_io_b; // @[Snxn100k.scala 15757:35]
  wire  inst_SnxnLv4Inst217_io_z; // @[Snxn100k.scala 15757:35]
  wire  inst_SnxnLv4Inst218_io_a; // @[Snxn100k.scala 15761:35]
  wire  inst_SnxnLv4Inst218_io_b; // @[Snxn100k.scala 15761:35]
  wire  inst_SnxnLv4Inst218_io_z; // @[Snxn100k.scala 15761:35]
  wire  inst_SnxnLv4Inst219_io_a; // @[Snxn100k.scala 15765:35]
  wire  inst_SnxnLv4Inst219_io_b; // @[Snxn100k.scala 15765:35]
  wire  inst_SnxnLv4Inst219_io_z; // @[Snxn100k.scala 15765:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst216_io_z + inst_SnxnLv4Inst217_io_z; // @[Snxn100k.scala 15769:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst218_io_z; // @[Snxn100k.scala 15769:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst219_io_z; // @[Snxn100k.scala 15769:92]
  SnxnLv4Inst0 inst_SnxnLv4Inst216 ( // @[Snxn100k.scala 15753:35]
    .io_a(inst_SnxnLv4Inst216_io_a),
    .io_b(inst_SnxnLv4Inst216_io_b),
    .io_z(inst_SnxnLv4Inst216_io_z)
  );
  SnxnLv4Inst55 inst_SnxnLv4Inst217 ( // @[Snxn100k.scala 15757:35]
    .io_a(inst_SnxnLv4Inst217_io_a),
    .io_b(inst_SnxnLv4Inst217_io_b),
    .io_z(inst_SnxnLv4Inst217_io_z)
  );
  SnxnLv4Inst218 inst_SnxnLv4Inst218 ( // @[Snxn100k.scala 15761:35]
    .io_a(inst_SnxnLv4Inst218_io_a),
    .io_b(inst_SnxnLv4Inst218_io_b),
    .io_z(inst_SnxnLv4Inst218_io_z)
  );
  SnxnLv4Inst219 inst_SnxnLv4Inst219 ( // @[Snxn100k.scala 15765:35]
    .io_a(inst_SnxnLv4Inst219_io_a),
    .io_b(inst_SnxnLv4Inst219_io_b),
    .io_z(inst_SnxnLv4Inst219_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 15770:15]
  assign inst_SnxnLv4Inst216_io_a = io_a; // @[Snxn100k.scala 15754:28]
  assign inst_SnxnLv4Inst216_io_b = io_b; // @[Snxn100k.scala 15755:28]
  assign inst_SnxnLv4Inst217_io_a = io_a; // @[Snxn100k.scala 15758:28]
  assign inst_SnxnLv4Inst217_io_b = io_b; // @[Snxn100k.scala 15759:28]
  assign inst_SnxnLv4Inst218_io_a = io_a; // @[Snxn100k.scala 15762:28]
  assign inst_SnxnLv4Inst218_io_b = io_b; // @[Snxn100k.scala 15763:28]
  assign inst_SnxnLv4Inst219_io_a = io_a; // @[Snxn100k.scala 15766:28]
  assign inst_SnxnLv4Inst219_io_b = io_b; // @[Snxn100k.scala 15767:28]
endmodule
module SnxnLv4Inst221(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 53919:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 53920:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 53921:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 53922:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 53923:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 53924:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 53925:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 53926:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 53927:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 53928:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 53929:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 53930:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 53931:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 53932:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 53933:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 53934:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 53935:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 53936:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 53937:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 53938:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 53939:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 53940:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 53941:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 53942:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 53943:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 53944:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 53945:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 53946:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 53947:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 53948:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 53949:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 53950:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 53951:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 53952:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 53953:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 53954:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 53955:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 53956:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 53957:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 53958:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 53959:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 53960:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 53961:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 53962:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 53963:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 53964:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 53965:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 53966:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 53967:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 53968:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 53969:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 53970:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 53971:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 53972:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 53973:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 53974:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 53975:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 53976:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 53977:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 53978:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 53979:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 53980:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 53981:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 53982:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 53983:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 53984:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 53985:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 53986:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 53987:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 53988:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 53989:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 53990:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 53991:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 53992:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 53993:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 53994:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 53995:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 53996:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 53997:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 53998:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 53999:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 54000:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 54001:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 54002:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 54003:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 54004:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 54005:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 54006:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 54007:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 54008:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 54009:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 54010:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 54011:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 54012:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 54013:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 54014:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 54015:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 54016:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 54017:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 54018:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 54019:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 54020:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 54021:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 54022:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 54023:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 54024:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 54025:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 54026:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 54027:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 54028:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 54029:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 54030:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 54031:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 54032:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 54033:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 54034:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 54035:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 54036:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 54037:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 54038:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 54039:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 54040:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 54041:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 54042:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 54043:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 54044:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 54045:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 54046:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 54047:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 54048:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 54049:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 54050:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 54051:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 54052:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 54053:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 54054:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 54055:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 54056:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 54057:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 54058:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 54059:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 54060:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 54061:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 54062:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 54063:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 54064:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 54065:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 54066:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 54067:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 54068:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 54069:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 54070:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 54071:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 54072:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 54073:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 54074:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 54075:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 54076:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 54077:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 54078:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 54079:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 54080:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 54081:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 54082:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 54083:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 54084:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 54085:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 54086:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 54087:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 54088:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 54089:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 54090:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 54091:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 54092:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 54093:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 54094:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 54095:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 54096:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 54097:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 54098:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 54099:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 54100:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 54101:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 54102:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 54103:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 54104:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 54105:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 54106:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 54107:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 54108:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 54109:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 54110:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 54111:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 54112:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 54113:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 54114:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 54115:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 54116:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 54117:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 54118:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 54119:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 54120:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 54121:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 54122:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 54123:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 54124:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 54125:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 54126:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 54127:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 54128:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 54129:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 54130:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 54131:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 54132:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 54133:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 54134:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 54135:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 54136:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 54137:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 54138:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 54139:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 54140:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 54141:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 54142:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 54143:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 54144:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 54145:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 54146:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 54147:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 54148:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 54149:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 54150:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 54151:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 54152:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 54153:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 54154:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 54155:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 54156:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 54157:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 54158:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 54159:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 54160:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 54161:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 54162:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 54163:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 54164:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 54165:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 54166:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 54167:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 54168:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 54169:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 54170:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 54171:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 54172:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 54173:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 54174:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 54175:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 54176:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 54177:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 54178:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 54179:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 54180:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 54181:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 54182:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 54183:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 54184:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 54185:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 54186:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 54187:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 54188:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 54189:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 54190:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 54191:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 54192:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 54193:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 54194:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 54195:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 54196:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 54197:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 54198:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 54199:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 54200:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 54201:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 54202:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 54203:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 54204:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 54205:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 54206:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 54207:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 54208:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 54209:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 54210:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 54211:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 54212:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 54213:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 54214:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 54215:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 54216:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 54217:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 54218:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 54219:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 54220:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 54221:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 54222:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 54223:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 54224:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 54225:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 54226:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 54227:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 54228:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 54229:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 54230:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 54231:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 54232:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 54233:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 54234:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 54235:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 54236:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 54237:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 54238:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 54239:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 54240:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 54241:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 54242:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 54243:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 54244:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 54245:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 54246:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 54247:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 54248:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 54249:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 54250:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 54251:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 54252:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 54253:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 54254:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 54255:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 54256:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 54257:20]
  wire  invx84 = ~x84; // @[Snxn100k.scala 54258:16]
  wire  t85 = x84 + invx84; // @[Snxn100k.scala 54259:20]
  wire  inv85 = ~t85; // @[Snxn100k.scala 54260:16]
  wire  x85 = t85 ^ inv85; // @[Snxn100k.scala 54261:20]
  wire  invx85 = ~x85; // @[Snxn100k.scala 54262:16]
  wire  t86 = x85 + invx85; // @[Snxn100k.scala 54263:20]
  wire  inv86 = ~t86; // @[Snxn100k.scala 54264:16]
  wire  x86 = t86 ^ inv86; // @[Snxn100k.scala 54265:20]
  wire  invx86 = ~x86; // @[Snxn100k.scala 54266:16]
  wire  t87 = x86 + invx86; // @[Snxn100k.scala 54267:20]
  wire  inv87 = ~t87; // @[Snxn100k.scala 54268:16]
  wire  x87 = t87 ^ inv87; // @[Snxn100k.scala 54269:20]
  wire  invx87 = ~x87; // @[Snxn100k.scala 54270:16]
  wire  t88 = x87 + invx87; // @[Snxn100k.scala 54271:20]
  wire  inv88 = ~t88; // @[Snxn100k.scala 54272:16]
  wire  x88 = t88 ^ inv88; // @[Snxn100k.scala 54273:20]
  wire  invx88 = ~x88; // @[Snxn100k.scala 54274:16]
  wire  t89 = x88 + invx88; // @[Snxn100k.scala 54275:20]
  wire  inv89 = ~t89; // @[Snxn100k.scala 54276:16]
  wire  x89 = t89 ^ inv89; // @[Snxn100k.scala 54277:20]
  wire  invx89 = ~x89; // @[Snxn100k.scala 54278:16]
  wire  t90 = x89 + invx89; // @[Snxn100k.scala 54279:20]
  wire  inv90 = ~t90; // @[Snxn100k.scala 54280:16]
  wire  x90 = t90 ^ inv90; // @[Snxn100k.scala 54281:20]
  wire  invx90 = ~x90; // @[Snxn100k.scala 54282:16]
  wire  t91 = x90 + invx90; // @[Snxn100k.scala 54283:20]
  wire  inv91 = ~t91; // @[Snxn100k.scala 54284:16]
  wire  x91 = t91 ^ inv91; // @[Snxn100k.scala 54285:20]
  wire  invx91 = ~x91; // @[Snxn100k.scala 54286:16]
  wire  t92 = x91 + invx91; // @[Snxn100k.scala 54287:20]
  wire  inv92 = ~t92; // @[Snxn100k.scala 54288:16]
  wire  x92 = t92 ^ inv92; // @[Snxn100k.scala 54289:20]
  wire  invx92 = ~x92; // @[Snxn100k.scala 54290:16]
  wire  t93 = x92 + invx92; // @[Snxn100k.scala 54291:20]
  wire  inv93 = ~t93; // @[Snxn100k.scala 54292:16]
  wire  x93 = t93 ^ inv93; // @[Snxn100k.scala 54293:20]
  wire  invx93 = ~x93; // @[Snxn100k.scala 54294:16]
  wire  t94 = x93 + invx93; // @[Snxn100k.scala 54295:20]
  wire  inv94 = ~t94; // @[Snxn100k.scala 54296:16]
  wire  x94 = t94 ^ inv94; // @[Snxn100k.scala 54297:20]
  wire  invx94 = ~x94; // @[Snxn100k.scala 54298:16]
  wire  t95 = x94 + invx94; // @[Snxn100k.scala 54299:20]
  wire  inv95 = ~t95; // @[Snxn100k.scala 54300:16]
  wire  x95 = t95 ^ inv95; // @[Snxn100k.scala 54301:20]
  wire  invx95 = ~x95; // @[Snxn100k.scala 54302:16]
  wire  t96 = x95 + invx95; // @[Snxn100k.scala 54303:20]
  wire  inv96 = ~t96; // @[Snxn100k.scala 54304:16]
  wire  x96 = t96 ^ inv96; // @[Snxn100k.scala 54305:20]
  wire  invx96 = ~x96; // @[Snxn100k.scala 54306:16]
  wire  t97 = x96 + invx96; // @[Snxn100k.scala 54307:20]
  wire  inv97 = ~t97; // @[Snxn100k.scala 54308:16]
  wire  x97 = t97 ^ inv97; // @[Snxn100k.scala 54309:20]
  wire  invx97 = ~x97; // @[Snxn100k.scala 54310:16]
  wire  t98 = x97 + invx97; // @[Snxn100k.scala 54311:20]
  wire  inv98 = ~t98; // @[Snxn100k.scala 54312:16]
  wire  x98 = t98 ^ inv98; // @[Snxn100k.scala 54313:20]
  wire  invx98 = ~x98; // @[Snxn100k.scala 54314:16]
  wire  t99 = x98 + invx98; // @[Snxn100k.scala 54315:20]
  wire  inv99 = ~t99; // @[Snxn100k.scala 54316:16]
  wire  x99 = t99 ^ inv99; // @[Snxn100k.scala 54317:20]
  wire  invx99 = ~x99; // @[Snxn100k.scala 54318:16]
  wire  t100 = x99 + invx99; // @[Snxn100k.scala 54319:21]
  wire  inv100 = ~t100; // @[Snxn100k.scala 54320:17]
  wire  x100 = t100 ^ inv100; // @[Snxn100k.scala 54321:22]
  wire  invx100 = ~x100; // @[Snxn100k.scala 54322:17]
  wire  t101 = x100 + invx100; // @[Snxn100k.scala 54323:22]
  wire  inv101 = ~t101; // @[Snxn100k.scala 54324:17]
  wire  x101 = t101 ^ inv101; // @[Snxn100k.scala 54325:22]
  wire  invx101 = ~x101; // @[Snxn100k.scala 54326:17]
  wire  t102 = x101 + invx101; // @[Snxn100k.scala 54327:22]
  wire  inv102 = ~t102; // @[Snxn100k.scala 54328:17]
  wire  x102 = t102 ^ inv102; // @[Snxn100k.scala 54329:22]
  wire  invx102 = ~x102; // @[Snxn100k.scala 54330:17]
  wire  t103 = x102 + invx102; // @[Snxn100k.scala 54331:22]
  wire  inv103 = ~t103; // @[Snxn100k.scala 54332:17]
  wire  x103 = t103 ^ inv103; // @[Snxn100k.scala 54333:22]
  wire  invx103 = ~x103; // @[Snxn100k.scala 54334:17]
  wire  t104 = x103 + invx103; // @[Snxn100k.scala 54335:22]
  wire  inv104 = ~t104; // @[Snxn100k.scala 54336:17]
  wire  x104 = t104 ^ inv104; // @[Snxn100k.scala 54337:22]
  wire  invx104 = ~x104; // @[Snxn100k.scala 54338:17]
  wire  t105 = x104 + invx104; // @[Snxn100k.scala 54339:22]
  wire  inv105 = ~t105; // @[Snxn100k.scala 54340:17]
  wire  x105 = t105 ^ inv105; // @[Snxn100k.scala 54341:22]
  wire  invx105 = ~x105; // @[Snxn100k.scala 54342:17]
  wire  t106 = x105 + invx105; // @[Snxn100k.scala 54343:22]
  wire  inv106 = ~t106; // @[Snxn100k.scala 54344:17]
  wire  x106 = t106 ^ inv106; // @[Snxn100k.scala 54345:22]
  wire  invx106 = ~x106; // @[Snxn100k.scala 54346:17]
  wire  t107 = x106 + invx106; // @[Snxn100k.scala 54347:22]
  wire  inv107 = ~t107; // @[Snxn100k.scala 54348:17]
  wire  x107 = t107 ^ inv107; // @[Snxn100k.scala 54349:22]
  wire  invx107 = ~x107; // @[Snxn100k.scala 54350:17]
  wire  t108 = x107 + invx107; // @[Snxn100k.scala 54351:22]
  wire  inv108 = ~t108; // @[Snxn100k.scala 54352:17]
  wire  x108 = t108 ^ inv108; // @[Snxn100k.scala 54353:22]
  wire  invx108 = ~x108; // @[Snxn100k.scala 54354:17]
  wire  t109 = x108 + invx108; // @[Snxn100k.scala 54355:22]
  wire  inv109 = ~t109; // @[Snxn100k.scala 54356:17]
  wire  x109 = t109 ^ inv109; // @[Snxn100k.scala 54357:22]
  wire  invx109 = ~x109; // @[Snxn100k.scala 54358:17]
  wire  t110 = x109 + invx109; // @[Snxn100k.scala 54359:22]
  wire  inv110 = ~t110; // @[Snxn100k.scala 54360:17]
  wire  x110 = t110 ^ inv110; // @[Snxn100k.scala 54361:22]
  wire  invx110 = ~x110; // @[Snxn100k.scala 54362:17]
  wire  t111 = x110 + invx110; // @[Snxn100k.scala 54363:22]
  wire  inv111 = ~t111; // @[Snxn100k.scala 54364:17]
  wire  x111 = t111 ^ inv111; // @[Snxn100k.scala 54365:22]
  wire  invx111 = ~x111; // @[Snxn100k.scala 54366:17]
  wire  t112 = x111 + invx111; // @[Snxn100k.scala 54367:22]
  wire  inv112 = ~t112; // @[Snxn100k.scala 54368:17]
  wire  x112 = t112 ^ inv112; // @[Snxn100k.scala 54369:22]
  wire  invx112 = ~x112; // @[Snxn100k.scala 54370:17]
  wire  t113 = x112 + invx112; // @[Snxn100k.scala 54371:22]
  wire  inv113 = ~t113; // @[Snxn100k.scala 54372:17]
  wire  x113 = t113 ^ inv113; // @[Snxn100k.scala 54373:22]
  wire  invx113 = ~x113; // @[Snxn100k.scala 54374:17]
  wire  t114 = x113 + invx113; // @[Snxn100k.scala 54375:22]
  wire  inv114 = ~t114; // @[Snxn100k.scala 54376:17]
  wire  x114 = t114 ^ inv114; // @[Snxn100k.scala 54377:22]
  wire  invx114 = ~x114; // @[Snxn100k.scala 54378:17]
  wire  t115 = x114 + invx114; // @[Snxn100k.scala 54379:22]
  wire  inv115 = ~t115; // @[Snxn100k.scala 54380:17]
  wire  x115 = t115 ^ inv115; // @[Snxn100k.scala 54381:22]
  wire  invx115 = ~x115; // @[Snxn100k.scala 54382:17]
  wire  t116 = x115 + invx115; // @[Snxn100k.scala 54383:22]
  wire  inv116 = ~t116; // @[Snxn100k.scala 54384:17]
  wire  x116 = t116 ^ inv116; // @[Snxn100k.scala 54385:22]
  wire  invx116 = ~x116; // @[Snxn100k.scala 54386:17]
  wire  t117 = x116 + invx116; // @[Snxn100k.scala 54387:22]
  wire  inv117 = ~t117; // @[Snxn100k.scala 54388:17]
  wire  x117 = t117 ^ inv117; // @[Snxn100k.scala 54389:22]
  wire  invx117 = ~x117; // @[Snxn100k.scala 54390:17]
  wire  t118 = x117 + invx117; // @[Snxn100k.scala 54391:22]
  wire  inv118 = ~t118; // @[Snxn100k.scala 54392:17]
  wire  x118 = t118 ^ inv118; // @[Snxn100k.scala 54393:22]
  wire  invx118 = ~x118; // @[Snxn100k.scala 54394:17]
  wire  t119 = x118 + invx118; // @[Snxn100k.scala 54395:22]
  wire  inv119 = ~t119; // @[Snxn100k.scala 54396:17]
  wire  x119 = t119 ^ inv119; // @[Snxn100k.scala 54397:22]
  wire  invx119 = ~x119; // @[Snxn100k.scala 54398:17]
  wire  t120 = x119 + invx119; // @[Snxn100k.scala 54399:22]
  wire  inv120 = ~t120; // @[Snxn100k.scala 54400:17]
  wire  x120 = t120 ^ inv120; // @[Snxn100k.scala 54401:22]
  wire  invx120 = ~x120; // @[Snxn100k.scala 54402:17]
  wire  t121 = x120 + invx120; // @[Snxn100k.scala 54403:22]
  wire  inv121 = ~t121; // @[Snxn100k.scala 54404:17]
  wire  x121 = t121 ^ inv121; // @[Snxn100k.scala 54405:22]
  assign io_z = ~x121; // @[Snxn100k.scala 54406:17]
endmodule
module SnxnLv4Inst223(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 53347:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 53348:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 53349:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 53350:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 53351:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 53352:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 53353:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 53354:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 53355:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 53356:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 53357:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 53358:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 53359:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 53360:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 53361:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 53362:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 53363:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 53364:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 53365:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 53366:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 53367:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 53368:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 53369:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 53370:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 53371:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 53372:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 53373:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 53374:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 53375:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 53376:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 53377:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 53378:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 53379:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 53380:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 53381:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 53382:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 53383:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 53384:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 53385:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 53386:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 53387:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 53388:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 53389:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 53390:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 53391:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 53392:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 53393:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 53394:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 53395:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 53396:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 53397:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 53398:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 53399:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 53400:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 53401:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 53402:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 53403:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 53404:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 53405:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 53406:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 53407:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 53408:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 53409:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 53410:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 53411:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 53412:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 53413:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 53414:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 53415:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 53416:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 53417:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 53418:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 53419:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 53420:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 53421:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 53422:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 53423:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 53424:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 53425:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 53426:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 53427:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 53428:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 53429:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 53430:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 53431:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 53432:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 53433:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 53434:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 53435:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 53436:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 53437:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 53438:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 53439:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 53440:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 53441:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 53442:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 53443:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 53444:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 53445:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 53446:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 53447:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 53448:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 53449:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 53450:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 53451:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 53452:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 53453:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 53454:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 53455:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 53456:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 53457:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 53458:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 53459:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 53460:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 53461:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 53462:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 53463:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 53464:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 53465:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 53466:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 53467:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 53468:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 53469:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 53470:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 53471:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 53472:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 53473:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 53474:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 53475:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 53476:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 53477:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 53478:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 53479:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 53480:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 53481:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 53482:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 53483:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 53484:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 53485:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 53486:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 53487:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 53488:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 53489:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 53490:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 53491:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 53492:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 53493:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 53494:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 53495:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 53496:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 53497:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 53498:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 53499:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 53500:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 53501:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 53502:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 53503:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 53504:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 53505:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 53506:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 53507:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 53508:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 53509:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 53510:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 53511:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 53512:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 53513:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 53514:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 53515:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 53516:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 53517:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 53518:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 53519:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 53520:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 53521:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 53522:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 53523:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 53524:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 53525:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 53526:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 53527:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 53528:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 53529:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 53530:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 53531:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 53532:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 53533:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 53534:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 53535:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 53536:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 53537:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 53538:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 53539:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 53540:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 53541:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 53542:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 53543:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 53544:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 53545:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 53546:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 53547:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 53548:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 53549:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 53550:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 53551:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 53552:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 53553:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 53554:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 53555:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 53556:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 53557:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 53558:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 53559:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 53560:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 53561:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 53562:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 53563:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 53564:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 53565:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 53566:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 53567:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 53568:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 53569:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 53570:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 53571:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 53572:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 53573:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 53574:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 53575:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 53576:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 53577:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 53578:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 53579:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 53580:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 53581:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 53582:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 53583:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 53584:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 53585:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 53586:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 53587:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 53588:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 53589:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 53590:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 53591:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 53592:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 53593:20]
  assign io_z = ~x61; // @[Snxn100k.scala 53594:16]
endmodule
module SnxnLv3Inst55(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst220_io_a; // @[Snxn100k.scala 15262:35]
  wire  inst_SnxnLv4Inst220_io_b; // @[Snxn100k.scala 15262:35]
  wire  inst_SnxnLv4Inst220_io_z; // @[Snxn100k.scala 15262:35]
  wire  inst_SnxnLv4Inst221_io_a; // @[Snxn100k.scala 15266:35]
  wire  inst_SnxnLv4Inst221_io_b; // @[Snxn100k.scala 15266:35]
  wire  inst_SnxnLv4Inst221_io_z; // @[Snxn100k.scala 15266:35]
  wire  inst_SnxnLv4Inst222_io_a; // @[Snxn100k.scala 15270:35]
  wire  inst_SnxnLv4Inst222_io_b; // @[Snxn100k.scala 15270:35]
  wire  inst_SnxnLv4Inst222_io_z; // @[Snxn100k.scala 15270:35]
  wire  inst_SnxnLv4Inst223_io_a; // @[Snxn100k.scala 15274:35]
  wire  inst_SnxnLv4Inst223_io_b; // @[Snxn100k.scala 15274:35]
  wire  inst_SnxnLv4Inst223_io_z; // @[Snxn100k.scala 15274:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst220_io_z + inst_SnxnLv4Inst221_io_z; // @[Snxn100k.scala 15278:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst222_io_z; // @[Snxn100k.scala 15278:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst223_io_z; // @[Snxn100k.scala 15278:92]
  SnxnLv4Inst211 inst_SnxnLv4Inst220 ( // @[Snxn100k.scala 15262:35]
    .io_a(inst_SnxnLv4Inst220_io_a),
    .io_b(inst_SnxnLv4Inst220_io_b),
    .io_z(inst_SnxnLv4Inst220_io_z)
  );
  SnxnLv4Inst221 inst_SnxnLv4Inst221 ( // @[Snxn100k.scala 15266:35]
    .io_a(inst_SnxnLv4Inst221_io_a),
    .io_b(inst_SnxnLv4Inst221_io_b),
    .io_z(inst_SnxnLv4Inst221_io_z)
  );
  SnxnLv4Inst77 inst_SnxnLv4Inst222 ( // @[Snxn100k.scala 15270:35]
    .io_a(inst_SnxnLv4Inst222_io_a),
    .io_b(inst_SnxnLv4Inst222_io_b),
    .io_z(inst_SnxnLv4Inst222_io_z)
  );
  SnxnLv4Inst223 inst_SnxnLv4Inst223 ( // @[Snxn100k.scala 15274:35]
    .io_a(inst_SnxnLv4Inst223_io_a),
    .io_b(inst_SnxnLv4Inst223_io_b),
    .io_z(inst_SnxnLv4Inst223_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 15279:15]
  assign inst_SnxnLv4Inst220_io_a = io_a; // @[Snxn100k.scala 15263:28]
  assign inst_SnxnLv4Inst220_io_b = io_b; // @[Snxn100k.scala 15264:28]
  assign inst_SnxnLv4Inst221_io_a = io_a; // @[Snxn100k.scala 15267:28]
  assign inst_SnxnLv4Inst221_io_b = io_b; // @[Snxn100k.scala 15268:28]
  assign inst_SnxnLv4Inst222_io_a = io_a; // @[Snxn100k.scala 15271:28]
  assign inst_SnxnLv4Inst222_io_b = io_b; // @[Snxn100k.scala 15272:28]
  assign inst_SnxnLv4Inst223_io_a = io_a; // @[Snxn100k.scala 15275:28]
  assign inst_SnxnLv4Inst223_io_b = io_b; // @[Snxn100k.scala 15276:28]
endmodule
module SnxnLv2Inst13(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst52_io_a; // @[Snxn100k.scala 3760:34]
  wire  inst_SnxnLv3Inst52_io_b; // @[Snxn100k.scala 3760:34]
  wire  inst_SnxnLv3Inst52_io_z; // @[Snxn100k.scala 3760:34]
  wire  inst_SnxnLv3Inst53_io_a; // @[Snxn100k.scala 3764:34]
  wire  inst_SnxnLv3Inst53_io_b; // @[Snxn100k.scala 3764:34]
  wire  inst_SnxnLv3Inst53_io_z; // @[Snxn100k.scala 3764:34]
  wire  inst_SnxnLv3Inst54_io_a; // @[Snxn100k.scala 3768:34]
  wire  inst_SnxnLv3Inst54_io_b; // @[Snxn100k.scala 3768:34]
  wire  inst_SnxnLv3Inst54_io_z; // @[Snxn100k.scala 3768:34]
  wire  inst_SnxnLv3Inst55_io_a; // @[Snxn100k.scala 3772:34]
  wire  inst_SnxnLv3Inst55_io_b; // @[Snxn100k.scala 3772:34]
  wire  inst_SnxnLv3Inst55_io_z; // @[Snxn100k.scala 3772:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst52_io_z + inst_SnxnLv3Inst53_io_z; // @[Snxn100k.scala 3776:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst54_io_z; // @[Snxn100k.scala 3776:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst55_io_z; // @[Snxn100k.scala 3776:89]
  SnxnLv3Inst52 inst_SnxnLv3Inst52 ( // @[Snxn100k.scala 3760:34]
    .io_a(inst_SnxnLv3Inst52_io_a),
    .io_b(inst_SnxnLv3Inst52_io_b),
    .io_z(inst_SnxnLv3Inst52_io_z)
  );
  SnxnLv3Inst53 inst_SnxnLv3Inst53 ( // @[Snxn100k.scala 3764:34]
    .io_a(inst_SnxnLv3Inst53_io_a),
    .io_b(inst_SnxnLv3Inst53_io_b),
    .io_z(inst_SnxnLv3Inst53_io_z)
  );
  SnxnLv3Inst54 inst_SnxnLv3Inst54 ( // @[Snxn100k.scala 3768:34]
    .io_a(inst_SnxnLv3Inst54_io_a),
    .io_b(inst_SnxnLv3Inst54_io_b),
    .io_z(inst_SnxnLv3Inst54_io_z)
  );
  SnxnLv3Inst55 inst_SnxnLv3Inst55 ( // @[Snxn100k.scala 3772:34]
    .io_a(inst_SnxnLv3Inst55_io_a),
    .io_b(inst_SnxnLv3Inst55_io_b),
    .io_z(inst_SnxnLv3Inst55_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 3777:15]
  assign inst_SnxnLv3Inst52_io_a = io_a; // @[Snxn100k.scala 3761:27]
  assign inst_SnxnLv3Inst52_io_b = io_b; // @[Snxn100k.scala 3762:27]
  assign inst_SnxnLv3Inst53_io_a = io_a; // @[Snxn100k.scala 3765:27]
  assign inst_SnxnLv3Inst53_io_b = io_b; // @[Snxn100k.scala 3766:27]
  assign inst_SnxnLv3Inst54_io_a = io_a; // @[Snxn100k.scala 3769:27]
  assign inst_SnxnLv3Inst54_io_b = io_b; // @[Snxn100k.scala 3770:27]
  assign inst_SnxnLv3Inst55_io_a = io_a; // @[Snxn100k.scala 3773:27]
  assign inst_SnxnLv3Inst55_io_b = io_b; // @[Snxn100k.scala 3774:27]
endmodule
module SnxnLv4Inst224(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  t0 = io_a + io_b; // @[Snxn100k.scala 61171:20]
  wire  inv0 = ~t0; // @[Snxn100k.scala 61172:15]
  wire  x0 = t0 ^ inv0; // @[Snxn100k.scala 61173:18]
  wire  invx0 = ~x0; // @[Snxn100k.scala 61174:15]
  wire  t1 = x0 + invx0; // @[Snxn100k.scala 61175:18]
  wire  inv1 = ~t1; // @[Snxn100k.scala 61176:15]
  wire  x1 = t1 ^ inv1; // @[Snxn100k.scala 61177:18]
  wire  invx1 = ~x1; // @[Snxn100k.scala 61178:15]
  wire  t2 = x1 + invx1; // @[Snxn100k.scala 61179:18]
  wire  inv2 = ~t2; // @[Snxn100k.scala 61180:15]
  wire  x2 = t2 ^ inv2; // @[Snxn100k.scala 61181:18]
  wire  invx2 = ~x2; // @[Snxn100k.scala 61182:15]
  wire  t3 = x2 + invx2; // @[Snxn100k.scala 61183:18]
  wire  inv3 = ~t3; // @[Snxn100k.scala 61184:15]
  wire  x3 = t3 ^ inv3; // @[Snxn100k.scala 61185:18]
  wire  invx3 = ~x3; // @[Snxn100k.scala 61186:15]
  wire  t4 = x3 + invx3; // @[Snxn100k.scala 61187:18]
  wire  inv4 = ~t4; // @[Snxn100k.scala 61188:15]
  wire  x4 = t4 ^ inv4; // @[Snxn100k.scala 61189:18]
  wire  invx4 = ~x4; // @[Snxn100k.scala 61190:15]
  wire  t5 = x4 + invx4; // @[Snxn100k.scala 61191:18]
  wire  inv5 = ~t5; // @[Snxn100k.scala 61192:15]
  wire  x5 = t5 ^ inv5; // @[Snxn100k.scala 61193:18]
  wire  invx5 = ~x5; // @[Snxn100k.scala 61194:15]
  wire  t6 = x5 + invx5; // @[Snxn100k.scala 61195:18]
  wire  inv6 = ~t6; // @[Snxn100k.scala 61196:15]
  wire  x6 = t6 ^ inv6; // @[Snxn100k.scala 61197:18]
  wire  invx6 = ~x6; // @[Snxn100k.scala 61198:15]
  wire  t7 = x6 + invx6; // @[Snxn100k.scala 61199:18]
  wire  inv7 = ~t7; // @[Snxn100k.scala 61200:15]
  wire  x7 = t7 ^ inv7; // @[Snxn100k.scala 61201:18]
  wire  invx7 = ~x7; // @[Snxn100k.scala 61202:15]
  wire  t8 = x7 + invx7; // @[Snxn100k.scala 61203:18]
  wire  inv8 = ~t8; // @[Snxn100k.scala 61204:15]
  wire  x8 = t8 ^ inv8; // @[Snxn100k.scala 61205:18]
  wire  invx8 = ~x8; // @[Snxn100k.scala 61206:15]
  wire  t9 = x8 + invx8; // @[Snxn100k.scala 61207:18]
  wire  inv9 = ~t9; // @[Snxn100k.scala 61208:15]
  wire  x9 = t9 ^ inv9; // @[Snxn100k.scala 61209:18]
  wire  invx9 = ~x9; // @[Snxn100k.scala 61210:15]
  wire  t10 = x9 + invx9; // @[Snxn100k.scala 61211:19]
  wire  inv10 = ~t10; // @[Snxn100k.scala 61212:16]
  wire  x10 = t10 ^ inv10; // @[Snxn100k.scala 61213:20]
  wire  invx10 = ~x10; // @[Snxn100k.scala 61214:16]
  wire  t11 = x10 + invx10; // @[Snxn100k.scala 61215:20]
  wire  inv11 = ~t11; // @[Snxn100k.scala 61216:16]
  wire  x11 = t11 ^ inv11; // @[Snxn100k.scala 61217:20]
  wire  invx11 = ~x11; // @[Snxn100k.scala 61218:16]
  wire  t12 = x11 + invx11; // @[Snxn100k.scala 61219:20]
  wire  inv12 = ~t12; // @[Snxn100k.scala 61220:16]
  wire  x12 = t12 ^ inv12; // @[Snxn100k.scala 61221:20]
  wire  invx12 = ~x12; // @[Snxn100k.scala 61222:16]
  wire  t13 = x12 + invx12; // @[Snxn100k.scala 61223:20]
  wire  inv13 = ~t13; // @[Snxn100k.scala 61224:16]
  wire  x13 = t13 ^ inv13; // @[Snxn100k.scala 61225:20]
  wire  invx13 = ~x13; // @[Snxn100k.scala 61226:16]
  wire  t14 = x13 + invx13; // @[Snxn100k.scala 61227:20]
  wire  inv14 = ~t14; // @[Snxn100k.scala 61228:16]
  wire  x14 = t14 ^ inv14; // @[Snxn100k.scala 61229:20]
  wire  invx14 = ~x14; // @[Snxn100k.scala 61230:16]
  wire  t15 = x14 + invx14; // @[Snxn100k.scala 61231:20]
  wire  inv15 = ~t15; // @[Snxn100k.scala 61232:16]
  wire  x15 = t15 ^ inv15; // @[Snxn100k.scala 61233:20]
  wire  invx15 = ~x15; // @[Snxn100k.scala 61234:16]
  wire  t16 = x15 + invx15; // @[Snxn100k.scala 61235:20]
  wire  inv16 = ~t16; // @[Snxn100k.scala 61236:16]
  wire  x16 = t16 ^ inv16; // @[Snxn100k.scala 61237:20]
  wire  invx16 = ~x16; // @[Snxn100k.scala 61238:16]
  wire  t17 = x16 + invx16; // @[Snxn100k.scala 61239:20]
  wire  inv17 = ~t17; // @[Snxn100k.scala 61240:16]
  wire  x17 = t17 ^ inv17; // @[Snxn100k.scala 61241:20]
  wire  invx17 = ~x17; // @[Snxn100k.scala 61242:16]
  wire  t18 = x17 + invx17; // @[Snxn100k.scala 61243:20]
  wire  inv18 = ~t18; // @[Snxn100k.scala 61244:16]
  wire  x18 = t18 ^ inv18; // @[Snxn100k.scala 61245:20]
  wire  invx18 = ~x18; // @[Snxn100k.scala 61246:16]
  wire  t19 = x18 + invx18; // @[Snxn100k.scala 61247:20]
  wire  inv19 = ~t19; // @[Snxn100k.scala 61248:16]
  wire  x19 = t19 ^ inv19; // @[Snxn100k.scala 61249:20]
  wire  invx19 = ~x19; // @[Snxn100k.scala 61250:16]
  wire  t20 = x19 + invx19; // @[Snxn100k.scala 61251:20]
  wire  inv20 = ~t20; // @[Snxn100k.scala 61252:16]
  wire  x20 = t20 ^ inv20; // @[Snxn100k.scala 61253:20]
  wire  invx20 = ~x20; // @[Snxn100k.scala 61254:16]
  wire  t21 = x20 + invx20; // @[Snxn100k.scala 61255:20]
  wire  inv21 = ~t21; // @[Snxn100k.scala 61256:16]
  wire  x21 = t21 ^ inv21; // @[Snxn100k.scala 61257:20]
  wire  invx21 = ~x21; // @[Snxn100k.scala 61258:16]
  wire  t22 = x21 + invx21; // @[Snxn100k.scala 61259:20]
  wire  inv22 = ~t22; // @[Snxn100k.scala 61260:16]
  wire  x22 = t22 ^ inv22; // @[Snxn100k.scala 61261:20]
  wire  invx22 = ~x22; // @[Snxn100k.scala 61262:16]
  wire  t23 = x22 + invx22; // @[Snxn100k.scala 61263:20]
  wire  inv23 = ~t23; // @[Snxn100k.scala 61264:16]
  wire  x23 = t23 ^ inv23; // @[Snxn100k.scala 61265:20]
  wire  invx23 = ~x23; // @[Snxn100k.scala 61266:16]
  wire  t24 = x23 + invx23; // @[Snxn100k.scala 61267:20]
  wire  inv24 = ~t24; // @[Snxn100k.scala 61268:16]
  wire  x24 = t24 ^ inv24; // @[Snxn100k.scala 61269:20]
  wire  invx24 = ~x24; // @[Snxn100k.scala 61270:16]
  wire  t25 = x24 + invx24; // @[Snxn100k.scala 61271:20]
  wire  inv25 = ~t25; // @[Snxn100k.scala 61272:16]
  wire  x25 = t25 ^ inv25; // @[Snxn100k.scala 61273:20]
  wire  invx25 = ~x25; // @[Snxn100k.scala 61274:16]
  wire  t26 = x25 + invx25; // @[Snxn100k.scala 61275:20]
  wire  inv26 = ~t26; // @[Snxn100k.scala 61276:16]
  wire  x26 = t26 ^ inv26; // @[Snxn100k.scala 61277:20]
  wire  invx26 = ~x26; // @[Snxn100k.scala 61278:16]
  wire  t27 = x26 + invx26; // @[Snxn100k.scala 61279:20]
  wire  inv27 = ~t27; // @[Snxn100k.scala 61280:16]
  wire  x27 = t27 ^ inv27; // @[Snxn100k.scala 61281:20]
  wire  invx27 = ~x27; // @[Snxn100k.scala 61282:16]
  wire  t28 = x27 + invx27; // @[Snxn100k.scala 61283:20]
  wire  inv28 = ~t28; // @[Snxn100k.scala 61284:16]
  wire  x28 = t28 ^ inv28; // @[Snxn100k.scala 61285:20]
  wire  invx28 = ~x28; // @[Snxn100k.scala 61286:16]
  wire  t29 = x28 + invx28; // @[Snxn100k.scala 61287:20]
  wire  inv29 = ~t29; // @[Snxn100k.scala 61288:16]
  wire  x29 = t29 ^ inv29; // @[Snxn100k.scala 61289:20]
  wire  invx29 = ~x29; // @[Snxn100k.scala 61290:16]
  wire  t30 = x29 + invx29; // @[Snxn100k.scala 61291:20]
  wire  inv30 = ~t30; // @[Snxn100k.scala 61292:16]
  wire  x30 = t30 ^ inv30; // @[Snxn100k.scala 61293:20]
  wire  invx30 = ~x30; // @[Snxn100k.scala 61294:16]
  wire  t31 = x30 + invx30; // @[Snxn100k.scala 61295:20]
  wire  inv31 = ~t31; // @[Snxn100k.scala 61296:16]
  wire  x31 = t31 ^ inv31; // @[Snxn100k.scala 61297:20]
  wire  invx31 = ~x31; // @[Snxn100k.scala 61298:16]
  wire  t32 = x31 + invx31; // @[Snxn100k.scala 61299:20]
  wire  inv32 = ~t32; // @[Snxn100k.scala 61300:16]
  wire  x32 = t32 ^ inv32; // @[Snxn100k.scala 61301:20]
  wire  invx32 = ~x32; // @[Snxn100k.scala 61302:16]
  wire  t33 = x32 + invx32; // @[Snxn100k.scala 61303:20]
  wire  inv33 = ~t33; // @[Snxn100k.scala 61304:16]
  wire  x33 = t33 ^ inv33; // @[Snxn100k.scala 61305:20]
  wire  invx33 = ~x33; // @[Snxn100k.scala 61306:16]
  wire  t34 = x33 + invx33; // @[Snxn100k.scala 61307:20]
  wire  inv34 = ~t34; // @[Snxn100k.scala 61308:16]
  wire  x34 = t34 ^ inv34; // @[Snxn100k.scala 61309:20]
  wire  invx34 = ~x34; // @[Snxn100k.scala 61310:16]
  wire  t35 = x34 + invx34; // @[Snxn100k.scala 61311:20]
  wire  inv35 = ~t35; // @[Snxn100k.scala 61312:16]
  wire  x35 = t35 ^ inv35; // @[Snxn100k.scala 61313:20]
  wire  invx35 = ~x35; // @[Snxn100k.scala 61314:16]
  wire  t36 = x35 + invx35; // @[Snxn100k.scala 61315:20]
  wire  inv36 = ~t36; // @[Snxn100k.scala 61316:16]
  wire  x36 = t36 ^ inv36; // @[Snxn100k.scala 61317:20]
  wire  invx36 = ~x36; // @[Snxn100k.scala 61318:16]
  wire  t37 = x36 + invx36; // @[Snxn100k.scala 61319:20]
  wire  inv37 = ~t37; // @[Snxn100k.scala 61320:16]
  wire  x37 = t37 ^ inv37; // @[Snxn100k.scala 61321:20]
  wire  invx37 = ~x37; // @[Snxn100k.scala 61322:16]
  wire  t38 = x37 + invx37; // @[Snxn100k.scala 61323:20]
  wire  inv38 = ~t38; // @[Snxn100k.scala 61324:16]
  wire  x38 = t38 ^ inv38; // @[Snxn100k.scala 61325:20]
  wire  invx38 = ~x38; // @[Snxn100k.scala 61326:16]
  wire  t39 = x38 + invx38; // @[Snxn100k.scala 61327:20]
  wire  inv39 = ~t39; // @[Snxn100k.scala 61328:16]
  wire  x39 = t39 ^ inv39; // @[Snxn100k.scala 61329:20]
  wire  invx39 = ~x39; // @[Snxn100k.scala 61330:16]
  wire  t40 = x39 + invx39; // @[Snxn100k.scala 61331:20]
  wire  inv40 = ~t40; // @[Snxn100k.scala 61332:16]
  wire  x40 = t40 ^ inv40; // @[Snxn100k.scala 61333:20]
  wire  invx40 = ~x40; // @[Snxn100k.scala 61334:16]
  wire  t41 = x40 + invx40; // @[Snxn100k.scala 61335:20]
  wire  inv41 = ~t41; // @[Snxn100k.scala 61336:16]
  wire  x41 = t41 ^ inv41; // @[Snxn100k.scala 61337:20]
  wire  invx41 = ~x41; // @[Snxn100k.scala 61338:16]
  wire  t42 = x41 + invx41; // @[Snxn100k.scala 61339:20]
  wire  inv42 = ~t42; // @[Snxn100k.scala 61340:16]
  wire  x42 = t42 ^ inv42; // @[Snxn100k.scala 61341:20]
  wire  invx42 = ~x42; // @[Snxn100k.scala 61342:16]
  wire  t43 = x42 + invx42; // @[Snxn100k.scala 61343:20]
  wire  inv43 = ~t43; // @[Snxn100k.scala 61344:16]
  wire  x43 = t43 ^ inv43; // @[Snxn100k.scala 61345:20]
  wire  invx43 = ~x43; // @[Snxn100k.scala 61346:16]
  wire  t44 = x43 + invx43; // @[Snxn100k.scala 61347:20]
  wire  inv44 = ~t44; // @[Snxn100k.scala 61348:16]
  wire  x44 = t44 ^ inv44; // @[Snxn100k.scala 61349:20]
  wire  invx44 = ~x44; // @[Snxn100k.scala 61350:16]
  wire  t45 = x44 + invx44; // @[Snxn100k.scala 61351:20]
  wire  inv45 = ~t45; // @[Snxn100k.scala 61352:16]
  wire  x45 = t45 ^ inv45; // @[Snxn100k.scala 61353:20]
  wire  invx45 = ~x45; // @[Snxn100k.scala 61354:16]
  wire  t46 = x45 + invx45; // @[Snxn100k.scala 61355:20]
  wire  inv46 = ~t46; // @[Snxn100k.scala 61356:16]
  wire  x46 = t46 ^ inv46; // @[Snxn100k.scala 61357:20]
  wire  invx46 = ~x46; // @[Snxn100k.scala 61358:16]
  wire  t47 = x46 + invx46; // @[Snxn100k.scala 61359:20]
  wire  inv47 = ~t47; // @[Snxn100k.scala 61360:16]
  wire  x47 = t47 ^ inv47; // @[Snxn100k.scala 61361:20]
  wire  invx47 = ~x47; // @[Snxn100k.scala 61362:16]
  wire  t48 = x47 + invx47; // @[Snxn100k.scala 61363:20]
  wire  inv48 = ~t48; // @[Snxn100k.scala 61364:16]
  wire  x48 = t48 ^ inv48; // @[Snxn100k.scala 61365:20]
  wire  invx48 = ~x48; // @[Snxn100k.scala 61366:16]
  wire  t49 = x48 + invx48; // @[Snxn100k.scala 61367:20]
  wire  inv49 = ~t49; // @[Snxn100k.scala 61368:16]
  wire  x49 = t49 ^ inv49; // @[Snxn100k.scala 61369:20]
  wire  invx49 = ~x49; // @[Snxn100k.scala 61370:16]
  wire  t50 = x49 + invx49; // @[Snxn100k.scala 61371:20]
  wire  inv50 = ~t50; // @[Snxn100k.scala 61372:16]
  wire  x50 = t50 ^ inv50; // @[Snxn100k.scala 61373:20]
  wire  invx50 = ~x50; // @[Snxn100k.scala 61374:16]
  wire  t51 = x50 + invx50; // @[Snxn100k.scala 61375:20]
  wire  inv51 = ~t51; // @[Snxn100k.scala 61376:16]
  wire  x51 = t51 ^ inv51; // @[Snxn100k.scala 61377:20]
  wire  invx51 = ~x51; // @[Snxn100k.scala 61378:16]
  wire  t52 = x51 + invx51; // @[Snxn100k.scala 61379:20]
  wire  inv52 = ~t52; // @[Snxn100k.scala 61380:16]
  wire  x52 = t52 ^ inv52; // @[Snxn100k.scala 61381:20]
  wire  invx52 = ~x52; // @[Snxn100k.scala 61382:16]
  wire  t53 = x52 + invx52; // @[Snxn100k.scala 61383:20]
  wire  inv53 = ~t53; // @[Snxn100k.scala 61384:16]
  wire  x53 = t53 ^ inv53; // @[Snxn100k.scala 61385:20]
  wire  invx53 = ~x53; // @[Snxn100k.scala 61386:16]
  wire  t54 = x53 + invx53; // @[Snxn100k.scala 61387:20]
  wire  inv54 = ~t54; // @[Snxn100k.scala 61388:16]
  wire  x54 = t54 ^ inv54; // @[Snxn100k.scala 61389:20]
  wire  invx54 = ~x54; // @[Snxn100k.scala 61390:16]
  wire  t55 = x54 + invx54; // @[Snxn100k.scala 61391:20]
  wire  inv55 = ~t55; // @[Snxn100k.scala 61392:16]
  wire  x55 = t55 ^ inv55; // @[Snxn100k.scala 61393:20]
  wire  invx55 = ~x55; // @[Snxn100k.scala 61394:16]
  wire  t56 = x55 + invx55; // @[Snxn100k.scala 61395:20]
  wire  inv56 = ~t56; // @[Snxn100k.scala 61396:16]
  wire  x56 = t56 ^ inv56; // @[Snxn100k.scala 61397:20]
  wire  invx56 = ~x56; // @[Snxn100k.scala 61398:16]
  wire  t57 = x56 + invx56; // @[Snxn100k.scala 61399:20]
  wire  inv57 = ~t57; // @[Snxn100k.scala 61400:16]
  wire  x57 = t57 ^ inv57; // @[Snxn100k.scala 61401:20]
  wire  invx57 = ~x57; // @[Snxn100k.scala 61402:16]
  wire  t58 = x57 + invx57; // @[Snxn100k.scala 61403:20]
  wire  inv58 = ~t58; // @[Snxn100k.scala 61404:16]
  wire  x58 = t58 ^ inv58; // @[Snxn100k.scala 61405:20]
  wire  invx58 = ~x58; // @[Snxn100k.scala 61406:16]
  wire  t59 = x58 + invx58; // @[Snxn100k.scala 61407:20]
  wire  inv59 = ~t59; // @[Snxn100k.scala 61408:16]
  wire  x59 = t59 ^ inv59; // @[Snxn100k.scala 61409:20]
  wire  invx59 = ~x59; // @[Snxn100k.scala 61410:16]
  wire  t60 = x59 + invx59; // @[Snxn100k.scala 61411:20]
  wire  inv60 = ~t60; // @[Snxn100k.scala 61412:16]
  wire  x60 = t60 ^ inv60; // @[Snxn100k.scala 61413:20]
  wire  invx60 = ~x60; // @[Snxn100k.scala 61414:16]
  wire  t61 = x60 + invx60; // @[Snxn100k.scala 61415:20]
  wire  inv61 = ~t61; // @[Snxn100k.scala 61416:16]
  wire  x61 = t61 ^ inv61; // @[Snxn100k.scala 61417:20]
  wire  invx61 = ~x61; // @[Snxn100k.scala 61418:16]
  wire  t62 = x61 + invx61; // @[Snxn100k.scala 61419:20]
  wire  inv62 = ~t62; // @[Snxn100k.scala 61420:16]
  wire  x62 = t62 ^ inv62; // @[Snxn100k.scala 61421:20]
  wire  invx62 = ~x62; // @[Snxn100k.scala 61422:16]
  wire  t63 = x62 + invx62; // @[Snxn100k.scala 61423:20]
  wire  inv63 = ~t63; // @[Snxn100k.scala 61424:16]
  wire  x63 = t63 ^ inv63; // @[Snxn100k.scala 61425:20]
  wire  invx63 = ~x63; // @[Snxn100k.scala 61426:16]
  wire  t64 = x63 + invx63; // @[Snxn100k.scala 61427:20]
  wire  inv64 = ~t64; // @[Snxn100k.scala 61428:16]
  wire  x64 = t64 ^ inv64; // @[Snxn100k.scala 61429:20]
  wire  invx64 = ~x64; // @[Snxn100k.scala 61430:16]
  wire  t65 = x64 + invx64; // @[Snxn100k.scala 61431:20]
  wire  inv65 = ~t65; // @[Snxn100k.scala 61432:16]
  wire  x65 = t65 ^ inv65; // @[Snxn100k.scala 61433:20]
  wire  invx65 = ~x65; // @[Snxn100k.scala 61434:16]
  wire  t66 = x65 + invx65; // @[Snxn100k.scala 61435:20]
  wire  inv66 = ~t66; // @[Snxn100k.scala 61436:16]
  wire  x66 = t66 ^ inv66; // @[Snxn100k.scala 61437:20]
  wire  invx66 = ~x66; // @[Snxn100k.scala 61438:16]
  wire  t67 = x66 + invx66; // @[Snxn100k.scala 61439:20]
  wire  inv67 = ~t67; // @[Snxn100k.scala 61440:16]
  wire  x67 = t67 ^ inv67; // @[Snxn100k.scala 61441:20]
  wire  invx67 = ~x67; // @[Snxn100k.scala 61442:16]
  wire  t68 = x67 + invx67; // @[Snxn100k.scala 61443:20]
  wire  inv68 = ~t68; // @[Snxn100k.scala 61444:16]
  wire  x68 = t68 ^ inv68; // @[Snxn100k.scala 61445:20]
  wire  invx68 = ~x68; // @[Snxn100k.scala 61446:16]
  wire  t69 = x68 + invx68; // @[Snxn100k.scala 61447:20]
  wire  inv69 = ~t69; // @[Snxn100k.scala 61448:16]
  wire  x69 = t69 ^ inv69; // @[Snxn100k.scala 61449:20]
  wire  invx69 = ~x69; // @[Snxn100k.scala 61450:16]
  wire  t70 = x69 + invx69; // @[Snxn100k.scala 61451:20]
  wire  inv70 = ~t70; // @[Snxn100k.scala 61452:16]
  wire  x70 = t70 ^ inv70; // @[Snxn100k.scala 61453:20]
  wire  invx70 = ~x70; // @[Snxn100k.scala 61454:16]
  wire  t71 = x70 + invx70; // @[Snxn100k.scala 61455:20]
  wire  inv71 = ~t71; // @[Snxn100k.scala 61456:16]
  wire  x71 = t71 ^ inv71; // @[Snxn100k.scala 61457:20]
  wire  invx71 = ~x71; // @[Snxn100k.scala 61458:16]
  wire  t72 = x71 + invx71; // @[Snxn100k.scala 61459:20]
  wire  inv72 = ~t72; // @[Snxn100k.scala 61460:16]
  wire  x72 = t72 ^ inv72; // @[Snxn100k.scala 61461:20]
  wire  invx72 = ~x72; // @[Snxn100k.scala 61462:16]
  wire  t73 = x72 + invx72; // @[Snxn100k.scala 61463:20]
  wire  inv73 = ~t73; // @[Snxn100k.scala 61464:16]
  wire  x73 = t73 ^ inv73; // @[Snxn100k.scala 61465:20]
  wire  invx73 = ~x73; // @[Snxn100k.scala 61466:16]
  wire  t74 = x73 + invx73; // @[Snxn100k.scala 61467:20]
  wire  inv74 = ~t74; // @[Snxn100k.scala 61468:16]
  wire  x74 = t74 ^ inv74; // @[Snxn100k.scala 61469:20]
  wire  invx74 = ~x74; // @[Snxn100k.scala 61470:16]
  wire  t75 = x74 + invx74; // @[Snxn100k.scala 61471:20]
  wire  inv75 = ~t75; // @[Snxn100k.scala 61472:16]
  wire  x75 = t75 ^ inv75; // @[Snxn100k.scala 61473:20]
  wire  invx75 = ~x75; // @[Snxn100k.scala 61474:16]
  wire  t76 = x75 + invx75; // @[Snxn100k.scala 61475:20]
  wire  inv76 = ~t76; // @[Snxn100k.scala 61476:16]
  wire  x76 = t76 ^ inv76; // @[Snxn100k.scala 61477:20]
  wire  invx76 = ~x76; // @[Snxn100k.scala 61478:16]
  wire  t77 = x76 + invx76; // @[Snxn100k.scala 61479:20]
  wire  inv77 = ~t77; // @[Snxn100k.scala 61480:16]
  wire  x77 = t77 ^ inv77; // @[Snxn100k.scala 61481:20]
  wire  invx77 = ~x77; // @[Snxn100k.scala 61482:16]
  wire  t78 = x77 + invx77; // @[Snxn100k.scala 61483:20]
  wire  inv78 = ~t78; // @[Snxn100k.scala 61484:16]
  wire  x78 = t78 ^ inv78; // @[Snxn100k.scala 61485:20]
  wire  invx78 = ~x78; // @[Snxn100k.scala 61486:16]
  wire  t79 = x78 + invx78; // @[Snxn100k.scala 61487:20]
  wire  inv79 = ~t79; // @[Snxn100k.scala 61488:16]
  wire  x79 = t79 ^ inv79; // @[Snxn100k.scala 61489:20]
  wire  invx79 = ~x79; // @[Snxn100k.scala 61490:16]
  wire  t80 = x79 + invx79; // @[Snxn100k.scala 61491:20]
  wire  inv80 = ~t80; // @[Snxn100k.scala 61492:16]
  wire  x80 = t80 ^ inv80; // @[Snxn100k.scala 61493:20]
  wire  invx80 = ~x80; // @[Snxn100k.scala 61494:16]
  wire  t81 = x80 + invx80; // @[Snxn100k.scala 61495:20]
  wire  inv81 = ~t81; // @[Snxn100k.scala 61496:16]
  wire  x81 = t81 ^ inv81; // @[Snxn100k.scala 61497:20]
  wire  invx81 = ~x81; // @[Snxn100k.scala 61498:16]
  wire  t82 = x81 + invx81; // @[Snxn100k.scala 61499:20]
  wire  inv82 = ~t82; // @[Snxn100k.scala 61500:16]
  wire  x82 = t82 ^ inv82; // @[Snxn100k.scala 61501:20]
  wire  invx82 = ~x82; // @[Snxn100k.scala 61502:16]
  wire  t83 = x82 + invx82; // @[Snxn100k.scala 61503:20]
  wire  inv83 = ~t83; // @[Snxn100k.scala 61504:16]
  wire  x83 = t83 ^ inv83; // @[Snxn100k.scala 61505:20]
  wire  invx83 = ~x83; // @[Snxn100k.scala 61506:16]
  wire  t84 = x83 + invx83; // @[Snxn100k.scala 61507:20]
  wire  inv84 = ~t84; // @[Snxn100k.scala 61508:16]
  wire  x84 = t84 ^ inv84; // @[Snxn100k.scala 61509:20]
  assign io_z = ~x84; // @[Snxn100k.scala 61510:16]
endmodule
module SnxnLv3Inst56(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst224_io_a; // @[Snxn100k.scala 17952:35]
  wire  inst_SnxnLv4Inst224_io_b; // @[Snxn100k.scala 17952:35]
  wire  inst_SnxnLv4Inst224_io_z; // @[Snxn100k.scala 17952:35]
  wire  inst_SnxnLv4Inst225_io_a; // @[Snxn100k.scala 17956:35]
  wire  inst_SnxnLv4Inst225_io_b; // @[Snxn100k.scala 17956:35]
  wire  inst_SnxnLv4Inst225_io_z; // @[Snxn100k.scala 17956:35]
  wire  inst_SnxnLv4Inst226_io_a; // @[Snxn100k.scala 17960:35]
  wire  inst_SnxnLv4Inst226_io_b; // @[Snxn100k.scala 17960:35]
  wire  inst_SnxnLv4Inst226_io_z; // @[Snxn100k.scala 17960:35]
  wire  inst_SnxnLv4Inst227_io_a; // @[Snxn100k.scala 17964:35]
  wire  inst_SnxnLv4Inst227_io_b; // @[Snxn100k.scala 17964:35]
  wire  inst_SnxnLv4Inst227_io_z; // @[Snxn100k.scala 17964:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst224_io_z + inst_SnxnLv4Inst225_io_z; // @[Snxn100k.scala 17968:38]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv4Inst226_io_z; // @[Snxn100k.scala 17968:65]
  wire  sum = _sum_T_3 + inst_SnxnLv4Inst227_io_z; // @[Snxn100k.scala 17968:92]
  SnxnLv4Inst224 inst_SnxnLv4Inst224 ( // @[Snxn100k.scala 17952:35]
    .io_a(inst_SnxnLv4Inst224_io_a),
    .io_b(inst_SnxnLv4Inst224_io_b),
    .io_z(inst_SnxnLv4Inst224_io_z)
  );
  SnxnLv4Inst95 inst_SnxnLv4Inst225 ( // @[Snxn100k.scala 17956:35]
    .io_a(inst_SnxnLv4Inst225_io_a),
    .io_b(inst_SnxnLv4Inst225_io_b),
    .io_z(inst_SnxnLv4Inst225_io_z)
  );
  SnxnLv4Inst33 inst_SnxnLv4Inst226 ( // @[Snxn100k.scala 17960:35]
    .io_a(inst_SnxnLv4Inst226_io_a),
    .io_b(inst_SnxnLv4Inst226_io_b),
    .io_z(inst_SnxnLv4Inst226_io_z)
  );
  SnxnLv4Inst101 inst_SnxnLv4Inst227 ( // @[Snxn100k.scala 17964:35]
    .io_a(inst_SnxnLv4Inst227_io_a),
    .io_b(inst_SnxnLv4Inst227_io_b),
    .io_z(inst_SnxnLv4Inst227_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 17969:15]
  assign inst_SnxnLv4Inst224_io_a = io_a; // @[Snxn100k.scala 17953:28]
  assign inst_SnxnLv4Inst224_io_b = io_b; // @[Snxn100k.scala 17954:28]
  assign inst_SnxnLv4Inst225_io_a = io_a; // @[Snxn100k.scala 17957:28]
  assign inst_SnxnLv4Inst225_io_b = io_b; // @[Snxn100k.scala 17958:28]
  assign inst_SnxnLv4Inst226_io_a = io_a; // @[Snxn100k.scala 17961:28]
  assign inst_SnxnLv4Inst226_io_b = io_b; // @[Snxn100k.scala 17962:28]
  assign inst_SnxnLv4Inst227_io_a = io_a; // @[Snxn100k.scala 17965:28]
  assign inst_SnxnLv4Inst227_io_b = io_b; // @[Snxn100k.scala 17966:28]
endmodule
module SnxnLv3Inst57(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv4Inst228_io_a; // @[Snxn100k.scala 18367:35]
  wire  inst_SnxnLv4Inst228_io_b; // @[Snxn100k.scala 18367:35]
  wire  inst_SnxnLv4Inst228_io_z; // @[Snxn100k.scala 18367:35]
  wire  inst_SnxnLv4Inst229_io_a; // @[Snxn100k.scala 18371:35]
  wire  inst_SnxnLv4Inst229_io_b; // @[Snxn100k.scala 18371:35]
  wire  inst_SnxnLv4Inst229_io_z; // @[Snxn100k.scala 18371:35]
  wire  inst_SnxnLv4Inst230_io_a; // @[Snxn100k.scala 18375:35]
  wire  inst_SnxnLv4Inst230_io_b; // @[Snxn100k.scala 18375:35]
  wire  inst_SnxnLv4Inst230_io_z; // @[Snxn100k.scala 18375:35]
  wire  _sum_T_1 = inst_SnxnLv4Inst228_io_z + inst_SnxnLv4Inst229_io_z; // @[Snxn100k.scala 18379:38]
  wire  sum = _sum_T_1 + inst_SnxnLv4Inst230_io_z; // @[Snxn100k.scala 18379:65]
  SnxnLv4Inst44 inst_SnxnLv4Inst228 ( // @[Snxn100k.scala 18367:35]
    .io_a(inst_SnxnLv4Inst228_io_a),
    .io_b(inst_SnxnLv4Inst228_io_b),
    .io_z(inst_SnxnLv4Inst228_io_z)
  );
  SnxnLv4Inst154 inst_SnxnLv4Inst229 ( // @[Snxn100k.scala 18371:35]
    .io_a(inst_SnxnLv4Inst229_io_a),
    .io_b(inst_SnxnLv4Inst229_io_b),
    .io_z(inst_SnxnLv4Inst229_io_z)
  );
  SnxnLv4Inst152 inst_SnxnLv4Inst230 ( // @[Snxn100k.scala 18375:35]
    .io_a(inst_SnxnLv4Inst230_io_a),
    .io_b(inst_SnxnLv4Inst230_io_b),
    .io_z(inst_SnxnLv4Inst230_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 18380:15]
  assign inst_SnxnLv4Inst228_io_a = io_a; // @[Snxn100k.scala 18368:28]
  assign inst_SnxnLv4Inst228_io_b = io_b; // @[Snxn100k.scala 18369:28]
  assign inst_SnxnLv4Inst229_io_a = io_a; // @[Snxn100k.scala 18372:28]
  assign inst_SnxnLv4Inst229_io_b = io_b; // @[Snxn100k.scala 18373:28]
  assign inst_SnxnLv4Inst230_io_a = io_a; // @[Snxn100k.scala 18376:28]
  assign inst_SnxnLv4Inst230_io_b = io_b; // @[Snxn100k.scala 18377:28]
endmodule
module SnxnLv2Inst14(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst56_io_a; // @[Snxn100k.scala 4806:34]
  wire  inst_SnxnLv3Inst56_io_b; // @[Snxn100k.scala 4806:34]
  wire  inst_SnxnLv3Inst56_io_z; // @[Snxn100k.scala 4806:34]
  wire  inst_SnxnLv3Inst57_io_a; // @[Snxn100k.scala 4810:34]
  wire  inst_SnxnLv3Inst57_io_b; // @[Snxn100k.scala 4810:34]
  wire  inst_SnxnLv3Inst57_io_z; // @[Snxn100k.scala 4810:34]
  wire  inst_SnxnLv3Inst58_io_a; // @[Snxn100k.scala 4814:34]
  wire  inst_SnxnLv3Inst58_io_b; // @[Snxn100k.scala 4814:34]
  wire  inst_SnxnLv3Inst58_io_z; // @[Snxn100k.scala 4814:34]
  wire  inst_SnxnLv3Inst59_io_a; // @[Snxn100k.scala 4818:34]
  wire  inst_SnxnLv3Inst59_io_b; // @[Snxn100k.scala 4818:34]
  wire  inst_SnxnLv3Inst59_io_z; // @[Snxn100k.scala 4818:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst56_io_z + inst_SnxnLv3Inst57_io_z; // @[Snxn100k.scala 4822:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst58_io_z; // @[Snxn100k.scala 4822:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst59_io_z; // @[Snxn100k.scala 4822:89]
  SnxnLv3Inst56 inst_SnxnLv3Inst56 ( // @[Snxn100k.scala 4806:34]
    .io_a(inst_SnxnLv3Inst56_io_a),
    .io_b(inst_SnxnLv3Inst56_io_b),
    .io_z(inst_SnxnLv3Inst56_io_z)
  );
  SnxnLv3Inst57 inst_SnxnLv3Inst57 ( // @[Snxn100k.scala 4810:34]
    .io_a(inst_SnxnLv3Inst57_io_a),
    .io_b(inst_SnxnLv3Inst57_io_b),
    .io_z(inst_SnxnLv3Inst57_io_z)
  );
  SnxnLv4Inst51 inst_SnxnLv3Inst58 ( // @[Snxn100k.scala 4814:34]
    .io_a(inst_SnxnLv3Inst58_io_a),
    .io_b(inst_SnxnLv3Inst58_io_b),
    .io_z(inst_SnxnLv3Inst58_io_z)
  );
  SnxnLv4Inst67 inst_SnxnLv3Inst59 ( // @[Snxn100k.scala 4818:34]
    .io_a(inst_SnxnLv3Inst59_io_a),
    .io_b(inst_SnxnLv3Inst59_io_b),
    .io_z(inst_SnxnLv3Inst59_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 4823:15]
  assign inst_SnxnLv3Inst56_io_a = io_a; // @[Snxn100k.scala 4807:27]
  assign inst_SnxnLv3Inst56_io_b = io_b; // @[Snxn100k.scala 4808:27]
  assign inst_SnxnLv3Inst57_io_a = io_a; // @[Snxn100k.scala 4811:27]
  assign inst_SnxnLv3Inst57_io_b = io_b; // @[Snxn100k.scala 4812:27]
  assign inst_SnxnLv3Inst58_io_a = io_a; // @[Snxn100k.scala 4815:27]
  assign inst_SnxnLv3Inst58_io_b = io_b; // @[Snxn100k.scala 4816:27]
  assign inst_SnxnLv3Inst59_io_a = io_a; // @[Snxn100k.scala 4819:27]
  assign inst_SnxnLv3Inst59_io_b = io_b; // @[Snxn100k.scala 4820:27]
endmodule
module SnxnLv2Inst15(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv3Inst60_io_a; // @[Snxn100k.scala 5361:34]
  wire  inst_SnxnLv3Inst60_io_b; // @[Snxn100k.scala 5361:34]
  wire  inst_SnxnLv3Inst60_io_z; // @[Snxn100k.scala 5361:34]
  wire  inst_SnxnLv3Inst61_io_a; // @[Snxn100k.scala 5365:34]
  wire  inst_SnxnLv3Inst61_io_b; // @[Snxn100k.scala 5365:34]
  wire  inst_SnxnLv3Inst61_io_z; // @[Snxn100k.scala 5365:34]
  wire  inst_SnxnLv3Inst62_io_a; // @[Snxn100k.scala 5369:34]
  wire  inst_SnxnLv3Inst62_io_b; // @[Snxn100k.scala 5369:34]
  wire  inst_SnxnLv3Inst62_io_z; // @[Snxn100k.scala 5369:34]
  wire  inst_SnxnLv3Inst63_io_a; // @[Snxn100k.scala 5373:34]
  wire  inst_SnxnLv3Inst63_io_b; // @[Snxn100k.scala 5373:34]
  wire  inst_SnxnLv3Inst63_io_z; // @[Snxn100k.scala 5373:34]
  wire  _sum_T_1 = inst_SnxnLv3Inst60_io_z + inst_SnxnLv3Inst61_io_z; // @[Snxn100k.scala 5377:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv3Inst62_io_z; // @[Snxn100k.scala 5377:63]
  wire  sum = _sum_T_3 + inst_SnxnLv3Inst63_io_z; // @[Snxn100k.scala 5377:89]
  SnxnLv4Inst67 inst_SnxnLv3Inst60 ( // @[Snxn100k.scala 5361:34]
    .io_a(inst_SnxnLv3Inst60_io_a),
    .io_b(inst_SnxnLv3Inst60_io_b),
    .io_z(inst_SnxnLv3Inst60_io_z)
  );
  SnxnLv4Inst8 inst_SnxnLv3Inst61 ( // @[Snxn100k.scala 5365:34]
    .io_a(inst_SnxnLv3Inst61_io_a),
    .io_b(inst_SnxnLv3Inst61_io_b),
    .io_z(inst_SnxnLv3Inst61_io_z)
  );
  SnxnLv4Inst72 inst_SnxnLv3Inst62 ( // @[Snxn100k.scala 5369:34]
    .io_a(inst_SnxnLv3Inst62_io_a),
    .io_b(inst_SnxnLv3Inst62_io_b),
    .io_z(inst_SnxnLv3Inst62_io_z)
  );
  SnxnLv4Inst59 inst_SnxnLv3Inst63 ( // @[Snxn100k.scala 5373:34]
    .io_a(inst_SnxnLv3Inst63_io_a),
    .io_b(inst_SnxnLv3Inst63_io_b),
    .io_z(inst_SnxnLv3Inst63_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 5378:15]
  assign inst_SnxnLv3Inst60_io_a = io_a; // @[Snxn100k.scala 5362:27]
  assign inst_SnxnLv3Inst60_io_b = io_b; // @[Snxn100k.scala 5363:27]
  assign inst_SnxnLv3Inst61_io_a = io_a; // @[Snxn100k.scala 5366:27]
  assign inst_SnxnLv3Inst61_io_b = io_b; // @[Snxn100k.scala 5367:27]
  assign inst_SnxnLv3Inst62_io_a = io_a; // @[Snxn100k.scala 5370:27]
  assign inst_SnxnLv3Inst62_io_b = io_b; // @[Snxn100k.scala 5371:27]
  assign inst_SnxnLv3Inst63_io_a = io_a; // @[Snxn100k.scala 5374:27]
  assign inst_SnxnLv3Inst63_io_b = io_b; // @[Snxn100k.scala 5375:27]
endmodule
module SnxnLv1Inst3(
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv2Inst12_io_a; // @[Snxn100k.scala 671:34]
  wire  inst_SnxnLv2Inst12_io_b; // @[Snxn100k.scala 671:34]
  wire  inst_SnxnLv2Inst12_io_z; // @[Snxn100k.scala 671:34]
  wire  inst_SnxnLv2Inst13_io_a; // @[Snxn100k.scala 675:34]
  wire  inst_SnxnLv2Inst13_io_b; // @[Snxn100k.scala 675:34]
  wire  inst_SnxnLv2Inst13_io_z; // @[Snxn100k.scala 675:34]
  wire  inst_SnxnLv2Inst14_io_a; // @[Snxn100k.scala 679:34]
  wire  inst_SnxnLv2Inst14_io_b; // @[Snxn100k.scala 679:34]
  wire  inst_SnxnLv2Inst14_io_z; // @[Snxn100k.scala 679:34]
  wire  inst_SnxnLv2Inst15_io_a; // @[Snxn100k.scala 683:34]
  wire  inst_SnxnLv2Inst15_io_b; // @[Snxn100k.scala 683:34]
  wire  inst_SnxnLv2Inst15_io_z; // @[Snxn100k.scala 683:34]
  wire  _sum_T_1 = inst_SnxnLv2Inst12_io_z + inst_SnxnLv2Inst13_io_z; // @[Snxn100k.scala 687:37]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv2Inst14_io_z; // @[Snxn100k.scala 687:63]
  wire  sum = _sum_T_3 + inst_SnxnLv2Inst15_io_z; // @[Snxn100k.scala 687:89]
  SnxnLv2Inst12 inst_SnxnLv2Inst12 ( // @[Snxn100k.scala 671:34]
    .io_a(inst_SnxnLv2Inst12_io_a),
    .io_b(inst_SnxnLv2Inst12_io_b),
    .io_z(inst_SnxnLv2Inst12_io_z)
  );
  SnxnLv2Inst13 inst_SnxnLv2Inst13 ( // @[Snxn100k.scala 675:34]
    .io_a(inst_SnxnLv2Inst13_io_a),
    .io_b(inst_SnxnLv2Inst13_io_b),
    .io_z(inst_SnxnLv2Inst13_io_z)
  );
  SnxnLv2Inst14 inst_SnxnLv2Inst14 ( // @[Snxn100k.scala 679:34]
    .io_a(inst_SnxnLv2Inst14_io_a),
    .io_b(inst_SnxnLv2Inst14_io_b),
    .io_z(inst_SnxnLv2Inst14_io_z)
  );
  SnxnLv2Inst15 inst_SnxnLv2Inst15 ( // @[Snxn100k.scala 683:34]
    .io_a(inst_SnxnLv2Inst15_io_a),
    .io_b(inst_SnxnLv2Inst15_io_b),
    .io_z(inst_SnxnLv2Inst15_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 688:15]
  assign inst_SnxnLv2Inst12_io_a = io_a; // @[Snxn100k.scala 672:27]
  assign inst_SnxnLv2Inst12_io_b = io_b; // @[Snxn100k.scala 673:27]
  assign inst_SnxnLv2Inst13_io_a = io_a; // @[Snxn100k.scala 676:27]
  assign inst_SnxnLv2Inst13_io_b = io_b; // @[Snxn100k.scala 677:27]
  assign inst_SnxnLv2Inst14_io_a = io_a; // @[Snxn100k.scala 680:27]
  assign inst_SnxnLv2Inst14_io_b = io_b; // @[Snxn100k.scala 681:27]
  assign inst_SnxnLv2Inst15_io_a = io_a; // @[Snxn100k.scala 684:27]
  assign inst_SnxnLv2Inst15_io_b = io_b; // @[Snxn100k.scala 685:27]
endmodule
module Snxn100k(
  input   clock,
  input   reset,
  input   io_a,
  input   io_b,
  output  io_z
);
  wire  inst_SnxnLv1Inst0_io_a; // @[Snxn100k.scala 473:33]
  wire  inst_SnxnLv1Inst0_io_b; // @[Snxn100k.scala 473:33]
  wire  inst_SnxnLv1Inst0_io_z; // @[Snxn100k.scala 473:33]
  wire  inst_SnxnLv1Inst1_io_a; // @[Snxn100k.scala 477:33]
  wire  inst_SnxnLv1Inst1_io_b; // @[Snxn100k.scala 477:33]
  wire  inst_SnxnLv1Inst1_io_z; // @[Snxn100k.scala 477:33]
  wire  inst_SnxnLv1Inst2_io_a; // @[Snxn100k.scala 481:33]
  wire  inst_SnxnLv1Inst2_io_b; // @[Snxn100k.scala 481:33]
  wire  inst_SnxnLv1Inst2_io_z; // @[Snxn100k.scala 481:33]
  wire  inst_SnxnLv1Inst3_io_a; // @[Snxn100k.scala 485:33]
  wire  inst_SnxnLv1Inst3_io_b; // @[Snxn100k.scala 485:33]
  wire  inst_SnxnLv1Inst3_io_z; // @[Snxn100k.scala 485:33]
  wire  _sum_T_1 = inst_SnxnLv1Inst0_io_z + inst_SnxnLv1Inst1_io_z; // @[Snxn100k.scala 489:36]
  wire  _sum_T_3 = _sum_T_1 + inst_SnxnLv1Inst2_io_z; // @[Snxn100k.scala 489:61]
  wire  sum = _sum_T_3 + inst_SnxnLv1Inst3_io_z; // @[Snxn100k.scala 489:86]
  SnxnLv1Inst0 inst_SnxnLv1Inst0 ( // @[Snxn100k.scala 473:33]
    .io_a(inst_SnxnLv1Inst0_io_a),
    .io_b(inst_SnxnLv1Inst0_io_b),
    .io_z(inst_SnxnLv1Inst0_io_z)
  );
  SnxnLv1Inst1 inst_SnxnLv1Inst1 ( // @[Snxn100k.scala 477:33]
    .io_a(inst_SnxnLv1Inst1_io_a),
    .io_b(inst_SnxnLv1Inst1_io_b),
    .io_z(inst_SnxnLv1Inst1_io_z)
  );
  SnxnLv1Inst2 inst_SnxnLv1Inst2 ( // @[Snxn100k.scala 481:33]
    .io_a(inst_SnxnLv1Inst2_io_a),
    .io_b(inst_SnxnLv1Inst2_io_b),
    .io_z(inst_SnxnLv1Inst2_io_z)
  );
  SnxnLv1Inst3 inst_SnxnLv1Inst3 ( // @[Snxn100k.scala 485:33]
    .io_a(inst_SnxnLv1Inst3_io_a),
    .io_b(inst_SnxnLv1Inst3_io_b),
    .io_z(inst_SnxnLv1Inst3_io_z)
  );
  assign io_z = sum ^ io_a; // @[Snxn100k.scala 490:15]
  assign inst_SnxnLv1Inst0_io_a = io_a; // @[Snxn100k.scala 474:26]
  assign inst_SnxnLv1Inst0_io_b = io_b; // @[Snxn100k.scala 475:26]
  assign inst_SnxnLv1Inst1_io_a = io_a; // @[Snxn100k.scala 478:26]
  assign inst_SnxnLv1Inst1_io_b = io_b; // @[Snxn100k.scala 479:26]
  assign inst_SnxnLv1Inst2_io_a = io_a; // @[Snxn100k.scala 482:26]
  assign inst_SnxnLv1Inst2_io_b = io_b; // @[Snxn100k.scala 483:26]
  assign inst_SnxnLv1Inst3_io_a = io_a; // @[Snxn100k.scala 486:26]
  assign inst_SnxnLv1Inst3_io_b = io_b; // @[Snxn100k.scala 487:26]
endmodule
