module RecFNToIN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [63:0] io_out,
  output [2:0]  io_intExceptionFlags
);
  wire  rawIn_isZero = io_in[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_in[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn_isNaN = _T_4 & io_in[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_isInf = _T_4 & ~io_in[61]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn_sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn_sExp = {1'b0,$signed(io_in[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_12 = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] rawIn_sig = {1'h0,_T_12,io_in[51:0]}; // @[Cat.scala 29:58]
  wire  magGeOne = rawIn_sExp[11]; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp = rawIn_sExp[10:0]; // @[RecFNToIN.scala 59:28]
  wire  magJustBelowOne = ~magGeOne & &posExp; // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  wire [52:0] _T_19 = {magGeOne,rawIn_sig[51:0]}; // @[Cat.scala 29:58]
  wire [5:0] _T_21 = magGeOne ? rawIn_sExp[5:0] : 6'h0; // @[RecFNToIN.scala 81:16]
  wire [115:0] _GEN_2 = {{63'd0}, _T_19}; // @[RecFNToIN.scala 80:50]
  wire [115:0] shiftedSig = _GEN_2 << _T_21; // @[RecFNToIN.scala 80:50]
  wire  _T_24 = |shiftedSig[50:0]; // @[RecFNToIN.scala 86:69]
  wire [65:0] alignedSig = {shiftedSig[115:51],_T_24}; // @[Cat.scala 29:58]
  wire [63:0] unroundedInt = alignedSig[65:2]; // @[RecFNToIN.scala 87:54]
  wire  _T_27 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57]
  wire  common_inexact = magGeOne ? |alignedSig[1:0] : _T_12; // @[RecFNToIN.scala 89:29]
  wire  _T_37 = magJustBelowOne & _T_27; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even = magGeOne & (&alignedSig[2:1] | &alignedSig[1:0]) | _T_37; // @[RecFNToIN.scala 91:78]
  wire  roundIncr_near_maxMag = magGeOne & alignedSig[1] | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  wire  _T_41 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  wire  _T_42 = roundingMode_near_even & roundIncr_near_even | _T_41; // @[RecFNToIN.scala 95:61]
  wire  _T_44 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:26]
  wire  _T_45 = (roundingMode_min | roundingMode_odd) & _T_44; // @[RecFNToIN.scala 97:49]
  wire  _T_46 = _T_42 | _T_45; // @[RecFNToIN.scala 96:61]
  wire  _T_49 = roundingMode_max & (~rawIn_sign & common_inexact); // @[RecFNToIN.scala 99:27]
  wire  roundIncr = _T_46 | _T_49; // @[RecFNToIN.scala 98:46]
  wire [63:0] _T_50 = ~unroundedInt; // @[RecFNToIN.scala 100:45]
  wire [63:0] complUnroundedInt = rawIn_sign ? _T_50 : unroundedInt; // @[RecFNToIN.scala 100:32]
  wire [63:0] _T_53 = complUnroundedInt + 64'h1; // @[RecFNToIN.scala 103:31]
  wire [63:0] _T_54 = roundIncr ^ rawIn_sign ? _T_53 : complUnroundedInt; // @[RecFNToIN.scala 102:12]
  wire  _T_55 = roundingMode_odd & common_inexact; // @[RecFNToIN.scala 105:31]
  wire [63:0] _GEN_0 = {{63'd0}, _T_55}; // @[RecFNToIN.scala 105:11]
  wire [63:0] roundedInt = _T_54 | _GEN_0; // @[RecFNToIN.scala 105:11]
  wire  magGeOne_atOverflowEdge = posExp == 11'h3f; // @[RecFNToIN.scala 107:43]
  wire  roundCarryBut2 = &unroundedInt[61:0] & roundIncr; // @[RecFNToIN.scala 110:61]
  wire  _T_61 = |unroundedInt[62:0] | roundIncr; // @[RecFNToIN.scala 117:64]
  wire  _T_62 = magGeOne_atOverflowEdge & _T_61; // @[RecFNToIN.scala 116:49]
  wire  _T_64 = posExp == 11'h3e & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  wire  _T_65 = magGeOne_atOverflowEdge | _T_64; // @[RecFNToIN.scala 118:49]
  wire  _T_66 = rawIn_sign ? _T_62 : _T_65; // @[RecFNToIN.scala 115:24]
  wire  _T_68 = magGeOne_atOverflowEdge & unroundedInt[62]; // @[RecFNToIN.scala 122:50]
  wire  _T_69 = _T_68 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  wire  _T_70 = rawIn_sign | _T_69; // @[RecFNToIN.scala 121:32]
  wire  _T_71 = io_signedOut ? _T_66 : _T_70; // @[RecFNToIN.scala 114:20]
  wire  _T_72 = posExp >= 11'h40 | _T_71; // @[RecFNToIN.scala 113:40]
  wire  _T_75 = ~io_signedOut & rawIn_sign & roundIncr; // @[RecFNToIN.scala 125:41]
  wire  common_overflow = magGeOne ? _T_72 : _T_75; // @[RecFNToIN.scala 112:12]
  wire  invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 130:34]
  wire  _T_76 = ~invalidExc; // @[RecFNToIN.scala 131:20]
  wire  overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 131:32]
  wire  inexact = _T_76 & ~common_overflow & common_inexact; // @[RecFNToIN.scala 132:52]
  wire  excSign = ~rawIn_isNaN & rawIn_sign; // @[RecFNToIN.scala 134:32]
  wire [63:0] _T_82 = io_signedOut == excSign ? 64'h8000000000000000 : 64'h0; // @[RecFNToIN.scala 136:12]
  wire [62:0] _T_84 = ~excSign ? 63'h7fffffffffffffff : 63'h0; // @[RecFNToIN.scala 140:12]
  wire [63:0] _GEN_1 = {{1'd0}, _T_84}; // @[RecFNToIN.scala 139:11]
  wire [63:0] excOut = _T_82 | _GEN_1; // @[RecFNToIN.scala 139:11]
  wire [1:0] _T_87 = {invalidExc,overflow}; // @[Cat.scala 29:58]
  assign io_out = invalidExc | common_overflow ? excOut : roundedInt; // @[RecFNToIN.scala 142:18]
  assign io_intExceptionFlags = {_T_87,inexact}; // @[Cat.scala 29:58]
endmodule
