module Adder_1(
  input         clock,
  input         reset,
  input  [31:0] io_inputx,
  input  [31:0] io_inputy,
  output [31:0] io_result
);
  assign io_result = io_inputx + io_inputy;
endmodule
