module drop ( input [3:0] a, output [1:0] b);
assign b = a;
endmodule
