module sum( input a, input b, output [2:0] c);
assign c = a + b;
endmodule

