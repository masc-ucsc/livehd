module xor_10000(
    input a,
    input b,
    output z
    );

wire temp0, temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14, temp15, temp16, temp17, temp18, temp19, temp20, temp21, temp22, temp23, temp24, temp25, temp26, temp27, temp28, temp29, temp30, temp31, temp32, temp33, temp34, temp35, temp36, temp37, temp38, temp39, temp40, temp41, temp42, temp43, temp44, temp45, temp46, temp47, temp48, temp49, temp50, temp51, temp52, temp53, temp54, temp55, temp56, temp57, temp58, temp59, temp60, temp61, temp62, temp63, temp64, temp65, temp66, temp67, temp68, temp69, temp70, temp71, temp72, temp73, temp74, temp75, temp76, temp77, temp78, temp79, temp80, temp81, temp82, temp83, temp84, temp85, temp86, temp87, temp88, temp89, temp90, temp91, temp92, temp93, temp94, temp95, temp96, temp97, temp98, temp99, temp100, temp101, temp102, temp103, temp104, temp105, temp106, temp107, temp108, temp109, temp110, temp111, temp112, temp113, temp114, temp115, temp116, temp117, temp118, temp119, temp120, temp121, temp122, temp123, temp124, temp125, temp126, temp127, temp128, temp129, temp130, temp131, temp132, temp133, temp134, temp135, temp136, temp137, temp138, temp139, temp140, temp141, temp142, temp143, temp144, temp145, temp146, temp147, temp148, temp149, temp150, temp151, temp152, temp153, temp154, temp155, temp156, temp157, temp158, temp159, temp160, temp161, temp162, temp163, temp164, temp165, temp166, temp167, temp168, temp169, temp170, temp171, temp172, temp173, temp174, temp175, temp176, temp177, temp178, temp179, temp180, temp181, temp182, temp183, temp184, temp185, temp186, temp187, temp188, temp189, temp190, temp191, temp192, temp193, temp194, temp195, temp196, temp197, temp198, temp199, temp200, temp201, temp202, temp203, temp204, temp205, temp206, temp207, temp208, temp209, temp210, temp211, temp212, temp213, temp214, temp215, temp216, temp217, temp218, temp219, temp220, temp221, temp222, temp223, temp224, temp225, temp226, temp227, temp228, temp229, temp230, temp231, temp232, temp233, temp234, temp235, temp236, temp237, temp238, temp239, temp240, temp241, temp242, temp243, temp244, temp245, temp246, temp247, temp248, temp249, temp250, temp251, temp252, temp253, temp254, temp255, temp256, temp257, temp258, temp259, temp260, temp261, temp262, temp263, temp264, temp265, temp266, temp267, temp268, temp269, temp270, temp271, temp272, temp273, temp274, temp275, temp276, temp277, temp278, temp279, temp280, temp281, temp282, temp283, temp284, temp285, temp286, temp287, temp288, temp289, temp290, temp291, temp292, temp293, temp294, temp295, temp296, temp297, temp298, temp299, temp300, temp301, temp302, temp303, temp304, temp305, temp306, temp307, temp308, temp309, temp310, temp311, temp312, temp313, temp314, temp315, temp316, temp317, temp318, temp319, temp320, temp321, temp322, temp323, temp324, temp325, temp326, temp327, temp328, temp329, temp330, temp331, temp332, temp333, temp334, temp335, temp336, temp337, temp338, temp339, temp340, temp341, temp342, temp343, temp344, temp345, temp346, temp347, temp348, temp349, temp350, temp351, temp352, temp353, temp354, temp355, temp356, temp357, temp358, temp359, temp360, temp361, temp362, temp363, temp364, temp365, temp366, temp367, temp368, temp369, temp370, temp371, temp372, temp373, temp374, temp375, temp376, temp377, temp378, temp379, temp380, temp381, temp382, temp383, temp384, temp385, temp386, temp387, temp388, temp389, temp390, temp391, temp392, temp393, temp394, temp395, temp396, temp397, temp398, temp399, temp400, temp401, temp402, temp403, temp404, temp405, temp406, temp407, temp408, temp409, temp410, temp411, temp412, temp413, temp414, temp415, temp416, temp417, temp418, temp419, temp420, temp421, temp422, temp423, temp424, temp425, temp426, temp427, temp428, temp429, temp430, temp431, temp432, temp433, temp434, temp435, temp436, temp437, temp438, temp439, temp440, temp441, temp442, temp443, temp444, temp445, temp446, temp447, temp448, temp449, temp450, temp451, temp452, temp453, temp454, temp455, temp456, temp457, temp458, temp459, temp460, temp461, temp462, temp463, temp464, temp465, temp466, temp467, temp468, temp469, temp470, temp471, temp472, temp473, temp474, temp475, temp476, temp477, temp478, temp479, temp480, temp481, temp482, temp483, temp484, temp485, temp486, temp487, temp488, temp489, temp490, temp491, temp492, temp493, temp494, temp495, temp496, temp497, temp498, temp499, temp500, temp501, temp502, temp503, temp504, temp505, temp506, temp507, temp508, temp509, temp510, temp511, temp512, temp513, temp514, temp515, temp516, temp517, temp518, temp519, temp520, temp521, temp522, temp523, temp524, temp525, temp526, temp527, temp528, temp529, temp530, temp531, temp532, temp533, temp534, temp535, temp536, temp537, temp538, temp539, temp540, temp541, temp542, temp543, temp544, temp545, temp546, temp547, temp548, temp549, temp550, temp551, temp552, temp553, temp554, temp555, temp556, temp557, temp558, temp559, temp560, temp561, temp562, temp563, temp564, temp565, temp566, temp567, temp568, temp569, temp570, temp571, temp572, temp573, temp574, temp575, temp576, temp577, temp578, temp579, temp580, temp581, temp582, temp583, temp584, temp585, temp586, temp587, temp588, temp589, temp590, temp591, temp592, temp593, temp594, temp595, temp596, temp597, temp598, temp599, temp600, temp601, temp602, temp603, temp604, temp605, temp606, temp607, temp608, temp609, temp610, temp611, temp612, temp613, temp614, temp615, temp616, temp617, temp618, temp619, temp620, temp621, temp622, temp623, temp624, temp625, temp626, temp627, temp628, temp629, temp630, temp631, temp632, temp633, temp634, temp635, temp636, temp637, temp638, temp639, temp640, temp641, temp642, temp643, temp644, temp645, temp646, temp647, temp648, temp649, temp650, temp651, temp652, temp653, temp654, temp655, temp656, temp657, temp658, temp659, temp660, temp661, temp662, temp663, temp664, temp665, temp666, temp667, temp668, temp669, temp670, temp671, temp672, temp673, temp674, temp675, temp676, temp677, temp678, temp679, temp680, temp681, temp682, temp683, temp684, temp685, temp686, temp687, temp688, temp689, temp690, temp691, temp692, temp693, temp694, temp695, temp696, temp697, temp698, temp699, temp700, temp701, temp702, temp703, temp704, temp705, temp706, temp707, temp708, temp709, temp710, temp711, temp712, temp713, temp714, temp715, temp716, temp717, temp718, temp719, temp720, temp721, temp722, temp723, temp724, temp725, temp726, temp727, temp728, temp729, temp730, temp731, temp732, temp733, temp734, temp735, temp736, temp737, temp738, temp739, temp740, temp741, temp742, temp743, temp744, temp745, temp746, temp747, temp748, temp749, temp750, temp751, temp752, temp753, temp754, temp755, temp756, temp757, temp758, temp759, temp760, temp761, temp762, temp763, temp764, temp765, temp766, temp767, temp768, temp769, temp770, temp771, temp772, temp773, temp774, temp775, temp776, temp777, temp778, temp779, temp780, temp781, temp782, temp783, temp784, temp785, temp786, temp787, temp788, temp789, temp790, temp791, temp792, temp793, temp794, temp795, temp796, temp797, temp798, temp799, temp800, temp801, temp802, temp803, temp804, temp805, temp806, temp807, temp808, temp809, temp810, temp811, temp812, temp813, temp814, temp815, temp816, temp817, temp818, temp819, temp820, temp821, temp822, temp823, temp824, temp825, temp826, temp827, temp828, temp829, temp830, temp831, temp832, temp833, temp834, temp835, temp836, temp837, temp838, temp839, temp840, temp841, temp842, temp843, temp844, temp845, temp846, temp847, temp848, temp849, temp850, temp851, temp852, temp853, temp854, temp855, temp856, temp857, temp858, temp859, temp860, temp861, temp862, temp863, temp864, temp865, temp866, temp867, temp868, temp869, temp870, temp871, temp872, temp873, temp874, temp875, temp876, temp877, temp878, temp879, temp880, temp881, temp882, temp883, temp884, temp885, temp886, temp887, temp888, temp889, temp890, temp891, temp892, temp893, temp894, temp895, temp896, temp897, temp898, temp899, temp900, temp901, temp902, temp903, temp904, temp905, temp906, temp907, temp908, temp909, temp910, temp911, temp912, temp913, temp914, temp915, temp916, temp917, temp918, temp919, temp920, temp921, temp922, temp923, temp924, temp925, temp926, temp927, temp928, temp929, temp930, temp931, temp932, temp933, temp934, temp935, temp936, temp937, temp938, temp939, temp940, temp941, temp942, temp943, temp944, temp945, temp946, temp947, temp948, temp949, temp950, temp951, temp952, temp953, temp954, temp955, temp956, temp957, temp958, temp959, temp960, temp961, temp962, temp963, temp964, temp965, temp966, temp967, temp968, temp969, temp970, temp971, temp972, temp973, temp974, temp975, temp976, temp977, temp978, temp979, temp980, temp981, temp982, temp983, temp984, temp985, temp986, temp987, temp988, temp989, temp990, temp991, temp992, temp993, temp994, temp995, temp996, temp997, temp998, temp999, temp1000, temp1001, temp1002, temp1003, temp1004, temp1005, temp1006, temp1007, temp1008, temp1009, temp1010, temp1011, temp1012, temp1013, temp1014, temp1015, temp1016, temp1017, temp1018, temp1019, temp1020, temp1021, temp1022, temp1023, temp1024, temp1025, temp1026, temp1027, temp1028, temp1029, temp1030, temp1031, temp1032, temp1033, temp1034, temp1035, temp1036, temp1037, temp1038, temp1039, temp1040, temp1041, temp1042, temp1043, temp1044, temp1045, temp1046, temp1047, temp1048, temp1049, temp1050, temp1051, temp1052, temp1053, temp1054, temp1055, temp1056, temp1057, temp1058, temp1059, temp1060, temp1061, temp1062, temp1063, temp1064, temp1065, temp1066, temp1067, temp1068, temp1069, temp1070, temp1071, temp1072, temp1073, temp1074, temp1075, temp1076, temp1077, temp1078, temp1079, temp1080, temp1081, temp1082, temp1083, temp1084, temp1085, temp1086, temp1087, temp1088, temp1089, temp1090, temp1091, temp1092, temp1093, temp1094, temp1095, temp1096, temp1097, temp1098, temp1099, temp1100, temp1101, temp1102, temp1103, temp1104, temp1105, temp1106, temp1107, temp1108, temp1109, temp1110, temp1111, temp1112, temp1113, temp1114, temp1115, temp1116, temp1117, temp1118, temp1119, temp1120, temp1121, temp1122, temp1123, temp1124, temp1125, temp1126, temp1127, temp1128, temp1129, temp1130, temp1131, temp1132, temp1133, temp1134, temp1135, temp1136, temp1137, temp1138, temp1139, temp1140, temp1141, temp1142, temp1143, temp1144, temp1145, temp1146, temp1147, temp1148, temp1149, temp1150, temp1151, temp1152, temp1153, temp1154, temp1155, temp1156, temp1157, temp1158, temp1159, temp1160, temp1161, temp1162, temp1163, temp1164, temp1165, temp1166, temp1167, temp1168, temp1169, temp1170, temp1171, temp1172, temp1173, temp1174, temp1175, temp1176, temp1177, temp1178, temp1179, temp1180, temp1181, temp1182, temp1183, temp1184, temp1185, temp1186, temp1187, temp1188, temp1189, temp1190, temp1191, temp1192, temp1193, temp1194, temp1195, temp1196, temp1197, temp1198, temp1199, temp1200, temp1201, temp1202, temp1203, temp1204, temp1205, temp1206, temp1207, temp1208, temp1209, temp1210, temp1211, temp1212, temp1213, temp1214, temp1215, temp1216, temp1217, temp1218, temp1219, temp1220, temp1221, temp1222, temp1223, temp1224, temp1225, temp1226, temp1227, temp1228, temp1229, temp1230, temp1231, temp1232, temp1233, temp1234, temp1235, temp1236, temp1237, temp1238, temp1239, temp1240, temp1241, temp1242, temp1243, temp1244, temp1245, temp1246, temp1247, temp1248, temp1249, temp1250, temp1251, temp1252, temp1253, temp1254, temp1255, temp1256, temp1257, temp1258, temp1259, temp1260, temp1261, temp1262, temp1263, temp1264, temp1265, temp1266, temp1267, temp1268, temp1269, temp1270, temp1271, temp1272, temp1273, temp1274, temp1275, temp1276, temp1277, temp1278, temp1279, temp1280, temp1281, temp1282, temp1283, temp1284, temp1285, temp1286, temp1287, temp1288, temp1289, temp1290, temp1291, temp1292, temp1293, temp1294, temp1295, temp1296, temp1297, temp1298, temp1299, temp1300, temp1301, temp1302, temp1303, temp1304, temp1305, temp1306, temp1307, temp1308, temp1309, temp1310, temp1311, temp1312, temp1313, temp1314, temp1315, temp1316, temp1317, temp1318, temp1319, temp1320, temp1321, temp1322, temp1323, temp1324, temp1325, temp1326, temp1327, temp1328, temp1329, temp1330, temp1331, temp1332, temp1333, temp1334, temp1335, temp1336, temp1337, temp1338, temp1339, temp1340, temp1341, temp1342, temp1343, temp1344, temp1345, temp1346, temp1347, temp1348, temp1349, temp1350, temp1351, temp1352, temp1353, temp1354, temp1355, temp1356, temp1357, temp1358, temp1359, temp1360, temp1361, temp1362, temp1363, temp1364, temp1365, temp1366, temp1367, temp1368, temp1369, temp1370, temp1371, temp1372, temp1373, temp1374, temp1375, temp1376, temp1377, temp1378, temp1379, temp1380, temp1381, temp1382, temp1383, temp1384, temp1385, temp1386, temp1387, temp1388, temp1389, temp1390, temp1391, temp1392, temp1393, temp1394, temp1395, temp1396, temp1397, temp1398, temp1399, temp1400, temp1401, temp1402, temp1403, temp1404, temp1405, temp1406, temp1407, temp1408, temp1409, temp1410, temp1411, temp1412, temp1413, temp1414, temp1415, temp1416, temp1417, temp1418, temp1419, temp1420, temp1421, temp1422, temp1423, temp1424, temp1425, temp1426, temp1427, temp1428, temp1429, temp1430, temp1431, temp1432, temp1433, temp1434, temp1435, temp1436, temp1437, temp1438, temp1439, temp1440, temp1441, temp1442, temp1443, temp1444, temp1445, temp1446, temp1447, temp1448, temp1449, temp1450, temp1451, temp1452, temp1453, temp1454, temp1455, temp1456, temp1457, temp1458, temp1459, temp1460, temp1461, temp1462, temp1463, temp1464, temp1465, temp1466, temp1467, temp1468, temp1469, temp1470, temp1471, temp1472, temp1473, temp1474, temp1475, temp1476, temp1477, temp1478, temp1479, temp1480, temp1481, temp1482, temp1483, temp1484, temp1485, temp1486, temp1487, temp1488, temp1489, temp1490, temp1491, temp1492, temp1493, temp1494, temp1495, temp1496, temp1497, temp1498, temp1499, temp1500, temp1501, temp1502, temp1503, temp1504, temp1505, temp1506, temp1507, temp1508, temp1509, temp1510, temp1511, temp1512, temp1513, temp1514, temp1515, temp1516, temp1517, temp1518, temp1519, temp1520, temp1521, temp1522, temp1523, temp1524, temp1525, temp1526, temp1527, temp1528, temp1529, temp1530, temp1531, temp1532, temp1533, temp1534, temp1535, temp1536, temp1537, temp1538, temp1539, temp1540, temp1541, temp1542, temp1543, temp1544, temp1545, temp1546, temp1547, temp1548, temp1549, temp1550, temp1551, temp1552, temp1553, temp1554, temp1555, temp1556, temp1557, temp1558, temp1559, temp1560, temp1561, temp1562, temp1563, temp1564, temp1565, temp1566, temp1567, temp1568, temp1569, temp1570, temp1571, temp1572, temp1573, temp1574, temp1575, temp1576, temp1577, temp1578, temp1579, temp1580, temp1581, temp1582, temp1583, temp1584, temp1585, temp1586, temp1587, temp1588, temp1589, temp1590, temp1591, temp1592, temp1593, temp1594, temp1595, temp1596, temp1597, temp1598, temp1599, temp1600, temp1601, temp1602, temp1603, temp1604, temp1605, temp1606, temp1607, temp1608, temp1609, temp1610, temp1611, temp1612, temp1613, temp1614, temp1615, temp1616, temp1617, temp1618, temp1619, temp1620, temp1621, temp1622, temp1623, temp1624, temp1625, temp1626, temp1627, temp1628, temp1629, temp1630, temp1631, temp1632, temp1633, temp1634, temp1635, temp1636, temp1637, temp1638, temp1639, temp1640, temp1641, temp1642, temp1643, temp1644, temp1645, temp1646, temp1647, temp1648, temp1649, temp1650, temp1651, temp1652, temp1653, temp1654, temp1655, temp1656, temp1657, temp1658, temp1659, temp1660, temp1661, temp1662, temp1663, temp1664, temp1665, temp1666, temp1667, temp1668, temp1669, temp1670, temp1671, temp1672, temp1673, temp1674, temp1675, temp1676, temp1677, temp1678, temp1679, temp1680, temp1681, temp1682, temp1683, temp1684, temp1685, temp1686, temp1687, temp1688, temp1689, temp1690, temp1691, temp1692, temp1693, temp1694, temp1695, temp1696, temp1697, temp1698, temp1699, temp1700, temp1701, temp1702, temp1703, temp1704, temp1705, temp1706, temp1707, temp1708, temp1709, temp1710, temp1711, temp1712, temp1713, temp1714, temp1715, temp1716, temp1717, temp1718, temp1719, temp1720, temp1721, temp1722, temp1723, temp1724, temp1725, temp1726, temp1727, temp1728, temp1729, temp1730, temp1731, temp1732, temp1733, temp1734, temp1735, temp1736, temp1737, temp1738, temp1739, temp1740, temp1741, temp1742, temp1743, temp1744, temp1745, temp1746, temp1747, temp1748, temp1749, temp1750, temp1751, temp1752, temp1753, temp1754, temp1755, temp1756, temp1757, temp1758, temp1759, temp1760, temp1761, temp1762, temp1763, temp1764, temp1765, temp1766, temp1767, temp1768, temp1769, temp1770, temp1771, temp1772, temp1773, temp1774, temp1775, temp1776, temp1777, temp1778, temp1779, temp1780, temp1781, temp1782, temp1783, temp1784, temp1785, temp1786, temp1787, temp1788, temp1789, temp1790, temp1791, temp1792, temp1793, temp1794, temp1795, temp1796, temp1797, temp1798, temp1799, temp1800, temp1801, temp1802, temp1803, temp1804, temp1805, temp1806, temp1807, temp1808, temp1809, temp1810, temp1811, temp1812, temp1813, temp1814, temp1815, temp1816, temp1817, temp1818, temp1819, temp1820, temp1821, temp1822, temp1823, temp1824, temp1825, temp1826, temp1827, temp1828, temp1829, temp1830, temp1831, temp1832, temp1833, temp1834, temp1835, temp1836, temp1837, temp1838, temp1839, temp1840, temp1841, temp1842, temp1843, temp1844, temp1845, temp1846, temp1847, temp1848, temp1849, temp1850, temp1851, temp1852, temp1853, temp1854, temp1855, temp1856, temp1857, temp1858, temp1859, temp1860, temp1861, temp1862, temp1863, temp1864, temp1865, temp1866, temp1867, temp1868, temp1869, temp1870, temp1871, temp1872, temp1873, temp1874, temp1875, temp1876, temp1877, temp1878, temp1879, temp1880, temp1881, temp1882, temp1883, temp1884, temp1885, temp1886, temp1887, temp1888, temp1889, temp1890, temp1891, temp1892, temp1893, temp1894, temp1895, temp1896, temp1897, temp1898, temp1899, temp1900, temp1901, temp1902, temp1903, temp1904, temp1905, temp1906, temp1907, temp1908, temp1909, temp1910, temp1911, temp1912, temp1913, temp1914, temp1915, temp1916, temp1917, temp1918, temp1919, temp1920, temp1921, temp1922, temp1923, temp1924, temp1925, temp1926, temp1927, temp1928, temp1929, temp1930, temp1931, temp1932, temp1933, temp1934, temp1935, temp1936, temp1937, temp1938, temp1939, temp1940, temp1941, temp1942, temp1943, temp1944, temp1945, temp1946, temp1947, temp1948, temp1949, temp1950, temp1951, temp1952, temp1953, temp1954, temp1955, temp1956, temp1957, temp1958, temp1959, temp1960, temp1961, temp1962, temp1963, temp1964, temp1965, temp1966, temp1967, temp1968, temp1969, temp1970, temp1971, temp1972, temp1973, temp1974, temp1975, temp1976, temp1977, temp1978, temp1979, temp1980, temp1981, temp1982, temp1983, temp1984, temp1985, temp1986, temp1987, temp1988, temp1989, temp1990, temp1991, temp1992, temp1993, temp1994, temp1995, temp1996, temp1997, temp1998, temp1999, temp2000, temp2001, temp2002, temp2003, temp2004, temp2005, temp2006, temp2007, temp2008, temp2009, temp2010, temp2011, temp2012, temp2013, temp2014, temp2015, temp2016, temp2017, temp2018, temp2019, temp2020, temp2021, temp2022, temp2023, temp2024, temp2025, temp2026, temp2027, temp2028, temp2029, temp2030, temp2031, temp2032, temp2033, temp2034, temp2035, temp2036, temp2037, temp2038, temp2039, temp2040, temp2041, temp2042, temp2043, temp2044, temp2045, temp2046, temp2047, temp2048, temp2049, temp2050, temp2051, temp2052, temp2053, temp2054, temp2055, temp2056, temp2057, temp2058, temp2059, temp2060, temp2061, temp2062, temp2063, temp2064, temp2065, temp2066, temp2067, temp2068, temp2069, temp2070, temp2071, temp2072, temp2073, temp2074, temp2075, temp2076, temp2077, temp2078, temp2079, temp2080, temp2081, temp2082, temp2083, temp2084, temp2085, temp2086, temp2087, temp2088, temp2089, temp2090, temp2091, temp2092, temp2093, temp2094, temp2095, temp2096, temp2097, temp2098, temp2099, temp2100, temp2101, temp2102, temp2103, temp2104, temp2105, temp2106, temp2107, temp2108, temp2109, temp2110, temp2111, temp2112, temp2113, temp2114, temp2115, temp2116, temp2117, temp2118, temp2119, temp2120, temp2121, temp2122, temp2123, temp2124, temp2125, temp2126, temp2127, temp2128, temp2129, temp2130, temp2131, temp2132, temp2133, temp2134, temp2135, temp2136, temp2137, temp2138, temp2139, temp2140, temp2141, temp2142, temp2143, temp2144, temp2145, temp2146, temp2147, temp2148, temp2149, temp2150, temp2151, temp2152, temp2153, temp2154, temp2155, temp2156, temp2157, temp2158, temp2159, temp2160, temp2161, temp2162, temp2163, temp2164, temp2165, temp2166, temp2167, temp2168, temp2169, temp2170, temp2171, temp2172, temp2173, temp2174, temp2175, temp2176, temp2177, temp2178, temp2179, temp2180, temp2181, temp2182, temp2183, temp2184, temp2185, temp2186, temp2187, temp2188, temp2189, temp2190, temp2191, temp2192, temp2193, temp2194, temp2195, temp2196, temp2197, temp2198, temp2199, temp2200, temp2201, temp2202, temp2203, temp2204, temp2205, temp2206, temp2207, temp2208, temp2209, temp2210, temp2211, temp2212, temp2213, temp2214, temp2215, temp2216, temp2217, temp2218, temp2219, temp2220, temp2221, temp2222, temp2223, temp2224, temp2225, temp2226, temp2227, temp2228, temp2229, temp2230, temp2231, temp2232, temp2233, temp2234, temp2235, temp2236, temp2237, temp2238, temp2239, temp2240, temp2241, temp2242, temp2243, temp2244, temp2245, temp2246, temp2247, temp2248, temp2249, temp2250, temp2251, temp2252, temp2253, temp2254, temp2255, temp2256, temp2257, temp2258, temp2259, temp2260, temp2261, temp2262, temp2263, temp2264, temp2265, temp2266, temp2267, temp2268, temp2269, temp2270, temp2271, temp2272, temp2273, temp2274, temp2275, temp2276, temp2277, temp2278, temp2279, temp2280, temp2281, temp2282, temp2283, temp2284, temp2285, temp2286, temp2287, temp2288, temp2289, temp2290, temp2291, temp2292, temp2293, temp2294, temp2295, temp2296, temp2297, temp2298, temp2299, temp2300, temp2301, temp2302, temp2303, temp2304, temp2305, temp2306, temp2307, temp2308, temp2309, temp2310, temp2311, temp2312, temp2313, temp2314, temp2315, temp2316, temp2317, temp2318, temp2319, temp2320, temp2321, temp2322, temp2323, temp2324, temp2325, temp2326, temp2327, temp2328, temp2329, temp2330, temp2331, temp2332, temp2333, temp2334, temp2335, temp2336, temp2337, temp2338, temp2339, temp2340, temp2341, temp2342, temp2343, temp2344, temp2345, temp2346, temp2347, temp2348, temp2349, temp2350, temp2351, temp2352, temp2353, temp2354, temp2355, temp2356, temp2357, temp2358, temp2359, temp2360, temp2361, temp2362, temp2363, temp2364, temp2365, temp2366, temp2367, temp2368, temp2369, temp2370, temp2371, temp2372, temp2373, temp2374, temp2375, temp2376, temp2377, temp2378, temp2379, temp2380, temp2381, temp2382, temp2383, temp2384, temp2385, temp2386, temp2387, temp2388, temp2389, temp2390, temp2391, temp2392, temp2393, temp2394, temp2395, temp2396, temp2397, temp2398, temp2399, temp2400, temp2401, temp2402, temp2403, temp2404, temp2405, temp2406, temp2407, temp2408, temp2409, temp2410, temp2411, temp2412, temp2413, temp2414, temp2415, temp2416, temp2417, temp2418, temp2419, temp2420, temp2421, temp2422, temp2423, temp2424, temp2425, temp2426, temp2427, temp2428, temp2429, temp2430, temp2431, temp2432, temp2433, temp2434, temp2435, temp2436, temp2437, temp2438, temp2439, temp2440, temp2441, temp2442, temp2443, temp2444, temp2445, temp2446, temp2447, temp2448, temp2449, temp2450, temp2451, temp2452, temp2453, temp2454, temp2455, temp2456, temp2457, temp2458, temp2459, temp2460, temp2461, temp2462, temp2463, temp2464, temp2465, temp2466, temp2467, temp2468, temp2469, temp2470, temp2471, temp2472, temp2473, temp2474, temp2475, temp2476, temp2477, temp2478, temp2479, temp2480, temp2481, temp2482, temp2483, temp2484, temp2485, temp2486, temp2487, temp2488, temp2489, temp2490, temp2491, temp2492, temp2493, temp2494, temp2495, temp2496, temp2497, temp2498, temp2499, temp2500, temp2501, temp2502, temp2503, temp2504, temp2505, temp2506, temp2507, temp2508, temp2509, temp2510, temp2511, temp2512, temp2513, temp2514, temp2515, temp2516, temp2517, temp2518, temp2519, temp2520, temp2521, temp2522, temp2523, temp2524, temp2525, temp2526, temp2527, temp2528, temp2529, temp2530, temp2531, temp2532, temp2533, temp2534, temp2535, temp2536, temp2537, temp2538, temp2539, temp2540, temp2541, temp2542, temp2543, temp2544, temp2545, temp2546, temp2547, temp2548, temp2549, temp2550, temp2551, temp2552, temp2553, temp2554, temp2555, temp2556, temp2557, temp2558, temp2559, temp2560, temp2561, temp2562, temp2563, temp2564, temp2565, temp2566, temp2567, temp2568, temp2569, temp2570, temp2571, temp2572, temp2573, temp2574, temp2575, temp2576, temp2577, temp2578, temp2579, temp2580, temp2581, temp2582, temp2583, temp2584, temp2585, temp2586, temp2587, temp2588, temp2589, temp2590, temp2591, temp2592, temp2593, temp2594, temp2595, temp2596, temp2597, temp2598, temp2599, temp2600, temp2601, temp2602, temp2603, temp2604, temp2605, temp2606, temp2607, temp2608, temp2609, temp2610, temp2611, temp2612, temp2613, temp2614, temp2615, temp2616, temp2617, temp2618, temp2619, temp2620, temp2621, temp2622, temp2623, temp2624, temp2625, temp2626, temp2627, temp2628, temp2629, temp2630, temp2631, temp2632, temp2633, temp2634, temp2635, temp2636, temp2637, temp2638, temp2639, temp2640, temp2641, temp2642, temp2643, temp2644, temp2645, temp2646, temp2647, temp2648, temp2649, temp2650, temp2651, temp2652, temp2653, temp2654, temp2655, temp2656, temp2657, temp2658, temp2659, temp2660, temp2661, temp2662, temp2663, temp2664, temp2665, temp2666, temp2667, temp2668, temp2669, temp2670, temp2671, temp2672, temp2673, temp2674, temp2675, temp2676, temp2677, temp2678, temp2679, temp2680, temp2681, temp2682, temp2683, temp2684, temp2685, temp2686, temp2687, temp2688, temp2689, temp2690, temp2691, temp2692, temp2693, temp2694, temp2695, temp2696, temp2697, temp2698, temp2699, temp2700, temp2701, temp2702, temp2703, temp2704, temp2705, temp2706, temp2707, temp2708, temp2709, temp2710, temp2711, temp2712, temp2713, temp2714, temp2715, temp2716, temp2717, temp2718, temp2719, temp2720, temp2721, temp2722, temp2723, temp2724, temp2725, temp2726, temp2727, temp2728, temp2729, temp2730, temp2731, temp2732, temp2733, temp2734, temp2735, temp2736, temp2737, temp2738, temp2739, temp2740, temp2741, temp2742, temp2743, temp2744, temp2745, temp2746, temp2747, temp2748, temp2749, temp2750, temp2751, temp2752, temp2753, temp2754, temp2755, temp2756, temp2757, temp2758, temp2759, temp2760, temp2761, temp2762, temp2763, temp2764, temp2765, temp2766, temp2767, temp2768, temp2769, temp2770, temp2771, temp2772, temp2773, temp2774, temp2775, temp2776, temp2777, temp2778, temp2779, temp2780, temp2781, temp2782, temp2783, temp2784, temp2785, temp2786, temp2787, temp2788, temp2789, temp2790, temp2791, temp2792, temp2793, temp2794, temp2795, temp2796, temp2797, temp2798, temp2799, temp2800, temp2801, temp2802, temp2803, temp2804, temp2805, temp2806, temp2807, temp2808, temp2809, temp2810, temp2811, temp2812, temp2813, temp2814, temp2815, temp2816, temp2817, temp2818, temp2819, temp2820, temp2821, temp2822, temp2823, temp2824, temp2825, temp2826, temp2827, temp2828, temp2829, temp2830, temp2831, temp2832, temp2833, temp2834, temp2835, temp2836, temp2837, temp2838, temp2839, temp2840, temp2841, temp2842, temp2843, temp2844, temp2845, temp2846, temp2847, temp2848, temp2849, temp2850, temp2851, temp2852, temp2853, temp2854, temp2855, temp2856, temp2857, temp2858, temp2859, temp2860, temp2861, temp2862, temp2863, temp2864, temp2865, temp2866, temp2867, temp2868, temp2869, temp2870, temp2871, temp2872, temp2873, temp2874, temp2875, temp2876, temp2877, temp2878, temp2879, temp2880, temp2881, temp2882, temp2883, temp2884, temp2885, temp2886, temp2887, temp2888, temp2889, temp2890, temp2891, temp2892, temp2893, temp2894, temp2895, temp2896, temp2897, temp2898, temp2899, temp2900, temp2901, temp2902, temp2903, temp2904, temp2905, temp2906, temp2907, temp2908, temp2909, temp2910, temp2911, temp2912, temp2913, temp2914, temp2915, temp2916, temp2917, temp2918, temp2919, temp2920, temp2921, temp2922, temp2923, temp2924, temp2925, temp2926, temp2927, temp2928, temp2929, temp2930, temp2931, temp2932, temp2933, temp2934, temp2935, temp2936, temp2937, temp2938, temp2939, temp2940, temp2941, temp2942, temp2943, temp2944, temp2945, temp2946, temp2947, temp2948, temp2949, temp2950, temp2951, temp2952, temp2953, temp2954, temp2955, temp2956, temp2957, temp2958, temp2959, temp2960, temp2961, temp2962, temp2963, temp2964, temp2965, temp2966, temp2967, temp2968, temp2969, temp2970, temp2971, temp2972, temp2973, temp2974, temp2975, temp2976, temp2977, temp2978, temp2979, temp2980, temp2981, temp2982, temp2983, temp2984, temp2985, temp2986, temp2987, temp2988, temp2989, temp2990, temp2991, temp2992, temp2993, temp2994, temp2995, temp2996, temp2997, temp2998, temp2999, temp3000, temp3001, temp3002, temp3003, temp3004, temp3005, temp3006, temp3007, temp3008, temp3009, temp3010, temp3011, temp3012, temp3013, temp3014, temp3015, temp3016, temp3017, temp3018, temp3019, temp3020, temp3021, temp3022, temp3023, temp3024, temp3025, temp3026, temp3027, temp3028, temp3029, temp3030, temp3031, temp3032, temp3033, temp3034, temp3035, temp3036, temp3037, temp3038, temp3039, temp3040, temp3041, temp3042, temp3043, temp3044, temp3045, temp3046, temp3047, temp3048, temp3049, temp3050, temp3051, temp3052, temp3053, temp3054, temp3055, temp3056, temp3057, temp3058, temp3059, temp3060, temp3061, temp3062, temp3063, temp3064, temp3065, temp3066, temp3067, temp3068, temp3069, temp3070, temp3071, temp3072, temp3073, temp3074, temp3075, temp3076, temp3077, temp3078, temp3079, temp3080, temp3081, temp3082, temp3083, temp3084, temp3085, temp3086, temp3087, temp3088, temp3089, temp3090, temp3091, temp3092, temp3093, temp3094, temp3095, temp3096, temp3097, temp3098, temp3099, temp3100, temp3101, temp3102, temp3103, temp3104, temp3105, temp3106, temp3107, temp3108, temp3109, temp3110, temp3111, temp3112, temp3113, temp3114, temp3115, temp3116, temp3117, temp3118, temp3119, temp3120, temp3121, temp3122, temp3123, temp3124, temp3125, temp3126, temp3127, temp3128, temp3129, temp3130, temp3131, temp3132, temp3133, temp3134, temp3135, temp3136, temp3137, temp3138, temp3139, temp3140, temp3141, temp3142, temp3143, temp3144, temp3145, temp3146, temp3147, temp3148, temp3149, temp3150, temp3151, temp3152, temp3153, temp3154, temp3155, temp3156, temp3157, temp3158, temp3159, temp3160, temp3161, temp3162, temp3163, temp3164, temp3165, temp3166, temp3167, temp3168, temp3169, temp3170, temp3171, temp3172, temp3173, temp3174, temp3175, temp3176, temp3177, temp3178, temp3179, temp3180, temp3181, temp3182, temp3183, temp3184, temp3185, temp3186, temp3187, temp3188, temp3189, temp3190, temp3191, temp3192, temp3193, temp3194, temp3195, temp3196, temp3197, temp3198, temp3199, temp3200, temp3201, temp3202, temp3203, temp3204, temp3205, temp3206, temp3207, temp3208, temp3209, temp3210, temp3211, temp3212, temp3213, temp3214, temp3215, temp3216, temp3217, temp3218, temp3219, temp3220, temp3221, temp3222, temp3223, temp3224, temp3225, temp3226, temp3227, temp3228, temp3229, temp3230, temp3231, temp3232, temp3233, temp3234, temp3235, temp3236, temp3237, temp3238, temp3239, temp3240, temp3241, temp3242, temp3243, temp3244, temp3245, temp3246, temp3247, temp3248, temp3249, temp3250, temp3251, temp3252, temp3253, temp3254, temp3255, temp3256, temp3257, temp3258, temp3259, temp3260, temp3261, temp3262, temp3263, temp3264, temp3265, temp3266, temp3267, temp3268, temp3269, temp3270, temp3271, temp3272, temp3273, temp3274, temp3275, temp3276, temp3277, temp3278, temp3279, temp3280, temp3281, temp3282, temp3283, temp3284, temp3285, temp3286, temp3287, temp3288, temp3289, temp3290, temp3291, temp3292, temp3293, temp3294, temp3295, temp3296, temp3297, temp3298, temp3299, temp3300, temp3301, temp3302, temp3303, temp3304, temp3305, temp3306, temp3307, temp3308, temp3309, temp3310, temp3311, temp3312, temp3313, temp3314, temp3315, temp3316, temp3317, temp3318, temp3319, temp3320, temp3321, temp3322, temp3323, temp3324, temp3325, temp3326, temp3327, temp3328, temp3329, temp3330, temp3331, temp3332, temp3333, temp3334, temp3335, temp3336, temp3337, temp3338, temp3339, temp3340, temp3341, temp3342, temp3343, temp3344, temp3345, temp3346, temp3347, temp3348, temp3349, temp3350, temp3351, temp3352, temp3353, temp3354, temp3355, temp3356, temp3357, temp3358, temp3359, temp3360, temp3361, temp3362, temp3363, temp3364, temp3365, temp3366, temp3367, temp3368, temp3369, temp3370, temp3371, temp3372, temp3373, temp3374, temp3375, temp3376, temp3377, temp3378, temp3379, temp3380, temp3381, temp3382, temp3383, temp3384, temp3385, temp3386, temp3387, temp3388, temp3389, temp3390, temp3391, temp3392, temp3393, temp3394, temp3395, temp3396, temp3397, temp3398, temp3399, temp3400, temp3401, temp3402, temp3403, temp3404, temp3405, temp3406, temp3407, temp3408, temp3409, temp3410, temp3411, temp3412, temp3413, temp3414, temp3415, temp3416, temp3417, temp3418, temp3419, temp3420, temp3421, temp3422, temp3423, temp3424, temp3425, temp3426, temp3427, temp3428, temp3429, temp3430, temp3431, temp3432, temp3433, temp3434, temp3435, temp3436, temp3437, temp3438, temp3439, temp3440, temp3441, temp3442, temp3443, temp3444, temp3445, temp3446, temp3447, temp3448, temp3449, temp3450, temp3451, temp3452, temp3453, temp3454, temp3455, temp3456, temp3457, temp3458, temp3459, temp3460, temp3461, temp3462, temp3463, temp3464, temp3465, temp3466, temp3467, temp3468, temp3469, temp3470, temp3471, temp3472, temp3473, temp3474, temp3475, temp3476, temp3477, temp3478, temp3479, temp3480, temp3481, temp3482, temp3483, temp3484, temp3485, temp3486, temp3487, temp3488, temp3489, temp3490, temp3491, temp3492, temp3493, temp3494, temp3495, temp3496, temp3497, temp3498, temp3499, temp3500, temp3501, temp3502, temp3503, temp3504, temp3505, temp3506, temp3507, temp3508, temp3509, temp3510, temp3511, temp3512, temp3513, temp3514, temp3515, temp3516, temp3517, temp3518, temp3519, temp3520, temp3521, temp3522, temp3523, temp3524, temp3525, temp3526, temp3527, temp3528, temp3529, temp3530, temp3531, temp3532, temp3533, temp3534, temp3535, temp3536, temp3537, temp3538, temp3539, temp3540, temp3541, temp3542, temp3543, temp3544, temp3545, temp3546, temp3547, temp3548, temp3549, temp3550, temp3551, temp3552, temp3553, temp3554, temp3555, temp3556, temp3557, temp3558, temp3559, temp3560, temp3561, temp3562, temp3563, temp3564, temp3565, temp3566, temp3567, temp3568, temp3569, temp3570, temp3571, temp3572, temp3573, temp3574, temp3575, temp3576, temp3577, temp3578, temp3579, temp3580, temp3581, temp3582, temp3583, temp3584, temp3585, temp3586, temp3587, temp3588, temp3589, temp3590, temp3591, temp3592, temp3593, temp3594, temp3595, temp3596, temp3597, temp3598, temp3599, temp3600, temp3601, temp3602, temp3603, temp3604, temp3605, temp3606, temp3607, temp3608, temp3609, temp3610, temp3611, temp3612, temp3613, temp3614, temp3615, temp3616, temp3617, temp3618, temp3619, temp3620, temp3621, temp3622, temp3623, temp3624, temp3625, temp3626, temp3627, temp3628, temp3629, temp3630, temp3631, temp3632, temp3633, temp3634, temp3635, temp3636, temp3637, temp3638, temp3639, temp3640, temp3641, temp3642, temp3643, temp3644, temp3645, temp3646, temp3647, temp3648, temp3649, temp3650, temp3651, temp3652, temp3653, temp3654, temp3655, temp3656, temp3657, temp3658, temp3659, temp3660, temp3661, temp3662, temp3663, temp3664, temp3665, temp3666, temp3667, temp3668, temp3669, temp3670, temp3671, temp3672, temp3673, temp3674, temp3675, temp3676, temp3677, temp3678, temp3679, temp3680, temp3681, temp3682, temp3683, temp3684, temp3685, temp3686, temp3687, temp3688, temp3689, temp3690, temp3691, temp3692, temp3693, temp3694, temp3695, temp3696, temp3697, temp3698, temp3699, temp3700, temp3701, temp3702, temp3703, temp3704, temp3705, temp3706, temp3707, temp3708, temp3709, temp3710, temp3711, temp3712, temp3713, temp3714, temp3715, temp3716, temp3717, temp3718, temp3719, temp3720, temp3721, temp3722, temp3723, temp3724, temp3725, temp3726, temp3727, temp3728, temp3729, temp3730, temp3731, temp3732, temp3733, temp3734, temp3735, temp3736, temp3737, temp3738, temp3739, temp3740, temp3741, temp3742, temp3743, temp3744, temp3745, temp3746, temp3747, temp3748, temp3749, temp3750, temp3751, temp3752, temp3753, temp3754, temp3755, temp3756, temp3757, temp3758, temp3759, temp3760, temp3761, temp3762, temp3763, temp3764, temp3765, temp3766, temp3767, temp3768, temp3769, temp3770, temp3771, temp3772, temp3773, temp3774, temp3775, temp3776, temp3777, temp3778, temp3779, temp3780, temp3781, temp3782, temp3783, temp3784, temp3785, temp3786, temp3787, temp3788, temp3789, temp3790, temp3791, temp3792, temp3793, temp3794, temp3795, temp3796, temp3797, temp3798, temp3799, temp3800, temp3801, temp3802, temp3803, temp3804, temp3805, temp3806, temp3807, temp3808, temp3809, temp3810, temp3811, temp3812, temp3813, temp3814, temp3815, temp3816, temp3817, temp3818, temp3819, temp3820, temp3821, temp3822, temp3823, temp3824, temp3825, temp3826, temp3827, temp3828, temp3829, temp3830, temp3831, temp3832, temp3833, temp3834, temp3835, temp3836, temp3837, temp3838, temp3839, temp3840, temp3841, temp3842, temp3843, temp3844, temp3845, temp3846, temp3847, temp3848, temp3849, temp3850, temp3851, temp3852, temp3853, temp3854, temp3855, temp3856, temp3857, temp3858, temp3859, temp3860, temp3861, temp3862, temp3863, temp3864, temp3865, temp3866, temp3867, temp3868, temp3869, temp3870, temp3871, temp3872, temp3873, temp3874, temp3875, temp3876, temp3877, temp3878, temp3879, temp3880, temp3881, temp3882, temp3883, temp3884, temp3885, temp3886, temp3887, temp3888, temp3889, temp3890, temp3891, temp3892, temp3893, temp3894, temp3895, temp3896, temp3897, temp3898, temp3899, temp3900, temp3901, temp3902, temp3903, temp3904, temp3905, temp3906, temp3907, temp3908, temp3909, temp3910, temp3911, temp3912, temp3913, temp3914, temp3915, temp3916, temp3917, temp3918, temp3919, temp3920, temp3921, temp3922, temp3923, temp3924, temp3925, temp3926, temp3927, temp3928, temp3929, temp3930, temp3931, temp3932, temp3933, temp3934, temp3935, temp3936, temp3937, temp3938, temp3939, temp3940, temp3941, temp3942, temp3943, temp3944, temp3945, temp3946, temp3947, temp3948, temp3949, temp3950, temp3951, temp3952, temp3953, temp3954, temp3955, temp3956, temp3957, temp3958, temp3959, temp3960, temp3961, temp3962, temp3963, temp3964, temp3965, temp3966, temp3967, temp3968, temp3969, temp3970, temp3971, temp3972, temp3973, temp3974, temp3975, temp3976, temp3977, temp3978, temp3979, temp3980, temp3981, temp3982, temp3983, temp3984, temp3985, temp3986, temp3987, temp3988, temp3989, temp3990, temp3991, temp3992, temp3993, temp3994, temp3995, temp3996, temp3997, temp3998, temp3999, temp4000, temp4001, temp4002, temp4003, temp4004, temp4005, temp4006, temp4007, temp4008, temp4009, temp4010, temp4011, temp4012, temp4013, temp4014, temp4015, temp4016, temp4017, temp4018, temp4019, temp4020, temp4021, temp4022, temp4023, temp4024, temp4025, temp4026, temp4027, temp4028, temp4029, temp4030, temp4031, temp4032, temp4033, temp4034, temp4035, temp4036, temp4037, temp4038, temp4039, temp4040, temp4041, temp4042, temp4043, temp4044, temp4045, temp4046, temp4047, temp4048, temp4049, temp4050, temp4051, temp4052, temp4053, temp4054, temp4055, temp4056, temp4057, temp4058, temp4059, temp4060, temp4061, temp4062, temp4063, temp4064, temp4065, temp4066, temp4067, temp4068, temp4069, temp4070, temp4071, temp4072, temp4073, temp4074, temp4075, temp4076, temp4077, temp4078, temp4079, temp4080, temp4081, temp4082, temp4083, temp4084, temp4085, temp4086, temp4087, temp4088, temp4089, temp4090, temp4091, temp4092, temp4093, temp4094, temp4095, temp4096, temp4097, temp4098, temp4099, temp4100, temp4101, temp4102, temp4103, temp4104, temp4105, temp4106, temp4107, temp4108, temp4109, temp4110, temp4111, temp4112, temp4113, temp4114, temp4115, temp4116, temp4117, temp4118, temp4119, temp4120, temp4121, temp4122, temp4123, temp4124, temp4125, temp4126, temp4127, temp4128, temp4129, temp4130, temp4131, temp4132, temp4133, temp4134, temp4135, temp4136, temp4137, temp4138, temp4139, temp4140, temp4141, temp4142, temp4143, temp4144, temp4145, temp4146, temp4147, temp4148, temp4149, temp4150, temp4151, temp4152, temp4153, temp4154, temp4155, temp4156, temp4157, temp4158, temp4159, temp4160, temp4161, temp4162, temp4163, temp4164, temp4165, temp4166, temp4167, temp4168, temp4169, temp4170, temp4171, temp4172, temp4173, temp4174, temp4175, temp4176, temp4177, temp4178, temp4179, temp4180, temp4181, temp4182, temp4183, temp4184, temp4185, temp4186, temp4187, temp4188, temp4189, temp4190, temp4191, temp4192, temp4193, temp4194, temp4195, temp4196, temp4197, temp4198, temp4199, temp4200, temp4201, temp4202, temp4203, temp4204, temp4205, temp4206, temp4207, temp4208, temp4209, temp4210, temp4211, temp4212, temp4213, temp4214, temp4215, temp4216, temp4217, temp4218, temp4219, temp4220, temp4221, temp4222, temp4223, temp4224, temp4225, temp4226, temp4227, temp4228, temp4229, temp4230, temp4231, temp4232, temp4233, temp4234, temp4235, temp4236, temp4237, temp4238, temp4239, temp4240, temp4241, temp4242, temp4243, temp4244, temp4245, temp4246, temp4247, temp4248, temp4249, temp4250, temp4251, temp4252, temp4253, temp4254, temp4255, temp4256, temp4257, temp4258, temp4259, temp4260, temp4261, temp4262, temp4263, temp4264, temp4265, temp4266, temp4267, temp4268, temp4269, temp4270, temp4271, temp4272, temp4273, temp4274, temp4275, temp4276, temp4277, temp4278, temp4279, temp4280, temp4281, temp4282, temp4283, temp4284, temp4285, temp4286, temp4287, temp4288, temp4289, temp4290, temp4291, temp4292, temp4293, temp4294, temp4295, temp4296, temp4297, temp4298, temp4299, temp4300, temp4301, temp4302, temp4303, temp4304, temp4305, temp4306, temp4307, temp4308, temp4309, temp4310, temp4311, temp4312, temp4313, temp4314, temp4315, temp4316, temp4317, temp4318, temp4319, temp4320, temp4321, temp4322, temp4323, temp4324, temp4325, temp4326, temp4327, temp4328, temp4329, temp4330, temp4331, temp4332, temp4333, temp4334, temp4335, temp4336, temp4337, temp4338, temp4339, temp4340, temp4341, temp4342, temp4343, temp4344, temp4345, temp4346, temp4347, temp4348, temp4349, temp4350, temp4351, temp4352, temp4353, temp4354, temp4355, temp4356, temp4357, temp4358, temp4359, temp4360, temp4361, temp4362, temp4363, temp4364, temp4365, temp4366, temp4367, temp4368, temp4369, temp4370, temp4371, temp4372, temp4373, temp4374, temp4375, temp4376, temp4377, temp4378, temp4379, temp4380, temp4381, temp4382, temp4383, temp4384, temp4385, temp4386, temp4387, temp4388, temp4389, temp4390, temp4391, temp4392, temp4393, temp4394, temp4395, temp4396, temp4397, temp4398, temp4399, temp4400, temp4401, temp4402, temp4403, temp4404, temp4405, temp4406, temp4407, temp4408, temp4409, temp4410, temp4411, temp4412, temp4413, temp4414, temp4415, temp4416, temp4417, temp4418, temp4419, temp4420, temp4421, temp4422, temp4423, temp4424, temp4425, temp4426, temp4427, temp4428, temp4429, temp4430, temp4431, temp4432, temp4433, temp4434, temp4435, temp4436, temp4437, temp4438, temp4439, temp4440, temp4441, temp4442, temp4443, temp4444, temp4445, temp4446, temp4447, temp4448, temp4449, temp4450, temp4451, temp4452, temp4453, temp4454, temp4455, temp4456, temp4457, temp4458, temp4459, temp4460, temp4461, temp4462, temp4463, temp4464, temp4465, temp4466, temp4467, temp4468, temp4469, temp4470, temp4471, temp4472, temp4473, temp4474, temp4475, temp4476, temp4477, temp4478, temp4479, temp4480, temp4481, temp4482, temp4483, temp4484, temp4485, temp4486, temp4487, temp4488, temp4489, temp4490, temp4491, temp4492, temp4493, temp4494, temp4495, temp4496, temp4497, temp4498, temp4499, temp4500, temp4501, temp4502, temp4503, temp4504, temp4505, temp4506, temp4507, temp4508, temp4509, temp4510, temp4511, temp4512, temp4513, temp4514, temp4515, temp4516, temp4517, temp4518, temp4519, temp4520, temp4521, temp4522, temp4523, temp4524, temp4525, temp4526, temp4527, temp4528, temp4529, temp4530, temp4531, temp4532, temp4533, temp4534, temp4535, temp4536, temp4537, temp4538, temp4539, temp4540, temp4541, temp4542, temp4543, temp4544, temp4545, temp4546, temp4547, temp4548, temp4549, temp4550, temp4551, temp4552, temp4553, temp4554, temp4555, temp4556, temp4557, temp4558, temp4559, temp4560, temp4561, temp4562, temp4563, temp4564, temp4565, temp4566, temp4567, temp4568, temp4569, temp4570, temp4571, temp4572, temp4573, temp4574, temp4575, temp4576, temp4577, temp4578, temp4579, temp4580, temp4581, temp4582, temp4583, temp4584, temp4585, temp4586, temp4587, temp4588, temp4589, temp4590, temp4591, temp4592, temp4593, temp4594, temp4595, temp4596, temp4597, temp4598, temp4599, temp4600, temp4601, temp4602, temp4603, temp4604, temp4605, temp4606, temp4607, temp4608, temp4609, temp4610, temp4611, temp4612, temp4613, temp4614, temp4615, temp4616, temp4617, temp4618, temp4619, temp4620, temp4621, temp4622, temp4623, temp4624, temp4625, temp4626, temp4627, temp4628, temp4629, temp4630, temp4631, temp4632, temp4633, temp4634, temp4635, temp4636, temp4637, temp4638, temp4639, temp4640, temp4641, temp4642, temp4643, temp4644, temp4645, temp4646, temp4647, temp4648, temp4649, temp4650, temp4651, temp4652, temp4653, temp4654, temp4655, temp4656, temp4657, temp4658, temp4659, temp4660, temp4661, temp4662, temp4663, temp4664, temp4665, temp4666, temp4667, temp4668, temp4669, temp4670, temp4671, temp4672, temp4673, temp4674, temp4675, temp4676, temp4677, temp4678, temp4679, temp4680, temp4681, temp4682, temp4683, temp4684, temp4685, temp4686, temp4687, temp4688, temp4689, temp4690, temp4691, temp4692, temp4693, temp4694, temp4695, temp4696, temp4697, temp4698, temp4699, temp4700, temp4701, temp4702, temp4703, temp4704, temp4705, temp4706, temp4707, temp4708, temp4709, temp4710, temp4711, temp4712, temp4713, temp4714, temp4715, temp4716, temp4717, temp4718, temp4719, temp4720, temp4721, temp4722, temp4723, temp4724, temp4725, temp4726, temp4727, temp4728, temp4729, temp4730, temp4731, temp4732, temp4733, temp4734, temp4735, temp4736, temp4737, temp4738, temp4739, temp4740, temp4741, temp4742, temp4743, temp4744, temp4745, temp4746, temp4747, temp4748, temp4749, temp4750, temp4751, temp4752, temp4753, temp4754, temp4755, temp4756, temp4757, temp4758, temp4759, temp4760, temp4761, temp4762, temp4763, temp4764, temp4765, temp4766, temp4767, temp4768, temp4769, temp4770, temp4771, temp4772, temp4773, temp4774, temp4775, temp4776, temp4777, temp4778, temp4779, temp4780, temp4781, temp4782, temp4783, temp4784, temp4785, temp4786, temp4787, temp4788, temp4789, temp4790, temp4791, temp4792, temp4793, temp4794, temp4795, temp4796, temp4797, temp4798, temp4799, temp4800, temp4801, temp4802, temp4803, temp4804, temp4805, temp4806, temp4807, temp4808, temp4809, temp4810, temp4811, temp4812, temp4813, temp4814, temp4815, temp4816, temp4817, temp4818, temp4819, temp4820, temp4821, temp4822, temp4823, temp4824, temp4825, temp4826, temp4827, temp4828, temp4829, temp4830, temp4831, temp4832, temp4833, temp4834, temp4835, temp4836, temp4837, temp4838, temp4839, temp4840, temp4841, temp4842, temp4843, temp4844, temp4845, temp4846, temp4847, temp4848, temp4849, temp4850, temp4851, temp4852, temp4853, temp4854, temp4855, temp4856, temp4857, temp4858, temp4859, temp4860, temp4861, temp4862, temp4863, temp4864, temp4865, temp4866, temp4867, temp4868, temp4869, temp4870, temp4871, temp4872, temp4873, temp4874, temp4875, temp4876, temp4877, temp4878, temp4879, temp4880, temp4881, temp4882, temp4883, temp4884, temp4885, temp4886, temp4887, temp4888, temp4889, temp4890, temp4891, temp4892, temp4893, temp4894, temp4895, temp4896, temp4897, temp4898, temp4899, temp4900, temp4901, temp4902, temp4903, temp4904, temp4905, temp4906, temp4907, temp4908, temp4909, temp4910, temp4911, temp4912, temp4913, temp4914, temp4915, temp4916, temp4917, temp4918, temp4919, temp4920, temp4921, temp4922, temp4923, temp4924, temp4925, temp4926, temp4927, temp4928, temp4929, temp4930, temp4931, temp4932, temp4933, temp4934, temp4935, temp4936, temp4937, temp4938, temp4939, temp4940, temp4941, temp4942, temp4943, temp4944, temp4945, temp4946, temp4947, temp4948, temp4949, temp4950, temp4951, temp4952, temp4953, temp4954, temp4955, temp4956, temp4957, temp4958, temp4959, temp4960, temp4961, temp4962, temp4963, temp4964, temp4965, temp4966, temp4967, temp4968, temp4969, temp4970, temp4971, temp4972, temp4973, temp4974, temp4975, temp4976, temp4977, temp4978, temp4979, temp4980, temp4981, temp4982, temp4983, temp4984, temp4985, temp4986, temp4987, temp4988, temp4989, temp4990, temp4991, temp4992, temp4993, temp4994, temp4995, temp4996, temp4997, temp4998, temp4999, temp5000, temp5001, temp5002, temp5003, temp5004, temp5005, temp5006, temp5007, temp5008, temp5009, temp5010, temp5011, temp5012, temp5013, temp5014, temp5015, temp5016, temp5017, temp5018, temp5019, temp5020, temp5021, temp5022, temp5023, temp5024, temp5025, temp5026, temp5027, temp5028, temp5029, temp5030, temp5031, temp5032, temp5033, temp5034, temp5035, temp5036, temp5037, temp5038, temp5039, temp5040, temp5041, temp5042, temp5043, temp5044, temp5045, temp5046, temp5047, temp5048, temp5049, temp5050, temp5051, temp5052, temp5053, temp5054, temp5055, temp5056, temp5057, temp5058, temp5059, temp5060, temp5061, temp5062, temp5063, temp5064, temp5065, temp5066, temp5067, temp5068, temp5069, temp5070, temp5071, temp5072, temp5073, temp5074, temp5075, temp5076, temp5077, temp5078, temp5079, temp5080, temp5081, temp5082, temp5083, temp5084, temp5085, temp5086, temp5087, temp5088, temp5089, temp5090, temp5091, temp5092, temp5093, temp5094, temp5095, temp5096, temp5097, temp5098, temp5099, temp5100, temp5101, temp5102, temp5103, temp5104, temp5105, temp5106, temp5107, temp5108, temp5109, temp5110, temp5111, temp5112, temp5113, temp5114, temp5115, temp5116, temp5117, temp5118, temp5119, temp5120, temp5121, temp5122, temp5123, temp5124, temp5125, temp5126, temp5127, temp5128, temp5129, temp5130, temp5131, temp5132, temp5133, temp5134, temp5135, temp5136, temp5137, temp5138, temp5139, temp5140, temp5141, temp5142, temp5143, temp5144, temp5145, temp5146, temp5147, temp5148, temp5149, temp5150, temp5151, temp5152, temp5153, temp5154, temp5155, temp5156, temp5157, temp5158, temp5159, temp5160, temp5161, temp5162, temp5163, temp5164, temp5165, temp5166, temp5167, temp5168, temp5169, temp5170, temp5171, temp5172, temp5173, temp5174, temp5175, temp5176, temp5177, temp5178, temp5179, temp5180, temp5181, temp5182, temp5183, temp5184, temp5185, temp5186, temp5187, temp5188, temp5189, temp5190, temp5191, temp5192, temp5193, temp5194, temp5195, temp5196, temp5197, temp5198, temp5199, temp5200, temp5201, temp5202, temp5203, temp5204, temp5205, temp5206, temp5207, temp5208, temp5209, temp5210, temp5211, temp5212, temp5213, temp5214, temp5215, temp5216, temp5217, temp5218, temp5219, temp5220, temp5221, temp5222, temp5223, temp5224, temp5225, temp5226, temp5227, temp5228, temp5229, temp5230, temp5231, temp5232, temp5233, temp5234, temp5235, temp5236, temp5237, temp5238, temp5239, temp5240, temp5241, temp5242, temp5243, temp5244, temp5245, temp5246, temp5247, temp5248, temp5249, temp5250, temp5251, temp5252, temp5253, temp5254, temp5255, temp5256, temp5257, temp5258, temp5259, temp5260, temp5261, temp5262, temp5263, temp5264, temp5265, temp5266, temp5267, temp5268, temp5269, temp5270, temp5271, temp5272, temp5273, temp5274, temp5275, temp5276, temp5277, temp5278, temp5279, temp5280, temp5281, temp5282, temp5283, temp5284, temp5285, temp5286, temp5287, temp5288, temp5289, temp5290, temp5291, temp5292, temp5293, temp5294, temp5295, temp5296, temp5297, temp5298, temp5299, temp5300, temp5301, temp5302, temp5303, temp5304, temp5305, temp5306, temp5307, temp5308, temp5309, temp5310, temp5311, temp5312, temp5313, temp5314, temp5315, temp5316, temp5317, temp5318, temp5319, temp5320, temp5321, temp5322, temp5323, temp5324, temp5325, temp5326, temp5327, temp5328, temp5329, temp5330, temp5331, temp5332, temp5333, temp5334, temp5335, temp5336, temp5337, temp5338, temp5339, temp5340, temp5341, temp5342, temp5343, temp5344, temp5345, temp5346, temp5347, temp5348, temp5349, temp5350, temp5351, temp5352, temp5353, temp5354, temp5355, temp5356, temp5357, temp5358, temp5359, temp5360, temp5361, temp5362, temp5363, temp5364, temp5365, temp5366, temp5367, temp5368, temp5369, temp5370, temp5371, temp5372, temp5373, temp5374, temp5375, temp5376, temp5377, temp5378, temp5379, temp5380, temp5381, temp5382, temp5383, temp5384, temp5385, temp5386, temp5387, temp5388, temp5389, temp5390, temp5391, temp5392, temp5393, temp5394, temp5395, temp5396, temp5397, temp5398, temp5399, temp5400, temp5401, temp5402, temp5403, temp5404, temp5405, temp5406, temp5407, temp5408, temp5409, temp5410, temp5411, temp5412, temp5413, temp5414, temp5415, temp5416, temp5417, temp5418, temp5419, temp5420, temp5421, temp5422, temp5423, temp5424, temp5425, temp5426, temp5427, temp5428, temp5429, temp5430, temp5431, temp5432, temp5433, temp5434, temp5435, temp5436, temp5437, temp5438, temp5439, temp5440, temp5441, temp5442, temp5443, temp5444, temp5445, temp5446, temp5447, temp5448, temp5449, temp5450, temp5451, temp5452, temp5453, temp5454, temp5455, temp5456, temp5457, temp5458, temp5459, temp5460, temp5461, temp5462, temp5463, temp5464, temp5465, temp5466, temp5467, temp5468, temp5469, temp5470, temp5471, temp5472, temp5473, temp5474, temp5475, temp5476, temp5477, temp5478, temp5479, temp5480, temp5481, temp5482, temp5483, temp5484, temp5485, temp5486, temp5487, temp5488, temp5489, temp5490, temp5491, temp5492, temp5493, temp5494, temp5495, temp5496, temp5497, temp5498, temp5499, temp5500, temp5501, temp5502, temp5503, temp5504, temp5505, temp5506, temp5507, temp5508, temp5509, temp5510, temp5511, temp5512, temp5513, temp5514, temp5515, temp5516, temp5517, temp5518, temp5519, temp5520, temp5521, temp5522, temp5523, temp5524, temp5525, temp5526, temp5527, temp5528, temp5529, temp5530, temp5531, temp5532, temp5533, temp5534, temp5535, temp5536, temp5537, temp5538, temp5539, temp5540, temp5541, temp5542, temp5543, temp5544, temp5545, temp5546, temp5547, temp5548, temp5549, temp5550, temp5551, temp5552, temp5553, temp5554, temp5555, temp5556, temp5557, temp5558, temp5559, temp5560, temp5561, temp5562, temp5563, temp5564, temp5565, temp5566, temp5567, temp5568, temp5569, temp5570, temp5571, temp5572, temp5573, temp5574, temp5575, temp5576, temp5577, temp5578, temp5579, temp5580, temp5581, temp5582, temp5583, temp5584, temp5585, temp5586, temp5587, temp5588, temp5589, temp5590, temp5591, temp5592, temp5593, temp5594, temp5595, temp5596, temp5597, temp5598, temp5599, temp5600, temp5601, temp5602, temp5603, temp5604, temp5605, temp5606, temp5607, temp5608, temp5609, temp5610, temp5611, temp5612, temp5613, temp5614, temp5615, temp5616, temp5617, temp5618, temp5619, temp5620, temp5621, temp5622, temp5623, temp5624, temp5625, temp5626, temp5627, temp5628, temp5629, temp5630, temp5631, temp5632, temp5633, temp5634, temp5635, temp5636, temp5637, temp5638, temp5639, temp5640, temp5641, temp5642, temp5643, temp5644, temp5645, temp5646, temp5647, temp5648, temp5649, temp5650, temp5651, temp5652, temp5653, temp5654, temp5655, temp5656, temp5657, temp5658, temp5659, temp5660, temp5661, temp5662, temp5663, temp5664, temp5665, temp5666, temp5667, temp5668, temp5669, temp5670, temp5671, temp5672, temp5673, temp5674, temp5675, temp5676, temp5677, temp5678, temp5679, temp5680, temp5681, temp5682, temp5683, temp5684, temp5685, temp5686, temp5687, temp5688, temp5689, temp5690, temp5691, temp5692, temp5693, temp5694, temp5695, temp5696, temp5697, temp5698, temp5699, temp5700, temp5701, temp5702, temp5703, temp5704, temp5705, temp5706, temp5707, temp5708, temp5709, temp5710, temp5711, temp5712, temp5713, temp5714, temp5715, temp5716, temp5717, temp5718, temp5719, temp5720, temp5721, temp5722, temp5723, temp5724, temp5725, temp5726, temp5727, temp5728, temp5729, temp5730, temp5731, temp5732, temp5733, temp5734, temp5735, temp5736, temp5737, temp5738, temp5739, temp5740, temp5741, temp5742, temp5743, temp5744, temp5745, temp5746, temp5747, temp5748, temp5749, temp5750, temp5751, temp5752, temp5753, temp5754, temp5755, temp5756, temp5757, temp5758, temp5759, temp5760, temp5761, temp5762, temp5763, temp5764, temp5765, temp5766, temp5767, temp5768, temp5769, temp5770, temp5771, temp5772, temp5773, temp5774, temp5775, temp5776, temp5777, temp5778, temp5779, temp5780, temp5781, temp5782, temp5783, temp5784, temp5785, temp5786, temp5787, temp5788, temp5789, temp5790, temp5791, temp5792, temp5793, temp5794, temp5795, temp5796, temp5797, temp5798, temp5799, temp5800, temp5801, temp5802, temp5803, temp5804, temp5805, temp5806, temp5807, temp5808, temp5809, temp5810, temp5811, temp5812, temp5813, temp5814, temp5815, temp5816, temp5817, temp5818, temp5819, temp5820, temp5821, temp5822, temp5823, temp5824, temp5825, temp5826, temp5827, temp5828, temp5829, temp5830, temp5831, temp5832, temp5833, temp5834, temp5835, temp5836, temp5837, temp5838, temp5839, temp5840, temp5841, temp5842, temp5843, temp5844, temp5845, temp5846, temp5847, temp5848, temp5849, temp5850, temp5851, temp5852, temp5853, temp5854, temp5855, temp5856, temp5857, temp5858, temp5859, temp5860, temp5861, temp5862, temp5863, temp5864, temp5865, temp5866, temp5867, temp5868, temp5869, temp5870, temp5871, temp5872, temp5873, temp5874, temp5875, temp5876, temp5877, temp5878, temp5879, temp5880, temp5881, temp5882, temp5883, temp5884, temp5885, temp5886, temp5887, temp5888, temp5889, temp5890, temp5891, temp5892, temp5893, temp5894, temp5895, temp5896, temp5897, temp5898, temp5899, temp5900, temp5901, temp5902, temp5903, temp5904, temp5905, temp5906, temp5907, temp5908, temp5909, temp5910, temp5911, temp5912, temp5913, temp5914, temp5915, temp5916, temp5917, temp5918, temp5919, temp5920, temp5921, temp5922, temp5923, temp5924, temp5925, temp5926, temp5927, temp5928, temp5929, temp5930, temp5931, temp5932, temp5933, temp5934, temp5935, temp5936, temp5937, temp5938, temp5939, temp5940, temp5941, temp5942, temp5943, temp5944, temp5945, temp5946, temp5947, temp5948, temp5949, temp5950, temp5951, temp5952, temp5953, temp5954, temp5955, temp5956, temp5957, temp5958, temp5959, temp5960, temp5961, temp5962, temp5963, temp5964, temp5965, temp5966, temp5967, temp5968, temp5969, temp5970, temp5971, temp5972, temp5973, temp5974, temp5975, temp5976, temp5977, temp5978, temp5979, temp5980, temp5981, temp5982, temp5983, temp5984, temp5985, temp5986, temp5987, temp5988, temp5989, temp5990, temp5991, temp5992, temp5993, temp5994, temp5995, temp5996, temp5997, temp5998, temp5999, temp6000, temp6001, temp6002, temp6003, temp6004, temp6005, temp6006, temp6007, temp6008, temp6009, temp6010, temp6011, temp6012, temp6013, temp6014, temp6015, temp6016, temp6017, temp6018, temp6019, temp6020, temp6021, temp6022, temp6023, temp6024, temp6025, temp6026, temp6027, temp6028, temp6029, temp6030, temp6031, temp6032, temp6033, temp6034, temp6035, temp6036, temp6037, temp6038, temp6039, temp6040, temp6041, temp6042, temp6043, temp6044, temp6045, temp6046, temp6047, temp6048, temp6049, temp6050, temp6051, temp6052, temp6053, temp6054, temp6055, temp6056, temp6057, temp6058, temp6059, temp6060, temp6061, temp6062, temp6063, temp6064, temp6065, temp6066, temp6067, temp6068, temp6069, temp6070, temp6071, temp6072, temp6073, temp6074, temp6075, temp6076, temp6077, temp6078, temp6079, temp6080, temp6081, temp6082, temp6083, temp6084, temp6085, temp6086, temp6087, temp6088, temp6089, temp6090, temp6091, temp6092, temp6093, temp6094, temp6095, temp6096, temp6097, temp6098, temp6099, temp6100, temp6101, temp6102, temp6103, temp6104, temp6105, temp6106, temp6107, temp6108, temp6109, temp6110, temp6111, temp6112, temp6113, temp6114, temp6115, temp6116, temp6117, temp6118, temp6119, temp6120, temp6121, temp6122, temp6123, temp6124, temp6125, temp6126, temp6127, temp6128, temp6129, temp6130, temp6131, temp6132, temp6133, temp6134, temp6135, temp6136, temp6137, temp6138, temp6139, temp6140, temp6141, temp6142, temp6143, temp6144, temp6145, temp6146, temp6147, temp6148, temp6149, temp6150, temp6151, temp6152, temp6153, temp6154, temp6155, temp6156, temp6157, temp6158, temp6159, temp6160, temp6161, temp6162, temp6163, temp6164, temp6165, temp6166, temp6167, temp6168, temp6169, temp6170, temp6171, temp6172, temp6173, temp6174, temp6175, temp6176, temp6177, temp6178, temp6179, temp6180, temp6181, temp6182, temp6183, temp6184, temp6185, temp6186, temp6187, temp6188, temp6189, temp6190, temp6191, temp6192, temp6193, temp6194, temp6195, temp6196, temp6197, temp6198, temp6199, temp6200, temp6201, temp6202, temp6203, temp6204, temp6205, temp6206, temp6207, temp6208, temp6209, temp6210, temp6211, temp6212, temp6213, temp6214, temp6215, temp6216, temp6217, temp6218, temp6219, temp6220, temp6221, temp6222, temp6223, temp6224, temp6225, temp6226, temp6227, temp6228, temp6229, temp6230, temp6231, temp6232, temp6233, temp6234, temp6235, temp6236, temp6237, temp6238, temp6239, temp6240, temp6241, temp6242, temp6243, temp6244, temp6245, temp6246, temp6247, temp6248, temp6249, temp6250, temp6251, temp6252, temp6253, temp6254, temp6255, temp6256, temp6257, temp6258, temp6259, temp6260, temp6261, temp6262, temp6263, temp6264, temp6265, temp6266, temp6267, temp6268, temp6269, temp6270, temp6271, temp6272, temp6273, temp6274, temp6275, temp6276, temp6277, temp6278, temp6279, temp6280, temp6281, temp6282, temp6283, temp6284, temp6285, temp6286, temp6287, temp6288, temp6289, temp6290, temp6291, temp6292, temp6293, temp6294, temp6295, temp6296, temp6297, temp6298, temp6299, temp6300, temp6301, temp6302, temp6303, temp6304, temp6305, temp6306, temp6307, temp6308, temp6309, temp6310, temp6311, temp6312, temp6313, temp6314, temp6315, temp6316, temp6317, temp6318, temp6319, temp6320, temp6321, temp6322, temp6323, temp6324, temp6325, temp6326, temp6327, temp6328, temp6329, temp6330, temp6331, temp6332, temp6333, temp6334, temp6335, temp6336, temp6337, temp6338, temp6339, temp6340, temp6341, temp6342, temp6343, temp6344, temp6345, temp6346, temp6347, temp6348, temp6349, temp6350, temp6351, temp6352, temp6353, temp6354, temp6355, temp6356, temp6357, temp6358, temp6359, temp6360, temp6361, temp6362, temp6363, temp6364, temp6365, temp6366, temp6367, temp6368, temp6369, temp6370, temp6371, temp6372, temp6373, temp6374, temp6375, temp6376, temp6377, temp6378, temp6379, temp6380, temp6381, temp6382, temp6383, temp6384, temp6385, temp6386, temp6387, temp6388, temp6389, temp6390, temp6391, temp6392, temp6393, temp6394, temp6395, temp6396, temp6397, temp6398, temp6399, temp6400, temp6401, temp6402, temp6403, temp6404, temp6405, temp6406, temp6407, temp6408, temp6409, temp6410, temp6411, temp6412, temp6413, temp6414, temp6415, temp6416, temp6417, temp6418, temp6419, temp6420, temp6421, temp6422, temp6423, temp6424, temp6425, temp6426, temp6427, temp6428, temp6429, temp6430, temp6431, temp6432, temp6433, temp6434, temp6435, temp6436, temp6437, temp6438, temp6439, temp6440, temp6441, temp6442, temp6443, temp6444, temp6445, temp6446, temp6447, temp6448, temp6449, temp6450, temp6451, temp6452, temp6453, temp6454, temp6455, temp6456, temp6457, temp6458, temp6459, temp6460, temp6461, temp6462, temp6463, temp6464, temp6465, temp6466, temp6467, temp6468, temp6469, temp6470, temp6471, temp6472, temp6473, temp6474, temp6475, temp6476, temp6477, temp6478, temp6479, temp6480, temp6481, temp6482, temp6483, temp6484, temp6485, temp6486, temp6487, temp6488, temp6489, temp6490, temp6491, temp6492, temp6493, temp6494, temp6495, temp6496, temp6497, temp6498, temp6499, temp6500, temp6501, temp6502, temp6503, temp6504, temp6505, temp6506, temp6507, temp6508, temp6509, temp6510, temp6511, temp6512, temp6513, temp6514, temp6515, temp6516, temp6517, temp6518, temp6519, temp6520, temp6521, temp6522, temp6523, temp6524, temp6525, temp6526, temp6527, temp6528, temp6529, temp6530, temp6531, temp6532, temp6533, temp6534, temp6535, temp6536, temp6537, temp6538, temp6539, temp6540, temp6541, temp6542, temp6543, temp6544, temp6545, temp6546, temp6547, temp6548, temp6549, temp6550, temp6551, temp6552, temp6553, temp6554, temp6555, temp6556, temp6557, temp6558, temp6559, temp6560, temp6561, temp6562, temp6563, temp6564, temp6565, temp6566, temp6567, temp6568, temp6569, temp6570, temp6571, temp6572, temp6573, temp6574, temp6575, temp6576, temp6577, temp6578, temp6579, temp6580, temp6581, temp6582, temp6583, temp6584, temp6585, temp6586, temp6587, temp6588, temp6589, temp6590, temp6591, temp6592, temp6593, temp6594, temp6595, temp6596, temp6597, temp6598, temp6599, temp6600, temp6601, temp6602, temp6603, temp6604, temp6605, temp6606, temp6607, temp6608, temp6609, temp6610, temp6611, temp6612, temp6613, temp6614, temp6615, temp6616, temp6617, temp6618, temp6619, temp6620, temp6621, temp6622, temp6623, temp6624, temp6625, temp6626, temp6627, temp6628, temp6629, temp6630, temp6631, temp6632, temp6633, temp6634, temp6635, temp6636, temp6637, temp6638, temp6639, temp6640, temp6641, temp6642, temp6643, temp6644, temp6645, temp6646, temp6647, temp6648, temp6649, temp6650, temp6651, temp6652, temp6653, temp6654, temp6655, temp6656, temp6657, temp6658, temp6659, temp6660, temp6661, temp6662, temp6663, temp6664, temp6665, temp6666, temp6667, temp6668, temp6669, temp6670, temp6671, temp6672, temp6673, temp6674, temp6675, temp6676, temp6677, temp6678, temp6679, temp6680, temp6681, temp6682, temp6683, temp6684, temp6685, temp6686, temp6687, temp6688, temp6689, temp6690, temp6691, temp6692, temp6693, temp6694, temp6695, temp6696, temp6697, temp6698, temp6699, temp6700, temp6701, temp6702, temp6703, temp6704, temp6705, temp6706, temp6707, temp6708, temp6709, temp6710, temp6711, temp6712, temp6713, temp6714, temp6715, temp6716, temp6717, temp6718, temp6719, temp6720, temp6721, temp6722, temp6723, temp6724, temp6725, temp6726, temp6727, temp6728, temp6729, temp6730, temp6731, temp6732, temp6733, temp6734, temp6735, temp6736, temp6737, temp6738, temp6739, temp6740, temp6741, temp6742, temp6743, temp6744, temp6745, temp6746, temp6747, temp6748, temp6749, temp6750, temp6751, temp6752, temp6753, temp6754, temp6755, temp6756, temp6757, temp6758, temp6759, temp6760, temp6761, temp6762, temp6763, temp6764, temp6765, temp6766, temp6767, temp6768, temp6769, temp6770, temp6771, temp6772, temp6773, temp6774, temp6775, temp6776, temp6777, temp6778, temp6779, temp6780, temp6781, temp6782, temp6783, temp6784, temp6785, temp6786, temp6787, temp6788, temp6789, temp6790, temp6791, temp6792, temp6793, temp6794, temp6795, temp6796, temp6797, temp6798, temp6799, temp6800, temp6801, temp6802, temp6803, temp6804, temp6805, temp6806, temp6807, temp6808, temp6809, temp6810, temp6811, temp6812, temp6813, temp6814, temp6815, temp6816, temp6817, temp6818, temp6819, temp6820, temp6821, temp6822, temp6823, temp6824, temp6825, temp6826, temp6827, temp6828, temp6829, temp6830, temp6831, temp6832, temp6833, temp6834, temp6835, temp6836, temp6837, temp6838, temp6839, temp6840, temp6841, temp6842, temp6843, temp6844, temp6845, temp6846, temp6847, temp6848, temp6849, temp6850, temp6851, temp6852, temp6853, temp6854, temp6855, temp6856, temp6857, temp6858, temp6859, temp6860, temp6861, temp6862, temp6863, temp6864, temp6865, temp6866, temp6867, temp6868, temp6869, temp6870, temp6871, temp6872, temp6873, temp6874, temp6875, temp6876, temp6877, temp6878, temp6879, temp6880, temp6881, temp6882, temp6883, temp6884, temp6885, temp6886, temp6887, temp6888, temp6889, temp6890, temp6891, temp6892, temp6893, temp6894, temp6895, temp6896, temp6897, temp6898, temp6899, temp6900, temp6901, temp6902, temp6903, temp6904, temp6905, temp6906, temp6907, temp6908, temp6909, temp6910, temp6911, temp6912, temp6913, temp6914, temp6915, temp6916, temp6917, temp6918, temp6919, temp6920, temp6921, temp6922, temp6923, temp6924, temp6925, temp6926, temp6927, temp6928, temp6929, temp6930, temp6931, temp6932, temp6933, temp6934, temp6935, temp6936, temp6937, temp6938, temp6939, temp6940, temp6941, temp6942, temp6943, temp6944, temp6945, temp6946, temp6947, temp6948, temp6949, temp6950, temp6951, temp6952, temp6953, temp6954, temp6955, temp6956, temp6957, temp6958, temp6959, temp6960, temp6961, temp6962, temp6963, temp6964, temp6965, temp6966, temp6967, temp6968, temp6969, temp6970, temp6971, temp6972, temp6973, temp6974, temp6975, temp6976, temp6977, temp6978, temp6979, temp6980, temp6981, temp6982, temp6983, temp6984, temp6985, temp6986, temp6987, temp6988, temp6989, temp6990, temp6991, temp6992, temp6993, temp6994, temp6995, temp6996, temp6997, temp6998, temp6999, temp7000, temp7001, temp7002, temp7003, temp7004, temp7005, temp7006, temp7007, temp7008, temp7009, temp7010, temp7011, temp7012, temp7013, temp7014, temp7015, temp7016, temp7017, temp7018, temp7019, temp7020, temp7021, temp7022, temp7023, temp7024, temp7025, temp7026, temp7027, temp7028, temp7029, temp7030, temp7031, temp7032, temp7033, temp7034, temp7035, temp7036, temp7037, temp7038, temp7039, temp7040, temp7041, temp7042, temp7043, temp7044, temp7045, temp7046, temp7047, temp7048, temp7049, temp7050, temp7051, temp7052, temp7053, temp7054, temp7055, temp7056, temp7057, temp7058, temp7059, temp7060, temp7061, temp7062, temp7063, temp7064, temp7065, temp7066, temp7067, temp7068, temp7069, temp7070, temp7071, temp7072, temp7073, temp7074, temp7075, temp7076, temp7077, temp7078, temp7079, temp7080, temp7081, temp7082, temp7083, temp7084, temp7085, temp7086, temp7087, temp7088, temp7089, temp7090, temp7091, temp7092, temp7093, temp7094, temp7095, temp7096, temp7097, temp7098, temp7099, temp7100, temp7101, temp7102, temp7103, temp7104, temp7105, temp7106, temp7107, temp7108, temp7109, temp7110, temp7111, temp7112, temp7113, temp7114, temp7115, temp7116, temp7117, temp7118, temp7119, temp7120, temp7121, temp7122, temp7123, temp7124, temp7125, temp7126, temp7127, temp7128, temp7129, temp7130, temp7131, temp7132, temp7133, temp7134, temp7135, temp7136, temp7137, temp7138, temp7139, temp7140, temp7141, temp7142, temp7143, temp7144, temp7145, temp7146, temp7147, temp7148, temp7149, temp7150, temp7151, temp7152, temp7153, temp7154, temp7155, temp7156, temp7157, temp7158, temp7159, temp7160, temp7161, temp7162, temp7163, temp7164, temp7165, temp7166, temp7167, temp7168, temp7169, temp7170, temp7171, temp7172, temp7173, temp7174, temp7175, temp7176, temp7177, temp7178, temp7179, temp7180, temp7181, temp7182, temp7183, temp7184, temp7185, temp7186, temp7187, temp7188, temp7189, temp7190, temp7191, temp7192, temp7193, temp7194, temp7195, temp7196, temp7197, temp7198, temp7199, temp7200, temp7201, temp7202, temp7203, temp7204, temp7205, temp7206, temp7207, temp7208, temp7209, temp7210, temp7211, temp7212, temp7213, temp7214, temp7215, temp7216, temp7217, temp7218, temp7219, temp7220, temp7221, temp7222, temp7223, temp7224, temp7225, temp7226, temp7227, temp7228, temp7229, temp7230, temp7231, temp7232, temp7233, temp7234, temp7235, temp7236, temp7237, temp7238, temp7239, temp7240, temp7241, temp7242, temp7243, temp7244, temp7245, temp7246, temp7247, temp7248, temp7249, temp7250, temp7251, temp7252, temp7253, temp7254, temp7255, temp7256, temp7257, temp7258, temp7259, temp7260, temp7261, temp7262, temp7263, temp7264, temp7265, temp7266, temp7267, temp7268, temp7269, temp7270, temp7271, temp7272, temp7273, temp7274, temp7275, temp7276, temp7277, temp7278, temp7279, temp7280, temp7281, temp7282, temp7283, temp7284, temp7285, temp7286, temp7287, temp7288, temp7289, temp7290, temp7291, temp7292, temp7293, temp7294, temp7295, temp7296, temp7297, temp7298, temp7299, temp7300, temp7301, temp7302, temp7303, temp7304, temp7305, temp7306, temp7307, temp7308, temp7309, temp7310, temp7311, temp7312, temp7313, temp7314, temp7315, temp7316, temp7317, temp7318, temp7319, temp7320, temp7321, temp7322, temp7323, temp7324, temp7325, temp7326, temp7327, temp7328, temp7329, temp7330, temp7331, temp7332, temp7333, temp7334, temp7335, temp7336, temp7337, temp7338, temp7339, temp7340, temp7341, temp7342, temp7343, temp7344, temp7345, temp7346, temp7347, temp7348, temp7349, temp7350, temp7351, temp7352, temp7353, temp7354, temp7355, temp7356, temp7357, temp7358, temp7359, temp7360, temp7361, temp7362, temp7363, temp7364, temp7365, temp7366, temp7367, temp7368, temp7369, temp7370, temp7371, temp7372, temp7373, temp7374, temp7375, temp7376, temp7377, temp7378, temp7379, temp7380, temp7381, temp7382, temp7383, temp7384, temp7385, temp7386, temp7387, temp7388, temp7389, temp7390, temp7391, temp7392, temp7393, temp7394, temp7395, temp7396, temp7397, temp7398, temp7399, temp7400, temp7401, temp7402, temp7403, temp7404, temp7405, temp7406, temp7407, temp7408, temp7409, temp7410, temp7411, temp7412, temp7413, temp7414, temp7415, temp7416, temp7417, temp7418, temp7419, temp7420, temp7421, temp7422, temp7423, temp7424, temp7425, temp7426, temp7427, temp7428, temp7429, temp7430, temp7431, temp7432, temp7433, temp7434, temp7435, temp7436, temp7437, temp7438, temp7439, temp7440, temp7441, temp7442, temp7443, temp7444, temp7445, temp7446, temp7447, temp7448, temp7449, temp7450, temp7451, temp7452, temp7453, temp7454, temp7455, temp7456, temp7457, temp7458, temp7459, temp7460, temp7461, temp7462, temp7463, temp7464, temp7465, temp7466, temp7467, temp7468, temp7469, temp7470, temp7471, temp7472, temp7473, temp7474, temp7475, temp7476, temp7477, temp7478, temp7479, temp7480, temp7481, temp7482, temp7483, temp7484, temp7485, temp7486, temp7487, temp7488, temp7489, temp7490, temp7491, temp7492, temp7493, temp7494, temp7495, temp7496, temp7497, temp7498, temp7499, temp7500, temp7501, temp7502, temp7503, temp7504, temp7505, temp7506, temp7507, temp7508, temp7509, temp7510, temp7511, temp7512, temp7513, temp7514, temp7515, temp7516, temp7517, temp7518, temp7519, temp7520, temp7521, temp7522, temp7523, temp7524, temp7525, temp7526, temp7527, temp7528, temp7529, temp7530, temp7531, temp7532, temp7533, temp7534, temp7535, temp7536, temp7537, temp7538, temp7539, temp7540, temp7541, temp7542, temp7543, temp7544, temp7545, temp7546, temp7547, temp7548, temp7549, temp7550, temp7551, temp7552, temp7553, temp7554, temp7555, temp7556, temp7557, temp7558, temp7559, temp7560, temp7561, temp7562, temp7563, temp7564, temp7565, temp7566, temp7567, temp7568, temp7569, temp7570, temp7571, temp7572, temp7573, temp7574, temp7575, temp7576, temp7577, temp7578, temp7579, temp7580, temp7581, temp7582, temp7583, temp7584, temp7585, temp7586, temp7587, temp7588, temp7589, temp7590, temp7591, temp7592, temp7593, temp7594, temp7595, temp7596, temp7597, temp7598, temp7599, temp7600, temp7601, temp7602, temp7603, temp7604, temp7605, temp7606, temp7607, temp7608, temp7609, temp7610, temp7611, temp7612, temp7613, temp7614, temp7615, temp7616, temp7617, temp7618, temp7619, temp7620, temp7621, temp7622, temp7623, temp7624, temp7625, temp7626, temp7627, temp7628, temp7629, temp7630, temp7631, temp7632, temp7633, temp7634, temp7635, temp7636, temp7637, temp7638, temp7639, temp7640, temp7641, temp7642, temp7643, temp7644, temp7645, temp7646, temp7647, temp7648, temp7649, temp7650, temp7651, temp7652, temp7653, temp7654, temp7655, temp7656, temp7657, temp7658, temp7659, temp7660, temp7661, temp7662, temp7663, temp7664, temp7665, temp7666, temp7667, temp7668, temp7669, temp7670, temp7671, temp7672, temp7673, temp7674, temp7675, temp7676, temp7677, temp7678, temp7679, temp7680, temp7681, temp7682, temp7683, temp7684, temp7685, temp7686, temp7687, temp7688, temp7689, temp7690, temp7691, temp7692, temp7693, temp7694, temp7695, temp7696, temp7697, temp7698, temp7699, temp7700, temp7701, temp7702, temp7703, temp7704, temp7705, temp7706, temp7707, temp7708, temp7709, temp7710, temp7711, temp7712, temp7713, temp7714, temp7715, temp7716, temp7717, temp7718, temp7719, temp7720, temp7721, temp7722, temp7723, temp7724, temp7725, temp7726, temp7727, temp7728, temp7729, temp7730, temp7731, temp7732, temp7733, temp7734, temp7735, temp7736, temp7737, temp7738, temp7739, temp7740, temp7741, temp7742, temp7743, temp7744, temp7745, temp7746, temp7747, temp7748, temp7749, temp7750, temp7751, temp7752, temp7753, temp7754, temp7755, temp7756, temp7757, temp7758, temp7759, temp7760, temp7761, temp7762, temp7763, temp7764, temp7765, temp7766, temp7767, temp7768, temp7769, temp7770, temp7771, temp7772, temp7773, temp7774, temp7775, temp7776, temp7777, temp7778, temp7779, temp7780, temp7781, temp7782, temp7783, temp7784, temp7785, temp7786, temp7787, temp7788, temp7789, temp7790, temp7791, temp7792, temp7793, temp7794, temp7795, temp7796, temp7797, temp7798, temp7799, temp7800, temp7801, temp7802, temp7803, temp7804, temp7805, temp7806, temp7807, temp7808, temp7809, temp7810, temp7811, temp7812, temp7813, temp7814, temp7815, temp7816, temp7817, temp7818, temp7819, temp7820, temp7821, temp7822, temp7823, temp7824, temp7825, temp7826, temp7827, temp7828, temp7829, temp7830, temp7831, temp7832, temp7833, temp7834, temp7835, temp7836, temp7837, temp7838, temp7839, temp7840, temp7841, temp7842, temp7843, temp7844, temp7845, temp7846, temp7847, temp7848, temp7849, temp7850, temp7851, temp7852, temp7853, temp7854, temp7855, temp7856, temp7857, temp7858, temp7859, temp7860, temp7861, temp7862, temp7863, temp7864, temp7865, temp7866, temp7867, temp7868, temp7869, temp7870, temp7871, temp7872, temp7873, temp7874, temp7875, temp7876, temp7877, temp7878, temp7879, temp7880, temp7881, temp7882, temp7883, temp7884, temp7885, temp7886, temp7887, temp7888, temp7889, temp7890, temp7891, temp7892, temp7893, temp7894, temp7895, temp7896, temp7897, temp7898, temp7899, temp7900, temp7901, temp7902, temp7903, temp7904, temp7905, temp7906, temp7907, temp7908, temp7909, temp7910, temp7911, temp7912, temp7913, temp7914, temp7915, temp7916, temp7917, temp7918, temp7919, temp7920, temp7921, temp7922, temp7923, temp7924, temp7925, temp7926, temp7927, temp7928, temp7929, temp7930, temp7931, temp7932, temp7933, temp7934, temp7935, temp7936, temp7937, temp7938, temp7939, temp7940, temp7941, temp7942, temp7943, temp7944, temp7945, temp7946, temp7947, temp7948, temp7949, temp7950, temp7951, temp7952, temp7953, temp7954, temp7955, temp7956, temp7957, temp7958, temp7959, temp7960, temp7961, temp7962, temp7963, temp7964, temp7965, temp7966, temp7967, temp7968, temp7969, temp7970, temp7971, temp7972, temp7973, temp7974, temp7975, temp7976, temp7977, temp7978, temp7979, temp7980, temp7981, temp7982, temp7983, temp7984, temp7985, temp7986, temp7987, temp7988, temp7989, temp7990, temp7991, temp7992, temp7993, temp7994, temp7995, temp7996, temp7997, temp7998, temp7999, temp8000, temp8001, temp8002, temp8003, temp8004, temp8005, temp8006, temp8007, temp8008, temp8009, temp8010, temp8011, temp8012, temp8013, temp8014, temp8015, temp8016, temp8017, temp8018, temp8019, temp8020, temp8021, temp8022, temp8023, temp8024, temp8025, temp8026, temp8027, temp8028, temp8029, temp8030, temp8031, temp8032, temp8033, temp8034, temp8035, temp8036, temp8037, temp8038, temp8039, temp8040, temp8041, temp8042, temp8043, temp8044, temp8045, temp8046, temp8047, temp8048, temp8049, temp8050, temp8051, temp8052, temp8053, temp8054, temp8055, temp8056, temp8057, temp8058, temp8059, temp8060, temp8061, temp8062, temp8063, temp8064, temp8065, temp8066, temp8067, temp8068, temp8069, temp8070, temp8071, temp8072, temp8073, temp8074, temp8075, temp8076, temp8077, temp8078, temp8079, temp8080, temp8081, temp8082, temp8083, temp8084, temp8085, temp8086, temp8087, temp8088, temp8089, temp8090, temp8091, temp8092, temp8093, temp8094, temp8095, temp8096, temp8097, temp8098, temp8099, temp8100, temp8101, temp8102, temp8103, temp8104, temp8105, temp8106, temp8107, temp8108, temp8109, temp8110, temp8111, temp8112, temp8113, temp8114, temp8115, temp8116, temp8117, temp8118, temp8119, temp8120, temp8121, temp8122, temp8123, temp8124, temp8125, temp8126, temp8127, temp8128, temp8129, temp8130, temp8131, temp8132, temp8133, temp8134, temp8135, temp8136, temp8137, temp8138, temp8139, temp8140, temp8141, temp8142, temp8143, temp8144, temp8145, temp8146, temp8147, temp8148, temp8149, temp8150, temp8151, temp8152, temp8153, temp8154, temp8155, temp8156, temp8157, temp8158, temp8159, temp8160, temp8161, temp8162, temp8163, temp8164, temp8165, temp8166, temp8167, temp8168, temp8169, temp8170, temp8171, temp8172, temp8173, temp8174, temp8175, temp8176, temp8177, temp8178, temp8179, temp8180, temp8181, temp8182, temp8183, temp8184, temp8185, temp8186, temp8187, temp8188, temp8189, temp8190, temp8191, temp8192, temp8193, temp8194, temp8195, temp8196, temp8197, temp8198, temp8199, temp8200, temp8201, temp8202, temp8203, temp8204, temp8205, temp8206, temp8207, temp8208, temp8209, temp8210, temp8211, temp8212, temp8213, temp8214, temp8215, temp8216, temp8217, temp8218, temp8219, temp8220, temp8221, temp8222, temp8223, temp8224, temp8225, temp8226, temp8227, temp8228, temp8229, temp8230, temp8231, temp8232, temp8233, temp8234, temp8235, temp8236, temp8237, temp8238, temp8239, temp8240, temp8241, temp8242, temp8243, temp8244, temp8245, temp8246, temp8247, temp8248, temp8249, temp8250, temp8251, temp8252, temp8253, temp8254, temp8255, temp8256, temp8257, temp8258, temp8259, temp8260, temp8261, temp8262, temp8263, temp8264, temp8265, temp8266, temp8267, temp8268, temp8269, temp8270, temp8271, temp8272, temp8273, temp8274, temp8275, temp8276, temp8277, temp8278, temp8279, temp8280, temp8281, temp8282, temp8283, temp8284, temp8285, temp8286, temp8287, temp8288, temp8289, temp8290, temp8291, temp8292, temp8293, temp8294, temp8295, temp8296, temp8297, temp8298, temp8299, temp8300, temp8301, temp8302, temp8303, temp8304, temp8305, temp8306, temp8307, temp8308, temp8309, temp8310, temp8311, temp8312, temp8313, temp8314, temp8315, temp8316, temp8317, temp8318, temp8319, temp8320, temp8321, temp8322, temp8323, temp8324, temp8325, temp8326, temp8327, temp8328, temp8329, temp8330, temp8331, temp8332, temp8333, temp8334, temp8335, temp8336, temp8337, temp8338, temp8339, temp8340, temp8341, temp8342, temp8343, temp8344, temp8345, temp8346, temp8347, temp8348, temp8349, temp8350, temp8351, temp8352, temp8353, temp8354, temp8355, temp8356, temp8357, temp8358, temp8359, temp8360, temp8361, temp8362, temp8363, temp8364, temp8365, temp8366, temp8367, temp8368, temp8369, temp8370, temp8371, temp8372, temp8373, temp8374, temp8375, temp8376, temp8377, temp8378, temp8379, temp8380, temp8381, temp8382, temp8383, temp8384, temp8385, temp8386, temp8387, temp8388, temp8389, temp8390, temp8391, temp8392, temp8393, temp8394, temp8395, temp8396, temp8397, temp8398, temp8399, temp8400, temp8401, temp8402, temp8403, temp8404, temp8405, temp8406, temp8407, temp8408, temp8409, temp8410, temp8411, temp8412, temp8413, temp8414, temp8415, temp8416, temp8417, temp8418, temp8419, temp8420, temp8421, temp8422, temp8423, temp8424, temp8425, temp8426, temp8427, temp8428, temp8429, temp8430, temp8431, temp8432, temp8433, temp8434, temp8435, temp8436, temp8437, temp8438, temp8439, temp8440, temp8441, temp8442, temp8443, temp8444, temp8445, temp8446, temp8447, temp8448, temp8449, temp8450, temp8451, temp8452, temp8453, temp8454, temp8455, temp8456, temp8457, temp8458, temp8459, temp8460, temp8461, temp8462, temp8463, temp8464, temp8465, temp8466, temp8467, temp8468, temp8469, temp8470, temp8471, temp8472, temp8473, temp8474, temp8475, temp8476, temp8477, temp8478, temp8479, temp8480, temp8481, temp8482, temp8483, temp8484, temp8485, temp8486, temp8487, temp8488, temp8489, temp8490, temp8491, temp8492, temp8493, temp8494, temp8495, temp8496, temp8497, temp8498, temp8499, temp8500, temp8501, temp8502, temp8503, temp8504, temp8505, temp8506, temp8507, temp8508, temp8509, temp8510, temp8511, temp8512, temp8513, temp8514, temp8515, temp8516, temp8517, temp8518, temp8519, temp8520, temp8521, temp8522, temp8523, temp8524, temp8525, temp8526, temp8527, temp8528, temp8529, temp8530, temp8531, temp8532, temp8533, temp8534, temp8535, temp8536, temp8537, temp8538, temp8539, temp8540, temp8541, temp8542, temp8543, temp8544, temp8545, temp8546, temp8547, temp8548, temp8549, temp8550, temp8551, temp8552, temp8553, temp8554, temp8555, temp8556, temp8557, temp8558, temp8559, temp8560, temp8561, temp8562, temp8563, temp8564, temp8565, temp8566, temp8567, temp8568, temp8569, temp8570, temp8571, temp8572, temp8573, temp8574, temp8575, temp8576, temp8577, temp8578, temp8579, temp8580, temp8581, temp8582, temp8583, temp8584, temp8585, temp8586, temp8587, temp8588, temp8589, temp8590, temp8591, temp8592, temp8593, temp8594, temp8595, temp8596, temp8597, temp8598, temp8599, temp8600, temp8601, temp8602, temp8603, temp8604, temp8605, temp8606, temp8607, temp8608, temp8609, temp8610, temp8611, temp8612, temp8613, temp8614, temp8615, temp8616, temp8617, temp8618, temp8619, temp8620, temp8621, temp8622, temp8623, temp8624, temp8625, temp8626, temp8627, temp8628, temp8629, temp8630, temp8631, temp8632, temp8633, temp8634, temp8635, temp8636, temp8637, temp8638, temp8639, temp8640, temp8641, temp8642, temp8643, temp8644, temp8645, temp8646, temp8647, temp8648, temp8649, temp8650, temp8651, temp8652, temp8653, temp8654, temp8655, temp8656, temp8657, temp8658, temp8659, temp8660, temp8661, temp8662, temp8663, temp8664, temp8665, temp8666, temp8667, temp8668, temp8669, temp8670, temp8671, temp8672, temp8673, temp8674, temp8675, temp8676, temp8677, temp8678, temp8679, temp8680, temp8681, temp8682, temp8683, temp8684, temp8685, temp8686, temp8687, temp8688, temp8689, temp8690, temp8691, temp8692, temp8693, temp8694, temp8695, temp8696, temp8697, temp8698, temp8699, temp8700, temp8701, temp8702, temp8703, temp8704, temp8705, temp8706, temp8707, temp8708, temp8709, temp8710, temp8711, temp8712, temp8713, temp8714, temp8715, temp8716, temp8717, temp8718, temp8719, temp8720, temp8721, temp8722, temp8723, temp8724, temp8725, temp8726, temp8727, temp8728, temp8729, temp8730, temp8731, temp8732, temp8733, temp8734, temp8735, temp8736, temp8737, temp8738, temp8739, temp8740, temp8741, temp8742, temp8743, temp8744, temp8745, temp8746, temp8747, temp8748, temp8749, temp8750, temp8751, temp8752, temp8753, temp8754, temp8755, temp8756, temp8757, temp8758, temp8759, temp8760, temp8761, temp8762, temp8763, temp8764, temp8765, temp8766, temp8767, temp8768, temp8769, temp8770, temp8771, temp8772, temp8773, temp8774, temp8775, temp8776, temp8777, temp8778, temp8779, temp8780, temp8781, temp8782, temp8783, temp8784, temp8785, temp8786, temp8787, temp8788, temp8789, temp8790, temp8791, temp8792, temp8793, temp8794, temp8795, temp8796, temp8797, temp8798, temp8799, temp8800, temp8801, temp8802, temp8803, temp8804, temp8805, temp8806, temp8807, temp8808, temp8809, temp8810, temp8811, temp8812, temp8813, temp8814, temp8815, temp8816, temp8817, temp8818, temp8819, temp8820, temp8821, temp8822, temp8823, temp8824, temp8825, temp8826, temp8827, temp8828, temp8829, temp8830, temp8831, temp8832, temp8833, temp8834, temp8835, temp8836, temp8837, temp8838, temp8839, temp8840, temp8841, temp8842, temp8843, temp8844, temp8845, temp8846, temp8847, temp8848, temp8849, temp8850, temp8851, temp8852, temp8853, temp8854, temp8855, temp8856, temp8857, temp8858, temp8859, temp8860, temp8861, temp8862, temp8863, temp8864, temp8865, temp8866, temp8867, temp8868, temp8869, temp8870, temp8871, temp8872, temp8873, temp8874, temp8875, temp8876, temp8877, temp8878, temp8879, temp8880, temp8881, temp8882, temp8883, temp8884, temp8885, temp8886, temp8887, temp8888, temp8889, temp8890, temp8891, temp8892, temp8893, temp8894, temp8895, temp8896, temp8897, temp8898, temp8899, temp8900, temp8901, temp8902, temp8903, temp8904, temp8905, temp8906, temp8907, temp8908, temp8909, temp8910, temp8911, temp8912, temp8913, temp8914, temp8915, temp8916, temp8917, temp8918, temp8919, temp8920, temp8921, temp8922, temp8923, temp8924, temp8925, temp8926, temp8927, temp8928, temp8929, temp8930, temp8931, temp8932, temp8933, temp8934, temp8935, temp8936, temp8937, temp8938, temp8939, temp8940, temp8941, temp8942, temp8943, temp8944, temp8945, temp8946, temp8947, temp8948, temp8949, temp8950, temp8951, temp8952, temp8953, temp8954, temp8955, temp8956, temp8957, temp8958, temp8959, temp8960, temp8961, temp8962, temp8963, temp8964, temp8965, temp8966, temp8967, temp8968, temp8969, temp8970, temp8971, temp8972, temp8973, temp8974, temp8975, temp8976, temp8977, temp8978, temp8979, temp8980, temp8981, temp8982, temp8983, temp8984, temp8985, temp8986, temp8987, temp8988, temp8989, temp8990, temp8991, temp8992, temp8993, temp8994, temp8995, temp8996, temp8997, temp8998, temp8999, temp9000, temp9001, temp9002, temp9003, temp9004, temp9005, temp9006, temp9007, temp9008, temp9009, temp9010, temp9011, temp9012, temp9013, temp9014, temp9015, temp9016, temp9017, temp9018, temp9019, temp9020, temp9021, temp9022, temp9023, temp9024, temp9025, temp9026, temp9027, temp9028, temp9029, temp9030, temp9031, temp9032, temp9033, temp9034, temp9035, temp9036, temp9037, temp9038, temp9039, temp9040, temp9041, temp9042, temp9043, temp9044, temp9045, temp9046, temp9047, temp9048, temp9049, temp9050, temp9051, temp9052, temp9053, temp9054, temp9055, temp9056, temp9057, temp9058, temp9059, temp9060, temp9061, temp9062, temp9063, temp9064, temp9065, temp9066, temp9067, temp9068, temp9069, temp9070, temp9071, temp9072, temp9073, temp9074, temp9075, temp9076, temp9077, temp9078, temp9079, temp9080, temp9081, temp9082, temp9083, temp9084, temp9085, temp9086, temp9087, temp9088, temp9089, temp9090, temp9091, temp9092, temp9093, temp9094, temp9095, temp9096, temp9097, temp9098, temp9099, temp9100, temp9101, temp9102, temp9103, temp9104, temp9105, temp9106, temp9107, temp9108, temp9109, temp9110, temp9111, temp9112, temp9113, temp9114, temp9115, temp9116, temp9117, temp9118, temp9119, temp9120, temp9121, temp9122, temp9123, temp9124, temp9125, temp9126, temp9127, temp9128, temp9129, temp9130, temp9131, temp9132, temp9133, temp9134, temp9135, temp9136, temp9137, temp9138, temp9139, temp9140, temp9141, temp9142, temp9143, temp9144, temp9145, temp9146, temp9147, temp9148, temp9149, temp9150, temp9151, temp9152, temp9153, temp9154, temp9155, temp9156, temp9157, temp9158, temp9159, temp9160, temp9161, temp9162, temp9163, temp9164, temp9165, temp9166, temp9167, temp9168, temp9169, temp9170, temp9171, temp9172, temp9173, temp9174, temp9175, temp9176, temp9177, temp9178, temp9179, temp9180, temp9181, temp9182, temp9183, temp9184, temp9185, temp9186, temp9187, temp9188, temp9189, temp9190, temp9191, temp9192, temp9193, temp9194, temp9195, temp9196, temp9197, temp9198, temp9199, temp9200, temp9201, temp9202, temp9203, temp9204, temp9205, temp9206, temp9207, temp9208, temp9209, temp9210, temp9211, temp9212, temp9213, temp9214, temp9215, temp9216, temp9217, temp9218, temp9219, temp9220, temp9221, temp9222, temp9223, temp9224, temp9225, temp9226, temp9227, temp9228, temp9229, temp9230, temp9231, temp9232, temp9233, temp9234, temp9235, temp9236, temp9237, temp9238, temp9239, temp9240, temp9241, temp9242, temp9243, temp9244, temp9245, temp9246, temp9247, temp9248, temp9249, temp9250, temp9251, temp9252, temp9253, temp9254, temp9255, temp9256, temp9257, temp9258, temp9259, temp9260, temp9261, temp9262, temp9263, temp9264, temp9265, temp9266, temp9267, temp9268, temp9269, temp9270, temp9271, temp9272, temp9273, temp9274, temp9275, temp9276, temp9277, temp9278, temp9279, temp9280, temp9281, temp9282, temp9283, temp9284, temp9285, temp9286, temp9287, temp9288, temp9289, temp9290, temp9291, temp9292, temp9293, temp9294, temp9295, temp9296, temp9297, temp9298, temp9299, temp9300, temp9301, temp9302, temp9303, temp9304, temp9305, temp9306, temp9307, temp9308, temp9309, temp9310, temp9311, temp9312, temp9313, temp9314, temp9315, temp9316, temp9317, temp9318, temp9319, temp9320, temp9321, temp9322, temp9323, temp9324, temp9325, temp9326, temp9327, temp9328, temp9329, temp9330, temp9331, temp9332, temp9333, temp9334, temp9335, temp9336, temp9337, temp9338, temp9339, temp9340, temp9341, temp9342, temp9343, temp9344, temp9345, temp9346, temp9347, temp9348, temp9349, temp9350, temp9351, temp9352, temp9353, temp9354, temp9355, temp9356, temp9357, temp9358, temp9359, temp9360, temp9361, temp9362, temp9363, temp9364, temp9365, temp9366, temp9367, temp9368, temp9369, temp9370, temp9371, temp9372, temp9373, temp9374, temp9375, temp9376, temp9377, temp9378, temp9379, temp9380, temp9381, temp9382, temp9383, temp9384, temp9385, temp9386, temp9387, temp9388, temp9389, temp9390, temp9391, temp9392, temp9393, temp9394, temp9395, temp9396, temp9397, temp9398, temp9399, temp9400, temp9401, temp9402, temp9403, temp9404, temp9405, temp9406, temp9407, temp9408, temp9409, temp9410, temp9411, temp9412, temp9413, temp9414, temp9415, temp9416, temp9417, temp9418, temp9419, temp9420, temp9421, temp9422, temp9423, temp9424, temp9425, temp9426, temp9427, temp9428, temp9429, temp9430, temp9431, temp9432, temp9433, temp9434, temp9435, temp9436, temp9437, temp9438, temp9439, temp9440, temp9441, temp9442, temp9443, temp9444, temp9445, temp9446, temp9447, temp9448, temp9449, temp9450, temp9451, temp9452, temp9453, temp9454, temp9455, temp9456, temp9457, temp9458, temp9459, temp9460, temp9461, temp9462, temp9463, temp9464, temp9465, temp9466, temp9467, temp9468, temp9469, temp9470, temp9471, temp9472, temp9473, temp9474, temp9475, temp9476, temp9477, temp9478, temp9479, temp9480, temp9481, temp9482, temp9483, temp9484, temp9485, temp9486, temp9487, temp9488, temp9489, temp9490, temp9491, temp9492, temp9493, temp9494, temp9495, temp9496, temp9497, temp9498, temp9499, temp9500, temp9501, temp9502, temp9503, temp9504, temp9505, temp9506, temp9507, temp9508, temp9509, temp9510, temp9511, temp9512, temp9513, temp9514, temp9515, temp9516, temp9517, temp9518, temp9519, temp9520, temp9521, temp9522, temp9523, temp9524, temp9525, temp9526, temp9527, temp9528, temp9529, temp9530, temp9531, temp9532, temp9533, temp9534, temp9535, temp9536, temp9537, temp9538, temp9539, temp9540, temp9541, temp9542, temp9543, temp9544, temp9545, temp9546, temp9547, temp9548, temp9549, temp9550, temp9551, temp9552, temp9553, temp9554, temp9555, temp9556, temp9557, temp9558, temp9559, temp9560, temp9561, temp9562, temp9563, temp9564, temp9565, temp9566, temp9567, temp9568, temp9569, temp9570, temp9571, temp9572, temp9573, temp9574, temp9575, temp9576, temp9577, temp9578, temp9579, temp9580, temp9581, temp9582, temp9583, temp9584, temp9585, temp9586, temp9587, temp9588, temp9589, temp9590, temp9591, temp9592, temp9593, temp9594, temp9595, temp9596, temp9597, temp9598, temp9599, temp9600, temp9601, temp9602, temp9603, temp9604, temp9605, temp9606, temp9607, temp9608, temp9609, temp9610, temp9611, temp9612, temp9613, temp9614, temp9615, temp9616, temp9617, temp9618, temp9619, temp9620, temp9621, temp9622, temp9623, temp9624, temp9625, temp9626, temp9627, temp9628, temp9629, temp9630, temp9631, temp9632, temp9633, temp9634, temp9635, temp9636, temp9637, temp9638, temp9639, temp9640, temp9641, temp9642, temp9643, temp9644, temp9645, temp9646, temp9647, temp9648, temp9649, temp9650, temp9651, temp9652, temp9653, temp9654, temp9655, temp9656, temp9657, temp9658, temp9659, temp9660, temp9661, temp9662, temp9663, temp9664, temp9665, temp9666, temp9667, temp9668, temp9669, temp9670, temp9671, temp9672, temp9673, temp9674, temp9675, temp9676, temp9677, temp9678, temp9679, temp9680, temp9681, temp9682, temp9683, temp9684, temp9685, temp9686, temp9687, temp9688, temp9689, temp9690, temp9691, temp9692, temp9693, temp9694, temp9695, temp9696, temp9697, temp9698, temp9699, temp9700, temp9701, temp9702, temp9703, temp9704, temp9705, temp9706, temp9707, temp9708, temp9709, temp9710, temp9711, temp9712, temp9713, temp9714, temp9715, temp9716, temp9717, temp9718, temp9719, temp9720, temp9721, temp9722, temp9723, temp9724, temp9725, temp9726, temp9727, temp9728, temp9729, temp9730, temp9731, temp9732, temp9733, temp9734, temp9735, temp9736, temp9737, temp9738, temp9739, temp9740, temp9741, temp9742, temp9743, temp9744, temp9745, temp9746, temp9747, temp9748, temp9749, temp9750, temp9751, temp9752, temp9753, temp9754, temp9755, temp9756, temp9757, temp9758, temp9759, temp9760, temp9761, temp9762, temp9763, temp9764, temp9765, temp9766, temp9767, temp9768, temp9769, temp9770, temp9771, temp9772, temp9773, temp9774, temp9775, temp9776, temp9777, temp9778, temp9779, temp9780, temp9781, temp9782, temp9783, temp9784, temp9785, temp9786, temp9787, temp9788, temp9789, temp9790, temp9791, temp9792, temp9793, temp9794, temp9795, temp9796, temp9797, temp9798, temp9799, temp9800, temp9801, temp9802, temp9803, temp9804, temp9805, temp9806, temp9807, temp9808, temp9809, temp9810, temp9811, temp9812, temp9813, temp9814, temp9815, temp9816, temp9817, temp9818, temp9819, temp9820, temp9821, temp9822, temp9823, temp9824, temp9825, temp9826, temp9827, temp9828, temp9829, temp9830, temp9831, temp9832, temp9833, temp9834, temp9835, temp9836, temp9837, temp9838, temp9839, temp9840, temp9841, temp9842, temp9843, temp9844, temp9845, temp9846, temp9847, temp9848, temp9849, temp9850, temp9851, temp9852, temp9853, temp9854, temp9855, temp9856, temp9857, temp9858, temp9859, temp9860, temp9861, temp9862, temp9863, temp9864, temp9865, temp9866, temp9867, temp9868, temp9869, temp9870, temp9871, temp9872, temp9873, temp9874, temp9875, temp9876, temp9877, temp9878, temp9879, temp9880, temp9881, temp9882, temp9883, temp9884, temp9885, temp9886, temp9887, temp9888, temp9889, temp9890, temp9891, temp9892, temp9893, temp9894, temp9895, temp9896, temp9897, temp9898, temp9899, temp9900, temp9901, temp9902, temp9903, temp9904, temp9905, temp9906, temp9907, temp9908, temp9909, temp9910, temp9911, temp9912, temp9913, temp9914, temp9915, temp9916, temp9917, temp9918, temp9919, temp9920, temp9921, temp9922, temp9923, temp9924, temp9925, temp9926, temp9927, temp9928, temp9929, temp9930, temp9931, temp9932, temp9933, temp9934, temp9935, temp9936, temp9937, temp9938, temp9939, temp9940, temp9941, temp9942, temp9943, temp9944, temp9945, temp9946, temp9947, temp9948, temp9949, temp9950, temp9951, temp9952, temp9953, temp9954, temp9955, temp9956, temp9957, temp9958, temp9959, temp9960, temp9961, temp9962, temp9963, temp9964, temp9965, temp9966, temp9967, temp9968, temp9969, temp9970, temp9971, temp9972, temp9973, temp9974, temp9975, temp9976, temp9977, temp9978, temp9979, temp9980, temp9981, temp9982, temp9983, temp9984, temp9985, temp9986, temp9987, temp9988, temp9989, temp9990, temp9991, temp9992, temp9993, temp9994, temp9995, temp9996, temp9997, temp9998;
    assign temp0 = a ^ b;
    assign temp1 = temp0 ^ temp0;
    assign temp2 = temp1 ^ temp1;
    assign temp3 = temp2 ^ temp2;
    assign temp4 = temp3 ^ temp3;
    assign temp5 = temp4 ^ temp4;
    assign temp6 = temp5 ^ temp5;
    assign temp7 = temp6 ^ temp6;
    assign temp8 = temp7 ^ temp7;
    assign temp9 = temp8 ^ temp8;
    assign temp10 = temp9 ^ temp9;
    assign temp11 = temp10 ^ temp10;
    assign temp12 = temp11 ^ temp11;
    assign temp13 = temp12 ^ temp12;
    assign temp14 = temp13 ^ temp13;
    assign temp15 = temp14 ^ temp14;
    assign temp16 = temp15 ^ temp15;
    assign temp17 = temp16 ^ temp16;
    assign temp18 = temp17 ^ temp17;
    assign temp19 = temp18 ^ temp18;
    assign temp20 = temp19 ^ temp19;
    assign temp21 = temp20 ^ temp20;
    assign temp22 = temp21 ^ temp21;
    assign temp23 = temp22 ^ temp22;
    assign temp24 = temp23 ^ temp23;
    assign temp25 = temp24 ^ temp24;
    assign temp26 = temp25 ^ temp25;
    assign temp27 = temp26 ^ temp26;
    assign temp28 = temp27 ^ temp27;
    assign temp29 = temp28 ^ temp28;
    assign temp30 = temp29 ^ temp29;
    assign temp31 = temp30 ^ temp30;
    assign temp32 = temp31 ^ temp31;
    assign temp33 = temp32 ^ temp32;
    assign temp34 = temp33 ^ temp33;
    assign temp35 = temp34 ^ temp34;
    assign temp36 = temp35 ^ temp35;
    assign temp37 = temp36 ^ temp36;
    assign temp38 = temp37 ^ temp37;
    assign temp39 = temp38 ^ temp38;
    assign temp40 = temp39 ^ temp39;
    assign temp41 = temp40 ^ temp40;
    assign temp42 = temp41 ^ temp41;
    assign temp43 = temp42 ^ temp42;
    assign temp44 = temp43 ^ temp43;
    assign temp45 = temp44 ^ temp44;
    assign temp46 = temp45 ^ temp45;
    assign temp47 = temp46 ^ temp46;
    assign temp48 = temp47 ^ temp47;
    assign temp49 = temp48 ^ temp48;
    assign temp50 = temp49 ^ temp49;
    assign temp51 = temp50 ^ temp50;
    assign temp52 = temp51 ^ temp51;
    assign temp53 = temp52 ^ temp52;
    assign temp54 = temp53 ^ temp53;
    assign temp55 = temp54 ^ temp54;
    assign temp56 = temp55 ^ temp55;
    assign temp57 = temp56 ^ temp56;
    assign temp58 = temp57 ^ temp57;
    assign temp59 = temp58 ^ temp58;
    assign temp60 = temp59 ^ temp59;
    assign temp61 = temp60 ^ temp60;
    assign temp62 = temp61 ^ temp61;
    assign temp63 = temp62 ^ temp62;
    assign temp64 = temp63 ^ temp63;
    assign temp65 = temp64 ^ temp64;
    assign temp66 = temp65 ^ temp65;
    assign temp67 = temp66 ^ temp66;
    assign temp68 = temp67 ^ temp67;
    assign temp69 = temp68 ^ temp68;
    assign temp70 = temp69 ^ temp69;
    assign temp71 = temp70 ^ temp70;
    assign temp72 = temp71 ^ temp71;
    assign temp73 = temp72 ^ temp72;
    assign temp74 = temp73 ^ temp73;
    assign temp75 = temp74 ^ temp74;
    assign temp76 = temp75 ^ temp75;
    assign temp77 = temp76 ^ temp76;
    assign temp78 = temp77 ^ temp77;
    assign temp79 = temp78 ^ temp78;
    assign temp80 = temp79 ^ temp79;
    assign temp81 = temp80 ^ temp80;
    assign temp82 = temp81 ^ temp81;
    assign temp83 = temp82 ^ temp82;
    assign temp84 = temp83 ^ temp83;
    assign temp85 = temp84 ^ temp84;
    assign temp86 = temp85 ^ temp85;
    assign temp87 = temp86 ^ temp86;
    assign temp88 = temp87 ^ temp87;
    assign temp89 = temp88 ^ temp88;
    assign temp90 = temp89 ^ temp89;
    assign temp91 = temp90 ^ temp90;
    assign temp92 = temp91 ^ temp91;
    assign temp93 = temp92 ^ temp92;
    assign temp94 = temp93 ^ temp93;
    assign temp95 = temp94 ^ temp94;
    assign temp96 = temp95 ^ temp95;
    assign temp97 = temp96 ^ temp96;
    assign temp98 = temp97 ^ temp97;
    assign temp99 = temp98 ^ temp98;
    assign temp100 = temp99 ^ temp99;
    assign temp101 = temp100 ^ temp100;
    assign temp102 = temp101 ^ temp101;
    assign temp103 = temp102 ^ temp102;
    assign temp104 = temp103 ^ temp103;
    assign temp105 = temp104 ^ temp104;
    assign temp106 = temp105 ^ temp105;
    assign temp107 = temp106 ^ temp106;
    assign temp108 = temp107 ^ temp107;
    assign temp109 = temp108 ^ temp108;
    assign temp110 = temp109 ^ temp109;
    assign temp111 = temp110 ^ temp110;
    assign temp112 = temp111 ^ temp111;
    assign temp113 = temp112 ^ temp112;
    assign temp114 = temp113 ^ temp113;
    assign temp115 = temp114 ^ temp114;
    assign temp116 = temp115 ^ temp115;
    assign temp117 = temp116 ^ temp116;
    assign temp118 = temp117 ^ temp117;
    assign temp119 = temp118 ^ temp118;
    assign temp120 = temp119 ^ temp119;
    assign temp121 = temp120 ^ temp120;
    assign temp122 = temp121 ^ temp121;
    assign temp123 = temp122 ^ temp122;
    assign temp124 = temp123 ^ temp123;
    assign temp125 = temp124 ^ temp124;
    assign temp126 = temp125 ^ temp125;
    assign temp127 = temp126 ^ temp126;
    assign temp128 = temp127 ^ temp127;
    assign temp129 = temp128 ^ temp128;
    assign temp130 = temp129 ^ temp129;
    assign temp131 = temp130 ^ temp130;
    assign temp132 = temp131 ^ temp131;
    assign temp133 = temp132 ^ temp132;
    assign temp134 = temp133 ^ temp133;
    assign temp135 = temp134 ^ temp134;
    assign temp136 = temp135 ^ temp135;
    assign temp137 = temp136 ^ temp136;
    assign temp138 = temp137 ^ temp137;
    assign temp139 = temp138 ^ temp138;
    assign temp140 = temp139 ^ temp139;
    assign temp141 = temp140 ^ temp140;
    assign temp142 = temp141 ^ temp141;
    assign temp143 = temp142 ^ temp142;
    assign temp144 = temp143 ^ temp143;
    assign temp145 = temp144 ^ temp144;
    assign temp146 = temp145 ^ temp145;
    assign temp147 = temp146 ^ temp146;
    assign temp148 = temp147 ^ temp147;
    assign temp149 = temp148 ^ temp148;
    assign temp150 = temp149 ^ temp149;
    assign temp151 = temp150 ^ temp150;
    assign temp152 = temp151 ^ temp151;
    assign temp153 = temp152 ^ temp152;
    assign temp154 = temp153 ^ temp153;
    assign temp155 = temp154 ^ temp154;
    assign temp156 = temp155 ^ temp155;
    assign temp157 = temp156 ^ temp156;
    assign temp158 = temp157 ^ temp157;
    assign temp159 = temp158 ^ temp158;
    assign temp160 = temp159 ^ temp159;
    assign temp161 = temp160 ^ temp160;
    assign temp162 = temp161 ^ temp161;
    assign temp163 = temp162 ^ temp162;
    assign temp164 = temp163 ^ temp163;
    assign temp165 = temp164 ^ temp164;
    assign temp166 = temp165 ^ temp165;
    assign temp167 = temp166 ^ temp166;
    assign temp168 = temp167 ^ temp167;
    assign temp169 = temp168 ^ temp168;
    assign temp170 = temp169 ^ temp169;
    assign temp171 = temp170 ^ temp170;
    assign temp172 = temp171 ^ temp171;
    assign temp173 = temp172 ^ temp172;
    assign temp174 = temp173 ^ temp173;
    assign temp175 = temp174 ^ temp174;
    assign temp176 = temp175 ^ temp175;
    assign temp177 = temp176 ^ temp176;
    assign temp178 = temp177 ^ temp177;
    assign temp179 = temp178 ^ temp178;
    assign temp180 = temp179 ^ temp179;
    assign temp181 = temp180 ^ temp180;
    assign temp182 = temp181 ^ temp181;
    assign temp183 = temp182 ^ temp182;
    assign temp184 = temp183 ^ temp183;
    assign temp185 = temp184 ^ temp184;
    assign temp186 = temp185 ^ temp185;
    assign temp187 = temp186 ^ temp186;
    assign temp188 = temp187 ^ temp187;
    assign temp189 = temp188 ^ temp188;
    assign temp190 = temp189 ^ temp189;
    assign temp191 = temp190 ^ temp190;
    assign temp192 = temp191 ^ temp191;
    assign temp193 = temp192 ^ temp192;
    assign temp194 = temp193 ^ temp193;
    assign temp195 = temp194 ^ temp194;
    assign temp196 = temp195 ^ temp195;
    assign temp197 = temp196 ^ temp196;
    assign temp198 = temp197 ^ temp197;
    assign temp199 = temp198 ^ temp198;
    assign temp200 = temp199 ^ temp199;
    assign temp201 = temp200 ^ temp200;
    assign temp202 = temp201 ^ temp201;
    assign temp203 = temp202 ^ temp202;
    assign temp204 = temp203 ^ temp203;
    assign temp205 = temp204 ^ temp204;
    assign temp206 = temp205 ^ temp205;
    assign temp207 = temp206 ^ temp206;
    assign temp208 = temp207 ^ temp207;
    assign temp209 = temp208 ^ temp208;
    assign temp210 = temp209 ^ temp209;
    assign temp211 = temp210 ^ temp210;
    assign temp212 = temp211 ^ temp211;
    assign temp213 = temp212 ^ temp212;
    assign temp214 = temp213 ^ temp213;
    assign temp215 = temp214 ^ temp214;
    assign temp216 = temp215 ^ temp215;
    assign temp217 = temp216 ^ temp216;
    assign temp218 = temp217 ^ temp217;
    assign temp219 = temp218 ^ temp218;
    assign temp220 = temp219 ^ temp219;
    assign temp221 = temp220 ^ temp220;
    assign temp222 = temp221 ^ temp221;
    assign temp223 = temp222 ^ temp222;
    assign temp224 = temp223 ^ temp223;
    assign temp225 = temp224 ^ temp224;
    assign temp226 = temp225 ^ temp225;
    assign temp227 = temp226 ^ temp226;
    assign temp228 = temp227 ^ temp227;
    assign temp229 = temp228 ^ temp228;
    assign temp230 = temp229 ^ temp229;
    assign temp231 = temp230 ^ temp230;
    assign temp232 = temp231 ^ temp231;
    assign temp233 = temp232 ^ temp232;
    assign temp234 = temp233 ^ temp233;
    assign temp235 = temp234 ^ temp234;
    assign temp236 = temp235 ^ temp235;
    assign temp237 = temp236 ^ temp236;
    assign temp238 = temp237 ^ temp237;
    assign temp239 = temp238 ^ temp238;
    assign temp240 = temp239 ^ temp239;
    assign temp241 = temp240 ^ temp240;
    assign temp242 = temp241 ^ temp241;
    assign temp243 = temp242 ^ temp242;
    assign temp244 = temp243 ^ temp243;
    assign temp245 = temp244 ^ temp244;
    assign temp246 = temp245 ^ temp245;
    assign temp247 = temp246 ^ temp246;
    assign temp248 = temp247 ^ temp247;
    assign temp249 = temp248 ^ temp248;
    assign temp250 = temp249 ^ temp249;
    assign temp251 = temp250 ^ temp250;
    assign temp252 = temp251 ^ temp251;
    assign temp253 = temp252 ^ temp252;
    assign temp254 = temp253 ^ temp253;
    assign temp255 = temp254 ^ temp254;
    assign temp256 = temp255 ^ temp255;
    assign temp257 = temp256 ^ temp256;
    assign temp258 = temp257 ^ temp257;
    assign temp259 = temp258 ^ temp258;
    assign temp260 = temp259 ^ temp259;
    assign temp261 = temp260 ^ temp260;
    assign temp262 = temp261 ^ temp261;
    assign temp263 = temp262 ^ temp262;
    assign temp264 = temp263 ^ temp263;
    assign temp265 = temp264 ^ temp264;
    assign temp266 = temp265 ^ temp265;
    assign temp267 = temp266 ^ temp266;
    assign temp268 = temp267 ^ temp267;
    assign temp269 = temp268 ^ temp268;
    assign temp270 = temp269 ^ temp269;
    assign temp271 = temp270 ^ temp270;
    assign temp272 = temp271 ^ temp271;
    assign temp273 = temp272 ^ temp272;
    assign temp274 = temp273 ^ temp273;
    assign temp275 = temp274 ^ temp274;
    assign temp276 = temp275 ^ temp275;
    assign temp277 = temp276 ^ temp276;
    assign temp278 = temp277 ^ temp277;
    assign temp279 = temp278 ^ temp278;
    assign temp280 = temp279 ^ temp279;
    assign temp281 = temp280 ^ temp280;
    assign temp282 = temp281 ^ temp281;
    assign temp283 = temp282 ^ temp282;
    assign temp284 = temp283 ^ temp283;
    assign temp285 = temp284 ^ temp284;
    assign temp286 = temp285 ^ temp285;
    assign temp287 = temp286 ^ temp286;
    assign temp288 = temp287 ^ temp287;
    assign temp289 = temp288 ^ temp288;
    assign temp290 = temp289 ^ temp289;
    assign temp291 = temp290 ^ temp290;
    assign temp292 = temp291 ^ temp291;
    assign temp293 = temp292 ^ temp292;
    assign temp294 = temp293 ^ temp293;
    assign temp295 = temp294 ^ temp294;
    assign temp296 = temp295 ^ temp295;
    assign temp297 = temp296 ^ temp296;
    assign temp298 = temp297 ^ temp297;
    assign temp299 = temp298 ^ temp298;
    assign temp300 = temp299 ^ temp299;
    assign temp301 = temp300 ^ temp300;
    assign temp302 = temp301 ^ temp301;
    assign temp303 = temp302 ^ temp302;
    assign temp304 = temp303 ^ temp303;
    assign temp305 = temp304 ^ temp304;
    assign temp306 = temp305 ^ temp305;
    assign temp307 = temp306 ^ temp306;
    assign temp308 = temp307 ^ temp307;
    assign temp309 = temp308 ^ temp308;
    assign temp310 = temp309 ^ temp309;
    assign temp311 = temp310 ^ temp310;
    assign temp312 = temp311 ^ temp311;
    assign temp313 = temp312 ^ temp312;
    assign temp314 = temp313 ^ temp313;
    assign temp315 = temp314 ^ temp314;
    assign temp316 = temp315 ^ temp315;
    assign temp317 = temp316 ^ temp316;
    assign temp318 = temp317 ^ temp317;
    assign temp319 = temp318 ^ temp318;
    assign temp320 = temp319 ^ temp319;
    assign temp321 = temp320 ^ temp320;
    assign temp322 = temp321 ^ temp321;
    assign temp323 = temp322 ^ temp322;
    assign temp324 = temp323 ^ temp323;
    assign temp325 = temp324 ^ temp324;
    assign temp326 = temp325 ^ temp325;
    assign temp327 = temp326 ^ temp326;
    assign temp328 = temp327 ^ temp327;
    assign temp329 = temp328 ^ temp328;
    assign temp330 = temp329 ^ temp329;
    assign temp331 = temp330 ^ temp330;
    assign temp332 = temp331 ^ temp331;
    assign temp333 = temp332 ^ temp332;
    assign temp334 = temp333 ^ temp333;
    assign temp335 = temp334 ^ temp334;
    assign temp336 = temp335 ^ temp335;
    assign temp337 = temp336 ^ temp336;
    assign temp338 = temp337 ^ temp337;
    assign temp339 = temp338 ^ temp338;
    assign temp340 = temp339 ^ temp339;
    assign temp341 = temp340 ^ temp340;
    assign temp342 = temp341 ^ temp341;
    assign temp343 = temp342 ^ temp342;
    assign temp344 = temp343 ^ temp343;
    assign temp345 = temp344 ^ temp344;
    assign temp346 = temp345 ^ temp345;
    assign temp347 = temp346 ^ temp346;
    assign temp348 = temp347 ^ temp347;
    assign temp349 = temp348 ^ temp348;
    assign temp350 = temp349 ^ temp349;
    assign temp351 = temp350 ^ temp350;
    assign temp352 = temp351 ^ temp351;
    assign temp353 = temp352 ^ temp352;
    assign temp354 = temp353 ^ temp353;
    assign temp355 = temp354 ^ temp354;
    assign temp356 = temp355 ^ temp355;
    assign temp357 = temp356 ^ temp356;
    assign temp358 = temp357 ^ temp357;
    assign temp359 = temp358 ^ temp358;
    assign temp360 = temp359 ^ temp359;
    assign temp361 = temp360 ^ temp360;
    assign temp362 = temp361 ^ temp361;
    assign temp363 = temp362 ^ temp362;
    assign temp364 = temp363 ^ temp363;
    assign temp365 = temp364 ^ temp364;
    assign temp366 = temp365 ^ temp365;
    assign temp367 = temp366 ^ temp366;
    assign temp368 = temp367 ^ temp367;
    assign temp369 = temp368 ^ temp368;
    assign temp370 = temp369 ^ temp369;
    assign temp371 = temp370 ^ temp370;
    assign temp372 = temp371 ^ temp371;
    assign temp373 = temp372 ^ temp372;
    assign temp374 = temp373 ^ temp373;
    assign temp375 = temp374 ^ temp374;
    assign temp376 = temp375 ^ temp375;
    assign temp377 = temp376 ^ temp376;
    assign temp378 = temp377 ^ temp377;
    assign temp379 = temp378 ^ temp378;
    assign temp380 = temp379 ^ temp379;
    assign temp381 = temp380 ^ temp380;
    assign temp382 = temp381 ^ temp381;
    assign temp383 = temp382 ^ temp382;
    assign temp384 = temp383 ^ temp383;
    assign temp385 = temp384 ^ temp384;
    assign temp386 = temp385 ^ temp385;
    assign temp387 = temp386 ^ temp386;
    assign temp388 = temp387 ^ temp387;
    assign temp389 = temp388 ^ temp388;
    assign temp390 = temp389 ^ temp389;
    assign temp391 = temp390 ^ temp390;
    assign temp392 = temp391 ^ temp391;
    assign temp393 = temp392 ^ temp392;
    assign temp394 = temp393 ^ temp393;
    assign temp395 = temp394 ^ temp394;
    assign temp396 = temp395 ^ temp395;
    assign temp397 = temp396 ^ temp396;
    assign temp398 = temp397 ^ temp397;
    assign temp399 = temp398 ^ temp398;
    assign temp400 = temp399 ^ temp399;
    assign temp401 = temp400 ^ temp400;
    assign temp402 = temp401 ^ temp401;
    assign temp403 = temp402 ^ temp402;
    assign temp404 = temp403 ^ temp403;
    assign temp405 = temp404 ^ temp404;
    assign temp406 = temp405 ^ temp405;
    assign temp407 = temp406 ^ temp406;
    assign temp408 = temp407 ^ temp407;
    assign temp409 = temp408 ^ temp408;
    assign temp410 = temp409 ^ temp409;
    assign temp411 = temp410 ^ temp410;
    assign temp412 = temp411 ^ temp411;
    assign temp413 = temp412 ^ temp412;
    assign temp414 = temp413 ^ temp413;
    assign temp415 = temp414 ^ temp414;
    assign temp416 = temp415 ^ temp415;
    assign temp417 = temp416 ^ temp416;
    assign temp418 = temp417 ^ temp417;
    assign temp419 = temp418 ^ temp418;
    assign temp420 = temp419 ^ temp419;
    assign temp421 = temp420 ^ temp420;
    assign temp422 = temp421 ^ temp421;
    assign temp423 = temp422 ^ temp422;
    assign temp424 = temp423 ^ temp423;
    assign temp425 = temp424 ^ temp424;
    assign temp426 = temp425 ^ temp425;
    assign temp427 = temp426 ^ temp426;
    assign temp428 = temp427 ^ temp427;
    assign temp429 = temp428 ^ temp428;
    assign temp430 = temp429 ^ temp429;
    assign temp431 = temp430 ^ temp430;
    assign temp432 = temp431 ^ temp431;
    assign temp433 = temp432 ^ temp432;
    assign temp434 = temp433 ^ temp433;
    assign temp435 = temp434 ^ temp434;
    assign temp436 = temp435 ^ temp435;
    assign temp437 = temp436 ^ temp436;
    assign temp438 = temp437 ^ temp437;
    assign temp439 = temp438 ^ temp438;
    assign temp440 = temp439 ^ temp439;
    assign temp441 = temp440 ^ temp440;
    assign temp442 = temp441 ^ temp441;
    assign temp443 = temp442 ^ temp442;
    assign temp444 = temp443 ^ temp443;
    assign temp445 = temp444 ^ temp444;
    assign temp446 = temp445 ^ temp445;
    assign temp447 = temp446 ^ temp446;
    assign temp448 = temp447 ^ temp447;
    assign temp449 = temp448 ^ temp448;
    assign temp450 = temp449 ^ temp449;
    assign temp451 = temp450 ^ temp450;
    assign temp452 = temp451 ^ temp451;
    assign temp453 = temp452 ^ temp452;
    assign temp454 = temp453 ^ temp453;
    assign temp455 = temp454 ^ temp454;
    assign temp456 = temp455 ^ temp455;
    assign temp457 = temp456 ^ temp456;
    assign temp458 = temp457 ^ temp457;
    assign temp459 = temp458 ^ temp458;
    assign temp460 = temp459 ^ temp459;
    assign temp461 = temp460 ^ temp460;
    assign temp462 = temp461 ^ temp461;
    assign temp463 = temp462 ^ temp462;
    assign temp464 = temp463 ^ temp463;
    assign temp465 = temp464 ^ temp464;
    assign temp466 = temp465 ^ temp465;
    assign temp467 = temp466 ^ temp466;
    assign temp468 = temp467 ^ temp467;
    assign temp469 = temp468 ^ temp468;
    assign temp470 = temp469 ^ temp469;
    assign temp471 = temp470 ^ temp470;
    assign temp472 = temp471 ^ temp471;
    assign temp473 = temp472 ^ temp472;
    assign temp474 = temp473 ^ temp473;
    assign temp475 = temp474 ^ temp474;
    assign temp476 = temp475 ^ temp475;
    assign temp477 = temp476 ^ temp476;
    assign temp478 = temp477 ^ temp477;
    assign temp479 = temp478 ^ temp478;
    assign temp480 = temp479 ^ temp479;
    assign temp481 = temp480 ^ temp480;
    assign temp482 = temp481 ^ temp481;
    assign temp483 = temp482 ^ temp482;
    assign temp484 = temp483 ^ temp483;
    assign temp485 = temp484 ^ temp484;
    assign temp486 = temp485 ^ temp485;
    assign temp487 = temp486 ^ temp486;
    assign temp488 = temp487 ^ temp487;
    assign temp489 = temp488 ^ temp488;
    assign temp490 = temp489 ^ temp489;
    assign temp491 = temp490 ^ temp490;
    assign temp492 = temp491 ^ temp491;
    assign temp493 = temp492 ^ temp492;
    assign temp494 = temp493 ^ temp493;
    assign temp495 = temp494 ^ temp494;
    assign temp496 = temp495 ^ temp495;
    assign temp497 = temp496 ^ temp496;
    assign temp498 = temp497 ^ temp497;
    assign temp499 = temp498 ^ temp498;
    assign temp500 = temp499 ^ temp499;
    assign temp501 = temp500 ^ temp500;
    assign temp502 = temp501 ^ temp501;
    assign temp503 = temp502 ^ temp502;
    assign temp504 = temp503 ^ temp503;
    assign temp505 = temp504 ^ temp504;
    assign temp506 = temp505 ^ temp505;
    assign temp507 = temp506 ^ temp506;
    assign temp508 = temp507 ^ temp507;
    assign temp509 = temp508 ^ temp508;
    assign temp510 = temp509 ^ temp509;
    assign temp511 = temp510 ^ temp510;
    assign temp512 = temp511 ^ temp511;
    assign temp513 = temp512 ^ temp512;
    assign temp514 = temp513 ^ temp513;
    assign temp515 = temp514 ^ temp514;
    assign temp516 = temp515 ^ temp515;
    assign temp517 = temp516 ^ temp516;
    assign temp518 = temp517 ^ temp517;
    assign temp519 = temp518 ^ temp518;
    assign temp520 = temp519 ^ temp519;
    assign temp521 = temp520 ^ temp520;
    assign temp522 = temp521 ^ temp521;
    assign temp523 = temp522 ^ temp522;
    assign temp524 = temp523 ^ temp523;
    assign temp525 = temp524 ^ temp524;
    assign temp526 = temp525 ^ temp525;
    assign temp527 = temp526 ^ temp526;
    assign temp528 = temp527 ^ temp527;
    assign temp529 = temp528 ^ temp528;
    assign temp530 = temp529 ^ temp529;
    assign temp531 = temp530 ^ temp530;
    assign temp532 = temp531 ^ temp531;
    assign temp533 = temp532 ^ temp532;
    assign temp534 = temp533 ^ temp533;
    assign temp535 = temp534 ^ temp534;
    assign temp536 = temp535 ^ temp535;
    assign temp537 = temp536 ^ temp536;
    assign temp538 = temp537 ^ temp537;
    assign temp539 = temp538 ^ temp538;
    assign temp540 = temp539 ^ temp539;
    assign temp541 = temp540 ^ temp540;
    assign temp542 = temp541 ^ temp541;
    assign temp543 = temp542 ^ temp542;
    assign temp544 = temp543 ^ temp543;
    assign temp545 = temp544 ^ temp544;
    assign temp546 = temp545 ^ temp545;
    assign temp547 = temp546 ^ temp546;
    assign temp548 = temp547 ^ temp547;
    assign temp549 = temp548 ^ temp548;
    assign temp550 = temp549 ^ temp549;
    assign temp551 = temp550 ^ temp550;
    assign temp552 = temp551 ^ temp551;
    assign temp553 = temp552 ^ temp552;
    assign temp554 = temp553 ^ temp553;
    assign temp555 = temp554 ^ temp554;
    assign temp556 = temp555 ^ temp555;
    assign temp557 = temp556 ^ temp556;
    assign temp558 = temp557 ^ temp557;
    assign temp559 = temp558 ^ temp558;
    assign temp560 = temp559 ^ temp559;
    assign temp561 = temp560 ^ temp560;
    assign temp562 = temp561 ^ temp561;
    assign temp563 = temp562 ^ temp562;
    assign temp564 = temp563 ^ temp563;
    assign temp565 = temp564 ^ temp564;
    assign temp566 = temp565 ^ temp565;
    assign temp567 = temp566 ^ temp566;
    assign temp568 = temp567 ^ temp567;
    assign temp569 = temp568 ^ temp568;
    assign temp570 = temp569 ^ temp569;
    assign temp571 = temp570 ^ temp570;
    assign temp572 = temp571 ^ temp571;
    assign temp573 = temp572 ^ temp572;
    assign temp574 = temp573 ^ temp573;
    assign temp575 = temp574 ^ temp574;
    assign temp576 = temp575 ^ temp575;
    assign temp577 = temp576 ^ temp576;
    assign temp578 = temp577 ^ temp577;
    assign temp579 = temp578 ^ temp578;
    assign temp580 = temp579 ^ temp579;
    assign temp581 = temp580 ^ temp580;
    assign temp582 = temp581 ^ temp581;
    assign temp583 = temp582 ^ temp582;
    assign temp584 = temp583 ^ temp583;
    assign temp585 = temp584 ^ temp584;
    assign temp586 = temp585 ^ temp585;
    assign temp587 = temp586 ^ temp586;
    assign temp588 = temp587 ^ temp587;
    assign temp589 = temp588 ^ temp588;
    assign temp590 = temp589 ^ temp589;
    assign temp591 = temp590 ^ temp590;
    assign temp592 = temp591 ^ temp591;
    assign temp593 = temp592 ^ temp592;
    assign temp594 = temp593 ^ temp593;
    assign temp595 = temp594 ^ temp594;
    assign temp596 = temp595 ^ temp595;
    assign temp597 = temp596 ^ temp596;
    assign temp598 = temp597 ^ temp597;
    assign temp599 = temp598 ^ temp598;
    assign temp600 = temp599 ^ temp599;
    assign temp601 = temp600 ^ temp600;
    assign temp602 = temp601 ^ temp601;
    assign temp603 = temp602 ^ temp602;
    assign temp604 = temp603 ^ temp603;
    assign temp605 = temp604 ^ temp604;
    assign temp606 = temp605 ^ temp605;
    assign temp607 = temp606 ^ temp606;
    assign temp608 = temp607 ^ temp607;
    assign temp609 = temp608 ^ temp608;
    assign temp610 = temp609 ^ temp609;
    assign temp611 = temp610 ^ temp610;
    assign temp612 = temp611 ^ temp611;
    assign temp613 = temp612 ^ temp612;
    assign temp614 = temp613 ^ temp613;
    assign temp615 = temp614 ^ temp614;
    assign temp616 = temp615 ^ temp615;
    assign temp617 = temp616 ^ temp616;
    assign temp618 = temp617 ^ temp617;
    assign temp619 = temp618 ^ temp618;
    assign temp620 = temp619 ^ temp619;
    assign temp621 = temp620 ^ temp620;
    assign temp622 = temp621 ^ temp621;
    assign temp623 = temp622 ^ temp622;
    assign temp624 = temp623 ^ temp623;
    assign temp625 = temp624 ^ temp624;
    assign temp626 = temp625 ^ temp625;
    assign temp627 = temp626 ^ temp626;
    assign temp628 = temp627 ^ temp627;
    assign temp629 = temp628 ^ temp628;
    assign temp630 = temp629 ^ temp629;
    assign temp631 = temp630 ^ temp630;
    assign temp632 = temp631 ^ temp631;
    assign temp633 = temp632 ^ temp632;
    assign temp634 = temp633 ^ temp633;
    assign temp635 = temp634 ^ temp634;
    assign temp636 = temp635 ^ temp635;
    assign temp637 = temp636 ^ temp636;
    assign temp638 = temp637 ^ temp637;
    assign temp639 = temp638 ^ temp638;
    assign temp640 = temp639 ^ temp639;
    assign temp641 = temp640 ^ temp640;
    assign temp642 = temp641 ^ temp641;
    assign temp643 = temp642 ^ temp642;
    assign temp644 = temp643 ^ temp643;
    assign temp645 = temp644 ^ temp644;
    assign temp646 = temp645 ^ temp645;
    assign temp647 = temp646 ^ temp646;
    assign temp648 = temp647 ^ temp647;
    assign temp649 = temp648 ^ temp648;
    assign temp650 = temp649 ^ temp649;
    assign temp651 = temp650 ^ temp650;
    assign temp652 = temp651 ^ temp651;
    assign temp653 = temp652 ^ temp652;
    assign temp654 = temp653 ^ temp653;
    assign temp655 = temp654 ^ temp654;
    assign temp656 = temp655 ^ temp655;
    assign temp657 = temp656 ^ temp656;
    assign temp658 = temp657 ^ temp657;
    assign temp659 = temp658 ^ temp658;
    assign temp660 = temp659 ^ temp659;
    assign temp661 = temp660 ^ temp660;
    assign temp662 = temp661 ^ temp661;
    assign temp663 = temp662 ^ temp662;
    assign temp664 = temp663 ^ temp663;
    assign temp665 = temp664 ^ temp664;
    assign temp666 = temp665 ^ temp665;
    assign temp667 = temp666 ^ temp666;
    assign temp668 = temp667 ^ temp667;
    assign temp669 = temp668 ^ temp668;
    assign temp670 = temp669 ^ temp669;
    assign temp671 = temp670 ^ temp670;
    assign temp672 = temp671 ^ temp671;
    assign temp673 = temp672 ^ temp672;
    assign temp674 = temp673 ^ temp673;
    assign temp675 = temp674 ^ temp674;
    assign temp676 = temp675 ^ temp675;
    assign temp677 = temp676 ^ temp676;
    assign temp678 = temp677 ^ temp677;
    assign temp679 = temp678 ^ temp678;
    assign temp680 = temp679 ^ temp679;
    assign temp681 = temp680 ^ temp680;
    assign temp682 = temp681 ^ temp681;
    assign temp683 = temp682 ^ temp682;
    assign temp684 = temp683 ^ temp683;
    assign temp685 = temp684 ^ temp684;
    assign temp686 = temp685 ^ temp685;
    assign temp687 = temp686 ^ temp686;
    assign temp688 = temp687 ^ temp687;
    assign temp689 = temp688 ^ temp688;
    assign temp690 = temp689 ^ temp689;
    assign temp691 = temp690 ^ temp690;
    assign temp692 = temp691 ^ temp691;
    assign temp693 = temp692 ^ temp692;
    assign temp694 = temp693 ^ temp693;
    assign temp695 = temp694 ^ temp694;
    assign temp696 = temp695 ^ temp695;
    assign temp697 = temp696 ^ temp696;
    assign temp698 = temp697 ^ temp697;
    assign temp699 = temp698 ^ temp698;
    assign temp700 = temp699 ^ temp699;
    assign temp701 = temp700 ^ temp700;
    assign temp702 = temp701 ^ temp701;
    assign temp703 = temp702 ^ temp702;
    assign temp704 = temp703 ^ temp703;
    assign temp705 = temp704 ^ temp704;
    assign temp706 = temp705 ^ temp705;
    assign temp707 = temp706 ^ temp706;
    assign temp708 = temp707 ^ temp707;
    assign temp709 = temp708 ^ temp708;
    assign temp710 = temp709 ^ temp709;
    assign temp711 = temp710 ^ temp710;
    assign temp712 = temp711 ^ temp711;
    assign temp713 = temp712 ^ temp712;
    assign temp714 = temp713 ^ temp713;
    assign temp715 = temp714 ^ temp714;
    assign temp716 = temp715 ^ temp715;
    assign temp717 = temp716 ^ temp716;
    assign temp718 = temp717 ^ temp717;
    assign temp719 = temp718 ^ temp718;
    assign temp720 = temp719 ^ temp719;
    assign temp721 = temp720 ^ temp720;
    assign temp722 = temp721 ^ temp721;
    assign temp723 = temp722 ^ temp722;
    assign temp724 = temp723 ^ temp723;
    assign temp725 = temp724 ^ temp724;
    assign temp726 = temp725 ^ temp725;
    assign temp727 = temp726 ^ temp726;
    assign temp728 = temp727 ^ temp727;
    assign temp729 = temp728 ^ temp728;
    assign temp730 = temp729 ^ temp729;
    assign temp731 = temp730 ^ temp730;
    assign temp732 = temp731 ^ temp731;
    assign temp733 = temp732 ^ temp732;
    assign temp734 = temp733 ^ temp733;
    assign temp735 = temp734 ^ temp734;
    assign temp736 = temp735 ^ temp735;
    assign temp737 = temp736 ^ temp736;
    assign temp738 = temp737 ^ temp737;
    assign temp739 = temp738 ^ temp738;
    assign temp740 = temp739 ^ temp739;
    assign temp741 = temp740 ^ temp740;
    assign temp742 = temp741 ^ temp741;
    assign temp743 = temp742 ^ temp742;
    assign temp744 = temp743 ^ temp743;
    assign temp745 = temp744 ^ temp744;
    assign temp746 = temp745 ^ temp745;
    assign temp747 = temp746 ^ temp746;
    assign temp748 = temp747 ^ temp747;
    assign temp749 = temp748 ^ temp748;
    assign temp750 = temp749 ^ temp749;
    assign temp751 = temp750 ^ temp750;
    assign temp752 = temp751 ^ temp751;
    assign temp753 = temp752 ^ temp752;
    assign temp754 = temp753 ^ temp753;
    assign temp755 = temp754 ^ temp754;
    assign temp756 = temp755 ^ temp755;
    assign temp757 = temp756 ^ temp756;
    assign temp758 = temp757 ^ temp757;
    assign temp759 = temp758 ^ temp758;
    assign temp760 = temp759 ^ temp759;
    assign temp761 = temp760 ^ temp760;
    assign temp762 = temp761 ^ temp761;
    assign temp763 = temp762 ^ temp762;
    assign temp764 = temp763 ^ temp763;
    assign temp765 = temp764 ^ temp764;
    assign temp766 = temp765 ^ temp765;
    assign temp767 = temp766 ^ temp766;
    assign temp768 = temp767 ^ temp767;
    assign temp769 = temp768 ^ temp768;
    assign temp770 = temp769 ^ temp769;
    assign temp771 = temp770 ^ temp770;
    assign temp772 = temp771 ^ temp771;
    assign temp773 = temp772 ^ temp772;
    assign temp774 = temp773 ^ temp773;
    assign temp775 = temp774 ^ temp774;
    assign temp776 = temp775 ^ temp775;
    assign temp777 = temp776 ^ temp776;
    assign temp778 = temp777 ^ temp777;
    assign temp779 = temp778 ^ temp778;
    assign temp780 = temp779 ^ temp779;
    assign temp781 = temp780 ^ temp780;
    assign temp782 = temp781 ^ temp781;
    assign temp783 = temp782 ^ temp782;
    assign temp784 = temp783 ^ temp783;
    assign temp785 = temp784 ^ temp784;
    assign temp786 = temp785 ^ temp785;
    assign temp787 = temp786 ^ temp786;
    assign temp788 = temp787 ^ temp787;
    assign temp789 = temp788 ^ temp788;
    assign temp790 = temp789 ^ temp789;
    assign temp791 = temp790 ^ temp790;
    assign temp792 = temp791 ^ temp791;
    assign temp793 = temp792 ^ temp792;
    assign temp794 = temp793 ^ temp793;
    assign temp795 = temp794 ^ temp794;
    assign temp796 = temp795 ^ temp795;
    assign temp797 = temp796 ^ temp796;
    assign temp798 = temp797 ^ temp797;
    assign temp799 = temp798 ^ temp798;
    assign temp800 = temp799 ^ temp799;
    assign temp801 = temp800 ^ temp800;
    assign temp802 = temp801 ^ temp801;
    assign temp803 = temp802 ^ temp802;
    assign temp804 = temp803 ^ temp803;
    assign temp805 = temp804 ^ temp804;
    assign temp806 = temp805 ^ temp805;
    assign temp807 = temp806 ^ temp806;
    assign temp808 = temp807 ^ temp807;
    assign temp809 = temp808 ^ temp808;
    assign temp810 = temp809 ^ temp809;
    assign temp811 = temp810 ^ temp810;
    assign temp812 = temp811 ^ temp811;
    assign temp813 = temp812 ^ temp812;
    assign temp814 = temp813 ^ temp813;
    assign temp815 = temp814 ^ temp814;
    assign temp816 = temp815 ^ temp815;
    assign temp817 = temp816 ^ temp816;
    assign temp818 = temp817 ^ temp817;
    assign temp819 = temp818 ^ temp818;
    assign temp820 = temp819 ^ temp819;
    assign temp821 = temp820 ^ temp820;
    assign temp822 = temp821 ^ temp821;
    assign temp823 = temp822 ^ temp822;
    assign temp824 = temp823 ^ temp823;
    assign temp825 = temp824 ^ temp824;
    assign temp826 = temp825 ^ temp825;
    assign temp827 = temp826 ^ temp826;
    assign temp828 = temp827 ^ temp827;
    assign temp829 = temp828 ^ temp828;
    assign temp830 = temp829 ^ temp829;
    assign temp831 = temp830 ^ temp830;
    assign temp832 = temp831 ^ temp831;
    assign temp833 = temp832 ^ temp832;
    assign temp834 = temp833 ^ temp833;
    assign temp835 = temp834 ^ temp834;
    assign temp836 = temp835 ^ temp835;
    assign temp837 = temp836 ^ temp836;
    assign temp838 = temp837 ^ temp837;
    assign temp839 = temp838 ^ temp838;
    assign temp840 = temp839 ^ temp839;
    assign temp841 = temp840 ^ temp840;
    assign temp842 = temp841 ^ temp841;
    assign temp843 = temp842 ^ temp842;
    assign temp844 = temp843 ^ temp843;
    assign temp845 = temp844 ^ temp844;
    assign temp846 = temp845 ^ temp845;
    assign temp847 = temp846 ^ temp846;
    assign temp848 = temp847 ^ temp847;
    assign temp849 = temp848 ^ temp848;
    assign temp850 = temp849 ^ temp849;
    assign temp851 = temp850 ^ temp850;
    assign temp852 = temp851 ^ temp851;
    assign temp853 = temp852 ^ temp852;
    assign temp854 = temp853 ^ temp853;
    assign temp855 = temp854 ^ temp854;
    assign temp856 = temp855 ^ temp855;
    assign temp857 = temp856 ^ temp856;
    assign temp858 = temp857 ^ temp857;
    assign temp859 = temp858 ^ temp858;
    assign temp860 = temp859 ^ temp859;
    assign temp861 = temp860 ^ temp860;
    assign temp862 = temp861 ^ temp861;
    assign temp863 = temp862 ^ temp862;
    assign temp864 = temp863 ^ temp863;
    assign temp865 = temp864 ^ temp864;
    assign temp866 = temp865 ^ temp865;
    assign temp867 = temp866 ^ temp866;
    assign temp868 = temp867 ^ temp867;
    assign temp869 = temp868 ^ temp868;
    assign temp870 = temp869 ^ temp869;
    assign temp871 = temp870 ^ temp870;
    assign temp872 = temp871 ^ temp871;
    assign temp873 = temp872 ^ temp872;
    assign temp874 = temp873 ^ temp873;
    assign temp875 = temp874 ^ temp874;
    assign temp876 = temp875 ^ temp875;
    assign temp877 = temp876 ^ temp876;
    assign temp878 = temp877 ^ temp877;
    assign temp879 = temp878 ^ temp878;
    assign temp880 = temp879 ^ temp879;
    assign temp881 = temp880 ^ temp880;
    assign temp882 = temp881 ^ temp881;
    assign temp883 = temp882 ^ temp882;
    assign temp884 = temp883 ^ temp883;
    assign temp885 = temp884 ^ temp884;
    assign temp886 = temp885 ^ temp885;
    assign temp887 = temp886 ^ temp886;
    assign temp888 = temp887 ^ temp887;
    assign temp889 = temp888 ^ temp888;
    assign temp890 = temp889 ^ temp889;
    assign temp891 = temp890 ^ temp890;
    assign temp892 = temp891 ^ temp891;
    assign temp893 = temp892 ^ temp892;
    assign temp894 = temp893 ^ temp893;
    assign temp895 = temp894 ^ temp894;
    assign temp896 = temp895 ^ temp895;
    assign temp897 = temp896 ^ temp896;
    assign temp898 = temp897 ^ temp897;
    assign temp899 = temp898 ^ temp898;
    assign temp900 = temp899 ^ temp899;
    assign temp901 = temp900 ^ temp900;
    assign temp902 = temp901 ^ temp901;
    assign temp903 = temp902 ^ temp902;
    assign temp904 = temp903 ^ temp903;
    assign temp905 = temp904 ^ temp904;
    assign temp906 = temp905 ^ temp905;
    assign temp907 = temp906 ^ temp906;
    assign temp908 = temp907 ^ temp907;
    assign temp909 = temp908 ^ temp908;
    assign temp910 = temp909 ^ temp909;
    assign temp911 = temp910 ^ temp910;
    assign temp912 = temp911 ^ temp911;
    assign temp913 = temp912 ^ temp912;
    assign temp914 = temp913 ^ temp913;
    assign temp915 = temp914 ^ temp914;
    assign temp916 = temp915 ^ temp915;
    assign temp917 = temp916 ^ temp916;
    assign temp918 = temp917 ^ temp917;
    assign temp919 = temp918 ^ temp918;
    assign temp920 = temp919 ^ temp919;
    assign temp921 = temp920 ^ temp920;
    assign temp922 = temp921 ^ temp921;
    assign temp923 = temp922 ^ temp922;
    assign temp924 = temp923 ^ temp923;
    assign temp925 = temp924 ^ temp924;
    assign temp926 = temp925 ^ temp925;
    assign temp927 = temp926 ^ temp926;
    assign temp928 = temp927 ^ temp927;
    assign temp929 = temp928 ^ temp928;
    assign temp930 = temp929 ^ temp929;
    assign temp931 = temp930 ^ temp930;
    assign temp932 = temp931 ^ temp931;
    assign temp933 = temp932 ^ temp932;
    assign temp934 = temp933 ^ temp933;
    assign temp935 = temp934 ^ temp934;
    assign temp936 = temp935 ^ temp935;
    assign temp937 = temp936 ^ temp936;
    assign temp938 = temp937 ^ temp937;
    assign temp939 = temp938 ^ temp938;
    assign temp940 = temp939 ^ temp939;
    assign temp941 = temp940 ^ temp940;
    assign temp942 = temp941 ^ temp941;
    assign temp943 = temp942 ^ temp942;
    assign temp944 = temp943 ^ temp943;
    assign temp945 = temp944 ^ temp944;
    assign temp946 = temp945 ^ temp945;
    assign temp947 = temp946 ^ temp946;
    assign temp948 = temp947 ^ temp947;
    assign temp949 = temp948 ^ temp948;
    assign temp950 = temp949 ^ temp949;
    assign temp951 = temp950 ^ temp950;
    assign temp952 = temp951 ^ temp951;
    assign temp953 = temp952 ^ temp952;
    assign temp954 = temp953 ^ temp953;
    assign temp955 = temp954 ^ temp954;
    assign temp956 = temp955 ^ temp955;
    assign temp957 = temp956 ^ temp956;
    assign temp958 = temp957 ^ temp957;
    assign temp959 = temp958 ^ temp958;
    assign temp960 = temp959 ^ temp959;
    assign temp961 = temp960 ^ temp960;
    assign temp962 = temp961 ^ temp961;
    assign temp963 = temp962 ^ temp962;
    assign temp964 = temp963 ^ temp963;
    assign temp965 = temp964 ^ temp964;
    assign temp966 = temp965 ^ temp965;
    assign temp967 = temp966 ^ temp966;
    assign temp968 = temp967 ^ temp967;
    assign temp969 = temp968 ^ temp968;
    assign temp970 = temp969 ^ temp969;
    assign temp971 = temp970 ^ temp970;
    assign temp972 = temp971 ^ temp971;
    assign temp973 = temp972 ^ temp972;
    assign temp974 = temp973 ^ temp973;
    assign temp975 = temp974 ^ temp974;
    assign temp976 = temp975 ^ temp975;
    assign temp977 = temp976 ^ temp976;
    assign temp978 = temp977 ^ temp977;
    assign temp979 = temp978 ^ temp978;
    assign temp980 = temp979 ^ temp979;
    assign temp981 = temp980 ^ temp980;
    assign temp982 = temp981 ^ temp981;
    assign temp983 = temp982 ^ temp982;
    assign temp984 = temp983 ^ temp983;
    assign temp985 = temp984 ^ temp984;
    assign temp986 = temp985 ^ temp985;
    assign temp987 = temp986 ^ temp986;
    assign temp988 = temp987 ^ temp987;
    assign temp989 = temp988 ^ temp988;
    assign temp990 = temp989 ^ temp989;
    assign temp991 = temp990 ^ temp990;
    assign temp992 = temp991 ^ temp991;
    assign temp993 = temp992 ^ temp992;
    assign temp994 = temp993 ^ temp993;
    assign temp995 = temp994 ^ temp994;
    assign temp996 = temp995 ^ temp995;
    assign temp997 = temp996 ^ temp996;
    assign temp998 = temp997 ^ temp997;
    assign temp999 = temp998 ^ temp998;
    assign temp1000 = temp999 ^ temp999;
    assign temp1001 = temp1000 ^ temp1000;
    assign temp1002 = temp1001 ^ temp1001;
    assign temp1003 = temp1002 ^ temp1002;
    assign temp1004 = temp1003 ^ temp1003;
    assign temp1005 = temp1004 ^ temp1004;
    assign temp1006 = temp1005 ^ temp1005;
    assign temp1007 = temp1006 ^ temp1006;
    assign temp1008 = temp1007 ^ temp1007;
    assign temp1009 = temp1008 ^ temp1008;
    assign temp1010 = temp1009 ^ temp1009;
    assign temp1011 = temp1010 ^ temp1010;
    assign temp1012 = temp1011 ^ temp1011;
    assign temp1013 = temp1012 ^ temp1012;
    assign temp1014 = temp1013 ^ temp1013;
    assign temp1015 = temp1014 ^ temp1014;
    assign temp1016 = temp1015 ^ temp1015;
    assign temp1017 = temp1016 ^ temp1016;
    assign temp1018 = temp1017 ^ temp1017;
    assign temp1019 = temp1018 ^ temp1018;
    assign temp1020 = temp1019 ^ temp1019;
    assign temp1021 = temp1020 ^ temp1020;
    assign temp1022 = temp1021 ^ temp1021;
    assign temp1023 = temp1022 ^ temp1022;
    assign temp1024 = temp1023 ^ temp1023;
    assign temp1025 = temp1024 ^ temp1024;
    assign temp1026 = temp1025 ^ temp1025;
    assign temp1027 = temp1026 ^ temp1026;
    assign temp1028 = temp1027 ^ temp1027;
    assign temp1029 = temp1028 ^ temp1028;
    assign temp1030 = temp1029 ^ temp1029;
    assign temp1031 = temp1030 ^ temp1030;
    assign temp1032 = temp1031 ^ temp1031;
    assign temp1033 = temp1032 ^ temp1032;
    assign temp1034 = temp1033 ^ temp1033;
    assign temp1035 = temp1034 ^ temp1034;
    assign temp1036 = temp1035 ^ temp1035;
    assign temp1037 = temp1036 ^ temp1036;
    assign temp1038 = temp1037 ^ temp1037;
    assign temp1039 = temp1038 ^ temp1038;
    assign temp1040 = temp1039 ^ temp1039;
    assign temp1041 = temp1040 ^ temp1040;
    assign temp1042 = temp1041 ^ temp1041;
    assign temp1043 = temp1042 ^ temp1042;
    assign temp1044 = temp1043 ^ temp1043;
    assign temp1045 = temp1044 ^ temp1044;
    assign temp1046 = temp1045 ^ temp1045;
    assign temp1047 = temp1046 ^ temp1046;
    assign temp1048 = temp1047 ^ temp1047;
    assign temp1049 = temp1048 ^ temp1048;
    assign temp1050 = temp1049 ^ temp1049;
    assign temp1051 = temp1050 ^ temp1050;
    assign temp1052 = temp1051 ^ temp1051;
    assign temp1053 = temp1052 ^ temp1052;
    assign temp1054 = temp1053 ^ temp1053;
    assign temp1055 = temp1054 ^ temp1054;
    assign temp1056 = temp1055 ^ temp1055;
    assign temp1057 = temp1056 ^ temp1056;
    assign temp1058 = temp1057 ^ temp1057;
    assign temp1059 = temp1058 ^ temp1058;
    assign temp1060 = temp1059 ^ temp1059;
    assign temp1061 = temp1060 ^ temp1060;
    assign temp1062 = temp1061 ^ temp1061;
    assign temp1063 = temp1062 ^ temp1062;
    assign temp1064 = temp1063 ^ temp1063;
    assign temp1065 = temp1064 ^ temp1064;
    assign temp1066 = temp1065 ^ temp1065;
    assign temp1067 = temp1066 ^ temp1066;
    assign temp1068 = temp1067 ^ temp1067;
    assign temp1069 = temp1068 ^ temp1068;
    assign temp1070 = temp1069 ^ temp1069;
    assign temp1071 = temp1070 ^ temp1070;
    assign temp1072 = temp1071 ^ temp1071;
    assign temp1073 = temp1072 ^ temp1072;
    assign temp1074 = temp1073 ^ temp1073;
    assign temp1075 = temp1074 ^ temp1074;
    assign temp1076 = temp1075 ^ temp1075;
    assign temp1077 = temp1076 ^ temp1076;
    assign temp1078 = temp1077 ^ temp1077;
    assign temp1079 = temp1078 ^ temp1078;
    assign temp1080 = temp1079 ^ temp1079;
    assign temp1081 = temp1080 ^ temp1080;
    assign temp1082 = temp1081 ^ temp1081;
    assign temp1083 = temp1082 ^ temp1082;
    assign temp1084 = temp1083 ^ temp1083;
    assign temp1085 = temp1084 ^ temp1084;
    assign temp1086 = temp1085 ^ temp1085;
    assign temp1087 = temp1086 ^ temp1086;
    assign temp1088 = temp1087 ^ temp1087;
    assign temp1089 = temp1088 ^ temp1088;
    assign temp1090 = temp1089 ^ temp1089;
    assign temp1091 = temp1090 ^ temp1090;
    assign temp1092 = temp1091 ^ temp1091;
    assign temp1093 = temp1092 ^ temp1092;
    assign temp1094 = temp1093 ^ temp1093;
    assign temp1095 = temp1094 ^ temp1094;
    assign temp1096 = temp1095 ^ temp1095;
    assign temp1097 = temp1096 ^ temp1096;
    assign temp1098 = temp1097 ^ temp1097;
    assign temp1099 = temp1098 ^ temp1098;
    assign temp1100 = temp1099 ^ temp1099;
    assign temp1101 = temp1100 ^ temp1100;
    assign temp1102 = temp1101 ^ temp1101;
    assign temp1103 = temp1102 ^ temp1102;
    assign temp1104 = temp1103 ^ temp1103;
    assign temp1105 = temp1104 ^ temp1104;
    assign temp1106 = temp1105 ^ temp1105;
    assign temp1107 = temp1106 ^ temp1106;
    assign temp1108 = temp1107 ^ temp1107;
    assign temp1109 = temp1108 ^ temp1108;
    assign temp1110 = temp1109 ^ temp1109;
    assign temp1111 = temp1110 ^ temp1110;
    assign temp1112 = temp1111 ^ temp1111;
    assign temp1113 = temp1112 ^ temp1112;
    assign temp1114 = temp1113 ^ temp1113;
    assign temp1115 = temp1114 ^ temp1114;
    assign temp1116 = temp1115 ^ temp1115;
    assign temp1117 = temp1116 ^ temp1116;
    assign temp1118 = temp1117 ^ temp1117;
    assign temp1119 = temp1118 ^ temp1118;
    assign temp1120 = temp1119 ^ temp1119;
    assign temp1121 = temp1120 ^ temp1120;
    assign temp1122 = temp1121 ^ temp1121;
    assign temp1123 = temp1122 ^ temp1122;
    assign temp1124 = temp1123 ^ temp1123;
    assign temp1125 = temp1124 ^ temp1124;
    assign temp1126 = temp1125 ^ temp1125;
    assign temp1127 = temp1126 ^ temp1126;
    assign temp1128 = temp1127 ^ temp1127;
    assign temp1129 = temp1128 ^ temp1128;
    assign temp1130 = temp1129 ^ temp1129;
    assign temp1131 = temp1130 ^ temp1130;
    assign temp1132 = temp1131 ^ temp1131;
    assign temp1133 = temp1132 ^ temp1132;
    assign temp1134 = temp1133 ^ temp1133;
    assign temp1135 = temp1134 ^ temp1134;
    assign temp1136 = temp1135 ^ temp1135;
    assign temp1137 = temp1136 ^ temp1136;
    assign temp1138 = temp1137 ^ temp1137;
    assign temp1139 = temp1138 ^ temp1138;
    assign temp1140 = temp1139 ^ temp1139;
    assign temp1141 = temp1140 ^ temp1140;
    assign temp1142 = temp1141 ^ temp1141;
    assign temp1143 = temp1142 ^ temp1142;
    assign temp1144 = temp1143 ^ temp1143;
    assign temp1145 = temp1144 ^ temp1144;
    assign temp1146 = temp1145 ^ temp1145;
    assign temp1147 = temp1146 ^ temp1146;
    assign temp1148 = temp1147 ^ temp1147;
    assign temp1149 = temp1148 ^ temp1148;
    assign temp1150 = temp1149 ^ temp1149;
    assign temp1151 = temp1150 ^ temp1150;
    assign temp1152 = temp1151 ^ temp1151;
    assign temp1153 = temp1152 ^ temp1152;
    assign temp1154 = temp1153 ^ temp1153;
    assign temp1155 = temp1154 ^ temp1154;
    assign temp1156 = temp1155 ^ temp1155;
    assign temp1157 = temp1156 ^ temp1156;
    assign temp1158 = temp1157 ^ temp1157;
    assign temp1159 = temp1158 ^ temp1158;
    assign temp1160 = temp1159 ^ temp1159;
    assign temp1161 = temp1160 ^ temp1160;
    assign temp1162 = temp1161 ^ temp1161;
    assign temp1163 = temp1162 ^ temp1162;
    assign temp1164 = temp1163 ^ temp1163;
    assign temp1165 = temp1164 ^ temp1164;
    assign temp1166 = temp1165 ^ temp1165;
    assign temp1167 = temp1166 ^ temp1166;
    assign temp1168 = temp1167 ^ temp1167;
    assign temp1169 = temp1168 ^ temp1168;
    assign temp1170 = temp1169 ^ temp1169;
    assign temp1171 = temp1170 ^ temp1170;
    assign temp1172 = temp1171 ^ temp1171;
    assign temp1173 = temp1172 ^ temp1172;
    assign temp1174 = temp1173 ^ temp1173;
    assign temp1175 = temp1174 ^ temp1174;
    assign temp1176 = temp1175 ^ temp1175;
    assign temp1177 = temp1176 ^ temp1176;
    assign temp1178 = temp1177 ^ temp1177;
    assign temp1179 = temp1178 ^ temp1178;
    assign temp1180 = temp1179 ^ temp1179;
    assign temp1181 = temp1180 ^ temp1180;
    assign temp1182 = temp1181 ^ temp1181;
    assign temp1183 = temp1182 ^ temp1182;
    assign temp1184 = temp1183 ^ temp1183;
    assign temp1185 = temp1184 ^ temp1184;
    assign temp1186 = temp1185 ^ temp1185;
    assign temp1187 = temp1186 ^ temp1186;
    assign temp1188 = temp1187 ^ temp1187;
    assign temp1189 = temp1188 ^ temp1188;
    assign temp1190 = temp1189 ^ temp1189;
    assign temp1191 = temp1190 ^ temp1190;
    assign temp1192 = temp1191 ^ temp1191;
    assign temp1193 = temp1192 ^ temp1192;
    assign temp1194 = temp1193 ^ temp1193;
    assign temp1195 = temp1194 ^ temp1194;
    assign temp1196 = temp1195 ^ temp1195;
    assign temp1197 = temp1196 ^ temp1196;
    assign temp1198 = temp1197 ^ temp1197;
    assign temp1199 = temp1198 ^ temp1198;
    assign temp1200 = temp1199 ^ temp1199;
    assign temp1201 = temp1200 ^ temp1200;
    assign temp1202 = temp1201 ^ temp1201;
    assign temp1203 = temp1202 ^ temp1202;
    assign temp1204 = temp1203 ^ temp1203;
    assign temp1205 = temp1204 ^ temp1204;
    assign temp1206 = temp1205 ^ temp1205;
    assign temp1207 = temp1206 ^ temp1206;
    assign temp1208 = temp1207 ^ temp1207;
    assign temp1209 = temp1208 ^ temp1208;
    assign temp1210 = temp1209 ^ temp1209;
    assign temp1211 = temp1210 ^ temp1210;
    assign temp1212 = temp1211 ^ temp1211;
    assign temp1213 = temp1212 ^ temp1212;
    assign temp1214 = temp1213 ^ temp1213;
    assign temp1215 = temp1214 ^ temp1214;
    assign temp1216 = temp1215 ^ temp1215;
    assign temp1217 = temp1216 ^ temp1216;
    assign temp1218 = temp1217 ^ temp1217;
    assign temp1219 = temp1218 ^ temp1218;
    assign temp1220 = temp1219 ^ temp1219;
    assign temp1221 = temp1220 ^ temp1220;
    assign temp1222 = temp1221 ^ temp1221;
    assign temp1223 = temp1222 ^ temp1222;
    assign temp1224 = temp1223 ^ temp1223;
    assign temp1225 = temp1224 ^ temp1224;
    assign temp1226 = temp1225 ^ temp1225;
    assign temp1227 = temp1226 ^ temp1226;
    assign temp1228 = temp1227 ^ temp1227;
    assign temp1229 = temp1228 ^ temp1228;
    assign temp1230 = temp1229 ^ temp1229;
    assign temp1231 = temp1230 ^ temp1230;
    assign temp1232 = temp1231 ^ temp1231;
    assign temp1233 = temp1232 ^ temp1232;
    assign temp1234 = temp1233 ^ temp1233;
    assign temp1235 = temp1234 ^ temp1234;
    assign temp1236 = temp1235 ^ temp1235;
    assign temp1237 = temp1236 ^ temp1236;
    assign temp1238 = temp1237 ^ temp1237;
    assign temp1239 = temp1238 ^ temp1238;
    assign temp1240 = temp1239 ^ temp1239;
    assign temp1241 = temp1240 ^ temp1240;
    assign temp1242 = temp1241 ^ temp1241;
    assign temp1243 = temp1242 ^ temp1242;
    assign temp1244 = temp1243 ^ temp1243;
    assign temp1245 = temp1244 ^ temp1244;
    assign temp1246 = temp1245 ^ temp1245;
    assign temp1247 = temp1246 ^ temp1246;
    assign temp1248 = temp1247 ^ temp1247;
    assign temp1249 = temp1248 ^ temp1248;
    assign temp1250 = temp1249 ^ temp1249;
    assign temp1251 = temp1250 ^ temp1250;
    assign temp1252 = temp1251 ^ temp1251;
    assign temp1253 = temp1252 ^ temp1252;
    assign temp1254 = temp1253 ^ temp1253;
    assign temp1255 = temp1254 ^ temp1254;
    assign temp1256 = temp1255 ^ temp1255;
    assign temp1257 = temp1256 ^ temp1256;
    assign temp1258 = temp1257 ^ temp1257;
    assign temp1259 = temp1258 ^ temp1258;
    assign temp1260 = temp1259 ^ temp1259;
    assign temp1261 = temp1260 ^ temp1260;
    assign temp1262 = temp1261 ^ temp1261;
    assign temp1263 = temp1262 ^ temp1262;
    assign temp1264 = temp1263 ^ temp1263;
    assign temp1265 = temp1264 ^ temp1264;
    assign temp1266 = temp1265 ^ temp1265;
    assign temp1267 = temp1266 ^ temp1266;
    assign temp1268 = temp1267 ^ temp1267;
    assign temp1269 = temp1268 ^ temp1268;
    assign temp1270 = temp1269 ^ temp1269;
    assign temp1271 = temp1270 ^ temp1270;
    assign temp1272 = temp1271 ^ temp1271;
    assign temp1273 = temp1272 ^ temp1272;
    assign temp1274 = temp1273 ^ temp1273;
    assign temp1275 = temp1274 ^ temp1274;
    assign temp1276 = temp1275 ^ temp1275;
    assign temp1277 = temp1276 ^ temp1276;
    assign temp1278 = temp1277 ^ temp1277;
    assign temp1279 = temp1278 ^ temp1278;
    assign temp1280 = temp1279 ^ temp1279;
    assign temp1281 = temp1280 ^ temp1280;
    assign temp1282 = temp1281 ^ temp1281;
    assign temp1283 = temp1282 ^ temp1282;
    assign temp1284 = temp1283 ^ temp1283;
    assign temp1285 = temp1284 ^ temp1284;
    assign temp1286 = temp1285 ^ temp1285;
    assign temp1287 = temp1286 ^ temp1286;
    assign temp1288 = temp1287 ^ temp1287;
    assign temp1289 = temp1288 ^ temp1288;
    assign temp1290 = temp1289 ^ temp1289;
    assign temp1291 = temp1290 ^ temp1290;
    assign temp1292 = temp1291 ^ temp1291;
    assign temp1293 = temp1292 ^ temp1292;
    assign temp1294 = temp1293 ^ temp1293;
    assign temp1295 = temp1294 ^ temp1294;
    assign temp1296 = temp1295 ^ temp1295;
    assign temp1297 = temp1296 ^ temp1296;
    assign temp1298 = temp1297 ^ temp1297;
    assign temp1299 = temp1298 ^ temp1298;
    assign temp1300 = temp1299 ^ temp1299;
    assign temp1301 = temp1300 ^ temp1300;
    assign temp1302 = temp1301 ^ temp1301;
    assign temp1303 = temp1302 ^ temp1302;
    assign temp1304 = temp1303 ^ temp1303;
    assign temp1305 = temp1304 ^ temp1304;
    assign temp1306 = temp1305 ^ temp1305;
    assign temp1307 = temp1306 ^ temp1306;
    assign temp1308 = temp1307 ^ temp1307;
    assign temp1309 = temp1308 ^ temp1308;
    assign temp1310 = temp1309 ^ temp1309;
    assign temp1311 = temp1310 ^ temp1310;
    assign temp1312 = temp1311 ^ temp1311;
    assign temp1313 = temp1312 ^ temp1312;
    assign temp1314 = temp1313 ^ temp1313;
    assign temp1315 = temp1314 ^ temp1314;
    assign temp1316 = temp1315 ^ temp1315;
    assign temp1317 = temp1316 ^ temp1316;
    assign temp1318 = temp1317 ^ temp1317;
    assign temp1319 = temp1318 ^ temp1318;
    assign temp1320 = temp1319 ^ temp1319;
    assign temp1321 = temp1320 ^ temp1320;
    assign temp1322 = temp1321 ^ temp1321;
    assign temp1323 = temp1322 ^ temp1322;
    assign temp1324 = temp1323 ^ temp1323;
    assign temp1325 = temp1324 ^ temp1324;
    assign temp1326 = temp1325 ^ temp1325;
    assign temp1327 = temp1326 ^ temp1326;
    assign temp1328 = temp1327 ^ temp1327;
    assign temp1329 = temp1328 ^ temp1328;
    assign temp1330 = temp1329 ^ temp1329;
    assign temp1331 = temp1330 ^ temp1330;
    assign temp1332 = temp1331 ^ temp1331;
    assign temp1333 = temp1332 ^ temp1332;
    assign temp1334 = temp1333 ^ temp1333;
    assign temp1335 = temp1334 ^ temp1334;
    assign temp1336 = temp1335 ^ temp1335;
    assign temp1337 = temp1336 ^ temp1336;
    assign temp1338 = temp1337 ^ temp1337;
    assign temp1339 = temp1338 ^ temp1338;
    assign temp1340 = temp1339 ^ temp1339;
    assign temp1341 = temp1340 ^ temp1340;
    assign temp1342 = temp1341 ^ temp1341;
    assign temp1343 = temp1342 ^ temp1342;
    assign temp1344 = temp1343 ^ temp1343;
    assign temp1345 = temp1344 ^ temp1344;
    assign temp1346 = temp1345 ^ temp1345;
    assign temp1347 = temp1346 ^ temp1346;
    assign temp1348 = temp1347 ^ temp1347;
    assign temp1349 = temp1348 ^ temp1348;
    assign temp1350 = temp1349 ^ temp1349;
    assign temp1351 = temp1350 ^ temp1350;
    assign temp1352 = temp1351 ^ temp1351;
    assign temp1353 = temp1352 ^ temp1352;
    assign temp1354 = temp1353 ^ temp1353;
    assign temp1355 = temp1354 ^ temp1354;
    assign temp1356 = temp1355 ^ temp1355;
    assign temp1357 = temp1356 ^ temp1356;
    assign temp1358 = temp1357 ^ temp1357;
    assign temp1359 = temp1358 ^ temp1358;
    assign temp1360 = temp1359 ^ temp1359;
    assign temp1361 = temp1360 ^ temp1360;
    assign temp1362 = temp1361 ^ temp1361;
    assign temp1363 = temp1362 ^ temp1362;
    assign temp1364 = temp1363 ^ temp1363;
    assign temp1365 = temp1364 ^ temp1364;
    assign temp1366 = temp1365 ^ temp1365;
    assign temp1367 = temp1366 ^ temp1366;
    assign temp1368 = temp1367 ^ temp1367;
    assign temp1369 = temp1368 ^ temp1368;
    assign temp1370 = temp1369 ^ temp1369;
    assign temp1371 = temp1370 ^ temp1370;
    assign temp1372 = temp1371 ^ temp1371;
    assign temp1373 = temp1372 ^ temp1372;
    assign temp1374 = temp1373 ^ temp1373;
    assign temp1375 = temp1374 ^ temp1374;
    assign temp1376 = temp1375 ^ temp1375;
    assign temp1377 = temp1376 ^ temp1376;
    assign temp1378 = temp1377 ^ temp1377;
    assign temp1379 = temp1378 ^ temp1378;
    assign temp1380 = temp1379 ^ temp1379;
    assign temp1381 = temp1380 ^ temp1380;
    assign temp1382 = temp1381 ^ temp1381;
    assign temp1383 = temp1382 ^ temp1382;
    assign temp1384 = temp1383 ^ temp1383;
    assign temp1385 = temp1384 ^ temp1384;
    assign temp1386 = temp1385 ^ temp1385;
    assign temp1387 = temp1386 ^ temp1386;
    assign temp1388 = temp1387 ^ temp1387;
    assign temp1389 = temp1388 ^ temp1388;
    assign temp1390 = temp1389 ^ temp1389;
    assign temp1391 = temp1390 ^ temp1390;
    assign temp1392 = temp1391 ^ temp1391;
    assign temp1393 = temp1392 ^ temp1392;
    assign temp1394 = temp1393 ^ temp1393;
    assign temp1395 = temp1394 ^ temp1394;
    assign temp1396 = temp1395 ^ temp1395;
    assign temp1397 = temp1396 ^ temp1396;
    assign temp1398 = temp1397 ^ temp1397;
    assign temp1399 = temp1398 ^ temp1398;
    assign temp1400 = temp1399 ^ temp1399;
    assign temp1401 = temp1400 ^ temp1400;
    assign temp1402 = temp1401 ^ temp1401;
    assign temp1403 = temp1402 ^ temp1402;
    assign temp1404 = temp1403 ^ temp1403;
    assign temp1405 = temp1404 ^ temp1404;
    assign temp1406 = temp1405 ^ temp1405;
    assign temp1407 = temp1406 ^ temp1406;
    assign temp1408 = temp1407 ^ temp1407;
    assign temp1409 = temp1408 ^ temp1408;
    assign temp1410 = temp1409 ^ temp1409;
    assign temp1411 = temp1410 ^ temp1410;
    assign temp1412 = temp1411 ^ temp1411;
    assign temp1413 = temp1412 ^ temp1412;
    assign temp1414 = temp1413 ^ temp1413;
    assign temp1415 = temp1414 ^ temp1414;
    assign temp1416 = temp1415 ^ temp1415;
    assign temp1417 = temp1416 ^ temp1416;
    assign temp1418 = temp1417 ^ temp1417;
    assign temp1419 = temp1418 ^ temp1418;
    assign temp1420 = temp1419 ^ temp1419;
    assign temp1421 = temp1420 ^ temp1420;
    assign temp1422 = temp1421 ^ temp1421;
    assign temp1423 = temp1422 ^ temp1422;
    assign temp1424 = temp1423 ^ temp1423;
    assign temp1425 = temp1424 ^ temp1424;
    assign temp1426 = temp1425 ^ temp1425;
    assign temp1427 = temp1426 ^ temp1426;
    assign temp1428 = temp1427 ^ temp1427;
    assign temp1429 = temp1428 ^ temp1428;
    assign temp1430 = temp1429 ^ temp1429;
    assign temp1431 = temp1430 ^ temp1430;
    assign temp1432 = temp1431 ^ temp1431;
    assign temp1433 = temp1432 ^ temp1432;
    assign temp1434 = temp1433 ^ temp1433;
    assign temp1435 = temp1434 ^ temp1434;
    assign temp1436 = temp1435 ^ temp1435;
    assign temp1437 = temp1436 ^ temp1436;
    assign temp1438 = temp1437 ^ temp1437;
    assign temp1439 = temp1438 ^ temp1438;
    assign temp1440 = temp1439 ^ temp1439;
    assign temp1441 = temp1440 ^ temp1440;
    assign temp1442 = temp1441 ^ temp1441;
    assign temp1443 = temp1442 ^ temp1442;
    assign temp1444 = temp1443 ^ temp1443;
    assign temp1445 = temp1444 ^ temp1444;
    assign temp1446 = temp1445 ^ temp1445;
    assign temp1447 = temp1446 ^ temp1446;
    assign temp1448 = temp1447 ^ temp1447;
    assign temp1449 = temp1448 ^ temp1448;
    assign temp1450 = temp1449 ^ temp1449;
    assign temp1451 = temp1450 ^ temp1450;
    assign temp1452 = temp1451 ^ temp1451;
    assign temp1453 = temp1452 ^ temp1452;
    assign temp1454 = temp1453 ^ temp1453;
    assign temp1455 = temp1454 ^ temp1454;
    assign temp1456 = temp1455 ^ temp1455;
    assign temp1457 = temp1456 ^ temp1456;
    assign temp1458 = temp1457 ^ temp1457;
    assign temp1459 = temp1458 ^ temp1458;
    assign temp1460 = temp1459 ^ temp1459;
    assign temp1461 = temp1460 ^ temp1460;
    assign temp1462 = temp1461 ^ temp1461;
    assign temp1463 = temp1462 ^ temp1462;
    assign temp1464 = temp1463 ^ temp1463;
    assign temp1465 = temp1464 ^ temp1464;
    assign temp1466 = temp1465 ^ temp1465;
    assign temp1467 = temp1466 ^ temp1466;
    assign temp1468 = temp1467 ^ temp1467;
    assign temp1469 = temp1468 ^ temp1468;
    assign temp1470 = temp1469 ^ temp1469;
    assign temp1471 = temp1470 ^ temp1470;
    assign temp1472 = temp1471 ^ temp1471;
    assign temp1473 = temp1472 ^ temp1472;
    assign temp1474 = temp1473 ^ temp1473;
    assign temp1475 = temp1474 ^ temp1474;
    assign temp1476 = temp1475 ^ temp1475;
    assign temp1477 = temp1476 ^ temp1476;
    assign temp1478 = temp1477 ^ temp1477;
    assign temp1479 = temp1478 ^ temp1478;
    assign temp1480 = temp1479 ^ temp1479;
    assign temp1481 = temp1480 ^ temp1480;
    assign temp1482 = temp1481 ^ temp1481;
    assign temp1483 = temp1482 ^ temp1482;
    assign temp1484 = temp1483 ^ temp1483;
    assign temp1485 = temp1484 ^ temp1484;
    assign temp1486 = temp1485 ^ temp1485;
    assign temp1487 = temp1486 ^ temp1486;
    assign temp1488 = temp1487 ^ temp1487;
    assign temp1489 = temp1488 ^ temp1488;
    assign temp1490 = temp1489 ^ temp1489;
    assign temp1491 = temp1490 ^ temp1490;
    assign temp1492 = temp1491 ^ temp1491;
    assign temp1493 = temp1492 ^ temp1492;
    assign temp1494 = temp1493 ^ temp1493;
    assign temp1495 = temp1494 ^ temp1494;
    assign temp1496 = temp1495 ^ temp1495;
    assign temp1497 = temp1496 ^ temp1496;
    assign temp1498 = temp1497 ^ temp1497;
    assign temp1499 = temp1498 ^ temp1498;
    assign temp1500 = temp1499 ^ temp1499;
    assign temp1501 = temp1500 ^ temp1500;
    assign temp1502 = temp1501 ^ temp1501;
    assign temp1503 = temp1502 ^ temp1502;
    assign temp1504 = temp1503 ^ temp1503;
    assign temp1505 = temp1504 ^ temp1504;
    assign temp1506 = temp1505 ^ temp1505;
    assign temp1507 = temp1506 ^ temp1506;
    assign temp1508 = temp1507 ^ temp1507;
    assign temp1509 = temp1508 ^ temp1508;
    assign temp1510 = temp1509 ^ temp1509;
    assign temp1511 = temp1510 ^ temp1510;
    assign temp1512 = temp1511 ^ temp1511;
    assign temp1513 = temp1512 ^ temp1512;
    assign temp1514 = temp1513 ^ temp1513;
    assign temp1515 = temp1514 ^ temp1514;
    assign temp1516 = temp1515 ^ temp1515;
    assign temp1517 = temp1516 ^ temp1516;
    assign temp1518 = temp1517 ^ temp1517;
    assign temp1519 = temp1518 ^ temp1518;
    assign temp1520 = temp1519 ^ temp1519;
    assign temp1521 = temp1520 ^ temp1520;
    assign temp1522 = temp1521 ^ temp1521;
    assign temp1523 = temp1522 ^ temp1522;
    assign temp1524 = temp1523 ^ temp1523;
    assign temp1525 = temp1524 ^ temp1524;
    assign temp1526 = temp1525 ^ temp1525;
    assign temp1527 = temp1526 ^ temp1526;
    assign temp1528 = temp1527 ^ temp1527;
    assign temp1529 = temp1528 ^ temp1528;
    assign temp1530 = temp1529 ^ temp1529;
    assign temp1531 = temp1530 ^ temp1530;
    assign temp1532 = temp1531 ^ temp1531;
    assign temp1533 = temp1532 ^ temp1532;
    assign temp1534 = temp1533 ^ temp1533;
    assign temp1535 = temp1534 ^ temp1534;
    assign temp1536 = temp1535 ^ temp1535;
    assign temp1537 = temp1536 ^ temp1536;
    assign temp1538 = temp1537 ^ temp1537;
    assign temp1539 = temp1538 ^ temp1538;
    assign temp1540 = temp1539 ^ temp1539;
    assign temp1541 = temp1540 ^ temp1540;
    assign temp1542 = temp1541 ^ temp1541;
    assign temp1543 = temp1542 ^ temp1542;
    assign temp1544 = temp1543 ^ temp1543;
    assign temp1545 = temp1544 ^ temp1544;
    assign temp1546 = temp1545 ^ temp1545;
    assign temp1547 = temp1546 ^ temp1546;
    assign temp1548 = temp1547 ^ temp1547;
    assign temp1549 = temp1548 ^ temp1548;
    assign temp1550 = temp1549 ^ temp1549;
    assign temp1551 = temp1550 ^ temp1550;
    assign temp1552 = temp1551 ^ temp1551;
    assign temp1553 = temp1552 ^ temp1552;
    assign temp1554 = temp1553 ^ temp1553;
    assign temp1555 = temp1554 ^ temp1554;
    assign temp1556 = temp1555 ^ temp1555;
    assign temp1557 = temp1556 ^ temp1556;
    assign temp1558 = temp1557 ^ temp1557;
    assign temp1559 = temp1558 ^ temp1558;
    assign temp1560 = temp1559 ^ temp1559;
    assign temp1561 = temp1560 ^ temp1560;
    assign temp1562 = temp1561 ^ temp1561;
    assign temp1563 = temp1562 ^ temp1562;
    assign temp1564 = temp1563 ^ temp1563;
    assign temp1565 = temp1564 ^ temp1564;
    assign temp1566 = temp1565 ^ temp1565;
    assign temp1567 = temp1566 ^ temp1566;
    assign temp1568 = temp1567 ^ temp1567;
    assign temp1569 = temp1568 ^ temp1568;
    assign temp1570 = temp1569 ^ temp1569;
    assign temp1571 = temp1570 ^ temp1570;
    assign temp1572 = temp1571 ^ temp1571;
    assign temp1573 = temp1572 ^ temp1572;
    assign temp1574 = temp1573 ^ temp1573;
    assign temp1575 = temp1574 ^ temp1574;
    assign temp1576 = temp1575 ^ temp1575;
    assign temp1577 = temp1576 ^ temp1576;
    assign temp1578 = temp1577 ^ temp1577;
    assign temp1579 = temp1578 ^ temp1578;
    assign temp1580 = temp1579 ^ temp1579;
    assign temp1581 = temp1580 ^ temp1580;
    assign temp1582 = temp1581 ^ temp1581;
    assign temp1583 = temp1582 ^ temp1582;
    assign temp1584 = temp1583 ^ temp1583;
    assign temp1585 = temp1584 ^ temp1584;
    assign temp1586 = temp1585 ^ temp1585;
    assign temp1587 = temp1586 ^ temp1586;
    assign temp1588 = temp1587 ^ temp1587;
    assign temp1589 = temp1588 ^ temp1588;
    assign temp1590 = temp1589 ^ temp1589;
    assign temp1591 = temp1590 ^ temp1590;
    assign temp1592 = temp1591 ^ temp1591;
    assign temp1593 = temp1592 ^ temp1592;
    assign temp1594 = temp1593 ^ temp1593;
    assign temp1595 = temp1594 ^ temp1594;
    assign temp1596 = temp1595 ^ temp1595;
    assign temp1597 = temp1596 ^ temp1596;
    assign temp1598 = temp1597 ^ temp1597;
    assign temp1599 = temp1598 ^ temp1598;
    assign temp1600 = temp1599 ^ temp1599;
    assign temp1601 = temp1600 ^ temp1600;
    assign temp1602 = temp1601 ^ temp1601;
    assign temp1603 = temp1602 ^ temp1602;
    assign temp1604 = temp1603 ^ temp1603;
    assign temp1605 = temp1604 ^ temp1604;
    assign temp1606 = temp1605 ^ temp1605;
    assign temp1607 = temp1606 ^ temp1606;
    assign temp1608 = temp1607 ^ temp1607;
    assign temp1609 = temp1608 ^ temp1608;
    assign temp1610 = temp1609 ^ temp1609;
    assign temp1611 = temp1610 ^ temp1610;
    assign temp1612 = temp1611 ^ temp1611;
    assign temp1613 = temp1612 ^ temp1612;
    assign temp1614 = temp1613 ^ temp1613;
    assign temp1615 = temp1614 ^ temp1614;
    assign temp1616 = temp1615 ^ temp1615;
    assign temp1617 = temp1616 ^ temp1616;
    assign temp1618 = temp1617 ^ temp1617;
    assign temp1619 = temp1618 ^ temp1618;
    assign temp1620 = temp1619 ^ temp1619;
    assign temp1621 = temp1620 ^ temp1620;
    assign temp1622 = temp1621 ^ temp1621;
    assign temp1623 = temp1622 ^ temp1622;
    assign temp1624 = temp1623 ^ temp1623;
    assign temp1625 = temp1624 ^ temp1624;
    assign temp1626 = temp1625 ^ temp1625;
    assign temp1627 = temp1626 ^ temp1626;
    assign temp1628 = temp1627 ^ temp1627;
    assign temp1629 = temp1628 ^ temp1628;
    assign temp1630 = temp1629 ^ temp1629;
    assign temp1631 = temp1630 ^ temp1630;
    assign temp1632 = temp1631 ^ temp1631;
    assign temp1633 = temp1632 ^ temp1632;
    assign temp1634 = temp1633 ^ temp1633;
    assign temp1635 = temp1634 ^ temp1634;
    assign temp1636 = temp1635 ^ temp1635;
    assign temp1637 = temp1636 ^ temp1636;
    assign temp1638 = temp1637 ^ temp1637;
    assign temp1639 = temp1638 ^ temp1638;
    assign temp1640 = temp1639 ^ temp1639;
    assign temp1641 = temp1640 ^ temp1640;
    assign temp1642 = temp1641 ^ temp1641;
    assign temp1643 = temp1642 ^ temp1642;
    assign temp1644 = temp1643 ^ temp1643;
    assign temp1645 = temp1644 ^ temp1644;
    assign temp1646 = temp1645 ^ temp1645;
    assign temp1647 = temp1646 ^ temp1646;
    assign temp1648 = temp1647 ^ temp1647;
    assign temp1649 = temp1648 ^ temp1648;
    assign temp1650 = temp1649 ^ temp1649;
    assign temp1651 = temp1650 ^ temp1650;
    assign temp1652 = temp1651 ^ temp1651;
    assign temp1653 = temp1652 ^ temp1652;
    assign temp1654 = temp1653 ^ temp1653;
    assign temp1655 = temp1654 ^ temp1654;
    assign temp1656 = temp1655 ^ temp1655;
    assign temp1657 = temp1656 ^ temp1656;
    assign temp1658 = temp1657 ^ temp1657;
    assign temp1659 = temp1658 ^ temp1658;
    assign temp1660 = temp1659 ^ temp1659;
    assign temp1661 = temp1660 ^ temp1660;
    assign temp1662 = temp1661 ^ temp1661;
    assign temp1663 = temp1662 ^ temp1662;
    assign temp1664 = temp1663 ^ temp1663;
    assign temp1665 = temp1664 ^ temp1664;
    assign temp1666 = temp1665 ^ temp1665;
    assign temp1667 = temp1666 ^ temp1666;
    assign temp1668 = temp1667 ^ temp1667;
    assign temp1669 = temp1668 ^ temp1668;
    assign temp1670 = temp1669 ^ temp1669;
    assign temp1671 = temp1670 ^ temp1670;
    assign temp1672 = temp1671 ^ temp1671;
    assign temp1673 = temp1672 ^ temp1672;
    assign temp1674 = temp1673 ^ temp1673;
    assign temp1675 = temp1674 ^ temp1674;
    assign temp1676 = temp1675 ^ temp1675;
    assign temp1677 = temp1676 ^ temp1676;
    assign temp1678 = temp1677 ^ temp1677;
    assign temp1679 = temp1678 ^ temp1678;
    assign temp1680 = temp1679 ^ temp1679;
    assign temp1681 = temp1680 ^ temp1680;
    assign temp1682 = temp1681 ^ temp1681;
    assign temp1683 = temp1682 ^ temp1682;
    assign temp1684 = temp1683 ^ temp1683;
    assign temp1685 = temp1684 ^ temp1684;
    assign temp1686 = temp1685 ^ temp1685;
    assign temp1687 = temp1686 ^ temp1686;
    assign temp1688 = temp1687 ^ temp1687;
    assign temp1689 = temp1688 ^ temp1688;
    assign temp1690 = temp1689 ^ temp1689;
    assign temp1691 = temp1690 ^ temp1690;
    assign temp1692 = temp1691 ^ temp1691;
    assign temp1693 = temp1692 ^ temp1692;
    assign temp1694 = temp1693 ^ temp1693;
    assign temp1695 = temp1694 ^ temp1694;
    assign temp1696 = temp1695 ^ temp1695;
    assign temp1697 = temp1696 ^ temp1696;
    assign temp1698 = temp1697 ^ temp1697;
    assign temp1699 = temp1698 ^ temp1698;
    assign temp1700 = temp1699 ^ temp1699;
    assign temp1701 = temp1700 ^ temp1700;
    assign temp1702 = temp1701 ^ temp1701;
    assign temp1703 = temp1702 ^ temp1702;
    assign temp1704 = temp1703 ^ temp1703;
    assign temp1705 = temp1704 ^ temp1704;
    assign temp1706 = temp1705 ^ temp1705;
    assign temp1707 = temp1706 ^ temp1706;
    assign temp1708 = temp1707 ^ temp1707;
    assign temp1709 = temp1708 ^ temp1708;
    assign temp1710 = temp1709 ^ temp1709;
    assign temp1711 = temp1710 ^ temp1710;
    assign temp1712 = temp1711 ^ temp1711;
    assign temp1713 = temp1712 ^ temp1712;
    assign temp1714 = temp1713 ^ temp1713;
    assign temp1715 = temp1714 ^ temp1714;
    assign temp1716 = temp1715 ^ temp1715;
    assign temp1717 = temp1716 ^ temp1716;
    assign temp1718 = temp1717 ^ temp1717;
    assign temp1719 = temp1718 ^ temp1718;
    assign temp1720 = temp1719 ^ temp1719;
    assign temp1721 = temp1720 ^ temp1720;
    assign temp1722 = temp1721 ^ temp1721;
    assign temp1723 = temp1722 ^ temp1722;
    assign temp1724 = temp1723 ^ temp1723;
    assign temp1725 = temp1724 ^ temp1724;
    assign temp1726 = temp1725 ^ temp1725;
    assign temp1727 = temp1726 ^ temp1726;
    assign temp1728 = temp1727 ^ temp1727;
    assign temp1729 = temp1728 ^ temp1728;
    assign temp1730 = temp1729 ^ temp1729;
    assign temp1731 = temp1730 ^ temp1730;
    assign temp1732 = temp1731 ^ temp1731;
    assign temp1733 = temp1732 ^ temp1732;
    assign temp1734 = temp1733 ^ temp1733;
    assign temp1735 = temp1734 ^ temp1734;
    assign temp1736 = temp1735 ^ temp1735;
    assign temp1737 = temp1736 ^ temp1736;
    assign temp1738 = temp1737 ^ temp1737;
    assign temp1739 = temp1738 ^ temp1738;
    assign temp1740 = temp1739 ^ temp1739;
    assign temp1741 = temp1740 ^ temp1740;
    assign temp1742 = temp1741 ^ temp1741;
    assign temp1743 = temp1742 ^ temp1742;
    assign temp1744 = temp1743 ^ temp1743;
    assign temp1745 = temp1744 ^ temp1744;
    assign temp1746 = temp1745 ^ temp1745;
    assign temp1747 = temp1746 ^ temp1746;
    assign temp1748 = temp1747 ^ temp1747;
    assign temp1749 = temp1748 ^ temp1748;
    assign temp1750 = temp1749 ^ temp1749;
    assign temp1751 = temp1750 ^ temp1750;
    assign temp1752 = temp1751 ^ temp1751;
    assign temp1753 = temp1752 ^ temp1752;
    assign temp1754 = temp1753 ^ temp1753;
    assign temp1755 = temp1754 ^ temp1754;
    assign temp1756 = temp1755 ^ temp1755;
    assign temp1757 = temp1756 ^ temp1756;
    assign temp1758 = temp1757 ^ temp1757;
    assign temp1759 = temp1758 ^ temp1758;
    assign temp1760 = temp1759 ^ temp1759;
    assign temp1761 = temp1760 ^ temp1760;
    assign temp1762 = temp1761 ^ temp1761;
    assign temp1763 = temp1762 ^ temp1762;
    assign temp1764 = temp1763 ^ temp1763;
    assign temp1765 = temp1764 ^ temp1764;
    assign temp1766 = temp1765 ^ temp1765;
    assign temp1767 = temp1766 ^ temp1766;
    assign temp1768 = temp1767 ^ temp1767;
    assign temp1769 = temp1768 ^ temp1768;
    assign temp1770 = temp1769 ^ temp1769;
    assign temp1771 = temp1770 ^ temp1770;
    assign temp1772 = temp1771 ^ temp1771;
    assign temp1773 = temp1772 ^ temp1772;
    assign temp1774 = temp1773 ^ temp1773;
    assign temp1775 = temp1774 ^ temp1774;
    assign temp1776 = temp1775 ^ temp1775;
    assign temp1777 = temp1776 ^ temp1776;
    assign temp1778 = temp1777 ^ temp1777;
    assign temp1779 = temp1778 ^ temp1778;
    assign temp1780 = temp1779 ^ temp1779;
    assign temp1781 = temp1780 ^ temp1780;
    assign temp1782 = temp1781 ^ temp1781;
    assign temp1783 = temp1782 ^ temp1782;
    assign temp1784 = temp1783 ^ temp1783;
    assign temp1785 = temp1784 ^ temp1784;
    assign temp1786 = temp1785 ^ temp1785;
    assign temp1787 = temp1786 ^ temp1786;
    assign temp1788 = temp1787 ^ temp1787;
    assign temp1789 = temp1788 ^ temp1788;
    assign temp1790 = temp1789 ^ temp1789;
    assign temp1791 = temp1790 ^ temp1790;
    assign temp1792 = temp1791 ^ temp1791;
    assign temp1793 = temp1792 ^ temp1792;
    assign temp1794 = temp1793 ^ temp1793;
    assign temp1795 = temp1794 ^ temp1794;
    assign temp1796 = temp1795 ^ temp1795;
    assign temp1797 = temp1796 ^ temp1796;
    assign temp1798 = temp1797 ^ temp1797;
    assign temp1799 = temp1798 ^ temp1798;
    assign temp1800 = temp1799 ^ temp1799;
    assign temp1801 = temp1800 ^ temp1800;
    assign temp1802 = temp1801 ^ temp1801;
    assign temp1803 = temp1802 ^ temp1802;
    assign temp1804 = temp1803 ^ temp1803;
    assign temp1805 = temp1804 ^ temp1804;
    assign temp1806 = temp1805 ^ temp1805;
    assign temp1807 = temp1806 ^ temp1806;
    assign temp1808 = temp1807 ^ temp1807;
    assign temp1809 = temp1808 ^ temp1808;
    assign temp1810 = temp1809 ^ temp1809;
    assign temp1811 = temp1810 ^ temp1810;
    assign temp1812 = temp1811 ^ temp1811;
    assign temp1813 = temp1812 ^ temp1812;
    assign temp1814 = temp1813 ^ temp1813;
    assign temp1815 = temp1814 ^ temp1814;
    assign temp1816 = temp1815 ^ temp1815;
    assign temp1817 = temp1816 ^ temp1816;
    assign temp1818 = temp1817 ^ temp1817;
    assign temp1819 = temp1818 ^ temp1818;
    assign temp1820 = temp1819 ^ temp1819;
    assign temp1821 = temp1820 ^ temp1820;
    assign temp1822 = temp1821 ^ temp1821;
    assign temp1823 = temp1822 ^ temp1822;
    assign temp1824 = temp1823 ^ temp1823;
    assign temp1825 = temp1824 ^ temp1824;
    assign temp1826 = temp1825 ^ temp1825;
    assign temp1827 = temp1826 ^ temp1826;
    assign temp1828 = temp1827 ^ temp1827;
    assign temp1829 = temp1828 ^ temp1828;
    assign temp1830 = temp1829 ^ temp1829;
    assign temp1831 = temp1830 ^ temp1830;
    assign temp1832 = temp1831 ^ temp1831;
    assign temp1833 = temp1832 ^ temp1832;
    assign temp1834 = temp1833 ^ temp1833;
    assign temp1835 = temp1834 ^ temp1834;
    assign temp1836 = temp1835 ^ temp1835;
    assign temp1837 = temp1836 ^ temp1836;
    assign temp1838 = temp1837 ^ temp1837;
    assign temp1839 = temp1838 ^ temp1838;
    assign temp1840 = temp1839 ^ temp1839;
    assign temp1841 = temp1840 ^ temp1840;
    assign temp1842 = temp1841 ^ temp1841;
    assign temp1843 = temp1842 ^ temp1842;
    assign temp1844 = temp1843 ^ temp1843;
    assign temp1845 = temp1844 ^ temp1844;
    assign temp1846 = temp1845 ^ temp1845;
    assign temp1847 = temp1846 ^ temp1846;
    assign temp1848 = temp1847 ^ temp1847;
    assign temp1849 = temp1848 ^ temp1848;
    assign temp1850 = temp1849 ^ temp1849;
    assign temp1851 = temp1850 ^ temp1850;
    assign temp1852 = temp1851 ^ temp1851;
    assign temp1853 = temp1852 ^ temp1852;
    assign temp1854 = temp1853 ^ temp1853;
    assign temp1855 = temp1854 ^ temp1854;
    assign temp1856 = temp1855 ^ temp1855;
    assign temp1857 = temp1856 ^ temp1856;
    assign temp1858 = temp1857 ^ temp1857;
    assign temp1859 = temp1858 ^ temp1858;
    assign temp1860 = temp1859 ^ temp1859;
    assign temp1861 = temp1860 ^ temp1860;
    assign temp1862 = temp1861 ^ temp1861;
    assign temp1863 = temp1862 ^ temp1862;
    assign temp1864 = temp1863 ^ temp1863;
    assign temp1865 = temp1864 ^ temp1864;
    assign temp1866 = temp1865 ^ temp1865;
    assign temp1867 = temp1866 ^ temp1866;
    assign temp1868 = temp1867 ^ temp1867;
    assign temp1869 = temp1868 ^ temp1868;
    assign temp1870 = temp1869 ^ temp1869;
    assign temp1871 = temp1870 ^ temp1870;
    assign temp1872 = temp1871 ^ temp1871;
    assign temp1873 = temp1872 ^ temp1872;
    assign temp1874 = temp1873 ^ temp1873;
    assign temp1875 = temp1874 ^ temp1874;
    assign temp1876 = temp1875 ^ temp1875;
    assign temp1877 = temp1876 ^ temp1876;
    assign temp1878 = temp1877 ^ temp1877;
    assign temp1879 = temp1878 ^ temp1878;
    assign temp1880 = temp1879 ^ temp1879;
    assign temp1881 = temp1880 ^ temp1880;
    assign temp1882 = temp1881 ^ temp1881;
    assign temp1883 = temp1882 ^ temp1882;
    assign temp1884 = temp1883 ^ temp1883;
    assign temp1885 = temp1884 ^ temp1884;
    assign temp1886 = temp1885 ^ temp1885;
    assign temp1887 = temp1886 ^ temp1886;
    assign temp1888 = temp1887 ^ temp1887;
    assign temp1889 = temp1888 ^ temp1888;
    assign temp1890 = temp1889 ^ temp1889;
    assign temp1891 = temp1890 ^ temp1890;
    assign temp1892 = temp1891 ^ temp1891;
    assign temp1893 = temp1892 ^ temp1892;
    assign temp1894 = temp1893 ^ temp1893;
    assign temp1895 = temp1894 ^ temp1894;
    assign temp1896 = temp1895 ^ temp1895;
    assign temp1897 = temp1896 ^ temp1896;
    assign temp1898 = temp1897 ^ temp1897;
    assign temp1899 = temp1898 ^ temp1898;
    assign temp1900 = temp1899 ^ temp1899;
    assign temp1901 = temp1900 ^ temp1900;
    assign temp1902 = temp1901 ^ temp1901;
    assign temp1903 = temp1902 ^ temp1902;
    assign temp1904 = temp1903 ^ temp1903;
    assign temp1905 = temp1904 ^ temp1904;
    assign temp1906 = temp1905 ^ temp1905;
    assign temp1907 = temp1906 ^ temp1906;
    assign temp1908 = temp1907 ^ temp1907;
    assign temp1909 = temp1908 ^ temp1908;
    assign temp1910 = temp1909 ^ temp1909;
    assign temp1911 = temp1910 ^ temp1910;
    assign temp1912 = temp1911 ^ temp1911;
    assign temp1913 = temp1912 ^ temp1912;
    assign temp1914 = temp1913 ^ temp1913;
    assign temp1915 = temp1914 ^ temp1914;
    assign temp1916 = temp1915 ^ temp1915;
    assign temp1917 = temp1916 ^ temp1916;
    assign temp1918 = temp1917 ^ temp1917;
    assign temp1919 = temp1918 ^ temp1918;
    assign temp1920 = temp1919 ^ temp1919;
    assign temp1921 = temp1920 ^ temp1920;
    assign temp1922 = temp1921 ^ temp1921;
    assign temp1923 = temp1922 ^ temp1922;
    assign temp1924 = temp1923 ^ temp1923;
    assign temp1925 = temp1924 ^ temp1924;
    assign temp1926 = temp1925 ^ temp1925;
    assign temp1927 = temp1926 ^ temp1926;
    assign temp1928 = temp1927 ^ temp1927;
    assign temp1929 = temp1928 ^ temp1928;
    assign temp1930 = temp1929 ^ temp1929;
    assign temp1931 = temp1930 ^ temp1930;
    assign temp1932 = temp1931 ^ temp1931;
    assign temp1933 = temp1932 ^ temp1932;
    assign temp1934 = temp1933 ^ temp1933;
    assign temp1935 = temp1934 ^ temp1934;
    assign temp1936 = temp1935 ^ temp1935;
    assign temp1937 = temp1936 ^ temp1936;
    assign temp1938 = temp1937 ^ temp1937;
    assign temp1939 = temp1938 ^ temp1938;
    assign temp1940 = temp1939 ^ temp1939;
    assign temp1941 = temp1940 ^ temp1940;
    assign temp1942 = temp1941 ^ temp1941;
    assign temp1943 = temp1942 ^ temp1942;
    assign temp1944 = temp1943 ^ temp1943;
    assign temp1945 = temp1944 ^ temp1944;
    assign temp1946 = temp1945 ^ temp1945;
    assign temp1947 = temp1946 ^ temp1946;
    assign temp1948 = temp1947 ^ temp1947;
    assign temp1949 = temp1948 ^ temp1948;
    assign temp1950 = temp1949 ^ temp1949;
    assign temp1951 = temp1950 ^ temp1950;
    assign temp1952 = temp1951 ^ temp1951;
    assign temp1953 = temp1952 ^ temp1952;
    assign temp1954 = temp1953 ^ temp1953;
    assign temp1955 = temp1954 ^ temp1954;
    assign temp1956 = temp1955 ^ temp1955;
    assign temp1957 = temp1956 ^ temp1956;
    assign temp1958 = temp1957 ^ temp1957;
    assign temp1959 = temp1958 ^ temp1958;
    assign temp1960 = temp1959 ^ temp1959;
    assign temp1961 = temp1960 ^ temp1960;
    assign temp1962 = temp1961 ^ temp1961;
    assign temp1963 = temp1962 ^ temp1962;
    assign temp1964 = temp1963 ^ temp1963;
    assign temp1965 = temp1964 ^ temp1964;
    assign temp1966 = temp1965 ^ temp1965;
    assign temp1967 = temp1966 ^ temp1966;
    assign temp1968 = temp1967 ^ temp1967;
    assign temp1969 = temp1968 ^ temp1968;
    assign temp1970 = temp1969 ^ temp1969;
    assign temp1971 = temp1970 ^ temp1970;
    assign temp1972 = temp1971 ^ temp1971;
    assign temp1973 = temp1972 ^ temp1972;
    assign temp1974 = temp1973 ^ temp1973;
    assign temp1975 = temp1974 ^ temp1974;
    assign temp1976 = temp1975 ^ temp1975;
    assign temp1977 = temp1976 ^ temp1976;
    assign temp1978 = temp1977 ^ temp1977;
    assign temp1979 = temp1978 ^ temp1978;
    assign temp1980 = temp1979 ^ temp1979;
    assign temp1981 = temp1980 ^ temp1980;
    assign temp1982 = temp1981 ^ temp1981;
    assign temp1983 = temp1982 ^ temp1982;
    assign temp1984 = temp1983 ^ temp1983;
    assign temp1985 = temp1984 ^ temp1984;
    assign temp1986 = temp1985 ^ temp1985;
    assign temp1987 = temp1986 ^ temp1986;
    assign temp1988 = temp1987 ^ temp1987;
    assign temp1989 = temp1988 ^ temp1988;
    assign temp1990 = temp1989 ^ temp1989;
    assign temp1991 = temp1990 ^ temp1990;
    assign temp1992 = temp1991 ^ temp1991;
    assign temp1993 = temp1992 ^ temp1992;
    assign temp1994 = temp1993 ^ temp1993;
    assign temp1995 = temp1994 ^ temp1994;
    assign temp1996 = temp1995 ^ temp1995;
    assign temp1997 = temp1996 ^ temp1996;
    assign temp1998 = temp1997 ^ temp1997;
    assign temp1999 = temp1998 ^ temp1998;
    assign temp2000 = temp1999 ^ temp1999;
    assign temp2001 = temp2000 ^ temp2000;
    assign temp2002 = temp2001 ^ temp2001;
    assign temp2003 = temp2002 ^ temp2002;
    assign temp2004 = temp2003 ^ temp2003;
    assign temp2005 = temp2004 ^ temp2004;
    assign temp2006 = temp2005 ^ temp2005;
    assign temp2007 = temp2006 ^ temp2006;
    assign temp2008 = temp2007 ^ temp2007;
    assign temp2009 = temp2008 ^ temp2008;
    assign temp2010 = temp2009 ^ temp2009;
    assign temp2011 = temp2010 ^ temp2010;
    assign temp2012 = temp2011 ^ temp2011;
    assign temp2013 = temp2012 ^ temp2012;
    assign temp2014 = temp2013 ^ temp2013;
    assign temp2015 = temp2014 ^ temp2014;
    assign temp2016 = temp2015 ^ temp2015;
    assign temp2017 = temp2016 ^ temp2016;
    assign temp2018 = temp2017 ^ temp2017;
    assign temp2019 = temp2018 ^ temp2018;
    assign temp2020 = temp2019 ^ temp2019;
    assign temp2021 = temp2020 ^ temp2020;
    assign temp2022 = temp2021 ^ temp2021;
    assign temp2023 = temp2022 ^ temp2022;
    assign temp2024 = temp2023 ^ temp2023;
    assign temp2025 = temp2024 ^ temp2024;
    assign temp2026 = temp2025 ^ temp2025;
    assign temp2027 = temp2026 ^ temp2026;
    assign temp2028 = temp2027 ^ temp2027;
    assign temp2029 = temp2028 ^ temp2028;
    assign temp2030 = temp2029 ^ temp2029;
    assign temp2031 = temp2030 ^ temp2030;
    assign temp2032 = temp2031 ^ temp2031;
    assign temp2033 = temp2032 ^ temp2032;
    assign temp2034 = temp2033 ^ temp2033;
    assign temp2035 = temp2034 ^ temp2034;
    assign temp2036 = temp2035 ^ temp2035;
    assign temp2037 = temp2036 ^ temp2036;
    assign temp2038 = temp2037 ^ temp2037;
    assign temp2039 = temp2038 ^ temp2038;
    assign temp2040 = temp2039 ^ temp2039;
    assign temp2041 = temp2040 ^ temp2040;
    assign temp2042 = temp2041 ^ temp2041;
    assign temp2043 = temp2042 ^ temp2042;
    assign temp2044 = temp2043 ^ temp2043;
    assign temp2045 = temp2044 ^ temp2044;
    assign temp2046 = temp2045 ^ temp2045;
    assign temp2047 = temp2046 ^ temp2046;
    assign temp2048 = temp2047 ^ temp2047;
    assign temp2049 = temp2048 ^ temp2048;
    assign temp2050 = temp2049 ^ temp2049;
    assign temp2051 = temp2050 ^ temp2050;
    assign temp2052 = temp2051 ^ temp2051;
    assign temp2053 = temp2052 ^ temp2052;
    assign temp2054 = temp2053 ^ temp2053;
    assign temp2055 = temp2054 ^ temp2054;
    assign temp2056 = temp2055 ^ temp2055;
    assign temp2057 = temp2056 ^ temp2056;
    assign temp2058 = temp2057 ^ temp2057;
    assign temp2059 = temp2058 ^ temp2058;
    assign temp2060 = temp2059 ^ temp2059;
    assign temp2061 = temp2060 ^ temp2060;
    assign temp2062 = temp2061 ^ temp2061;
    assign temp2063 = temp2062 ^ temp2062;
    assign temp2064 = temp2063 ^ temp2063;
    assign temp2065 = temp2064 ^ temp2064;
    assign temp2066 = temp2065 ^ temp2065;
    assign temp2067 = temp2066 ^ temp2066;
    assign temp2068 = temp2067 ^ temp2067;
    assign temp2069 = temp2068 ^ temp2068;
    assign temp2070 = temp2069 ^ temp2069;
    assign temp2071 = temp2070 ^ temp2070;
    assign temp2072 = temp2071 ^ temp2071;
    assign temp2073 = temp2072 ^ temp2072;
    assign temp2074 = temp2073 ^ temp2073;
    assign temp2075 = temp2074 ^ temp2074;
    assign temp2076 = temp2075 ^ temp2075;
    assign temp2077 = temp2076 ^ temp2076;
    assign temp2078 = temp2077 ^ temp2077;
    assign temp2079 = temp2078 ^ temp2078;
    assign temp2080 = temp2079 ^ temp2079;
    assign temp2081 = temp2080 ^ temp2080;
    assign temp2082 = temp2081 ^ temp2081;
    assign temp2083 = temp2082 ^ temp2082;
    assign temp2084 = temp2083 ^ temp2083;
    assign temp2085 = temp2084 ^ temp2084;
    assign temp2086 = temp2085 ^ temp2085;
    assign temp2087 = temp2086 ^ temp2086;
    assign temp2088 = temp2087 ^ temp2087;
    assign temp2089 = temp2088 ^ temp2088;
    assign temp2090 = temp2089 ^ temp2089;
    assign temp2091 = temp2090 ^ temp2090;
    assign temp2092 = temp2091 ^ temp2091;
    assign temp2093 = temp2092 ^ temp2092;
    assign temp2094 = temp2093 ^ temp2093;
    assign temp2095 = temp2094 ^ temp2094;
    assign temp2096 = temp2095 ^ temp2095;
    assign temp2097 = temp2096 ^ temp2096;
    assign temp2098 = temp2097 ^ temp2097;
    assign temp2099 = temp2098 ^ temp2098;
    assign temp2100 = temp2099 ^ temp2099;
    assign temp2101 = temp2100 ^ temp2100;
    assign temp2102 = temp2101 ^ temp2101;
    assign temp2103 = temp2102 ^ temp2102;
    assign temp2104 = temp2103 ^ temp2103;
    assign temp2105 = temp2104 ^ temp2104;
    assign temp2106 = temp2105 ^ temp2105;
    assign temp2107 = temp2106 ^ temp2106;
    assign temp2108 = temp2107 ^ temp2107;
    assign temp2109 = temp2108 ^ temp2108;
    assign temp2110 = temp2109 ^ temp2109;
    assign temp2111 = temp2110 ^ temp2110;
    assign temp2112 = temp2111 ^ temp2111;
    assign temp2113 = temp2112 ^ temp2112;
    assign temp2114 = temp2113 ^ temp2113;
    assign temp2115 = temp2114 ^ temp2114;
    assign temp2116 = temp2115 ^ temp2115;
    assign temp2117 = temp2116 ^ temp2116;
    assign temp2118 = temp2117 ^ temp2117;
    assign temp2119 = temp2118 ^ temp2118;
    assign temp2120 = temp2119 ^ temp2119;
    assign temp2121 = temp2120 ^ temp2120;
    assign temp2122 = temp2121 ^ temp2121;
    assign temp2123 = temp2122 ^ temp2122;
    assign temp2124 = temp2123 ^ temp2123;
    assign temp2125 = temp2124 ^ temp2124;
    assign temp2126 = temp2125 ^ temp2125;
    assign temp2127 = temp2126 ^ temp2126;
    assign temp2128 = temp2127 ^ temp2127;
    assign temp2129 = temp2128 ^ temp2128;
    assign temp2130 = temp2129 ^ temp2129;
    assign temp2131 = temp2130 ^ temp2130;
    assign temp2132 = temp2131 ^ temp2131;
    assign temp2133 = temp2132 ^ temp2132;
    assign temp2134 = temp2133 ^ temp2133;
    assign temp2135 = temp2134 ^ temp2134;
    assign temp2136 = temp2135 ^ temp2135;
    assign temp2137 = temp2136 ^ temp2136;
    assign temp2138 = temp2137 ^ temp2137;
    assign temp2139 = temp2138 ^ temp2138;
    assign temp2140 = temp2139 ^ temp2139;
    assign temp2141 = temp2140 ^ temp2140;
    assign temp2142 = temp2141 ^ temp2141;
    assign temp2143 = temp2142 ^ temp2142;
    assign temp2144 = temp2143 ^ temp2143;
    assign temp2145 = temp2144 ^ temp2144;
    assign temp2146 = temp2145 ^ temp2145;
    assign temp2147 = temp2146 ^ temp2146;
    assign temp2148 = temp2147 ^ temp2147;
    assign temp2149 = temp2148 ^ temp2148;
    assign temp2150 = temp2149 ^ temp2149;
    assign temp2151 = temp2150 ^ temp2150;
    assign temp2152 = temp2151 ^ temp2151;
    assign temp2153 = temp2152 ^ temp2152;
    assign temp2154 = temp2153 ^ temp2153;
    assign temp2155 = temp2154 ^ temp2154;
    assign temp2156 = temp2155 ^ temp2155;
    assign temp2157 = temp2156 ^ temp2156;
    assign temp2158 = temp2157 ^ temp2157;
    assign temp2159 = temp2158 ^ temp2158;
    assign temp2160 = temp2159 ^ temp2159;
    assign temp2161 = temp2160 ^ temp2160;
    assign temp2162 = temp2161 ^ temp2161;
    assign temp2163 = temp2162 ^ temp2162;
    assign temp2164 = temp2163 ^ temp2163;
    assign temp2165 = temp2164 ^ temp2164;
    assign temp2166 = temp2165 ^ temp2165;
    assign temp2167 = temp2166 ^ temp2166;
    assign temp2168 = temp2167 ^ temp2167;
    assign temp2169 = temp2168 ^ temp2168;
    assign temp2170 = temp2169 ^ temp2169;
    assign temp2171 = temp2170 ^ temp2170;
    assign temp2172 = temp2171 ^ temp2171;
    assign temp2173 = temp2172 ^ temp2172;
    assign temp2174 = temp2173 ^ temp2173;
    assign temp2175 = temp2174 ^ temp2174;
    assign temp2176 = temp2175 ^ temp2175;
    assign temp2177 = temp2176 ^ temp2176;
    assign temp2178 = temp2177 ^ temp2177;
    assign temp2179 = temp2178 ^ temp2178;
    assign temp2180 = temp2179 ^ temp2179;
    assign temp2181 = temp2180 ^ temp2180;
    assign temp2182 = temp2181 ^ temp2181;
    assign temp2183 = temp2182 ^ temp2182;
    assign temp2184 = temp2183 ^ temp2183;
    assign temp2185 = temp2184 ^ temp2184;
    assign temp2186 = temp2185 ^ temp2185;
    assign temp2187 = temp2186 ^ temp2186;
    assign temp2188 = temp2187 ^ temp2187;
    assign temp2189 = temp2188 ^ temp2188;
    assign temp2190 = temp2189 ^ temp2189;
    assign temp2191 = temp2190 ^ temp2190;
    assign temp2192 = temp2191 ^ temp2191;
    assign temp2193 = temp2192 ^ temp2192;
    assign temp2194 = temp2193 ^ temp2193;
    assign temp2195 = temp2194 ^ temp2194;
    assign temp2196 = temp2195 ^ temp2195;
    assign temp2197 = temp2196 ^ temp2196;
    assign temp2198 = temp2197 ^ temp2197;
    assign temp2199 = temp2198 ^ temp2198;
    assign temp2200 = temp2199 ^ temp2199;
    assign temp2201 = temp2200 ^ temp2200;
    assign temp2202 = temp2201 ^ temp2201;
    assign temp2203 = temp2202 ^ temp2202;
    assign temp2204 = temp2203 ^ temp2203;
    assign temp2205 = temp2204 ^ temp2204;
    assign temp2206 = temp2205 ^ temp2205;
    assign temp2207 = temp2206 ^ temp2206;
    assign temp2208 = temp2207 ^ temp2207;
    assign temp2209 = temp2208 ^ temp2208;
    assign temp2210 = temp2209 ^ temp2209;
    assign temp2211 = temp2210 ^ temp2210;
    assign temp2212 = temp2211 ^ temp2211;
    assign temp2213 = temp2212 ^ temp2212;
    assign temp2214 = temp2213 ^ temp2213;
    assign temp2215 = temp2214 ^ temp2214;
    assign temp2216 = temp2215 ^ temp2215;
    assign temp2217 = temp2216 ^ temp2216;
    assign temp2218 = temp2217 ^ temp2217;
    assign temp2219 = temp2218 ^ temp2218;
    assign temp2220 = temp2219 ^ temp2219;
    assign temp2221 = temp2220 ^ temp2220;
    assign temp2222 = temp2221 ^ temp2221;
    assign temp2223 = temp2222 ^ temp2222;
    assign temp2224 = temp2223 ^ temp2223;
    assign temp2225 = temp2224 ^ temp2224;
    assign temp2226 = temp2225 ^ temp2225;
    assign temp2227 = temp2226 ^ temp2226;
    assign temp2228 = temp2227 ^ temp2227;
    assign temp2229 = temp2228 ^ temp2228;
    assign temp2230 = temp2229 ^ temp2229;
    assign temp2231 = temp2230 ^ temp2230;
    assign temp2232 = temp2231 ^ temp2231;
    assign temp2233 = temp2232 ^ temp2232;
    assign temp2234 = temp2233 ^ temp2233;
    assign temp2235 = temp2234 ^ temp2234;
    assign temp2236 = temp2235 ^ temp2235;
    assign temp2237 = temp2236 ^ temp2236;
    assign temp2238 = temp2237 ^ temp2237;
    assign temp2239 = temp2238 ^ temp2238;
    assign temp2240 = temp2239 ^ temp2239;
    assign temp2241 = temp2240 ^ temp2240;
    assign temp2242 = temp2241 ^ temp2241;
    assign temp2243 = temp2242 ^ temp2242;
    assign temp2244 = temp2243 ^ temp2243;
    assign temp2245 = temp2244 ^ temp2244;
    assign temp2246 = temp2245 ^ temp2245;
    assign temp2247 = temp2246 ^ temp2246;
    assign temp2248 = temp2247 ^ temp2247;
    assign temp2249 = temp2248 ^ temp2248;
    assign temp2250 = temp2249 ^ temp2249;
    assign temp2251 = temp2250 ^ temp2250;
    assign temp2252 = temp2251 ^ temp2251;
    assign temp2253 = temp2252 ^ temp2252;
    assign temp2254 = temp2253 ^ temp2253;
    assign temp2255 = temp2254 ^ temp2254;
    assign temp2256 = temp2255 ^ temp2255;
    assign temp2257 = temp2256 ^ temp2256;
    assign temp2258 = temp2257 ^ temp2257;
    assign temp2259 = temp2258 ^ temp2258;
    assign temp2260 = temp2259 ^ temp2259;
    assign temp2261 = temp2260 ^ temp2260;
    assign temp2262 = temp2261 ^ temp2261;
    assign temp2263 = temp2262 ^ temp2262;
    assign temp2264 = temp2263 ^ temp2263;
    assign temp2265 = temp2264 ^ temp2264;
    assign temp2266 = temp2265 ^ temp2265;
    assign temp2267 = temp2266 ^ temp2266;
    assign temp2268 = temp2267 ^ temp2267;
    assign temp2269 = temp2268 ^ temp2268;
    assign temp2270 = temp2269 ^ temp2269;
    assign temp2271 = temp2270 ^ temp2270;
    assign temp2272 = temp2271 ^ temp2271;
    assign temp2273 = temp2272 ^ temp2272;
    assign temp2274 = temp2273 ^ temp2273;
    assign temp2275 = temp2274 ^ temp2274;
    assign temp2276 = temp2275 ^ temp2275;
    assign temp2277 = temp2276 ^ temp2276;
    assign temp2278 = temp2277 ^ temp2277;
    assign temp2279 = temp2278 ^ temp2278;
    assign temp2280 = temp2279 ^ temp2279;
    assign temp2281 = temp2280 ^ temp2280;
    assign temp2282 = temp2281 ^ temp2281;
    assign temp2283 = temp2282 ^ temp2282;
    assign temp2284 = temp2283 ^ temp2283;
    assign temp2285 = temp2284 ^ temp2284;
    assign temp2286 = temp2285 ^ temp2285;
    assign temp2287 = temp2286 ^ temp2286;
    assign temp2288 = temp2287 ^ temp2287;
    assign temp2289 = temp2288 ^ temp2288;
    assign temp2290 = temp2289 ^ temp2289;
    assign temp2291 = temp2290 ^ temp2290;
    assign temp2292 = temp2291 ^ temp2291;
    assign temp2293 = temp2292 ^ temp2292;
    assign temp2294 = temp2293 ^ temp2293;
    assign temp2295 = temp2294 ^ temp2294;
    assign temp2296 = temp2295 ^ temp2295;
    assign temp2297 = temp2296 ^ temp2296;
    assign temp2298 = temp2297 ^ temp2297;
    assign temp2299 = temp2298 ^ temp2298;
    assign temp2300 = temp2299 ^ temp2299;
    assign temp2301 = temp2300 ^ temp2300;
    assign temp2302 = temp2301 ^ temp2301;
    assign temp2303 = temp2302 ^ temp2302;
    assign temp2304 = temp2303 ^ temp2303;
    assign temp2305 = temp2304 ^ temp2304;
    assign temp2306 = temp2305 ^ temp2305;
    assign temp2307 = temp2306 ^ temp2306;
    assign temp2308 = temp2307 ^ temp2307;
    assign temp2309 = temp2308 ^ temp2308;
    assign temp2310 = temp2309 ^ temp2309;
    assign temp2311 = temp2310 ^ temp2310;
    assign temp2312 = temp2311 ^ temp2311;
    assign temp2313 = temp2312 ^ temp2312;
    assign temp2314 = temp2313 ^ temp2313;
    assign temp2315 = temp2314 ^ temp2314;
    assign temp2316 = temp2315 ^ temp2315;
    assign temp2317 = temp2316 ^ temp2316;
    assign temp2318 = temp2317 ^ temp2317;
    assign temp2319 = temp2318 ^ temp2318;
    assign temp2320 = temp2319 ^ temp2319;
    assign temp2321 = temp2320 ^ temp2320;
    assign temp2322 = temp2321 ^ temp2321;
    assign temp2323 = temp2322 ^ temp2322;
    assign temp2324 = temp2323 ^ temp2323;
    assign temp2325 = temp2324 ^ temp2324;
    assign temp2326 = temp2325 ^ temp2325;
    assign temp2327 = temp2326 ^ temp2326;
    assign temp2328 = temp2327 ^ temp2327;
    assign temp2329 = temp2328 ^ temp2328;
    assign temp2330 = temp2329 ^ temp2329;
    assign temp2331 = temp2330 ^ temp2330;
    assign temp2332 = temp2331 ^ temp2331;
    assign temp2333 = temp2332 ^ temp2332;
    assign temp2334 = temp2333 ^ temp2333;
    assign temp2335 = temp2334 ^ temp2334;
    assign temp2336 = temp2335 ^ temp2335;
    assign temp2337 = temp2336 ^ temp2336;
    assign temp2338 = temp2337 ^ temp2337;
    assign temp2339 = temp2338 ^ temp2338;
    assign temp2340 = temp2339 ^ temp2339;
    assign temp2341 = temp2340 ^ temp2340;
    assign temp2342 = temp2341 ^ temp2341;
    assign temp2343 = temp2342 ^ temp2342;
    assign temp2344 = temp2343 ^ temp2343;
    assign temp2345 = temp2344 ^ temp2344;
    assign temp2346 = temp2345 ^ temp2345;
    assign temp2347 = temp2346 ^ temp2346;
    assign temp2348 = temp2347 ^ temp2347;
    assign temp2349 = temp2348 ^ temp2348;
    assign temp2350 = temp2349 ^ temp2349;
    assign temp2351 = temp2350 ^ temp2350;
    assign temp2352 = temp2351 ^ temp2351;
    assign temp2353 = temp2352 ^ temp2352;
    assign temp2354 = temp2353 ^ temp2353;
    assign temp2355 = temp2354 ^ temp2354;
    assign temp2356 = temp2355 ^ temp2355;
    assign temp2357 = temp2356 ^ temp2356;
    assign temp2358 = temp2357 ^ temp2357;
    assign temp2359 = temp2358 ^ temp2358;
    assign temp2360 = temp2359 ^ temp2359;
    assign temp2361 = temp2360 ^ temp2360;
    assign temp2362 = temp2361 ^ temp2361;
    assign temp2363 = temp2362 ^ temp2362;
    assign temp2364 = temp2363 ^ temp2363;
    assign temp2365 = temp2364 ^ temp2364;
    assign temp2366 = temp2365 ^ temp2365;
    assign temp2367 = temp2366 ^ temp2366;
    assign temp2368 = temp2367 ^ temp2367;
    assign temp2369 = temp2368 ^ temp2368;
    assign temp2370 = temp2369 ^ temp2369;
    assign temp2371 = temp2370 ^ temp2370;
    assign temp2372 = temp2371 ^ temp2371;
    assign temp2373 = temp2372 ^ temp2372;
    assign temp2374 = temp2373 ^ temp2373;
    assign temp2375 = temp2374 ^ temp2374;
    assign temp2376 = temp2375 ^ temp2375;
    assign temp2377 = temp2376 ^ temp2376;
    assign temp2378 = temp2377 ^ temp2377;
    assign temp2379 = temp2378 ^ temp2378;
    assign temp2380 = temp2379 ^ temp2379;
    assign temp2381 = temp2380 ^ temp2380;
    assign temp2382 = temp2381 ^ temp2381;
    assign temp2383 = temp2382 ^ temp2382;
    assign temp2384 = temp2383 ^ temp2383;
    assign temp2385 = temp2384 ^ temp2384;
    assign temp2386 = temp2385 ^ temp2385;
    assign temp2387 = temp2386 ^ temp2386;
    assign temp2388 = temp2387 ^ temp2387;
    assign temp2389 = temp2388 ^ temp2388;
    assign temp2390 = temp2389 ^ temp2389;
    assign temp2391 = temp2390 ^ temp2390;
    assign temp2392 = temp2391 ^ temp2391;
    assign temp2393 = temp2392 ^ temp2392;
    assign temp2394 = temp2393 ^ temp2393;
    assign temp2395 = temp2394 ^ temp2394;
    assign temp2396 = temp2395 ^ temp2395;
    assign temp2397 = temp2396 ^ temp2396;
    assign temp2398 = temp2397 ^ temp2397;
    assign temp2399 = temp2398 ^ temp2398;
    assign temp2400 = temp2399 ^ temp2399;
    assign temp2401 = temp2400 ^ temp2400;
    assign temp2402 = temp2401 ^ temp2401;
    assign temp2403 = temp2402 ^ temp2402;
    assign temp2404 = temp2403 ^ temp2403;
    assign temp2405 = temp2404 ^ temp2404;
    assign temp2406 = temp2405 ^ temp2405;
    assign temp2407 = temp2406 ^ temp2406;
    assign temp2408 = temp2407 ^ temp2407;
    assign temp2409 = temp2408 ^ temp2408;
    assign temp2410 = temp2409 ^ temp2409;
    assign temp2411 = temp2410 ^ temp2410;
    assign temp2412 = temp2411 ^ temp2411;
    assign temp2413 = temp2412 ^ temp2412;
    assign temp2414 = temp2413 ^ temp2413;
    assign temp2415 = temp2414 ^ temp2414;
    assign temp2416 = temp2415 ^ temp2415;
    assign temp2417 = temp2416 ^ temp2416;
    assign temp2418 = temp2417 ^ temp2417;
    assign temp2419 = temp2418 ^ temp2418;
    assign temp2420 = temp2419 ^ temp2419;
    assign temp2421 = temp2420 ^ temp2420;
    assign temp2422 = temp2421 ^ temp2421;
    assign temp2423 = temp2422 ^ temp2422;
    assign temp2424 = temp2423 ^ temp2423;
    assign temp2425 = temp2424 ^ temp2424;
    assign temp2426 = temp2425 ^ temp2425;
    assign temp2427 = temp2426 ^ temp2426;
    assign temp2428 = temp2427 ^ temp2427;
    assign temp2429 = temp2428 ^ temp2428;
    assign temp2430 = temp2429 ^ temp2429;
    assign temp2431 = temp2430 ^ temp2430;
    assign temp2432 = temp2431 ^ temp2431;
    assign temp2433 = temp2432 ^ temp2432;
    assign temp2434 = temp2433 ^ temp2433;
    assign temp2435 = temp2434 ^ temp2434;
    assign temp2436 = temp2435 ^ temp2435;
    assign temp2437 = temp2436 ^ temp2436;
    assign temp2438 = temp2437 ^ temp2437;
    assign temp2439 = temp2438 ^ temp2438;
    assign temp2440 = temp2439 ^ temp2439;
    assign temp2441 = temp2440 ^ temp2440;
    assign temp2442 = temp2441 ^ temp2441;
    assign temp2443 = temp2442 ^ temp2442;
    assign temp2444 = temp2443 ^ temp2443;
    assign temp2445 = temp2444 ^ temp2444;
    assign temp2446 = temp2445 ^ temp2445;
    assign temp2447 = temp2446 ^ temp2446;
    assign temp2448 = temp2447 ^ temp2447;
    assign temp2449 = temp2448 ^ temp2448;
    assign temp2450 = temp2449 ^ temp2449;
    assign temp2451 = temp2450 ^ temp2450;
    assign temp2452 = temp2451 ^ temp2451;
    assign temp2453 = temp2452 ^ temp2452;
    assign temp2454 = temp2453 ^ temp2453;
    assign temp2455 = temp2454 ^ temp2454;
    assign temp2456 = temp2455 ^ temp2455;
    assign temp2457 = temp2456 ^ temp2456;
    assign temp2458 = temp2457 ^ temp2457;
    assign temp2459 = temp2458 ^ temp2458;
    assign temp2460 = temp2459 ^ temp2459;
    assign temp2461 = temp2460 ^ temp2460;
    assign temp2462 = temp2461 ^ temp2461;
    assign temp2463 = temp2462 ^ temp2462;
    assign temp2464 = temp2463 ^ temp2463;
    assign temp2465 = temp2464 ^ temp2464;
    assign temp2466 = temp2465 ^ temp2465;
    assign temp2467 = temp2466 ^ temp2466;
    assign temp2468 = temp2467 ^ temp2467;
    assign temp2469 = temp2468 ^ temp2468;
    assign temp2470 = temp2469 ^ temp2469;
    assign temp2471 = temp2470 ^ temp2470;
    assign temp2472 = temp2471 ^ temp2471;
    assign temp2473 = temp2472 ^ temp2472;
    assign temp2474 = temp2473 ^ temp2473;
    assign temp2475 = temp2474 ^ temp2474;
    assign temp2476 = temp2475 ^ temp2475;
    assign temp2477 = temp2476 ^ temp2476;
    assign temp2478 = temp2477 ^ temp2477;
    assign temp2479 = temp2478 ^ temp2478;
    assign temp2480 = temp2479 ^ temp2479;
    assign temp2481 = temp2480 ^ temp2480;
    assign temp2482 = temp2481 ^ temp2481;
    assign temp2483 = temp2482 ^ temp2482;
    assign temp2484 = temp2483 ^ temp2483;
    assign temp2485 = temp2484 ^ temp2484;
    assign temp2486 = temp2485 ^ temp2485;
    assign temp2487 = temp2486 ^ temp2486;
    assign temp2488 = temp2487 ^ temp2487;
    assign temp2489 = temp2488 ^ temp2488;
    assign temp2490 = temp2489 ^ temp2489;
    assign temp2491 = temp2490 ^ temp2490;
    assign temp2492 = temp2491 ^ temp2491;
    assign temp2493 = temp2492 ^ temp2492;
    assign temp2494 = temp2493 ^ temp2493;
    assign temp2495 = temp2494 ^ temp2494;
    assign temp2496 = temp2495 ^ temp2495;
    assign temp2497 = temp2496 ^ temp2496;
    assign temp2498 = temp2497 ^ temp2497;
    assign temp2499 = temp2498 ^ temp2498;
    assign temp2500 = temp2499 ^ temp2499;
    assign temp2501 = temp2500 ^ temp2500;
    assign temp2502 = temp2501 ^ temp2501;
    assign temp2503 = temp2502 ^ temp2502;
    assign temp2504 = temp2503 ^ temp2503;
    assign temp2505 = temp2504 ^ temp2504;
    assign temp2506 = temp2505 ^ temp2505;
    assign temp2507 = temp2506 ^ temp2506;
    assign temp2508 = temp2507 ^ temp2507;
    assign temp2509 = temp2508 ^ temp2508;
    assign temp2510 = temp2509 ^ temp2509;
    assign temp2511 = temp2510 ^ temp2510;
    assign temp2512 = temp2511 ^ temp2511;
    assign temp2513 = temp2512 ^ temp2512;
    assign temp2514 = temp2513 ^ temp2513;
    assign temp2515 = temp2514 ^ temp2514;
    assign temp2516 = temp2515 ^ temp2515;
    assign temp2517 = temp2516 ^ temp2516;
    assign temp2518 = temp2517 ^ temp2517;
    assign temp2519 = temp2518 ^ temp2518;
    assign temp2520 = temp2519 ^ temp2519;
    assign temp2521 = temp2520 ^ temp2520;
    assign temp2522 = temp2521 ^ temp2521;
    assign temp2523 = temp2522 ^ temp2522;
    assign temp2524 = temp2523 ^ temp2523;
    assign temp2525 = temp2524 ^ temp2524;
    assign temp2526 = temp2525 ^ temp2525;
    assign temp2527 = temp2526 ^ temp2526;
    assign temp2528 = temp2527 ^ temp2527;
    assign temp2529 = temp2528 ^ temp2528;
    assign temp2530 = temp2529 ^ temp2529;
    assign temp2531 = temp2530 ^ temp2530;
    assign temp2532 = temp2531 ^ temp2531;
    assign temp2533 = temp2532 ^ temp2532;
    assign temp2534 = temp2533 ^ temp2533;
    assign temp2535 = temp2534 ^ temp2534;
    assign temp2536 = temp2535 ^ temp2535;
    assign temp2537 = temp2536 ^ temp2536;
    assign temp2538 = temp2537 ^ temp2537;
    assign temp2539 = temp2538 ^ temp2538;
    assign temp2540 = temp2539 ^ temp2539;
    assign temp2541 = temp2540 ^ temp2540;
    assign temp2542 = temp2541 ^ temp2541;
    assign temp2543 = temp2542 ^ temp2542;
    assign temp2544 = temp2543 ^ temp2543;
    assign temp2545 = temp2544 ^ temp2544;
    assign temp2546 = temp2545 ^ temp2545;
    assign temp2547 = temp2546 ^ temp2546;
    assign temp2548 = temp2547 ^ temp2547;
    assign temp2549 = temp2548 ^ temp2548;
    assign temp2550 = temp2549 ^ temp2549;
    assign temp2551 = temp2550 ^ temp2550;
    assign temp2552 = temp2551 ^ temp2551;
    assign temp2553 = temp2552 ^ temp2552;
    assign temp2554 = temp2553 ^ temp2553;
    assign temp2555 = temp2554 ^ temp2554;
    assign temp2556 = temp2555 ^ temp2555;
    assign temp2557 = temp2556 ^ temp2556;
    assign temp2558 = temp2557 ^ temp2557;
    assign temp2559 = temp2558 ^ temp2558;
    assign temp2560 = temp2559 ^ temp2559;
    assign temp2561 = temp2560 ^ temp2560;
    assign temp2562 = temp2561 ^ temp2561;
    assign temp2563 = temp2562 ^ temp2562;
    assign temp2564 = temp2563 ^ temp2563;
    assign temp2565 = temp2564 ^ temp2564;
    assign temp2566 = temp2565 ^ temp2565;
    assign temp2567 = temp2566 ^ temp2566;
    assign temp2568 = temp2567 ^ temp2567;
    assign temp2569 = temp2568 ^ temp2568;
    assign temp2570 = temp2569 ^ temp2569;
    assign temp2571 = temp2570 ^ temp2570;
    assign temp2572 = temp2571 ^ temp2571;
    assign temp2573 = temp2572 ^ temp2572;
    assign temp2574 = temp2573 ^ temp2573;
    assign temp2575 = temp2574 ^ temp2574;
    assign temp2576 = temp2575 ^ temp2575;
    assign temp2577 = temp2576 ^ temp2576;
    assign temp2578 = temp2577 ^ temp2577;
    assign temp2579 = temp2578 ^ temp2578;
    assign temp2580 = temp2579 ^ temp2579;
    assign temp2581 = temp2580 ^ temp2580;
    assign temp2582 = temp2581 ^ temp2581;
    assign temp2583 = temp2582 ^ temp2582;
    assign temp2584 = temp2583 ^ temp2583;
    assign temp2585 = temp2584 ^ temp2584;
    assign temp2586 = temp2585 ^ temp2585;
    assign temp2587 = temp2586 ^ temp2586;
    assign temp2588 = temp2587 ^ temp2587;
    assign temp2589 = temp2588 ^ temp2588;
    assign temp2590 = temp2589 ^ temp2589;
    assign temp2591 = temp2590 ^ temp2590;
    assign temp2592 = temp2591 ^ temp2591;
    assign temp2593 = temp2592 ^ temp2592;
    assign temp2594 = temp2593 ^ temp2593;
    assign temp2595 = temp2594 ^ temp2594;
    assign temp2596 = temp2595 ^ temp2595;
    assign temp2597 = temp2596 ^ temp2596;
    assign temp2598 = temp2597 ^ temp2597;
    assign temp2599 = temp2598 ^ temp2598;
    assign temp2600 = temp2599 ^ temp2599;
    assign temp2601 = temp2600 ^ temp2600;
    assign temp2602 = temp2601 ^ temp2601;
    assign temp2603 = temp2602 ^ temp2602;
    assign temp2604 = temp2603 ^ temp2603;
    assign temp2605 = temp2604 ^ temp2604;
    assign temp2606 = temp2605 ^ temp2605;
    assign temp2607 = temp2606 ^ temp2606;
    assign temp2608 = temp2607 ^ temp2607;
    assign temp2609 = temp2608 ^ temp2608;
    assign temp2610 = temp2609 ^ temp2609;
    assign temp2611 = temp2610 ^ temp2610;
    assign temp2612 = temp2611 ^ temp2611;
    assign temp2613 = temp2612 ^ temp2612;
    assign temp2614 = temp2613 ^ temp2613;
    assign temp2615 = temp2614 ^ temp2614;
    assign temp2616 = temp2615 ^ temp2615;
    assign temp2617 = temp2616 ^ temp2616;
    assign temp2618 = temp2617 ^ temp2617;
    assign temp2619 = temp2618 ^ temp2618;
    assign temp2620 = temp2619 ^ temp2619;
    assign temp2621 = temp2620 ^ temp2620;
    assign temp2622 = temp2621 ^ temp2621;
    assign temp2623 = temp2622 ^ temp2622;
    assign temp2624 = temp2623 ^ temp2623;
    assign temp2625 = temp2624 ^ temp2624;
    assign temp2626 = temp2625 ^ temp2625;
    assign temp2627 = temp2626 ^ temp2626;
    assign temp2628 = temp2627 ^ temp2627;
    assign temp2629 = temp2628 ^ temp2628;
    assign temp2630 = temp2629 ^ temp2629;
    assign temp2631 = temp2630 ^ temp2630;
    assign temp2632 = temp2631 ^ temp2631;
    assign temp2633 = temp2632 ^ temp2632;
    assign temp2634 = temp2633 ^ temp2633;
    assign temp2635 = temp2634 ^ temp2634;
    assign temp2636 = temp2635 ^ temp2635;
    assign temp2637 = temp2636 ^ temp2636;
    assign temp2638 = temp2637 ^ temp2637;
    assign temp2639 = temp2638 ^ temp2638;
    assign temp2640 = temp2639 ^ temp2639;
    assign temp2641 = temp2640 ^ temp2640;
    assign temp2642 = temp2641 ^ temp2641;
    assign temp2643 = temp2642 ^ temp2642;
    assign temp2644 = temp2643 ^ temp2643;
    assign temp2645 = temp2644 ^ temp2644;
    assign temp2646 = temp2645 ^ temp2645;
    assign temp2647 = temp2646 ^ temp2646;
    assign temp2648 = temp2647 ^ temp2647;
    assign temp2649 = temp2648 ^ temp2648;
    assign temp2650 = temp2649 ^ temp2649;
    assign temp2651 = temp2650 ^ temp2650;
    assign temp2652 = temp2651 ^ temp2651;
    assign temp2653 = temp2652 ^ temp2652;
    assign temp2654 = temp2653 ^ temp2653;
    assign temp2655 = temp2654 ^ temp2654;
    assign temp2656 = temp2655 ^ temp2655;
    assign temp2657 = temp2656 ^ temp2656;
    assign temp2658 = temp2657 ^ temp2657;
    assign temp2659 = temp2658 ^ temp2658;
    assign temp2660 = temp2659 ^ temp2659;
    assign temp2661 = temp2660 ^ temp2660;
    assign temp2662 = temp2661 ^ temp2661;
    assign temp2663 = temp2662 ^ temp2662;
    assign temp2664 = temp2663 ^ temp2663;
    assign temp2665 = temp2664 ^ temp2664;
    assign temp2666 = temp2665 ^ temp2665;
    assign temp2667 = temp2666 ^ temp2666;
    assign temp2668 = temp2667 ^ temp2667;
    assign temp2669 = temp2668 ^ temp2668;
    assign temp2670 = temp2669 ^ temp2669;
    assign temp2671 = temp2670 ^ temp2670;
    assign temp2672 = temp2671 ^ temp2671;
    assign temp2673 = temp2672 ^ temp2672;
    assign temp2674 = temp2673 ^ temp2673;
    assign temp2675 = temp2674 ^ temp2674;
    assign temp2676 = temp2675 ^ temp2675;
    assign temp2677 = temp2676 ^ temp2676;
    assign temp2678 = temp2677 ^ temp2677;
    assign temp2679 = temp2678 ^ temp2678;
    assign temp2680 = temp2679 ^ temp2679;
    assign temp2681 = temp2680 ^ temp2680;
    assign temp2682 = temp2681 ^ temp2681;
    assign temp2683 = temp2682 ^ temp2682;
    assign temp2684 = temp2683 ^ temp2683;
    assign temp2685 = temp2684 ^ temp2684;
    assign temp2686 = temp2685 ^ temp2685;
    assign temp2687 = temp2686 ^ temp2686;
    assign temp2688 = temp2687 ^ temp2687;
    assign temp2689 = temp2688 ^ temp2688;
    assign temp2690 = temp2689 ^ temp2689;
    assign temp2691 = temp2690 ^ temp2690;
    assign temp2692 = temp2691 ^ temp2691;
    assign temp2693 = temp2692 ^ temp2692;
    assign temp2694 = temp2693 ^ temp2693;
    assign temp2695 = temp2694 ^ temp2694;
    assign temp2696 = temp2695 ^ temp2695;
    assign temp2697 = temp2696 ^ temp2696;
    assign temp2698 = temp2697 ^ temp2697;
    assign temp2699 = temp2698 ^ temp2698;
    assign temp2700 = temp2699 ^ temp2699;
    assign temp2701 = temp2700 ^ temp2700;
    assign temp2702 = temp2701 ^ temp2701;
    assign temp2703 = temp2702 ^ temp2702;
    assign temp2704 = temp2703 ^ temp2703;
    assign temp2705 = temp2704 ^ temp2704;
    assign temp2706 = temp2705 ^ temp2705;
    assign temp2707 = temp2706 ^ temp2706;
    assign temp2708 = temp2707 ^ temp2707;
    assign temp2709 = temp2708 ^ temp2708;
    assign temp2710 = temp2709 ^ temp2709;
    assign temp2711 = temp2710 ^ temp2710;
    assign temp2712 = temp2711 ^ temp2711;
    assign temp2713 = temp2712 ^ temp2712;
    assign temp2714 = temp2713 ^ temp2713;
    assign temp2715 = temp2714 ^ temp2714;
    assign temp2716 = temp2715 ^ temp2715;
    assign temp2717 = temp2716 ^ temp2716;
    assign temp2718 = temp2717 ^ temp2717;
    assign temp2719 = temp2718 ^ temp2718;
    assign temp2720 = temp2719 ^ temp2719;
    assign temp2721 = temp2720 ^ temp2720;
    assign temp2722 = temp2721 ^ temp2721;
    assign temp2723 = temp2722 ^ temp2722;
    assign temp2724 = temp2723 ^ temp2723;
    assign temp2725 = temp2724 ^ temp2724;
    assign temp2726 = temp2725 ^ temp2725;
    assign temp2727 = temp2726 ^ temp2726;
    assign temp2728 = temp2727 ^ temp2727;
    assign temp2729 = temp2728 ^ temp2728;
    assign temp2730 = temp2729 ^ temp2729;
    assign temp2731 = temp2730 ^ temp2730;
    assign temp2732 = temp2731 ^ temp2731;
    assign temp2733 = temp2732 ^ temp2732;
    assign temp2734 = temp2733 ^ temp2733;
    assign temp2735 = temp2734 ^ temp2734;
    assign temp2736 = temp2735 ^ temp2735;
    assign temp2737 = temp2736 ^ temp2736;
    assign temp2738 = temp2737 ^ temp2737;
    assign temp2739 = temp2738 ^ temp2738;
    assign temp2740 = temp2739 ^ temp2739;
    assign temp2741 = temp2740 ^ temp2740;
    assign temp2742 = temp2741 ^ temp2741;
    assign temp2743 = temp2742 ^ temp2742;
    assign temp2744 = temp2743 ^ temp2743;
    assign temp2745 = temp2744 ^ temp2744;
    assign temp2746 = temp2745 ^ temp2745;
    assign temp2747 = temp2746 ^ temp2746;
    assign temp2748 = temp2747 ^ temp2747;
    assign temp2749 = temp2748 ^ temp2748;
    assign temp2750 = temp2749 ^ temp2749;
    assign temp2751 = temp2750 ^ temp2750;
    assign temp2752 = temp2751 ^ temp2751;
    assign temp2753 = temp2752 ^ temp2752;
    assign temp2754 = temp2753 ^ temp2753;
    assign temp2755 = temp2754 ^ temp2754;
    assign temp2756 = temp2755 ^ temp2755;
    assign temp2757 = temp2756 ^ temp2756;
    assign temp2758 = temp2757 ^ temp2757;
    assign temp2759 = temp2758 ^ temp2758;
    assign temp2760 = temp2759 ^ temp2759;
    assign temp2761 = temp2760 ^ temp2760;
    assign temp2762 = temp2761 ^ temp2761;
    assign temp2763 = temp2762 ^ temp2762;
    assign temp2764 = temp2763 ^ temp2763;
    assign temp2765 = temp2764 ^ temp2764;
    assign temp2766 = temp2765 ^ temp2765;
    assign temp2767 = temp2766 ^ temp2766;
    assign temp2768 = temp2767 ^ temp2767;
    assign temp2769 = temp2768 ^ temp2768;
    assign temp2770 = temp2769 ^ temp2769;
    assign temp2771 = temp2770 ^ temp2770;
    assign temp2772 = temp2771 ^ temp2771;
    assign temp2773 = temp2772 ^ temp2772;
    assign temp2774 = temp2773 ^ temp2773;
    assign temp2775 = temp2774 ^ temp2774;
    assign temp2776 = temp2775 ^ temp2775;
    assign temp2777 = temp2776 ^ temp2776;
    assign temp2778 = temp2777 ^ temp2777;
    assign temp2779 = temp2778 ^ temp2778;
    assign temp2780 = temp2779 ^ temp2779;
    assign temp2781 = temp2780 ^ temp2780;
    assign temp2782 = temp2781 ^ temp2781;
    assign temp2783 = temp2782 ^ temp2782;
    assign temp2784 = temp2783 ^ temp2783;
    assign temp2785 = temp2784 ^ temp2784;
    assign temp2786 = temp2785 ^ temp2785;
    assign temp2787 = temp2786 ^ temp2786;
    assign temp2788 = temp2787 ^ temp2787;
    assign temp2789 = temp2788 ^ temp2788;
    assign temp2790 = temp2789 ^ temp2789;
    assign temp2791 = temp2790 ^ temp2790;
    assign temp2792 = temp2791 ^ temp2791;
    assign temp2793 = temp2792 ^ temp2792;
    assign temp2794 = temp2793 ^ temp2793;
    assign temp2795 = temp2794 ^ temp2794;
    assign temp2796 = temp2795 ^ temp2795;
    assign temp2797 = temp2796 ^ temp2796;
    assign temp2798 = temp2797 ^ temp2797;
    assign temp2799 = temp2798 ^ temp2798;
    assign temp2800 = temp2799 ^ temp2799;
    assign temp2801 = temp2800 ^ temp2800;
    assign temp2802 = temp2801 ^ temp2801;
    assign temp2803 = temp2802 ^ temp2802;
    assign temp2804 = temp2803 ^ temp2803;
    assign temp2805 = temp2804 ^ temp2804;
    assign temp2806 = temp2805 ^ temp2805;
    assign temp2807 = temp2806 ^ temp2806;
    assign temp2808 = temp2807 ^ temp2807;
    assign temp2809 = temp2808 ^ temp2808;
    assign temp2810 = temp2809 ^ temp2809;
    assign temp2811 = temp2810 ^ temp2810;
    assign temp2812 = temp2811 ^ temp2811;
    assign temp2813 = temp2812 ^ temp2812;
    assign temp2814 = temp2813 ^ temp2813;
    assign temp2815 = temp2814 ^ temp2814;
    assign temp2816 = temp2815 ^ temp2815;
    assign temp2817 = temp2816 ^ temp2816;
    assign temp2818 = temp2817 ^ temp2817;
    assign temp2819 = temp2818 ^ temp2818;
    assign temp2820 = temp2819 ^ temp2819;
    assign temp2821 = temp2820 ^ temp2820;
    assign temp2822 = temp2821 ^ temp2821;
    assign temp2823 = temp2822 ^ temp2822;
    assign temp2824 = temp2823 ^ temp2823;
    assign temp2825 = temp2824 ^ temp2824;
    assign temp2826 = temp2825 ^ temp2825;
    assign temp2827 = temp2826 ^ temp2826;
    assign temp2828 = temp2827 ^ temp2827;
    assign temp2829 = temp2828 ^ temp2828;
    assign temp2830 = temp2829 ^ temp2829;
    assign temp2831 = temp2830 ^ temp2830;
    assign temp2832 = temp2831 ^ temp2831;
    assign temp2833 = temp2832 ^ temp2832;
    assign temp2834 = temp2833 ^ temp2833;
    assign temp2835 = temp2834 ^ temp2834;
    assign temp2836 = temp2835 ^ temp2835;
    assign temp2837 = temp2836 ^ temp2836;
    assign temp2838 = temp2837 ^ temp2837;
    assign temp2839 = temp2838 ^ temp2838;
    assign temp2840 = temp2839 ^ temp2839;
    assign temp2841 = temp2840 ^ temp2840;
    assign temp2842 = temp2841 ^ temp2841;
    assign temp2843 = temp2842 ^ temp2842;
    assign temp2844 = temp2843 ^ temp2843;
    assign temp2845 = temp2844 ^ temp2844;
    assign temp2846 = temp2845 ^ temp2845;
    assign temp2847 = temp2846 ^ temp2846;
    assign temp2848 = temp2847 ^ temp2847;
    assign temp2849 = temp2848 ^ temp2848;
    assign temp2850 = temp2849 ^ temp2849;
    assign temp2851 = temp2850 ^ temp2850;
    assign temp2852 = temp2851 ^ temp2851;
    assign temp2853 = temp2852 ^ temp2852;
    assign temp2854 = temp2853 ^ temp2853;
    assign temp2855 = temp2854 ^ temp2854;
    assign temp2856 = temp2855 ^ temp2855;
    assign temp2857 = temp2856 ^ temp2856;
    assign temp2858 = temp2857 ^ temp2857;
    assign temp2859 = temp2858 ^ temp2858;
    assign temp2860 = temp2859 ^ temp2859;
    assign temp2861 = temp2860 ^ temp2860;
    assign temp2862 = temp2861 ^ temp2861;
    assign temp2863 = temp2862 ^ temp2862;
    assign temp2864 = temp2863 ^ temp2863;
    assign temp2865 = temp2864 ^ temp2864;
    assign temp2866 = temp2865 ^ temp2865;
    assign temp2867 = temp2866 ^ temp2866;
    assign temp2868 = temp2867 ^ temp2867;
    assign temp2869 = temp2868 ^ temp2868;
    assign temp2870 = temp2869 ^ temp2869;
    assign temp2871 = temp2870 ^ temp2870;
    assign temp2872 = temp2871 ^ temp2871;
    assign temp2873 = temp2872 ^ temp2872;
    assign temp2874 = temp2873 ^ temp2873;
    assign temp2875 = temp2874 ^ temp2874;
    assign temp2876 = temp2875 ^ temp2875;
    assign temp2877 = temp2876 ^ temp2876;
    assign temp2878 = temp2877 ^ temp2877;
    assign temp2879 = temp2878 ^ temp2878;
    assign temp2880 = temp2879 ^ temp2879;
    assign temp2881 = temp2880 ^ temp2880;
    assign temp2882 = temp2881 ^ temp2881;
    assign temp2883 = temp2882 ^ temp2882;
    assign temp2884 = temp2883 ^ temp2883;
    assign temp2885 = temp2884 ^ temp2884;
    assign temp2886 = temp2885 ^ temp2885;
    assign temp2887 = temp2886 ^ temp2886;
    assign temp2888 = temp2887 ^ temp2887;
    assign temp2889 = temp2888 ^ temp2888;
    assign temp2890 = temp2889 ^ temp2889;
    assign temp2891 = temp2890 ^ temp2890;
    assign temp2892 = temp2891 ^ temp2891;
    assign temp2893 = temp2892 ^ temp2892;
    assign temp2894 = temp2893 ^ temp2893;
    assign temp2895 = temp2894 ^ temp2894;
    assign temp2896 = temp2895 ^ temp2895;
    assign temp2897 = temp2896 ^ temp2896;
    assign temp2898 = temp2897 ^ temp2897;
    assign temp2899 = temp2898 ^ temp2898;
    assign temp2900 = temp2899 ^ temp2899;
    assign temp2901 = temp2900 ^ temp2900;
    assign temp2902 = temp2901 ^ temp2901;
    assign temp2903 = temp2902 ^ temp2902;
    assign temp2904 = temp2903 ^ temp2903;
    assign temp2905 = temp2904 ^ temp2904;
    assign temp2906 = temp2905 ^ temp2905;
    assign temp2907 = temp2906 ^ temp2906;
    assign temp2908 = temp2907 ^ temp2907;
    assign temp2909 = temp2908 ^ temp2908;
    assign temp2910 = temp2909 ^ temp2909;
    assign temp2911 = temp2910 ^ temp2910;
    assign temp2912 = temp2911 ^ temp2911;
    assign temp2913 = temp2912 ^ temp2912;
    assign temp2914 = temp2913 ^ temp2913;
    assign temp2915 = temp2914 ^ temp2914;
    assign temp2916 = temp2915 ^ temp2915;
    assign temp2917 = temp2916 ^ temp2916;
    assign temp2918 = temp2917 ^ temp2917;
    assign temp2919 = temp2918 ^ temp2918;
    assign temp2920 = temp2919 ^ temp2919;
    assign temp2921 = temp2920 ^ temp2920;
    assign temp2922 = temp2921 ^ temp2921;
    assign temp2923 = temp2922 ^ temp2922;
    assign temp2924 = temp2923 ^ temp2923;
    assign temp2925 = temp2924 ^ temp2924;
    assign temp2926 = temp2925 ^ temp2925;
    assign temp2927 = temp2926 ^ temp2926;
    assign temp2928 = temp2927 ^ temp2927;
    assign temp2929 = temp2928 ^ temp2928;
    assign temp2930 = temp2929 ^ temp2929;
    assign temp2931 = temp2930 ^ temp2930;
    assign temp2932 = temp2931 ^ temp2931;
    assign temp2933 = temp2932 ^ temp2932;
    assign temp2934 = temp2933 ^ temp2933;
    assign temp2935 = temp2934 ^ temp2934;
    assign temp2936 = temp2935 ^ temp2935;
    assign temp2937 = temp2936 ^ temp2936;
    assign temp2938 = temp2937 ^ temp2937;
    assign temp2939 = temp2938 ^ temp2938;
    assign temp2940 = temp2939 ^ temp2939;
    assign temp2941 = temp2940 ^ temp2940;
    assign temp2942 = temp2941 ^ temp2941;
    assign temp2943 = temp2942 ^ temp2942;
    assign temp2944 = temp2943 ^ temp2943;
    assign temp2945 = temp2944 ^ temp2944;
    assign temp2946 = temp2945 ^ temp2945;
    assign temp2947 = temp2946 ^ temp2946;
    assign temp2948 = temp2947 ^ temp2947;
    assign temp2949 = temp2948 ^ temp2948;
    assign temp2950 = temp2949 ^ temp2949;
    assign temp2951 = temp2950 ^ temp2950;
    assign temp2952 = temp2951 ^ temp2951;
    assign temp2953 = temp2952 ^ temp2952;
    assign temp2954 = temp2953 ^ temp2953;
    assign temp2955 = temp2954 ^ temp2954;
    assign temp2956 = temp2955 ^ temp2955;
    assign temp2957 = temp2956 ^ temp2956;
    assign temp2958 = temp2957 ^ temp2957;
    assign temp2959 = temp2958 ^ temp2958;
    assign temp2960 = temp2959 ^ temp2959;
    assign temp2961 = temp2960 ^ temp2960;
    assign temp2962 = temp2961 ^ temp2961;
    assign temp2963 = temp2962 ^ temp2962;
    assign temp2964 = temp2963 ^ temp2963;
    assign temp2965 = temp2964 ^ temp2964;
    assign temp2966 = temp2965 ^ temp2965;
    assign temp2967 = temp2966 ^ temp2966;
    assign temp2968 = temp2967 ^ temp2967;
    assign temp2969 = temp2968 ^ temp2968;
    assign temp2970 = temp2969 ^ temp2969;
    assign temp2971 = temp2970 ^ temp2970;
    assign temp2972 = temp2971 ^ temp2971;
    assign temp2973 = temp2972 ^ temp2972;
    assign temp2974 = temp2973 ^ temp2973;
    assign temp2975 = temp2974 ^ temp2974;
    assign temp2976 = temp2975 ^ temp2975;
    assign temp2977 = temp2976 ^ temp2976;
    assign temp2978 = temp2977 ^ temp2977;
    assign temp2979 = temp2978 ^ temp2978;
    assign temp2980 = temp2979 ^ temp2979;
    assign temp2981 = temp2980 ^ temp2980;
    assign temp2982 = temp2981 ^ temp2981;
    assign temp2983 = temp2982 ^ temp2982;
    assign temp2984 = temp2983 ^ temp2983;
    assign temp2985 = temp2984 ^ temp2984;
    assign temp2986 = temp2985 ^ temp2985;
    assign temp2987 = temp2986 ^ temp2986;
    assign temp2988 = temp2987 ^ temp2987;
    assign temp2989 = temp2988 ^ temp2988;
    assign temp2990 = temp2989 ^ temp2989;
    assign temp2991 = temp2990 ^ temp2990;
    assign temp2992 = temp2991 ^ temp2991;
    assign temp2993 = temp2992 ^ temp2992;
    assign temp2994 = temp2993 ^ temp2993;
    assign temp2995 = temp2994 ^ temp2994;
    assign temp2996 = temp2995 ^ temp2995;
    assign temp2997 = temp2996 ^ temp2996;
    assign temp2998 = temp2997 ^ temp2997;
    assign temp2999 = temp2998 ^ temp2998;
    assign temp3000 = temp2999 ^ temp2999;
    assign temp3001 = temp3000 ^ temp3000;
    assign temp3002 = temp3001 ^ temp3001;
    assign temp3003 = temp3002 ^ temp3002;
    assign temp3004 = temp3003 ^ temp3003;
    assign temp3005 = temp3004 ^ temp3004;
    assign temp3006 = temp3005 ^ temp3005;
    assign temp3007 = temp3006 ^ temp3006;
    assign temp3008 = temp3007 ^ temp3007;
    assign temp3009 = temp3008 ^ temp3008;
    assign temp3010 = temp3009 ^ temp3009;
    assign temp3011 = temp3010 ^ temp3010;
    assign temp3012 = temp3011 ^ temp3011;
    assign temp3013 = temp3012 ^ temp3012;
    assign temp3014 = temp3013 ^ temp3013;
    assign temp3015 = temp3014 ^ temp3014;
    assign temp3016 = temp3015 ^ temp3015;
    assign temp3017 = temp3016 ^ temp3016;
    assign temp3018 = temp3017 ^ temp3017;
    assign temp3019 = temp3018 ^ temp3018;
    assign temp3020 = temp3019 ^ temp3019;
    assign temp3021 = temp3020 ^ temp3020;
    assign temp3022 = temp3021 ^ temp3021;
    assign temp3023 = temp3022 ^ temp3022;
    assign temp3024 = temp3023 ^ temp3023;
    assign temp3025 = temp3024 ^ temp3024;
    assign temp3026 = temp3025 ^ temp3025;
    assign temp3027 = temp3026 ^ temp3026;
    assign temp3028 = temp3027 ^ temp3027;
    assign temp3029 = temp3028 ^ temp3028;
    assign temp3030 = temp3029 ^ temp3029;
    assign temp3031 = temp3030 ^ temp3030;
    assign temp3032 = temp3031 ^ temp3031;
    assign temp3033 = temp3032 ^ temp3032;
    assign temp3034 = temp3033 ^ temp3033;
    assign temp3035 = temp3034 ^ temp3034;
    assign temp3036 = temp3035 ^ temp3035;
    assign temp3037 = temp3036 ^ temp3036;
    assign temp3038 = temp3037 ^ temp3037;
    assign temp3039 = temp3038 ^ temp3038;
    assign temp3040 = temp3039 ^ temp3039;
    assign temp3041 = temp3040 ^ temp3040;
    assign temp3042 = temp3041 ^ temp3041;
    assign temp3043 = temp3042 ^ temp3042;
    assign temp3044 = temp3043 ^ temp3043;
    assign temp3045 = temp3044 ^ temp3044;
    assign temp3046 = temp3045 ^ temp3045;
    assign temp3047 = temp3046 ^ temp3046;
    assign temp3048 = temp3047 ^ temp3047;
    assign temp3049 = temp3048 ^ temp3048;
    assign temp3050 = temp3049 ^ temp3049;
    assign temp3051 = temp3050 ^ temp3050;
    assign temp3052 = temp3051 ^ temp3051;
    assign temp3053 = temp3052 ^ temp3052;
    assign temp3054 = temp3053 ^ temp3053;
    assign temp3055 = temp3054 ^ temp3054;
    assign temp3056 = temp3055 ^ temp3055;
    assign temp3057 = temp3056 ^ temp3056;
    assign temp3058 = temp3057 ^ temp3057;
    assign temp3059 = temp3058 ^ temp3058;
    assign temp3060 = temp3059 ^ temp3059;
    assign temp3061 = temp3060 ^ temp3060;
    assign temp3062 = temp3061 ^ temp3061;
    assign temp3063 = temp3062 ^ temp3062;
    assign temp3064 = temp3063 ^ temp3063;
    assign temp3065 = temp3064 ^ temp3064;
    assign temp3066 = temp3065 ^ temp3065;
    assign temp3067 = temp3066 ^ temp3066;
    assign temp3068 = temp3067 ^ temp3067;
    assign temp3069 = temp3068 ^ temp3068;
    assign temp3070 = temp3069 ^ temp3069;
    assign temp3071 = temp3070 ^ temp3070;
    assign temp3072 = temp3071 ^ temp3071;
    assign temp3073 = temp3072 ^ temp3072;
    assign temp3074 = temp3073 ^ temp3073;
    assign temp3075 = temp3074 ^ temp3074;
    assign temp3076 = temp3075 ^ temp3075;
    assign temp3077 = temp3076 ^ temp3076;
    assign temp3078 = temp3077 ^ temp3077;
    assign temp3079 = temp3078 ^ temp3078;
    assign temp3080 = temp3079 ^ temp3079;
    assign temp3081 = temp3080 ^ temp3080;
    assign temp3082 = temp3081 ^ temp3081;
    assign temp3083 = temp3082 ^ temp3082;
    assign temp3084 = temp3083 ^ temp3083;
    assign temp3085 = temp3084 ^ temp3084;
    assign temp3086 = temp3085 ^ temp3085;
    assign temp3087 = temp3086 ^ temp3086;
    assign temp3088 = temp3087 ^ temp3087;
    assign temp3089 = temp3088 ^ temp3088;
    assign temp3090 = temp3089 ^ temp3089;
    assign temp3091 = temp3090 ^ temp3090;
    assign temp3092 = temp3091 ^ temp3091;
    assign temp3093 = temp3092 ^ temp3092;
    assign temp3094 = temp3093 ^ temp3093;
    assign temp3095 = temp3094 ^ temp3094;
    assign temp3096 = temp3095 ^ temp3095;
    assign temp3097 = temp3096 ^ temp3096;
    assign temp3098 = temp3097 ^ temp3097;
    assign temp3099 = temp3098 ^ temp3098;
    assign temp3100 = temp3099 ^ temp3099;
    assign temp3101 = temp3100 ^ temp3100;
    assign temp3102 = temp3101 ^ temp3101;
    assign temp3103 = temp3102 ^ temp3102;
    assign temp3104 = temp3103 ^ temp3103;
    assign temp3105 = temp3104 ^ temp3104;
    assign temp3106 = temp3105 ^ temp3105;
    assign temp3107 = temp3106 ^ temp3106;
    assign temp3108 = temp3107 ^ temp3107;
    assign temp3109 = temp3108 ^ temp3108;
    assign temp3110 = temp3109 ^ temp3109;
    assign temp3111 = temp3110 ^ temp3110;
    assign temp3112 = temp3111 ^ temp3111;
    assign temp3113 = temp3112 ^ temp3112;
    assign temp3114 = temp3113 ^ temp3113;
    assign temp3115 = temp3114 ^ temp3114;
    assign temp3116 = temp3115 ^ temp3115;
    assign temp3117 = temp3116 ^ temp3116;
    assign temp3118 = temp3117 ^ temp3117;
    assign temp3119 = temp3118 ^ temp3118;
    assign temp3120 = temp3119 ^ temp3119;
    assign temp3121 = temp3120 ^ temp3120;
    assign temp3122 = temp3121 ^ temp3121;
    assign temp3123 = temp3122 ^ temp3122;
    assign temp3124 = temp3123 ^ temp3123;
    assign temp3125 = temp3124 ^ temp3124;
    assign temp3126 = temp3125 ^ temp3125;
    assign temp3127 = temp3126 ^ temp3126;
    assign temp3128 = temp3127 ^ temp3127;
    assign temp3129 = temp3128 ^ temp3128;
    assign temp3130 = temp3129 ^ temp3129;
    assign temp3131 = temp3130 ^ temp3130;
    assign temp3132 = temp3131 ^ temp3131;
    assign temp3133 = temp3132 ^ temp3132;
    assign temp3134 = temp3133 ^ temp3133;
    assign temp3135 = temp3134 ^ temp3134;
    assign temp3136 = temp3135 ^ temp3135;
    assign temp3137 = temp3136 ^ temp3136;
    assign temp3138 = temp3137 ^ temp3137;
    assign temp3139 = temp3138 ^ temp3138;
    assign temp3140 = temp3139 ^ temp3139;
    assign temp3141 = temp3140 ^ temp3140;
    assign temp3142 = temp3141 ^ temp3141;
    assign temp3143 = temp3142 ^ temp3142;
    assign temp3144 = temp3143 ^ temp3143;
    assign temp3145 = temp3144 ^ temp3144;
    assign temp3146 = temp3145 ^ temp3145;
    assign temp3147 = temp3146 ^ temp3146;
    assign temp3148 = temp3147 ^ temp3147;
    assign temp3149 = temp3148 ^ temp3148;
    assign temp3150 = temp3149 ^ temp3149;
    assign temp3151 = temp3150 ^ temp3150;
    assign temp3152 = temp3151 ^ temp3151;
    assign temp3153 = temp3152 ^ temp3152;
    assign temp3154 = temp3153 ^ temp3153;
    assign temp3155 = temp3154 ^ temp3154;
    assign temp3156 = temp3155 ^ temp3155;
    assign temp3157 = temp3156 ^ temp3156;
    assign temp3158 = temp3157 ^ temp3157;
    assign temp3159 = temp3158 ^ temp3158;
    assign temp3160 = temp3159 ^ temp3159;
    assign temp3161 = temp3160 ^ temp3160;
    assign temp3162 = temp3161 ^ temp3161;
    assign temp3163 = temp3162 ^ temp3162;
    assign temp3164 = temp3163 ^ temp3163;
    assign temp3165 = temp3164 ^ temp3164;
    assign temp3166 = temp3165 ^ temp3165;
    assign temp3167 = temp3166 ^ temp3166;
    assign temp3168 = temp3167 ^ temp3167;
    assign temp3169 = temp3168 ^ temp3168;
    assign temp3170 = temp3169 ^ temp3169;
    assign temp3171 = temp3170 ^ temp3170;
    assign temp3172 = temp3171 ^ temp3171;
    assign temp3173 = temp3172 ^ temp3172;
    assign temp3174 = temp3173 ^ temp3173;
    assign temp3175 = temp3174 ^ temp3174;
    assign temp3176 = temp3175 ^ temp3175;
    assign temp3177 = temp3176 ^ temp3176;
    assign temp3178 = temp3177 ^ temp3177;
    assign temp3179 = temp3178 ^ temp3178;
    assign temp3180 = temp3179 ^ temp3179;
    assign temp3181 = temp3180 ^ temp3180;
    assign temp3182 = temp3181 ^ temp3181;
    assign temp3183 = temp3182 ^ temp3182;
    assign temp3184 = temp3183 ^ temp3183;
    assign temp3185 = temp3184 ^ temp3184;
    assign temp3186 = temp3185 ^ temp3185;
    assign temp3187 = temp3186 ^ temp3186;
    assign temp3188 = temp3187 ^ temp3187;
    assign temp3189 = temp3188 ^ temp3188;
    assign temp3190 = temp3189 ^ temp3189;
    assign temp3191 = temp3190 ^ temp3190;
    assign temp3192 = temp3191 ^ temp3191;
    assign temp3193 = temp3192 ^ temp3192;
    assign temp3194 = temp3193 ^ temp3193;
    assign temp3195 = temp3194 ^ temp3194;
    assign temp3196 = temp3195 ^ temp3195;
    assign temp3197 = temp3196 ^ temp3196;
    assign temp3198 = temp3197 ^ temp3197;
    assign temp3199 = temp3198 ^ temp3198;
    assign temp3200 = temp3199 ^ temp3199;
    assign temp3201 = temp3200 ^ temp3200;
    assign temp3202 = temp3201 ^ temp3201;
    assign temp3203 = temp3202 ^ temp3202;
    assign temp3204 = temp3203 ^ temp3203;
    assign temp3205 = temp3204 ^ temp3204;
    assign temp3206 = temp3205 ^ temp3205;
    assign temp3207 = temp3206 ^ temp3206;
    assign temp3208 = temp3207 ^ temp3207;
    assign temp3209 = temp3208 ^ temp3208;
    assign temp3210 = temp3209 ^ temp3209;
    assign temp3211 = temp3210 ^ temp3210;
    assign temp3212 = temp3211 ^ temp3211;
    assign temp3213 = temp3212 ^ temp3212;
    assign temp3214 = temp3213 ^ temp3213;
    assign temp3215 = temp3214 ^ temp3214;
    assign temp3216 = temp3215 ^ temp3215;
    assign temp3217 = temp3216 ^ temp3216;
    assign temp3218 = temp3217 ^ temp3217;
    assign temp3219 = temp3218 ^ temp3218;
    assign temp3220 = temp3219 ^ temp3219;
    assign temp3221 = temp3220 ^ temp3220;
    assign temp3222 = temp3221 ^ temp3221;
    assign temp3223 = temp3222 ^ temp3222;
    assign temp3224 = temp3223 ^ temp3223;
    assign temp3225 = temp3224 ^ temp3224;
    assign temp3226 = temp3225 ^ temp3225;
    assign temp3227 = temp3226 ^ temp3226;
    assign temp3228 = temp3227 ^ temp3227;
    assign temp3229 = temp3228 ^ temp3228;
    assign temp3230 = temp3229 ^ temp3229;
    assign temp3231 = temp3230 ^ temp3230;
    assign temp3232 = temp3231 ^ temp3231;
    assign temp3233 = temp3232 ^ temp3232;
    assign temp3234 = temp3233 ^ temp3233;
    assign temp3235 = temp3234 ^ temp3234;
    assign temp3236 = temp3235 ^ temp3235;
    assign temp3237 = temp3236 ^ temp3236;
    assign temp3238 = temp3237 ^ temp3237;
    assign temp3239 = temp3238 ^ temp3238;
    assign temp3240 = temp3239 ^ temp3239;
    assign temp3241 = temp3240 ^ temp3240;
    assign temp3242 = temp3241 ^ temp3241;
    assign temp3243 = temp3242 ^ temp3242;
    assign temp3244 = temp3243 ^ temp3243;
    assign temp3245 = temp3244 ^ temp3244;
    assign temp3246 = temp3245 ^ temp3245;
    assign temp3247 = temp3246 ^ temp3246;
    assign temp3248 = temp3247 ^ temp3247;
    assign temp3249 = temp3248 ^ temp3248;
    assign temp3250 = temp3249 ^ temp3249;
    assign temp3251 = temp3250 ^ temp3250;
    assign temp3252 = temp3251 ^ temp3251;
    assign temp3253 = temp3252 ^ temp3252;
    assign temp3254 = temp3253 ^ temp3253;
    assign temp3255 = temp3254 ^ temp3254;
    assign temp3256 = temp3255 ^ temp3255;
    assign temp3257 = temp3256 ^ temp3256;
    assign temp3258 = temp3257 ^ temp3257;
    assign temp3259 = temp3258 ^ temp3258;
    assign temp3260 = temp3259 ^ temp3259;
    assign temp3261 = temp3260 ^ temp3260;
    assign temp3262 = temp3261 ^ temp3261;
    assign temp3263 = temp3262 ^ temp3262;
    assign temp3264 = temp3263 ^ temp3263;
    assign temp3265 = temp3264 ^ temp3264;
    assign temp3266 = temp3265 ^ temp3265;
    assign temp3267 = temp3266 ^ temp3266;
    assign temp3268 = temp3267 ^ temp3267;
    assign temp3269 = temp3268 ^ temp3268;
    assign temp3270 = temp3269 ^ temp3269;
    assign temp3271 = temp3270 ^ temp3270;
    assign temp3272 = temp3271 ^ temp3271;
    assign temp3273 = temp3272 ^ temp3272;
    assign temp3274 = temp3273 ^ temp3273;
    assign temp3275 = temp3274 ^ temp3274;
    assign temp3276 = temp3275 ^ temp3275;
    assign temp3277 = temp3276 ^ temp3276;
    assign temp3278 = temp3277 ^ temp3277;
    assign temp3279 = temp3278 ^ temp3278;
    assign temp3280 = temp3279 ^ temp3279;
    assign temp3281 = temp3280 ^ temp3280;
    assign temp3282 = temp3281 ^ temp3281;
    assign temp3283 = temp3282 ^ temp3282;
    assign temp3284 = temp3283 ^ temp3283;
    assign temp3285 = temp3284 ^ temp3284;
    assign temp3286 = temp3285 ^ temp3285;
    assign temp3287 = temp3286 ^ temp3286;
    assign temp3288 = temp3287 ^ temp3287;
    assign temp3289 = temp3288 ^ temp3288;
    assign temp3290 = temp3289 ^ temp3289;
    assign temp3291 = temp3290 ^ temp3290;
    assign temp3292 = temp3291 ^ temp3291;
    assign temp3293 = temp3292 ^ temp3292;
    assign temp3294 = temp3293 ^ temp3293;
    assign temp3295 = temp3294 ^ temp3294;
    assign temp3296 = temp3295 ^ temp3295;
    assign temp3297 = temp3296 ^ temp3296;
    assign temp3298 = temp3297 ^ temp3297;
    assign temp3299 = temp3298 ^ temp3298;
    assign temp3300 = temp3299 ^ temp3299;
    assign temp3301 = temp3300 ^ temp3300;
    assign temp3302 = temp3301 ^ temp3301;
    assign temp3303 = temp3302 ^ temp3302;
    assign temp3304 = temp3303 ^ temp3303;
    assign temp3305 = temp3304 ^ temp3304;
    assign temp3306 = temp3305 ^ temp3305;
    assign temp3307 = temp3306 ^ temp3306;
    assign temp3308 = temp3307 ^ temp3307;
    assign temp3309 = temp3308 ^ temp3308;
    assign temp3310 = temp3309 ^ temp3309;
    assign temp3311 = temp3310 ^ temp3310;
    assign temp3312 = temp3311 ^ temp3311;
    assign temp3313 = temp3312 ^ temp3312;
    assign temp3314 = temp3313 ^ temp3313;
    assign temp3315 = temp3314 ^ temp3314;
    assign temp3316 = temp3315 ^ temp3315;
    assign temp3317 = temp3316 ^ temp3316;
    assign temp3318 = temp3317 ^ temp3317;
    assign temp3319 = temp3318 ^ temp3318;
    assign temp3320 = temp3319 ^ temp3319;
    assign temp3321 = temp3320 ^ temp3320;
    assign temp3322 = temp3321 ^ temp3321;
    assign temp3323 = temp3322 ^ temp3322;
    assign temp3324 = temp3323 ^ temp3323;
    assign temp3325 = temp3324 ^ temp3324;
    assign temp3326 = temp3325 ^ temp3325;
    assign temp3327 = temp3326 ^ temp3326;
    assign temp3328 = temp3327 ^ temp3327;
    assign temp3329 = temp3328 ^ temp3328;
    assign temp3330 = temp3329 ^ temp3329;
    assign temp3331 = temp3330 ^ temp3330;
    assign temp3332 = temp3331 ^ temp3331;
    assign temp3333 = temp3332 ^ temp3332;
    assign temp3334 = temp3333 ^ temp3333;
    assign temp3335 = temp3334 ^ temp3334;
    assign temp3336 = temp3335 ^ temp3335;
    assign temp3337 = temp3336 ^ temp3336;
    assign temp3338 = temp3337 ^ temp3337;
    assign temp3339 = temp3338 ^ temp3338;
    assign temp3340 = temp3339 ^ temp3339;
    assign temp3341 = temp3340 ^ temp3340;
    assign temp3342 = temp3341 ^ temp3341;
    assign temp3343 = temp3342 ^ temp3342;
    assign temp3344 = temp3343 ^ temp3343;
    assign temp3345 = temp3344 ^ temp3344;
    assign temp3346 = temp3345 ^ temp3345;
    assign temp3347 = temp3346 ^ temp3346;
    assign temp3348 = temp3347 ^ temp3347;
    assign temp3349 = temp3348 ^ temp3348;
    assign temp3350 = temp3349 ^ temp3349;
    assign temp3351 = temp3350 ^ temp3350;
    assign temp3352 = temp3351 ^ temp3351;
    assign temp3353 = temp3352 ^ temp3352;
    assign temp3354 = temp3353 ^ temp3353;
    assign temp3355 = temp3354 ^ temp3354;
    assign temp3356 = temp3355 ^ temp3355;
    assign temp3357 = temp3356 ^ temp3356;
    assign temp3358 = temp3357 ^ temp3357;
    assign temp3359 = temp3358 ^ temp3358;
    assign temp3360 = temp3359 ^ temp3359;
    assign temp3361 = temp3360 ^ temp3360;
    assign temp3362 = temp3361 ^ temp3361;
    assign temp3363 = temp3362 ^ temp3362;
    assign temp3364 = temp3363 ^ temp3363;
    assign temp3365 = temp3364 ^ temp3364;
    assign temp3366 = temp3365 ^ temp3365;
    assign temp3367 = temp3366 ^ temp3366;
    assign temp3368 = temp3367 ^ temp3367;
    assign temp3369 = temp3368 ^ temp3368;
    assign temp3370 = temp3369 ^ temp3369;
    assign temp3371 = temp3370 ^ temp3370;
    assign temp3372 = temp3371 ^ temp3371;
    assign temp3373 = temp3372 ^ temp3372;
    assign temp3374 = temp3373 ^ temp3373;
    assign temp3375 = temp3374 ^ temp3374;
    assign temp3376 = temp3375 ^ temp3375;
    assign temp3377 = temp3376 ^ temp3376;
    assign temp3378 = temp3377 ^ temp3377;
    assign temp3379 = temp3378 ^ temp3378;
    assign temp3380 = temp3379 ^ temp3379;
    assign temp3381 = temp3380 ^ temp3380;
    assign temp3382 = temp3381 ^ temp3381;
    assign temp3383 = temp3382 ^ temp3382;
    assign temp3384 = temp3383 ^ temp3383;
    assign temp3385 = temp3384 ^ temp3384;
    assign temp3386 = temp3385 ^ temp3385;
    assign temp3387 = temp3386 ^ temp3386;
    assign temp3388 = temp3387 ^ temp3387;
    assign temp3389 = temp3388 ^ temp3388;
    assign temp3390 = temp3389 ^ temp3389;
    assign temp3391 = temp3390 ^ temp3390;
    assign temp3392 = temp3391 ^ temp3391;
    assign temp3393 = temp3392 ^ temp3392;
    assign temp3394 = temp3393 ^ temp3393;
    assign temp3395 = temp3394 ^ temp3394;
    assign temp3396 = temp3395 ^ temp3395;
    assign temp3397 = temp3396 ^ temp3396;
    assign temp3398 = temp3397 ^ temp3397;
    assign temp3399 = temp3398 ^ temp3398;
    assign temp3400 = temp3399 ^ temp3399;
    assign temp3401 = temp3400 ^ temp3400;
    assign temp3402 = temp3401 ^ temp3401;
    assign temp3403 = temp3402 ^ temp3402;
    assign temp3404 = temp3403 ^ temp3403;
    assign temp3405 = temp3404 ^ temp3404;
    assign temp3406 = temp3405 ^ temp3405;
    assign temp3407 = temp3406 ^ temp3406;
    assign temp3408 = temp3407 ^ temp3407;
    assign temp3409 = temp3408 ^ temp3408;
    assign temp3410 = temp3409 ^ temp3409;
    assign temp3411 = temp3410 ^ temp3410;
    assign temp3412 = temp3411 ^ temp3411;
    assign temp3413 = temp3412 ^ temp3412;
    assign temp3414 = temp3413 ^ temp3413;
    assign temp3415 = temp3414 ^ temp3414;
    assign temp3416 = temp3415 ^ temp3415;
    assign temp3417 = temp3416 ^ temp3416;
    assign temp3418 = temp3417 ^ temp3417;
    assign temp3419 = temp3418 ^ temp3418;
    assign temp3420 = temp3419 ^ temp3419;
    assign temp3421 = temp3420 ^ temp3420;
    assign temp3422 = temp3421 ^ temp3421;
    assign temp3423 = temp3422 ^ temp3422;
    assign temp3424 = temp3423 ^ temp3423;
    assign temp3425 = temp3424 ^ temp3424;
    assign temp3426 = temp3425 ^ temp3425;
    assign temp3427 = temp3426 ^ temp3426;
    assign temp3428 = temp3427 ^ temp3427;
    assign temp3429 = temp3428 ^ temp3428;
    assign temp3430 = temp3429 ^ temp3429;
    assign temp3431 = temp3430 ^ temp3430;
    assign temp3432 = temp3431 ^ temp3431;
    assign temp3433 = temp3432 ^ temp3432;
    assign temp3434 = temp3433 ^ temp3433;
    assign temp3435 = temp3434 ^ temp3434;
    assign temp3436 = temp3435 ^ temp3435;
    assign temp3437 = temp3436 ^ temp3436;
    assign temp3438 = temp3437 ^ temp3437;
    assign temp3439 = temp3438 ^ temp3438;
    assign temp3440 = temp3439 ^ temp3439;
    assign temp3441 = temp3440 ^ temp3440;
    assign temp3442 = temp3441 ^ temp3441;
    assign temp3443 = temp3442 ^ temp3442;
    assign temp3444 = temp3443 ^ temp3443;
    assign temp3445 = temp3444 ^ temp3444;
    assign temp3446 = temp3445 ^ temp3445;
    assign temp3447 = temp3446 ^ temp3446;
    assign temp3448 = temp3447 ^ temp3447;
    assign temp3449 = temp3448 ^ temp3448;
    assign temp3450 = temp3449 ^ temp3449;
    assign temp3451 = temp3450 ^ temp3450;
    assign temp3452 = temp3451 ^ temp3451;
    assign temp3453 = temp3452 ^ temp3452;
    assign temp3454 = temp3453 ^ temp3453;
    assign temp3455 = temp3454 ^ temp3454;
    assign temp3456 = temp3455 ^ temp3455;
    assign temp3457 = temp3456 ^ temp3456;
    assign temp3458 = temp3457 ^ temp3457;
    assign temp3459 = temp3458 ^ temp3458;
    assign temp3460 = temp3459 ^ temp3459;
    assign temp3461 = temp3460 ^ temp3460;
    assign temp3462 = temp3461 ^ temp3461;
    assign temp3463 = temp3462 ^ temp3462;
    assign temp3464 = temp3463 ^ temp3463;
    assign temp3465 = temp3464 ^ temp3464;
    assign temp3466 = temp3465 ^ temp3465;
    assign temp3467 = temp3466 ^ temp3466;
    assign temp3468 = temp3467 ^ temp3467;
    assign temp3469 = temp3468 ^ temp3468;
    assign temp3470 = temp3469 ^ temp3469;
    assign temp3471 = temp3470 ^ temp3470;
    assign temp3472 = temp3471 ^ temp3471;
    assign temp3473 = temp3472 ^ temp3472;
    assign temp3474 = temp3473 ^ temp3473;
    assign temp3475 = temp3474 ^ temp3474;
    assign temp3476 = temp3475 ^ temp3475;
    assign temp3477 = temp3476 ^ temp3476;
    assign temp3478 = temp3477 ^ temp3477;
    assign temp3479 = temp3478 ^ temp3478;
    assign temp3480 = temp3479 ^ temp3479;
    assign temp3481 = temp3480 ^ temp3480;
    assign temp3482 = temp3481 ^ temp3481;
    assign temp3483 = temp3482 ^ temp3482;
    assign temp3484 = temp3483 ^ temp3483;
    assign temp3485 = temp3484 ^ temp3484;
    assign temp3486 = temp3485 ^ temp3485;
    assign temp3487 = temp3486 ^ temp3486;
    assign temp3488 = temp3487 ^ temp3487;
    assign temp3489 = temp3488 ^ temp3488;
    assign temp3490 = temp3489 ^ temp3489;
    assign temp3491 = temp3490 ^ temp3490;
    assign temp3492 = temp3491 ^ temp3491;
    assign temp3493 = temp3492 ^ temp3492;
    assign temp3494 = temp3493 ^ temp3493;
    assign temp3495 = temp3494 ^ temp3494;
    assign temp3496 = temp3495 ^ temp3495;
    assign temp3497 = temp3496 ^ temp3496;
    assign temp3498 = temp3497 ^ temp3497;
    assign temp3499 = temp3498 ^ temp3498;
    assign temp3500 = temp3499 ^ temp3499;
    assign temp3501 = temp3500 ^ temp3500;
    assign temp3502 = temp3501 ^ temp3501;
    assign temp3503 = temp3502 ^ temp3502;
    assign temp3504 = temp3503 ^ temp3503;
    assign temp3505 = temp3504 ^ temp3504;
    assign temp3506 = temp3505 ^ temp3505;
    assign temp3507 = temp3506 ^ temp3506;
    assign temp3508 = temp3507 ^ temp3507;
    assign temp3509 = temp3508 ^ temp3508;
    assign temp3510 = temp3509 ^ temp3509;
    assign temp3511 = temp3510 ^ temp3510;
    assign temp3512 = temp3511 ^ temp3511;
    assign temp3513 = temp3512 ^ temp3512;
    assign temp3514 = temp3513 ^ temp3513;
    assign temp3515 = temp3514 ^ temp3514;
    assign temp3516 = temp3515 ^ temp3515;
    assign temp3517 = temp3516 ^ temp3516;
    assign temp3518 = temp3517 ^ temp3517;
    assign temp3519 = temp3518 ^ temp3518;
    assign temp3520 = temp3519 ^ temp3519;
    assign temp3521 = temp3520 ^ temp3520;
    assign temp3522 = temp3521 ^ temp3521;
    assign temp3523 = temp3522 ^ temp3522;
    assign temp3524 = temp3523 ^ temp3523;
    assign temp3525 = temp3524 ^ temp3524;
    assign temp3526 = temp3525 ^ temp3525;
    assign temp3527 = temp3526 ^ temp3526;
    assign temp3528 = temp3527 ^ temp3527;
    assign temp3529 = temp3528 ^ temp3528;
    assign temp3530 = temp3529 ^ temp3529;
    assign temp3531 = temp3530 ^ temp3530;
    assign temp3532 = temp3531 ^ temp3531;
    assign temp3533 = temp3532 ^ temp3532;
    assign temp3534 = temp3533 ^ temp3533;
    assign temp3535 = temp3534 ^ temp3534;
    assign temp3536 = temp3535 ^ temp3535;
    assign temp3537 = temp3536 ^ temp3536;
    assign temp3538 = temp3537 ^ temp3537;
    assign temp3539 = temp3538 ^ temp3538;
    assign temp3540 = temp3539 ^ temp3539;
    assign temp3541 = temp3540 ^ temp3540;
    assign temp3542 = temp3541 ^ temp3541;
    assign temp3543 = temp3542 ^ temp3542;
    assign temp3544 = temp3543 ^ temp3543;
    assign temp3545 = temp3544 ^ temp3544;
    assign temp3546 = temp3545 ^ temp3545;
    assign temp3547 = temp3546 ^ temp3546;
    assign temp3548 = temp3547 ^ temp3547;
    assign temp3549 = temp3548 ^ temp3548;
    assign temp3550 = temp3549 ^ temp3549;
    assign temp3551 = temp3550 ^ temp3550;
    assign temp3552 = temp3551 ^ temp3551;
    assign temp3553 = temp3552 ^ temp3552;
    assign temp3554 = temp3553 ^ temp3553;
    assign temp3555 = temp3554 ^ temp3554;
    assign temp3556 = temp3555 ^ temp3555;
    assign temp3557 = temp3556 ^ temp3556;
    assign temp3558 = temp3557 ^ temp3557;
    assign temp3559 = temp3558 ^ temp3558;
    assign temp3560 = temp3559 ^ temp3559;
    assign temp3561 = temp3560 ^ temp3560;
    assign temp3562 = temp3561 ^ temp3561;
    assign temp3563 = temp3562 ^ temp3562;
    assign temp3564 = temp3563 ^ temp3563;
    assign temp3565 = temp3564 ^ temp3564;
    assign temp3566 = temp3565 ^ temp3565;
    assign temp3567 = temp3566 ^ temp3566;
    assign temp3568 = temp3567 ^ temp3567;
    assign temp3569 = temp3568 ^ temp3568;
    assign temp3570 = temp3569 ^ temp3569;
    assign temp3571 = temp3570 ^ temp3570;
    assign temp3572 = temp3571 ^ temp3571;
    assign temp3573 = temp3572 ^ temp3572;
    assign temp3574 = temp3573 ^ temp3573;
    assign temp3575 = temp3574 ^ temp3574;
    assign temp3576 = temp3575 ^ temp3575;
    assign temp3577 = temp3576 ^ temp3576;
    assign temp3578 = temp3577 ^ temp3577;
    assign temp3579 = temp3578 ^ temp3578;
    assign temp3580 = temp3579 ^ temp3579;
    assign temp3581 = temp3580 ^ temp3580;
    assign temp3582 = temp3581 ^ temp3581;
    assign temp3583 = temp3582 ^ temp3582;
    assign temp3584 = temp3583 ^ temp3583;
    assign temp3585 = temp3584 ^ temp3584;
    assign temp3586 = temp3585 ^ temp3585;
    assign temp3587 = temp3586 ^ temp3586;
    assign temp3588 = temp3587 ^ temp3587;
    assign temp3589 = temp3588 ^ temp3588;
    assign temp3590 = temp3589 ^ temp3589;
    assign temp3591 = temp3590 ^ temp3590;
    assign temp3592 = temp3591 ^ temp3591;
    assign temp3593 = temp3592 ^ temp3592;
    assign temp3594 = temp3593 ^ temp3593;
    assign temp3595 = temp3594 ^ temp3594;
    assign temp3596 = temp3595 ^ temp3595;
    assign temp3597 = temp3596 ^ temp3596;
    assign temp3598 = temp3597 ^ temp3597;
    assign temp3599 = temp3598 ^ temp3598;
    assign temp3600 = temp3599 ^ temp3599;
    assign temp3601 = temp3600 ^ temp3600;
    assign temp3602 = temp3601 ^ temp3601;
    assign temp3603 = temp3602 ^ temp3602;
    assign temp3604 = temp3603 ^ temp3603;
    assign temp3605 = temp3604 ^ temp3604;
    assign temp3606 = temp3605 ^ temp3605;
    assign temp3607 = temp3606 ^ temp3606;
    assign temp3608 = temp3607 ^ temp3607;
    assign temp3609 = temp3608 ^ temp3608;
    assign temp3610 = temp3609 ^ temp3609;
    assign temp3611 = temp3610 ^ temp3610;
    assign temp3612 = temp3611 ^ temp3611;
    assign temp3613 = temp3612 ^ temp3612;
    assign temp3614 = temp3613 ^ temp3613;
    assign temp3615 = temp3614 ^ temp3614;
    assign temp3616 = temp3615 ^ temp3615;
    assign temp3617 = temp3616 ^ temp3616;
    assign temp3618 = temp3617 ^ temp3617;
    assign temp3619 = temp3618 ^ temp3618;
    assign temp3620 = temp3619 ^ temp3619;
    assign temp3621 = temp3620 ^ temp3620;
    assign temp3622 = temp3621 ^ temp3621;
    assign temp3623 = temp3622 ^ temp3622;
    assign temp3624 = temp3623 ^ temp3623;
    assign temp3625 = temp3624 ^ temp3624;
    assign temp3626 = temp3625 ^ temp3625;
    assign temp3627 = temp3626 ^ temp3626;
    assign temp3628 = temp3627 ^ temp3627;
    assign temp3629 = temp3628 ^ temp3628;
    assign temp3630 = temp3629 ^ temp3629;
    assign temp3631 = temp3630 ^ temp3630;
    assign temp3632 = temp3631 ^ temp3631;
    assign temp3633 = temp3632 ^ temp3632;
    assign temp3634 = temp3633 ^ temp3633;
    assign temp3635 = temp3634 ^ temp3634;
    assign temp3636 = temp3635 ^ temp3635;
    assign temp3637 = temp3636 ^ temp3636;
    assign temp3638 = temp3637 ^ temp3637;
    assign temp3639 = temp3638 ^ temp3638;
    assign temp3640 = temp3639 ^ temp3639;
    assign temp3641 = temp3640 ^ temp3640;
    assign temp3642 = temp3641 ^ temp3641;
    assign temp3643 = temp3642 ^ temp3642;
    assign temp3644 = temp3643 ^ temp3643;
    assign temp3645 = temp3644 ^ temp3644;
    assign temp3646 = temp3645 ^ temp3645;
    assign temp3647 = temp3646 ^ temp3646;
    assign temp3648 = temp3647 ^ temp3647;
    assign temp3649 = temp3648 ^ temp3648;
    assign temp3650 = temp3649 ^ temp3649;
    assign temp3651 = temp3650 ^ temp3650;
    assign temp3652 = temp3651 ^ temp3651;
    assign temp3653 = temp3652 ^ temp3652;
    assign temp3654 = temp3653 ^ temp3653;
    assign temp3655 = temp3654 ^ temp3654;
    assign temp3656 = temp3655 ^ temp3655;
    assign temp3657 = temp3656 ^ temp3656;
    assign temp3658 = temp3657 ^ temp3657;
    assign temp3659 = temp3658 ^ temp3658;
    assign temp3660 = temp3659 ^ temp3659;
    assign temp3661 = temp3660 ^ temp3660;
    assign temp3662 = temp3661 ^ temp3661;
    assign temp3663 = temp3662 ^ temp3662;
    assign temp3664 = temp3663 ^ temp3663;
    assign temp3665 = temp3664 ^ temp3664;
    assign temp3666 = temp3665 ^ temp3665;
    assign temp3667 = temp3666 ^ temp3666;
    assign temp3668 = temp3667 ^ temp3667;
    assign temp3669 = temp3668 ^ temp3668;
    assign temp3670 = temp3669 ^ temp3669;
    assign temp3671 = temp3670 ^ temp3670;
    assign temp3672 = temp3671 ^ temp3671;
    assign temp3673 = temp3672 ^ temp3672;
    assign temp3674 = temp3673 ^ temp3673;
    assign temp3675 = temp3674 ^ temp3674;
    assign temp3676 = temp3675 ^ temp3675;
    assign temp3677 = temp3676 ^ temp3676;
    assign temp3678 = temp3677 ^ temp3677;
    assign temp3679 = temp3678 ^ temp3678;
    assign temp3680 = temp3679 ^ temp3679;
    assign temp3681 = temp3680 ^ temp3680;
    assign temp3682 = temp3681 ^ temp3681;
    assign temp3683 = temp3682 ^ temp3682;
    assign temp3684 = temp3683 ^ temp3683;
    assign temp3685 = temp3684 ^ temp3684;
    assign temp3686 = temp3685 ^ temp3685;
    assign temp3687 = temp3686 ^ temp3686;
    assign temp3688 = temp3687 ^ temp3687;
    assign temp3689 = temp3688 ^ temp3688;
    assign temp3690 = temp3689 ^ temp3689;
    assign temp3691 = temp3690 ^ temp3690;
    assign temp3692 = temp3691 ^ temp3691;
    assign temp3693 = temp3692 ^ temp3692;
    assign temp3694 = temp3693 ^ temp3693;
    assign temp3695 = temp3694 ^ temp3694;
    assign temp3696 = temp3695 ^ temp3695;
    assign temp3697 = temp3696 ^ temp3696;
    assign temp3698 = temp3697 ^ temp3697;
    assign temp3699 = temp3698 ^ temp3698;
    assign temp3700 = temp3699 ^ temp3699;
    assign temp3701 = temp3700 ^ temp3700;
    assign temp3702 = temp3701 ^ temp3701;
    assign temp3703 = temp3702 ^ temp3702;
    assign temp3704 = temp3703 ^ temp3703;
    assign temp3705 = temp3704 ^ temp3704;
    assign temp3706 = temp3705 ^ temp3705;
    assign temp3707 = temp3706 ^ temp3706;
    assign temp3708 = temp3707 ^ temp3707;
    assign temp3709 = temp3708 ^ temp3708;
    assign temp3710 = temp3709 ^ temp3709;
    assign temp3711 = temp3710 ^ temp3710;
    assign temp3712 = temp3711 ^ temp3711;
    assign temp3713 = temp3712 ^ temp3712;
    assign temp3714 = temp3713 ^ temp3713;
    assign temp3715 = temp3714 ^ temp3714;
    assign temp3716 = temp3715 ^ temp3715;
    assign temp3717 = temp3716 ^ temp3716;
    assign temp3718 = temp3717 ^ temp3717;
    assign temp3719 = temp3718 ^ temp3718;
    assign temp3720 = temp3719 ^ temp3719;
    assign temp3721 = temp3720 ^ temp3720;
    assign temp3722 = temp3721 ^ temp3721;
    assign temp3723 = temp3722 ^ temp3722;
    assign temp3724 = temp3723 ^ temp3723;
    assign temp3725 = temp3724 ^ temp3724;
    assign temp3726 = temp3725 ^ temp3725;
    assign temp3727 = temp3726 ^ temp3726;
    assign temp3728 = temp3727 ^ temp3727;
    assign temp3729 = temp3728 ^ temp3728;
    assign temp3730 = temp3729 ^ temp3729;
    assign temp3731 = temp3730 ^ temp3730;
    assign temp3732 = temp3731 ^ temp3731;
    assign temp3733 = temp3732 ^ temp3732;
    assign temp3734 = temp3733 ^ temp3733;
    assign temp3735 = temp3734 ^ temp3734;
    assign temp3736 = temp3735 ^ temp3735;
    assign temp3737 = temp3736 ^ temp3736;
    assign temp3738 = temp3737 ^ temp3737;
    assign temp3739 = temp3738 ^ temp3738;
    assign temp3740 = temp3739 ^ temp3739;
    assign temp3741 = temp3740 ^ temp3740;
    assign temp3742 = temp3741 ^ temp3741;
    assign temp3743 = temp3742 ^ temp3742;
    assign temp3744 = temp3743 ^ temp3743;
    assign temp3745 = temp3744 ^ temp3744;
    assign temp3746 = temp3745 ^ temp3745;
    assign temp3747 = temp3746 ^ temp3746;
    assign temp3748 = temp3747 ^ temp3747;
    assign temp3749 = temp3748 ^ temp3748;
    assign temp3750 = temp3749 ^ temp3749;
    assign temp3751 = temp3750 ^ temp3750;
    assign temp3752 = temp3751 ^ temp3751;
    assign temp3753 = temp3752 ^ temp3752;
    assign temp3754 = temp3753 ^ temp3753;
    assign temp3755 = temp3754 ^ temp3754;
    assign temp3756 = temp3755 ^ temp3755;
    assign temp3757 = temp3756 ^ temp3756;
    assign temp3758 = temp3757 ^ temp3757;
    assign temp3759 = temp3758 ^ temp3758;
    assign temp3760 = temp3759 ^ temp3759;
    assign temp3761 = temp3760 ^ temp3760;
    assign temp3762 = temp3761 ^ temp3761;
    assign temp3763 = temp3762 ^ temp3762;
    assign temp3764 = temp3763 ^ temp3763;
    assign temp3765 = temp3764 ^ temp3764;
    assign temp3766 = temp3765 ^ temp3765;
    assign temp3767 = temp3766 ^ temp3766;
    assign temp3768 = temp3767 ^ temp3767;
    assign temp3769 = temp3768 ^ temp3768;
    assign temp3770 = temp3769 ^ temp3769;
    assign temp3771 = temp3770 ^ temp3770;
    assign temp3772 = temp3771 ^ temp3771;
    assign temp3773 = temp3772 ^ temp3772;
    assign temp3774 = temp3773 ^ temp3773;
    assign temp3775 = temp3774 ^ temp3774;
    assign temp3776 = temp3775 ^ temp3775;
    assign temp3777 = temp3776 ^ temp3776;
    assign temp3778 = temp3777 ^ temp3777;
    assign temp3779 = temp3778 ^ temp3778;
    assign temp3780 = temp3779 ^ temp3779;
    assign temp3781 = temp3780 ^ temp3780;
    assign temp3782 = temp3781 ^ temp3781;
    assign temp3783 = temp3782 ^ temp3782;
    assign temp3784 = temp3783 ^ temp3783;
    assign temp3785 = temp3784 ^ temp3784;
    assign temp3786 = temp3785 ^ temp3785;
    assign temp3787 = temp3786 ^ temp3786;
    assign temp3788 = temp3787 ^ temp3787;
    assign temp3789 = temp3788 ^ temp3788;
    assign temp3790 = temp3789 ^ temp3789;
    assign temp3791 = temp3790 ^ temp3790;
    assign temp3792 = temp3791 ^ temp3791;
    assign temp3793 = temp3792 ^ temp3792;
    assign temp3794 = temp3793 ^ temp3793;
    assign temp3795 = temp3794 ^ temp3794;
    assign temp3796 = temp3795 ^ temp3795;
    assign temp3797 = temp3796 ^ temp3796;
    assign temp3798 = temp3797 ^ temp3797;
    assign temp3799 = temp3798 ^ temp3798;
    assign temp3800 = temp3799 ^ temp3799;
    assign temp3801 = temp3800 ^ temp3800;
    assign temp3802 = temp3801 ^ temp3801;
    assign temp3803 = temp3802 ^ temp3802;
    assign temp3804 = temp3803 ^ temp3803;
    assign temp3805 = temp3804 ^ temp3804;
    assign temp3806 = temp3805 ^ temp3805;
    assign temp3807 = temp3806 ^ temp3806;
    assign temp3808 = temp3807 ^ temp3807;
    assign temp3809 = temp3808 ^ temp3808;
    assign temp3810 = temp3809 ^ temp3809;
    assign temp3811 = temp3810 ^ temp3810;
    assign temp3812 = temp3811 ^ temp3811;
    assign temp3813 = temp3812 ^ temp3812;
    assign temp3814 = temp3813 ^ temp3813;
    assign temp3815 = temp3814 ^ temp3814;
    assign temp3816 = temp3815 ^ temp3815;
    assign temp3817 = temp3816 ^ temp3816;
    assign temp3818 = temp3817 ^ temp3817;
    assign temp3819 = temp3818 ^ temp3818;
    assign temp3820 = temp3819 ^ temp3819;
    assign temp3821 = temp3820 ^ temp3820;
    assign temp3822 = temp3821 ^ temp3821;
    assign temp3823 = temp3822 ^ temp3822;
    assign temp3824 = temp3823 ^ temp3823;
    assign temp3825 = temp3824 ^ temp3824;
    assign temp3826 = temp3825 ^ temp3825;
    assign temp3827 = temp3826 ^ temp3826;
    assign temp3828 = temp3827 ^ temp3827;
    assign temp3829 = temp3828 ^ temp3828;
    assign temp3830 = temp3829 ^ temp3829;
    assign temp3831 = temp3830 ^ temp3830;
    assign temp3832 = temp3831 ^ temp3831;
    assign temp3833 = temp3832 ^ temp3832;
    assign temp3834 = temp3833 ^ temp3833;
    assign temp3835 = temp3834 ^ temp3834;
    assign temp3836 = temp3835 ^ temp3835;
    assign temp3837 = temp3836 ^ temp3836;
    assign temp3838 = temp3837 ^ temp3837;
    assign temp3839 = temp3838 ^ temp3838;
    assign temp3840 = temp3839 ^ temp3839;
    assign temp3841 = temp3840 ^ temp3840;
    assign temp3842 = temp3841 ^ temp3841;
    assign temp3843 = temp3842 ^ temp3842;
    assign temp3844 = temp3843 ^ temp3843;
    assign temp3845 = temp3844 ^ temp3844;
    assign temp3846 = temp3845 ^ temp3845;
    assign temp3847 = temp3846 ^ temp3846;
    assign temp3848 = temp3847 ^ temp3847;
    assign temp3849 = temp3848 ^ temp3848;
    assign temp3850 = temp3849 ^ temp3849;
    assign temp3851 = temp3850 ^ temp3850;
    assign temp3852 = temp3851 ^ temp3851;
    assign temp3853 = temp3852 ^ temp3852;
    assign temp3854 = temp3853 ^ temp3853;
    assign temp3855 = temp3854 ^ temp3854;
    assign temp3856 = temp3855 ^ temp3855;
    assign temp3857 = temp3856 ^ temp3856;
    assign temp3858 = temp3857 ^ temp3857;
    assign temp3859 = temp3858 ^ temp3858;
    assign temp3860 = temp3859 ^ temp3859;
    assign temp3861 = temp3860 ^ temp3860;
    assign temp3862 = temp3861 ^ temp3861;
    assign temp3863 = temp3862 ^ temp3862;
    assign temp3864 = temp3863 ^ temp3863;
    assign temp3865 = temp3864 ^ temp3864;
    assign temp3866 = temp3865 ^ temp3865;
    assign temp3867 = temp3866 ^ temp3866;
    assign temp3868 = temp3867 ^ temp3867;
    assign temp3869 = temp3868 ^ temp3868;
    assign temp3870 = temp3869 ^ temp3869;
    assign temp3871 = temp3870 ^ temp3870;
    assign temp3872 = temp3871 ^ temp3871;
    assign temp3873 = temp3872 ^ temp3872;
    assign temp3874 = temp3873 ^ temp3873;
    assign temp3875 = temp3874 ^ temp3874;
    assign temp3876 = temp3875 ^ temp3875;
    assign temp3877 = temp3876 ^ temp3876;
    assign temp3878 = temp3877 ^ temp3877;
    assign temp3879 = temp3878 ^ temp3878;
    assign temp3880 = temp3879 ^ temp3879;
    assign temp3881 = temp3880 ^ temp3880;
    assign temp3882 = temp3881 ^ temp3881;
    assign temp3883 = temp3882 ^ temp3882;
    assign temp3884 = temp3883 ^ temp3883;
    assign temp3885 = temp3884 ^ temp3884;
    assign temp3886 = temp3885 ^ temp3885;
    assign temp3887 = temp3886 ^ temp3886;
    assign temp3888 = temp3887 ^ temp3887;
    assign temp3889 = temp3888 ^ temp3888;
    assign temp3890 = temp3889 ^ temp3889;
    assign temp3891 = temp3890 ^ temp3890;
    assign temp3892 = temp3891 ^ temp3891;
    assign temp3893 = temp3892 ^ temp3892;
    assign temp3894 = temp3893 ^ temp3893;
    assign temp3895 = temp3894 ^ temp3894;
    assign temp3896 = temp3895 ^ temp3895;
    assign temp3897 = temp3896 ^ temp3896;
    assign temp3898 = temp3897 ^ temp3897;
    assign temp3899 = temp3898 ^ temp3898;
    assign temp3900 = temp3899 ^ temp3899;
    assign temp3901 = temp3900 ^ temp3900;
    assign temp3902 = temp3901 ^ temp3901;
    assign temp3903 = temp3902 ^ temp3902;
    assign temp3904 = temp3903 ^ temp3903;
    assign temp3905 = temp3904 ^ temp3904;
    assign temp3906 = temp3905 ^ temp3905;
    assign temp3907 = temp3906 ^ temp3906;
    assign temp3908 = temp3907 ^ temp3907;
    assign temp3909 = temp3908 ^ temp3908;
    assign temp3910 = temp3909 ^ temp3909;
    assign temp3911 = temp3910 ^ temp3910;
    assign temp3912 = temp3911 ^ temp3911;
    assign temp3913 = temp3912 ^ temp3912;
    assign temp3914 = temp3913 ^ temp3913;
    assign temp3915 = temp3914 ^ temp3914;
    assign temp3916 = temp3915 ^ temp3915;
    assign temp3917 = temp3916 ^ temp3916;
    assign temp3918 = temp3917 ^ temp3917;
    assign temp3919 = temp3918 ^ temp3918;
    assign temp3920 = temp3919 ^ temp3919;
    assign temp3921 = temp3920 ^ temp3920;
    assign temp3922 = temp3921 ^ temp3921;
    assign temp3923 = temp3922 ^ temp3922;
    assign temp3924 = temp3923 ^ temp3923;
    assign temp3925 = temp3924 ^ temp3924;
    assign temp3926 = temp3925 ^ temp3925;
    assign temp3927 = temp3926 ^ temp3926;
    assign temp3928 = temp3927 ^ temp3927;
    assign temp3929 = temp3928 ^ temp3928;
    assign temp3930 = temp3929 ^ temp3929;
    assign temp3931 = temp3930 ^ temp3930;
    assign temp3932 = temp3931 ^ temp3931;
    assign temp3933 = temp3932 ^ temp3932;
    assign temp3934 = temp3933 ^ temp3933;
    assign temp3935 = temp3934 ^ temp3934;
    assign temp3936 = temp3935 ^ temp3935;
    assign temp3937 = temp3936 ^ temp3936;
    assign temp3938 = temp3937 ^ temp3937;
    assign temp3939 = temp3938 ^ temp3938;
    assign temp3940 = temp3939 ^ temp3939;
    assign temp3941 = temp3940 ^ temp3940;
    assign temp3942 = temp3941 ^ temp3941;
    assign temp3943 = temp3942 ^ temp3942;
    assign temp3944 = temp3943 ^ temp3943;
    assign temp3945 = temp3944 ^ temp3944;
    assign temp3946 = temp3945 ^ temp3945;
    assign temp3947 = temp3946 ^ temp3946;
    assign temp3948 = temp3947 ^ temp3947;
    assign temp3949 = temp3948 ^ temp3948;
    assign temp3950 = temp3949 ^ temp3949;
    assign temp3951 = temp3950 ^ temp3950;
    assign temp3952 = temp3951 ^ temp3951;
    assign temp3953 = temp3952 ^ temp3952;
    assign temp3954 = temp3953 ^ temp3953;
    assign temp3955 = temp3954 ^ temp3954;
    assign temp3956 = temp3955 ^ temp3955;
    assign temp3957 = temp3956 ^ temp3956;
    assign temp3958 = temp3957 ^ temp3957;
    assign temp3959 = temp3958 ^ temp3958;
    assign temp3960 = temp3959 ^ temp3959;
    assign temp3961 = temp3960 ^ temp3960;
    assign temp3962 = temp3961 ^ temp3961;
    assign temp3963 = temp3962 ^ temp3962;
    assign temp3964 = temp3963 ^ temp3963;
    assign temp3965 = temp3964 ^ temp3964;
    assign temp3966 = temp3965 ^ temp3965;
    assign temp3967 = temp3966 ^ temp3966;
    assign temp3968 = temp3967 ^ temp3967;
    assign temp3969 = temp3968 ^ temp3968;
    assign temp3970 = temp3969 ^ temp3969;
    assign temp3971 = temp3970 ^ temp3970;
    assign temp3972 = temp3971 ^ temp3971;
    assign temp3973 = temp3972 ^ temp3972;
    assign temp3974 = temp3973 ^ temp3973;
    assign temp3975 = temp3974 ^ temp3974;
    assign temp3976 = temp3975 ^ temp3975;
    assign temp3977 = temp3976 ^ temp3976;
    assign temp3978 = temp3977 ^ temp3977;
    assign temp3979 = temp3978 ^ temp3978;
    assign temp3980 = temp3979 ^ temp3979;
    assign temp3981 = temp3980 ^ temp3980;
    assign temp3982 = temp3981 ^ temp3981;
    assign temp3983 = temp3982 ^ temp3982;
    assign temp3984 = temp3983 ^ temp3983;
    assign temp3985 = temp3984 ^ temp3984;
    assign temp3986 = temp3985 ^ temp3985;
    assign temp3987 = temp3986 ^ temp3986;
    assign temp3988 = temp3987 ^ temp3987;
    assign temp3989 = temp3988 ^ temp3988;
    assign temp3990 = temp3989 ^ temp3989;
    assign temp3991 = temp3990 ^ temp3990;
    assign temp3992 = temp3991 ^ temp3991;
    assign temp3993 = temp3992 ^ temp3992;
    assign temp3994 = temp3993 ^ temp3993;
    assign temp3995 = temp3994 ^ temp3994;
    assign temp3996 = temp3995 ^ temp3995;
    assign temp3997 = temp3996 ^ temp3996;
    assign temp3998 = temp3997 ^ temp3997;
    assign temp3999 = temp3998 ^ temp3998;
    assign temp4000 = temp3999 ^ temp3999;
    assign temp4001 = temp4000 ^ temp4000;
    assign temp4002 = temp4001 ^ temp4001;
    assign temp4003 = temp4002 ^ temp4002;
    assign temp4004 = temp4003 ^ temp4003;
    assign temp4005 = temp4004 ^ temp4004;
    assign temp4006 = temp4005 ^ temp4005;
    assign temp4007 = temp4006 ^ temp4006;
    assign temp4008 = temp4007 ^ temp4007;
    assign temp4009 = temp4008 ^ temp4008;
    assign temp4010 = temp4009 ^ temp4009;
    assign temp4011 = temp4010 ^ temp4010;
    assign temp4012 = temp4011 ^ temp4011;
    assign temp4013 = temp4012 ^ temp4012;
    assign temp4014 = temp4013 ^ temp4013;
    assign temp4015 = temp4014 ^ temp4014;
    assign temp4016 = temp4015 ^ temp4015;
    assign temp4017 = temp4016 ^ temp4016;
    assign temp4018 = temp4017 ^ temp4017;
    assign temp4019 = temp4018 ^ temp4018;
    assign temp4020 = temp4019 ^ temp4019;
    assign temp4021 = temp4020 ^ temp4020;
    assign temp4022 = temp4021 ^ temp4021;
    assign temp4023 = temp4022 ^ temp4022;
    assign temp4024 = temp4023 ^ temp4023;
    assign temp4025 = temp4024 ^ temp4024;
    assign temp4026 = temp4025 ^ temp4025;
    assign temp4027 = temp4026 ^ temp4026;
    assign temp4028 = temp4027 ^ temp4027;
    assign temp4029 = temp4028 ^ temp4028;
    assign temp4030 = temp4029 ^ temp4029;
    assign temp4031 = temp4030 ^ temp4030;
    assign temp4032 = temp4031 ^ temp4031;
    assign temp4033 = temp4032 ^ temp4032;
    assign temp4034 = temp4033 ^ temp4033;
    assign temp4035 = temp4034 ^ temp4034;
    assign temp4036 = temp4035 ^ temp4035;
    assign temp4037 = temp4036 ^ temp4036;
    assign temp4038 = temp4037 ^ temp4037;
    assign temp4039 = temp4038 ^ temp4038;
    assign temp4040 = temp4039 ^ temp4039;
    assign temp4041 = temp4040 ^ temp4040;
    assign temp4042 = temp4041 ^ temp4041;
    assign temp4043 = temp4042 ^ temp4042;
    assign temp4044 = temp4043 ^ temp4043;
    assign temp4045 = temp4044 ^ temp4044;
    assign temp4046 = temp4045 ^ temp4045;
    assign temp4047 = temp4046 ^ temp4046;
    assign temp4048 = temp4047 ^ temp4047;
    assign temp4049 = temp4048 ^ temp4048;
    assign temp4050 = temp4049 ^ temp4049;
    assign temp4051 = temp4050 ^ temp4050;
    assign temp4052 = temp4051 ^ temp4051;
    assign temp4053 = temp4052 ^ temp4052;
    assign temp4054 = temp4053 ^ temp4053;
    assign temp4055 = temp4054 ^ temp4054;
    assign temp4056 = temp4055 ^ temp4055;
    assign temp4057 = temp4056 ^ temp4056;
    assign temp4058 = temp4057 ^ temp4057;
    assign temp4059 = temp4058 ^ temp4058;
    assign temp4060 = temp4059 ^ temp4059;
    assign temp4061 = temp4060 ^ temp4060;
    assign temp4062 = temp4061 ^ temp4061;
    assign temp4063 = temp4062 ^ temp4062;
    assign temp4064 = temp4063 ^ temp4063;
    assign temp4065 = temp4064 ^ temp4064;
    assign temp4066 = temp4065 ^ temp4065;
    assign temp4067 = temp4066 ^ temp4066;
    assign temp4068 = temp4067 ^ temp4067;
    assign temp4069 = temp4068 ^ temp4068;
    assign temp4070 = temp4069 ^ temp4069;
    assign temp4071 = temp4070 ^ temp4070;
    assign temp4072 = temp4071 ^ temp4071;
    assign temp4073 = temp4072 ^ temp4072;
    assign temp4074 = temp4073 ^ temp4073;
    assign temp4075 = temp4074 ^ temp4074;
    assign temp4076 = temp4075 ^ temp4075;
    assign temp4077 = temp4076 ^ temp4076;
    assign temp4078 = temp4077 ^ temp4077;
    assign temp4079 = temp4078 ^ temp4078;
    assign temp4080 = temp4079 ^ temp4079;
    assign temp4081 = temp4080 ^ temp4080;
    assign temp4082 = temp4081 ^ temp4081;
    assign temp4083 = temp4082 ^ temp4082;
    assign temp4084 = temp4083 ^ temp4083;
    assign temp4085 = temp4084 ^ temp4084;
    assign temp4086 = temp4085 ^ temp4085;
    assign temp4087 = temp4086 ^ temp4086;
    assign temp4088 = temp4087 ^ temp4087;
    assign temp4089 = temp4088 ^ temp4088;
    assign temp4090 = temp4089 ^ temp4089;
    assign temp4091 = temp4090 ^ temp4090;
    assign temp4092 = temp4091 ^ temp4091;
    assign temp4093 = temp4092 ^ temp4092;
    assign temp4094 = temp4093 ^ temp4093;
    assign temp4095 = temp4094 ^ temp4094;
    assign temp4096 = temp4095 ^ temp4095;
    assign temp4097 = temp4096 ^ temp4096;
    assign temp4098 = temp4097 ^ temp4097;
    assign temp4099 = temp4098 ^ temp4098;
    assign temp4100 = temp4099 ^ temp4099;
    assign temp4101 = temp4100 ^ temp4100;
    assign temp4102 = temp4101 ^ temp4101;
    assign temp4103 = temp4102 ^ temp4102;
    assign temp4104 = temp4103 ^ temp4103;
    assign temp4105 = temp4104 ^ temp4104;
    assign temp4106 = temp4105 ^ temp4105;
    assign temp4107 = temp4106 ^ temp4106;
    assign temp4108 = temp4107 ^ temp4107;
    assign temp4109 = temp4108 ^ temp4108;
    assign temp4110 = temp4109 ^ temp4109;
    assign temp4111 = temp4110 ^ temp4110;
    assign temp4112 = temp4111 ^ temp4111;
    assign temp4113 = temp4112 ^ temp4112;
    assign temp4114 = temp4113 ^ temp4113;
    assign temp4115 = temp4114 ^ temp4114;
    assign temp4116 = temp4115 ^ temp4115;
    assign temp4117 = temp4116 ^ temp4116;
    assign temp4118 = temp4117 ^ temp4117;
    assign temp4119 = temp4118 ^ temp4118;
    assign temp4120 = temp4119 ^ temp4119;
    assign temp4121 = temp4120 ^ temp4120;
    assign temp4122 = temp4121 ^ temp4121;
    assign temp4123 = temp4122 ^ temp4122;
    assign temp4124 = temp4123 ^ temp4123;
    assign temp4125 = temp4124 ^ temp4124;
    assign temp4126 = temp4125 ^ temp4125;
    assign temp4127 = temp4126 ^ temp4126;
    assign temp4128 = temp4127 ^ temp4127;
    assign temp4129 = temp4128 ^ temp4128;
    assign temp4130 = temp4129 ^ temp4129;
    assign temp4131 = temp4130 ^ temp4130;
    assign temp4132 = temp4131 ^ temp4131;
    assign temp4133 = temp4132 ^ temp4132;
    assign temp4134 = temp4133 ^ temp4133;
    assign temp4135 = temp4134 ^ temp4134;
    assign temp4136 = temp4135 ^ temp4135;
    assign temp4137 = temp4136 ^ temp4136;
    assign temp4138 = temp4137 ^ temp4137;
    assign temp4139 = temp4138 ^ temp4138;
    assign temp4140 = temp4139 ^ temp4139;
    assign temp4141 = temp4140 ^ temp4140;
    assign temp4142 = temp4141 ^ temp4141;
    assign temp4143 = temp4142 ^ temp4142;
    assign temp4144 = temp4143 ^ temp4143;
    assign temp4145 = temp4144 ^ temp4144;
    assign temp4146 = temp4145 ^ temp4145;
    assign temp4147 = temp4146 ^ temp4146;
    assign temp4148 = temp4147 ^ temp4147;
    assign temp4149 = temp4148 ^ temp4148;
    assign temp4150 = temp4149 ^ temp4149;
    assign temp4151 = temp4150 ^ temp4150;
    assign temp4152 = temp4151 ^ temp4151;
    assign temp4153 = temp4152 ^ temp4152;
    assign temp4154 = temp4153 ^ temp4153;
    assign temp4155 = temp4154 ^ temp4154;
    assign temp4156 = temp4155 ^ temp4155;
    assign temp4157 = temp4156 ^ temp4156;
    assign temp4158 = temp4157 ^ temp4157;
    assign temp4159 = temp4158 ^ temp4158;
    assign temp4160 = temp4159 ^ temp4159;
    assign temp4161 = temp4160 ^ temp4160;
    assign temp4162 = temp4161 ^ temp4161;
    assign temp4163 = temp4162 ^ temp4162;
    assign temp4164 = temp4163 ^ temp4163;
    assign temp4165 = temp4164 ^ temp4164;
    assign temp4166 = temp4165 ^ temp4165;
    assign temp4167 = temp4166 ^ temp4166;
    assign temp4168 = temp4167 ^ temp4167;
    assign temp4169 = temp4168 ^ temp4168;
    assign temp4170 = temp4169 ^ temp4169;
    assign temp4171 = temp4170 ^ temp4170;
    assign temp4172 = temp4171 ^ temp4171;
    assign temp4173 = temp4172 ^ temp4172;
    assign temp4174 = temp4173 ^ temp4173;
    assign temp4175 = temp4174 ^ temp4174;
    assign temp4176 = temp4175 ^ temp4175;
    assign temp4177 = temp4176 ^ temp4176;
    assign temp4178 = temp4177 ^ temp4177;
    assign temp4179 = temp4178 ^ temp4178;
    assign temp4180 = temp4179 ^ temp4179;
    assign temp4181 = temp4180 ^ temp4180;
    assign temp4182 = temp4181 ^ temp4181;
    assign temp4183 = temp4182 ^ temp4182;
    assign temp4184 = temp4183 ^ temp4183;
    assign temp4185 = temp4184 ^ temp4184;
    assign temp4186 = temp4185 ^ temp4185;
    assign temp4187 = temp4186 ^ temp4186;
    assign temp4188 = temp4187 ^ temp4187;
    assign temp4189 = temp4188 ^ temp4188;
    assign temp4190 = temp4189 ^ temp4189;
    assign temp4191 = temp4190 ^ temp4190;
    assign temp4192 = temp4191 ^ temp4191;
    assign temp4193 = temp4192 ^ temp4192;
    assign temp4194 = temp4193 ^ temp4193;
    assign temp4195 = temp4194 ^ temp4194;
    assign temp4196 = temp4195 ^ temp4195;
    assign temp4197 = temp4196 ^ temp4196;
    assign temp4198 = temp4197 ^ temp4197;
    assign temp4199 = temp4198 ^ temp4198;
    assign temp4200 = temp4199 ^ temp4199;
    assign temp4201 = temp4200 ^ temp4200;
    assign temp4202 = temp4201 ^ temp4201;
    assign temp4203 = temp4202 ^ temp4202;
    assign temp4204 = temp4203 ^ temp4203;
    assign temp4205 = temp4204 ^ temp4204;
    assign temp4206 = temp4205 ^ temp4205;
    assign temp4207 = temp4206 ^ temp4206;
    assign temp4208 = temp4207 ^ temp4207;
    assign temp4209 = temp4208 ^ temp4208;
    assign temp4210 = temp4209 ^ temp4209;
    assign temp4211 = temp4210 ^ temp4210;
    assign temp4212 = temp4211 ^ temp4211;
    assign temp4213 = temp4212 ^ temp4212;
    assign temp4214 = temp4213 ^ temp4213;
    assign temp4215 = temp4214 ^ temp4214;
    assign temp4216 = temp4215 ^ temp4215;
    assign temp4217 = temp4216 ^ temp4216;
    assign temp4218 = temp4217 ^ temp4217;
    assign temp4219 = temp4218 ^ temp4218;
    assign temp4220 = temp4219 ^ temp4219;
    assign temp4221 = temp4220 ^ temp4220;
    assign temp4222 = temp4221 ^ temp4221;
    assign temp4223 = temp4222 ^ temp4222;
    assign temp4224 = temp4223 ^ temp4223;
    assign temp4225 = temp4224 ^ temp4224;
    assign temp4226 = temp4225 ^ temp4225;
    assign temp4227 = temp4226 ^ temp4226;
    assign temp4228 = temp4227 ^ temp4227;
    assign temp4229 = temp4228 ^ temp4228;
    assign temp4230 = temp4229 ^ temp4229;
    assign temp4231 = temp4230 ^ temp4230;
    assign temp4232 = temp4231 ^ temp4231;
    assign temp4233 = temp4232 ^ temp4232;
    assign temp4234 = temp4233 ^ temp4233;
    assign temp4235 = temp4234 ^ temp4234;
    assign temp4236 = temp4235 ^ temp4235;
    assign temp4237 = temp4236 ^ temp4236;
    assign temp4238 = temp4237 ^ temp4237;
    assign temp4239 = temp4238 ^ temp4238;
    assign temp4240 = temp4239 ^ temp4239;
    assign temp4241 = temp4240 ^ temp4240;
    assign temp4242 = temp4241 ^ temp4241;
    assign temp4243 = temp4242 ^ temp4242;
    assign temp4244 = temp4243 ^ temp4243;
    assign temp4245 = temp4244 ^ temp4244;
    assign temp4246 = temp4245 ^ temp4245;
    assign temp4247 = temp4246 ^ temp4246;
    assign temp4248 = temp4247 ^ temp4247;
    assign temp4249 = temp4248 ^ temp4248;
    assign temp4250 = temp4249 ^ temp4249;
    assign temp4251 = temp4250 ^ temp4250;
    assign temp4252 = temp4251 ^ temp4251;
    assign temp4253 = temp4252 ^ temp4252;
    assign temp4254 = temp4253 ^ temp4253;
    assign temp4255 = temp4254 ^ temp4254;
    assign temp4256 = temp4255 ^ temp4255;
    assign temp4257 = temp4256 ^ temp4256;
    assign temp4258 = temp4257 ^ temp4257;
    assign temp4259 = temp4258 ^ temp4258;
    assign temp4260 = temp4259 ^ temp4259;
    assign temp4261 = temp4260 ^ temp4260;
    assign temp4262 = temp4261 ^ temp4261;
    assign temp4263 = temp4262 ^ temp4262;
    assign temp4264 = temp4263 ^ temp4263;
    assign temp4265 = temp4264 ^ temp4264;
    assign temp4266 = temp4265 ^ temp4265;
    assign temp4267 = temp4266 ^ temp4266;
    assign temp4268 = temp4267 ^ temp4267;
    assign temp4269 = temp4268 ^ temp4268;
    assign temp4270 = temp4269 ^ temp4269;
    assign temp4271 = temp4270 ^ temp4270;
    assign temp4272 = temp4271 ^ temp4271;
    assign temp4273 = temp4272 ^ temp4272;
    assign temp4274 = temp4273 ^ temp4273;
    assign temp4275 = temp4274 ^ temp4274;
    assign temp4276 = temp4275 ^ temp4275;
    assign temp4277 = temp4276 ^ temp4276;
    assign temp4278 = temp4277 ^ temp4277;
    assign temp4279 = temp4278 ^ temp4278;
    assign temp4280 = temp4279 ^ temp4279;
    assign temp4281 = temp4280 ^ temp4280;
    assign temp4282 = temp4281 ^ temp4281;
    assign temp4283 = temp4282 ^ temp4282;
    assign temp4284 = temp4283 ^ temp4283;
    assign temp4285 = temp4284 ^ temp4284;
    assign temp4286 = temp4285 ^ temp4285;
    assign temp4287 = temp4286 ^ temp4286;
    assign temp4288 = temp4287 ^ temp4287;
    assign temp4289 = temp4288 ^ temp4288;
    assign temp4290 = temp4289 ^ temp4289;
    assign temp4291 = temp4290 ^ temp4290;
    assign temp4292 = temp4291 ^ temp4291;
    assign temp4293 = temp4292 ^ temp4292;
    assign temp4294 = temp4293 ^ temp4293;
    assign temp4295 = temp4294 ^ temp4294;
    assign temp4296 = temp4295 ^ temp4295;
    assign temp4297 = temp4296 ^ temp4296;
    assign temp4298 = temp4297 ^ temp4297;
    assign temp4299 = temp4298 ^ temp4298;
    assign temp4300 = temp4299 ^ temp4299;
    assign temp4301 = temp4300 ^ temp4300;
    assign temp4302 = temp4301 ^ temp4301;
    assign temp4303 = temp4302 ^ temp4302;
    assign temp4304 = temp4303 ^ temp4303;
    assign temp4305 = temp4304 ^ temp4304;
    assign temp4306 = temp4305 ^ temp4305;
    assign temp4307 = temp4306 ^ temp4306;
    assign temp4308 = temp4307 ^ temp4307;
    assign temp4309 = temp4308 ^ temp4308;
    assign temp4310 = temp4309 ^ temp4309;
    assign temp4311 = temp4310 ^ temp4310;
    assign temp4312 = temp4311 ^ temp4311;
    assign temp4313 = temp4312 ^ temp4312;
    assign temp4314 = temp4313 ^ temp4313;
    assign temp4315 = temp4314 ^ temp4314;
    assign temp4316 = temp4315 ^ temp4315;
    assign temp4317 = temp4316 ^ temp4316;
    assign temp4318 = temp4317 ^ temp4317;
    assign temp4319 = temp4318 ^ temp4318;
    assign temp4320 = temp4319 ^ temp4319;
    assign temp4321 = temp4320 ^ temp4320;
    assign temp4322 = temp4321 ^ temp4321;
    assign temp4323 = temp4322 ^ temp4322;
    assign temp4324 = temp4323 ^ temp4323;
    assign temp4325 = temp4324 ^ temp4324;
    assign temp4326 = temp4325 ^ temp4325;
    assign temp4327 = temp4326 ^ temp4326;
    assign temp4328 = temp4327 ^ temp4327;
    assign temp4329 = temp4328 ^ temp4328;
    assign temp4330 = temp4329 ^ temp4329;
    assign temp4331 = temp4330 ^ temp4330;
    assign temp4332 = temp4331 ^ temp4331;
    assign temp4333 = temp4332 ^ temp4332;
    assign temp4334 = temp4333 ^ temp4333;
    assign temp4335 = temp4334 ^ temp4334;
    assign temp4336 = temp4335 ^ temp4335;
    assign temp4337 = temp4336 ^ temp4336;
    assign temp4338 = temp4337 ^ temp4337;
    assign temp4339 = temp4338 ^ temp4338;
    assign temp4340 = temp4339 ^ temp4339;
    assign temp4341 = temp4340 ^ temp4340;
    assign temp4342 = temp4341 ^ temp4341;
    assign temp4343 = temp4342 ^ temp4342;
    assign temp4344 = temp4343 ^ temp4343;
    assign temp4345 = temp4344 ^ temp4344;
    assign temp4346 = temp4345 ^ temp4345;
    assign temp4347 = temp4346 ^ temp4346;
    assign temp4348 = temp4347 ^ temp4347;
    assign temp4349 = temp4348 ^ temp4348;
    assign temp4350 = temp4349 ^ temp4349;
    assign temp4351 = temp4350 ^ temp4350;
    assign temp4352 = temp4351 ^ temp4351;
    assign temp4353 = temp4352 ^ temp4352;
    assign temp4354 = temp4353 ^ temp4353;
    assign temp4355 = temp4354 ^ temp4354;
    assign temp4356 = temp4355 ^ temp4355;
    assign temp4357 = temp4356 ^ temp4356;
    assign temp4358 = temp4357 ^ temp4357;
    assign temp4359 = temp4358 ^ temp4358;
    assign temp4360 = temp4359 ^ temp4359;
    assign temp4361 = temp4360 ^ temp4360;
    assign temp4362 = temp4361 ^ temp4361;
    assign temp4363 = temp4362 ^ temp4362;
    assign temp4364 = temp4363 ^ temp4363;
    assign temp4365 = temp4364 ^ temp4364;
    assign temp4366 = temp4365 ^ temp4365;
    assign temp4367 = temp4366 ^ temp4366;
    assign temp4368 = temp4367 ^ temp4367;
    assign temp4369 = temp4368 ^ temp4368;
    assign temp4370 = temp4369 ^ temp4369;
    assign temp4371 = temp4370 ^ temp4370;
    assign temp4372 = temp4371 ^ temp4371;
    assign temp4373 = temp4372 ^ temp4372;
    assign temp4374 = temp4373 ^ temp4373;
    assign temp4375 = temp4374 ^ temp4374;
    assign temp4376 = temp4375 ^ temp4375;
    assign temp4377 = temp4376 ^ temp4376;
    assign temp4378 = temp4377 ^ temp4377;
    assign temp4379 = temp4378 ^ temp4378;
    assign temp4380 = temp4379 ^ temp4379;
    assign temp4381 = temp4380 ^ temp4380;
    assign temp4382 = temp4381 ^ temp4381;
    assign temp4383 = temp4382 ^ temp4382;
    assign temp4384 = temp4383 ^ temp4383;
    assign temp4385 = temp4384 ^ temp4384;
    assign temp4386 = temp4385 ^ temp4385;
    assign temp4387 = temp4386 ^ temp4386;
    assign temp4388 = temp4387 ^ temp4387;
    assign temp4389 = temp4388 ^ temp4388;
    assign temp4390 = temp4389 ^ temp4389;
    assign temp4391 = temp4390 ^ temp4390;
    assign temp4392 = temp4391 ^ temp4391;
    assign temp4393 = temp4392 ^ temp4392;
    assign temp4394 = temp4393 ^ temp4393;
    assign temp4395 = temp4394 ^ temp4394;
    assign temp4396 = temp4395 ^ temp4395;
    assign temp4397 = temp4396 ^ temp4396;
    assign temp4398 = temp4397 ^ temp4397;
    assign temp4399 = temp4398 ^ temp4398;
    assign temp4400 = temp4399 ^ temp4399;
    assign temp4401 = temp4400 ^ temp4400;
    assign temp4402 = temp4401 ^ temp4401;
    assign temp4403 = temp4402 ^ temp4402;
    assign temp4404 = temp4403 ^ temp4403;
    assign temp4405 = temp4404 ^ temp4404;
    assign temp4406 = temp4405 ^ temp4405;
    assign temp4407 = temp4406 ^ temp4406;
    assign temp4408 = temp4407 ^ temp4407;
    assign temp4409 = temp4408 ^ temp4408;
    assign temp4410 = temp4409 ^ temp4409;
    assign temp4411 = temp4410 ^ temp4410;
    assign temp4412 = temp4411 ^ temp4411;
    assign temp4413 = temp4412 ^ temp4412;
    assign temp4414 = temp4413 ^ temp4413;
    assign temp4415 = temp4414 ^ temp4414;
    assign temp4416 = temp4415 ^ temp4415;
    assign temp4417 = temp4416 ^ temp4416;
    assign temp4418 = temp4417 ^ temp4417;
    assign temp4419 = temp4418 ^ temp4418;
    assign temp4420 = temp4419 ^ temp4419;
    assign temp4421 = temp4420 ^ temp4420;
    assign temp4422 = temp4421 ^ temp4421;
    assign temp4423 = temp4422 ^ temp4422;
    assign temp4424 = temp4423 ^ temp4423;
    assign temp4425 = temp4424 ^ temp4424;
    assign temp4426 = temp4425 ^ temp4425;
    assign temp4427 = temp4426 ^ temp4426;
    assign temp4428 = temp4427 ^ temp4427;
    assign temp4429 = temp4428 ^ temp4428;
    assign temp4430 = temp4429 ^ temp4429;
    assign temp4431 = temp4430 ^ temp4430;
    assign temp4432 = temp4431 ^ temp4431;
    assign temp4433 = temp4432 ^ temp4432;
    assign temp4434 = temp4433 ^ temp4433;
    assign temp4435 = temp4434 ^ temp4434;
    assign temp4436 = temp4435 ^ temp4435;
    assign temp4437 = temp4436 ^ temp4436;
    assign temp4438 = temp4437 ^ temp4437;
    assign temp4439 = temp4438 ^ temp4438;
    assign temp4440 = temp4439 ^ temp4439;
    assign temp4441 = temp4440 ^ temp4440;
    assign temp4442 = temp4441 ^ temp4441;
    assign temp4443 = temp4442 ^ temp4442;
    assign temp4444 = temp4443 ^ temp4443;
    assign temp4445 = temp4444 ^ temp4444;
    assign temp4446 = temp4445 ^ temp4445;
    assign temp4447 = temp4446 ^ temp4446;
    assign temp4448 = temp4447 ^ temp4447;
    assign temp4449 = temp4448 ^ temp4448;
    assign temp4450 = temp4449 ^ temp4449;
    assign temp4451 = temp4450 ^ temp4450;
    assign temp4452 = temp4451 ^ temp4451;
    assign temp4453 = temp4452 ^ temp4452;
    assign temp4454 = temp4453 ^ temp4453;
    assign temp4455 = temp4454 ^ temp4454;
    assign temp4456 = temp4455 ^ temp4455;
    assign temp4457 = temp4456 ^ temp4456;
    assign temp4458 = temp4457 ^ temp4457;
    assign temp4459 = temp4458 ^ temp4458;
    assign temp4460 = temp4459 ^ temp4459;
    assign temp4461 = temp4460 ^ temp4460;
    assign temp4462 = temp4461 ^ temp4461;
    assign temp4463 = temp4462 ^ temp4462;
    assign temp4464 = temp4463 ^ temp4463;
    assign temp4465 = temp4464 ^ temp4464;
    assign temp4466 = temp4465 ^ temp4465;
    assign temp4467 = temp4466 ^ temp4466;
    assign temp4468 = temp4467 ^ temp4467;
    assign temp4469 = temp4468 ^ temp4468;
    assign temp4470 = temp4469 ^ temp4469;
    assign temp4471 = temp4470 ^ temp4470;
    assign temp4472 = temp4471 ^ temp4471;
    assign temp4473 = temp4472 ^ temp4472;
    assign temp4474 = temp4473 ^ temp4473;
    assign temp4475 = temp4474 ^ temp4474;
    assign temp4476 = temp4475 ^ temp4475;
    assign temp4477 = temp4476 ^ temp4476;
    assign temp4478 = temp4477 ^ temp4477;
    assign temp4479 = temp4478 ^ temp4478;
    assign temp4480 = temp4479 ^ temp4479;
    assign temp4481 = temp4480 ^ temp4480;
    assign temp4482 = temp4481 ^ temp4481;
    assign temp4483 = temp4482 ^ temp4482;
    assign temp4484 = temp4483 ^ temp4483;
    assign temp4485 = temp4484 ^ temp4484;
    assign temp4486 = temp4485 ^ temp4485;
    assign temp4487 = temp4486 ^ temp4486;
    assign temp4488 = temp4487 ^ temp4487;
    assign temp4489 = temp4488 ^ temp4488;
    assign temp4490 = temp4489 ^ temp4489;
    assign temp4491 = temp4490 ^ temp4490;
    assign temp4492 = temp4491 ^ temp4491;
    assign temp4493 = temp4492 ^ temp4492;
    assign temp4494 = temp4493 ^ temp4493;
    assign temp4495 = temp4494 ^ temp4494;
    assign temp4496 = temp4495 ^ temp4495;
    assign temp4497 = temp4496 ^ temp4496;
    assign temp4498 = temp4497 ^ temp4497;
    assign temp4499 = temp4498 ^ temp4498;
    assign temp4500 = temp4499 ^ temp4499;
    assign temp4501 = temp4500 ^ temp4500;
    assign temp4502 = temp4501 ^ temp4501;
    assign temp4503 = temp4502 ^ temp4502;
    assign temp4504 = temp4503 ^ temp4503;
    assign temp4505 = temp4504 ^ temp4504;
    assign temp4506 = temp4505 ^ temp4505;
    assign temp4507 = temp4506 ^ temp4506;
    assign temp4508 = temp4507 ^ temp4507;
    assign temp4509 = temp4508 ^ temp4508;
    assign temp4510 = temp4509 ^ temp4509;
    assign temp4511 = temp4510 ^ temp4510;
    assign temp4512 = temp4511 ^ temp4511;
    assign temp4513 = temp4512 ^ temp4512;
    assign temp4514 = temp4513 ^ temp4513;
    assign temp4515 = temp4514 ^ temp4514;
    assign temp4516 = temp4515 ^ temp4515;
    assign temp4517 = temp4516 ^ temp4516;
    assign temp4518 = temp4517 ^ temp4517;
    assign temp4519 = temp4518 ^ temp4518;
    assign temp4520 = temp4519 ^ temp4519;
    assign temp4521 = temp4520 ^ temp4520;
    assign temp4522 = temp4521 ^ temp4521;
    assign temp4523 = temp4522 ^ temp4522;
    assign temp4524 = temp4523 ^ temp4523;
    assign temp4525 = temp4524 ^ temp4524;
    assign temp4526 = temp4525 ^ temp4525;
    assign temp4527 = temp4526 ^ temp4526;
    assign temp4528 = temp4527 ^ temp4527;
    assign temp4529 = temp4528 ^ temp4528;
    assign temp4530 = temp4529 ^ temp4529;
    assign temp4531 = temp4530 ^ temp4530;
    assign temp4532 = temp4531 ^ temp4531;
    assign temp4533 = temp4532 ^ temp4532;
    assign temp4534 = temp4533 ^ temp4533;
    assign temp4535 = temp4534 ^ temp4534;
    assign temp4536 = temp4535 ^ temp4535;
    assign temp4537 = temp4536 ^ temp4536;
    assign temp4538 = temp4537 ^ temp4537;
    assign temp4539 = temp4538 ^ temp4538;
    assign temp4540 = temp4539 ^ temp4539;
    assign temp4541 = temp4540 ^ temp4540;
    assign temp4542 = temp4541 ^ temp4541;
    assign temp4543 = temp4542 ^ temp4542;
    assign temp4544 = temp4543 ^ temp4543;
    assign temp4545 = temp4544 ^ temp4544;
    assign temp4546 = temp4545 ^ temp4545;
    assign temp4547 = temp4546 ^ temp4546;
    assign temp4548 = temp4547 ^ temp4547;
    assign temp4549 = temp4548 ^ temp4548;
    assign temp4550 = temp4549 ^ temp4549;
    assign temp4551 = temp4550 ^ temp4550;
    assign temp4552 = temp4551 ^ temp4551;
    assign temp4553 = temp4552 ^ temp4552;
    assign temp4554 = temp4553 ^ temp4553;
    assign temp4555 = temp4554 ^ temp4554;
    assign temp4556 = temp4555 ^ temp4555;
    assign temp4557 = temp4556 ^ temp4556;
    assign temp4558 = temp4557 ^ temp4557;
    assign temp4559 = temp4558 ^ temp4558;
    assign temp4560 = temp4559 ^ temp4559;
    assign temp4561 = temp4560 ^ temp4560;
    assign temp4562 = temp4561 ^ temp4561;
    assign temp4563 = temp4562 ^ temp4562;
    assign temp4564 = temp4563 ^ temp4563;
    assign temp4565 = temp4564 ^ temp4564;
    assign temp4566 = temp4565 ^ temp4565;
    assign temp4567 = temp4566 ^ temp4566;
    assign temp4568 = temp4567 ^ temp4567;
    assign temp4569 = temp4568 ^ temp4568;
    assign temp4570 = temp4569 ^ temp4569;
    assign temp4571 = temp4570 ^ temp4570;
    assign temp4572 = temp4571 ^ temp4571;
    assign temp4573 = temp4572 ^ temp4572;
    assign temp4574 = temp4573 ^ temp4573;
    assign temp4575 = temp4574 ^ temp4574;
    assign temp4576 = temp4575 ^ temp4575;
    assign temp4577 = temp4576 ^ temp4576;
    assign temp4578 = temp4577 ^ temp4577;
    assign temp4579 = temp4578 ^ temp4578;
    assign temp4580 = temp4579 ^ temp4579;
    assign temp4581 = temp4580 ^ temp4580;
    assign temp4582 = temp4581 ^ temp4581;
    assign temp4583 = temp4582 ^ temp4582;
    assign temp4584 = temp4583 ^ temp4583;
    assign temp4585 = temp4584 ^ temp4584;
    assign temp4586 = temp4585 ^ temp4585;
    assign temp4587 = temp4586 ^ temp4586;
    assign temp4588 = temp4587 ^ temp4587;
    assign temp4589 = temp4588 ^ temp4588;
    assign temp4590 = temp4589 ^ temp4589;
    assign temp4591 = temp4590 ^ temp4590;
    assign temp4592 = temp4591 ^ temp4591;
    assign temp4593 = temp4592 ^ temp4592;
    assign temp4594 = temp4593 ^ temp4593;
    assign temp4595 = temp4594 ^ temp4594;
    assign temp4596 = temp4595 ^ temp4595;
    assign temp4597 = temp4596 ^ temp4596;
    assign temp4598 = temp4597 ^ temp4597;
    assign temp4599 = temp4598 ^ temp4598;
    assign temp4600 = temp4599 ^ temp4599;
    assign temp4601 = temp4600 ^ temp4600;
    assign temp4602 = temp4601 ^ temp4601;
    assign temp4603 = temp4602 ^ temp4602;
    assign temp4604 = temp4603 ^ temp4603;
    assign temp4605 = temp4604 ^ temp4604;
    assign temp4606 = temp4605 ^ temp4605;
    assign temp4607 = temp4606 ^ temp4606;
    assign temp4608 = temp4607 ^ temp4607;
    assign temp4609 = temp4608 ^ temp4608;
    assign temp4610 = temp4609 ^ temp4609;
    assign temp4611 = temp4610 ^ temp4610;
    assign temp4612 = temp4611 ^ temp4611;
    assign temp4613 = temp4612 ^ temp4612;
    assign temp4614 = temp4613 ^ temp4613;
    assign temp4615 = temp4614 ^ temp4614;
    assign temp4616 = temp4615 ^ temp4615;
    assign temp4617 = temp4616 ^ temp4616;
    assign temp4618 = temp4617 ^ temp4617;
    assign temp4619 = temp4618 ^ temp4618;
    assign temp4620 = temp4619 ^ temp4619;
    assign temp4621 = temp4620 ^ temp4620;
    assign temp4622 = temp4621 ^ temp4621;
    assign temp4623 = temp4622 ^ temp4622;
    assign temp4624 = temp4623 ^ temp4623;
    assign temp4625 = temp4624 ^ temp4624;
    assign temp4626 = temp4625 ^ temp4625;
    assign temp4627 = temp4626 ^ temp4626;
    assign temp4628 = temp4627 ^ temp4627;
    assign temp4629 = temp4628 ^ temp4628;
    assign temp4630 = temp4629 ^ temp4629;
    assign temp4631 = temp4630 ^ temp4630;
    assign temp4632 = temp4631 ^ temp4631;
    assign temp4633 = temp4632 ^ temp4632;
    assign temp4634 = temp4633 ^ temp4633;
    assign temp4635 = temp4634 ^ temp4634;
    assign temp4636 = temp4635 ^ temp4635;
    assign temp4637 = temp4636 ^ temp4636;
    assign temp4638 = temp4637 ^ temp4637;
    assign temp4639 = temp4638 ^ temp4638;
    assign temp4640 = temp4639 ^ temp4639;
    assign temp4641 = temp4640 ^ temp4640;
    assign temp4642 = temp4641 ^ temp4641;
    assign temp4643 = temp4642 ^ temp4642;
    assign temp4644 = temp4643 ^ temp4643;
    assign temp4645 = temp4644 ^ temp4644;
    assign temp4646 = temp4645 ^ temp4645;
    assign temp4647 = temp4646 ^ temp4646;
    assign temp4648 = temp4647 ^ temp4647;
    assign temp4649 = temp4648 ^ temp4648;
    assign temp4650 = temp4649 ^ temp4649;
    assign temp4651 = temp4650 ^ temp4650;
    assign temp4652 = temp4651 ^ temp4651;
    assign temp4653 = temp4652 ^ temp4652;
    assign temp4654 = temp4653 ^ temp4653;
    assign temp4655 = temp4654 ^ temp4654;
    assign temp4656 = temp4655 ^ temp4655;
    assign temp4657 = temp4656 ^ temp4656;
    assign temp4658 = temp4657 ^ temp4657;
    assign temp4659 = temp4658 ^ temp4658;
    assign temp4660 = temp4659 ^ temp4659;
    assign temp4661 = temp4660 ^ temp4660;
    assign temp4662 = temp4661 ^ temp4661;
    assign temp4663 = temp4662 ^ temp4662;
    assign temp4664 = temp4663 ^ temp4663;
    assign temp4665 = temp4664 ^ temp4664;
    assign temp4666 = temp4665 ^ temp4665;
    assign temp4667 = temp4666 ^ temp4666;
    assign temp4668 = temp4667 ^ temp4667;
    assign temp4669 = temp4668 ^ temp4668;
    assign temp4670 = temp4669 ^ temp4669;
    assign temp4671 = temp4670 ^ temp4670;
    assign temp4672 = temp4671 ^ temp4671;
    assign temp4673 = temp4672 ^ temp4672;
    assign temp4674 = temp4673 ^ temp4673;
    assign temp4675 = temp4674 ^ temp4674;
    assign temp4676 = temp4675 ^ temp4675;
    assign temp4677 = temp4676 ^ temp4676;
    assign temp4678 = temp4677 ^ temp4677;
    assign temp4679 = temp4678 ^ temp4678;
    assign temp4680 = temp4679 ^ temp4679;
    assign temp4681 = temp4680 ^ temp4680;
    assign temp4682 = temp4681 ^ temp4681;
    assign temp4683 = temp4682 ^ temp4682;
    assign temp4684 = temp4683 ^ temp4683;
    assign temp4685 = temp4684 ^ temp4684;
    assign temp4686 = temp4685 ^ temp4685;
    assign temp4687 = temp4686 ^ temp4686;
    assign temp4688 = temp4687 ^ temp4687;
    assign temp4689 = temp4688 ^ temp4688;
    assign temp4690 = temp4689 ^ temp4689;
    assign temp4691 = temp4690 ^ temp4690;
    assign temp4692 = temp4691 ^ temp4691;
    assign temp4693 = temp4692 ^ temp4692;
    assign temp4694 = temp4693 ^ temp4693;
    assign temp4695 = temp4694 ^ temp4694;
    assign temp4696 = temp4695 ^ temp4695;
    assign temp4697 = temp4696 ^ temp4696;
    assign temp4698 = temp4697 ^ temp4697;
    assign temp4699 = temp4698 ^ temp4698;
    assign temp4700 = temp4699 ^ temp4699;
    assign temp4701 = temp4700 ^ temp4700;
    assign temp4702 = temp4701 ^ temp4701;
    assign temp4703 = temp4702 ^ temp4702;
    assign temp4704 = temp4703 ^ temp4703;
    assign temp4705 = temp4704 ^ temp4704;
    assign temp4706 = temp4705 ^ temp4705;
    assign temp4707 = temp4706 ^ temp4706;
    assign temp4708 = temp4707 ^ temp4707;
    assign temp4709 = temp4708 ^ temp4708;
    assign temp4710 = temp4709 ^ temp4709;
    assign temp4711 = temp4710 ^ temp4710;
    assign temp4712 = temp4711 ^ temp4711;
    assign temp4713 = temp4712 ^ temp4712;
    assign temp4714 = temp4713 ^ temp4713;
    assign temp4715 = temp4714 ^ temp4714;
    assign temp4716 = temp4715 ^ temp4715;
    assign temp4717 = temp4716 ^ temp4716;
    assign temp4718 = temp4717 ^ temp4717;
    assign temp4719 = temp4718 ^ temp4718;
    assign temp4720 = temp4719 ^ temp4719;
    assign temp4721 = temp4720 ^ temp4720;
    assign temp4722 = temp4721 ^ temp4721;
    assign temp4723 = temp4722 ^ temp4722;
    assign temp4724 = temp4723 ^ temp4723;
    assign temp4725 = temp4724 ^ temp4724;
    assign temp4726 = temp4725 ^ temp4725;
    assign temp4727 = temp4726 ^ temp4726;
    assign temp4728 = temp4727 ^ temp4727;
    assign temp4729 = temp4728 ^ temp4728;
    assign temp4730 = temp4729 ^ temp4729;
    assign temp4731 = temp4730 ^ temp4730;
    assign temp4732 = temp4731 ^ temp4731;
    assign temp4733 = temp4732 ^ temp4732;
    assign temp4734 = temp4733 ^ temp4733;
    assign temp4735 = temp4734 ^ temp4734;
    assign temp4736 = temp4735 ^ temp4735;
    assign temp4737 = temp4736 ^ temp4736;
    assign temp4738 = temp4737 ^ temp4737;
    assign temp4739 = temp4738 ^ temp4738;
    assign temp4740 = temp4739 ^ temp4739;
    assign temp4741 = temp4740 ^ temp4740;
    assign temp4742 = temp4741 ^ temp4741;
    assign temp4743 = temp4742 ^ temp4742;
    assign temp4744 = temp4743 ^ temp4743;
    assign temp4745 = temp4744 ^ temp4744;
    assign temp4746 = temp4745 ^ temp4745;
    assign temp4747 = temp4746 ^ temp4746;
    assign temp4748 = temp4747 ^ temp4747;
    assign temp4749 = temp4748 ^ temp4748;
    assign temp4750 = temp4749 ^ temp4749;
    assign temp4751 = temp4750 ^ temp4750;
    assign temp4752 = temp4751 ^ temp4751;
    assign temp4753 = temp4752 ^ temp4752;
    assign temp4754 = temp4753 ^ temp4753;
    assign temp4755 = temp4754 ^ temp4754;
    assign temp4756 = temp4755 ^ temp4755;
    assign temp4757 = temp4756 ^ temp4756;
    assign temp4758 = temp4757 ^ temp4757;
    assign temp4759 = temp4758 ^ temp4758;
    assign temp4760 = temp4759 ^ temp4759;
    assign temp4761 = temp4760 ^ temp4760;
    assign temp4762 = temp4761 ^ temp4761;
    assign temp4763 = temp4762 ^ temp4762;
    assign temp4764 = temp4763 ^ temp4763;
    assign temp4765 = temp4764 ^ temp4764;
    assign temp4766 = temp4765 ^ temp4765;
    assign temp4767 = temp4766 ^ temp4766;
    assign temp4768 = temp4767 ^ temp4767;
    assign temp4769 = temp4768 ^ temp4768;
    assign temp4770 = temp4769 ^ temp4769;
    assign temp4771 = temp4770 ^ temp4770;
    assign temp4772 = temp4771 ^ temp4771;
    assign temp4773 = temp4772 ^ temp4772;
    assign temp4774 = temp4773 ^ temp4773;
    assign temp4775 = temp4774 ^ temp4774;
    assign temp4776 = temp4775 ^ temp4775;
    assign temp4777 = temp4776 ^ temp4776;
    assign temp4778 = temp4777 ^ temp4777;
    assign temp4779 = temp4778 ^ temp4778;
    assign temp4780 = temp4779 ^ temp4779;
    assign temp4781 = temp4780 ^ temp4780;
    assign temp4782 = temp4781 ^ temp4781;
    assign temp4783 = temp4782 ^ temp4782;
    assign temp4784 = temp4783 ^ temp4783;
    assign temp4785 = temp4784 ^ temp4784;
    assign temp4786 = temp4785 ^ temp4785;
    assign temp4787 = temp4786 ^ temp4786;
    assign temp4788 = temp4787 ^ temp4787;
    assign temp4789 = temp4788 ^ temp4788;
    assign temp4790 = temp4789 ^ temp4789;
    assign temp4791 = temp4790 ^ temp4790;
    assign temp4792 = temp4791 ^ temp4791;
    assign temp4793 = temp4792 ^ temp4792;
    assign temp4794 = temp4793 ^ temp4793;
    assign temp4795 = temp4794 ^ temp4794;
    assign temp4796 = temp4795 ^ temp4795;
    assign temp4797 = temp4796 ^ temp4796;
    assign temp4798 = temp4797 ^ temp4797;
    assign temp4799 = temp4798 ^ temp4798;
    assign temp4800 = temp4799 ^ temp4799;
    assign temp4801 = temp4800 ^ temp4800;
    assign temp4802 = temp4801 ^ temp4801;
    assign temp4803 = temp4802 ^ temp4802;
    assign temp4804 = temp4803 ^ temp4803;
    assign temp4805 = temp4804 ^ temp4804;
    assign temp4806 = temp4805 ^ temp4805;
    assign temp4807 = temp4806 ^ temp4806;
    assign temp4808 = temp4807 ^ temp4807;
    assign temp4809 = temp4808 ^ temp4808;
    assign temp4810 = temp4809 ^ temp4809;
    assign temp4811 = temp4810 ^ temp4810;
    assign temp4812 = temp4811 ^ temp4811;
    assign temp4813 = temp4812 ^ temp4812;
    assign temp4814 = temp4813 ^ temp4813;
    assign temp4815 = temp4814 ^ temp4814;
    assign temp4816 = temp4815 ^ temp4815;
    assign temp4817 = temp4816 ^ temp4816;
    assign temp4818 = temp4817 ^ temp4817;
    assign temp4819 = temp4818 ^ temp4818;
    assign temp4820 = temp4819 ^ temp4819;
    assign temp4821 = temp4820 ^ temp4820;
    assign temp4822 = temp4821 ^ temp4821;
    assign temp4823 = temp4822 ^ temp4822;
    assign temp4824 = temp4823 ^ temp4823;
    assign temp4825 = temp4824 ^ temp4824;
    assign temp4826 = temp4825 ^ temp4825;
    assign temp4827 = temp4826 ^ temp4826;
    assign temp4828 = temp4827 ^ temp4827;
    assign temp4829 = temp4828 ^ temp4828;
    assign temp4830 = temp4829 ^ temp4829;
    assign temp4831 = temp4830 ^ temp4830;
    assign temp4832 = temp4831 ^ temp4831;
    assign temp4833 = temp4832 ^ temp4832;
    assign temp4834 = temp4833 ^ temp4833;
    assign temp4835 = temp4834 ^ temp4834;
    assign temp4836 = temp4835 ^ temp4835;
    assign temp4837 = temp4836 ^ temp4836;
    assign temp4838 = temp4837 ^ temp4837;
    assign temp4839 = temp4838 ^ temp4838;
    assign temp4840 = temp4839 ^ temp4839;
    assign temp4841 = temp4840 ^ temp4840;
    assign temp4842 = temp4841 ^ temp4841;
    assign temp4843 = temp4842 ^ temp4842;
    assign temp4844 = temp4843 ^ temp4843;
    assign temp4845 = temp4844 ^ temp4844;
    assign temp4846 = temp4845 ^ temp4845;
    assign temp4847 = temp4846 ^ temp4846;
    assign temp4848 = temp4847 ^ temp4847;
    assign temp4849 = temp4848 ^ temp4848;
    assign temp4850 = temp4849 ^ temp4849;
    assign temp4851 = temp4850 ^ temp4850;
    assign temp4852 = temp4851 ^ temp4851;
    assign temp4853 = temp4852 ^ temp4852;
    assign temp4854 = temp4853 ^ temp4853;
    assign temp4855 = temp4854 ^ temp4854;
    assign temp4856 = temp4855 ^ temp4855;
    assign temp4857 = temp4856 ^ temp4856;
    assign temp4858 = temp4857 ^ temp4857;
    assign temp4859 = temp4858 ^ temp4858;
    assign temp4860 = temp4859 ^ temp4859;
    assign temp4861 = temp4860 ^ temp4860;
    assign temp4862 = temp4861 ^ temp4861;
    assign temp4863 = temp4862 ^ temp4862;
    assign temp4864 = temp4863 ^ temp4863;
    assign temp4865 = temp4864 ^ temp4864;
    assign temp4866 = temp4865 ^ temp4865;
    assign temp4867 = temp4866 ^ temp4866;
    assign temp4868 = temp4867 ^ temp4867;
    assign temp4869 = temp4868 ^ temp4868;
    assign temp4870 = temp4869 ^ temp4869;
    assign temp4871 = temp4870 ^ temp4870;
    assign temp4872 = temp4871 ^ temp4871;
    assign temp4873 = temp4872 ^ temp4872;
    assign temp4874 = temp4873 ^ temp4873;
    assign temp4875 = temp4874 ^ temp4874;
    assign temp4876 = temp4875 ^ temp4875;
    assign temp4877 = temp4876 ^ temp4876;
    assign temp4878 = temp4877 ^ temp4877;
    assign temp4879 = temp4878 ^ temp4878;
    assign temp4880 = temp4879 ^ temp4879;
    assign temp4881 = temp4880 ^ temp4880;
    assign temp4882 = temp4881 ^ temp4881;
    assign temp4883 = temp4882 ^ temp4882;
    assign temp4884 = temp4883 ^ temp4883;
    assign temp4885 = temp4884 ^ temp4884;
    assign temp4886 = temp4885 ^ temp4885;
    assign temp4887 = temp4886 ^ temp4886;
    assign temp4888 = temp4887 ^ temp4887;
    assign temp4889 = temp4888 ^ temp4888;
    assign temp4890 = temp4889 ^ temp4889;
    assign temp4891 = temp4890 ^ temp4890;
    assign temp4892 = temp4891 ^ temp4891;
    assign temp4893 = temp4892 ^ temp4892;
    assign temp4894 = temp4893 ^ temp4893;
    assign temp4895 = temp4894 ^ temp4894;
    assign temp4896 = temp4895 ^ temp4895;
    assign temp4897 = temp4896 ^ temp4896;
    assign temp4898 = temp4897 ^ temp4897;
    assign temp4899 = temp4898 ^ temp4898;
    assign temp4900 = temp4899 ^ temp4899;
    assign temp4901 = temp4900 ^ temp4900;
    assign temp4902 = temp4901 ^ temp4901;
    assign temp4903 = temp4902 ^ temp4902;
    assign temp4904 = temp4903 ^ temp4903;
    assign temp4905 = temp4904 ^ temp4904;
    assign temp4906 = temp4905 ^ temp4905;
    assign temp4907 = temp4906 ^ temp4906;
    assign temp4908 = temp4907 ^ temp4907;
    assign temp4909 = temp4908 ^ temp4908;
    assign temp4910 = temp4909 ^ temp4909;
    assign temp4911 = temp4910 ^ temp4910;
    assign temp4912 = temp4911 ^ temp4911;
    assign temp4913 = temp4912 ^ temp4912;
    assign temp4914 = temp4913 ^ temp4913;
    assign temp4915 = temp4914 ^ temp4914;
    assign temp4916 = temp4915 ^ temp4915;
    assign temp4917 = temp4916 ^ temp4916;
    assign temp4918 = temp4917 ^ temp4917;
    assign temp4919 = temp4918 ^ temp4918;
    assign temp4920 = temp4919 ^ temp4919;
    assign temp4921 = temp4920 ^ temp4920;
    assign temp4922 = temp4921 ^ temp4921;
    assign temp4923 = temp4922 ^ temp4922;
    assign temp4924 = temp4923 ^ temp4923;
    assign temp4925 = temp4924 ^ temp4924;
    assign temp4926 = temp4925 ^ temp4925;
    assign temp4927 = temp4926 ^ temp4926;
    assign temp4928 = temp4927 ^ temp4927;
    assign temp4929 = temp4928 ^ temp4928;
    assign temp4930 = temp4929 ^ temp4929;
    assign temp4931 = temp4930 ^ temp4930;
    assign temp4932 = temp4931 ^ temp4931;
    assign temp4933 = temp4932 ^ temp4932;
    assign temp4934 = temp4933 ^ temp4933;
    assign temp4935 = temp4934 ^ temp4934;
    assign temp4936 = temp4935 ^ temp4935;
    assign temp4937 = temp4936 ^ temp4936;
    assign temp4938 = temp4937 ^ temp4937;
    assign temp4939 = temp4938 ^ temp4938;
    assign temp4940 = temp4939 ^ temp4939;
    assign temp4941 = temp4940 ^ temp4940;
    assign temp4942 = temp4941 ^ temp4941;
    assign temp4943 = temp4942 ^ temp4942;
    assign temp4944 = temp4943 ^ temp4943;
    assign temp4945 = temp4944 ^ temp4944;
    assign temp4946 = temp4945 ^ temp4945;
    assign temp4947 = temp4946 ^ temp4946;
    assign temp4948 = temp4947 ^ temp4947;
    assign temp4949 = temp4948 ^ temp4948;
    assign temp4950 = temp4949 ^ temp4949;
    assign temp4951 = temp4950 ^ temp4950;
    assign temp4952 = temp4951 ^ temp4951;
    assign temp4953 = temp4952 ^ temp4952;
    assign temp4954 = temp4953 ^ temp4953;
    assign temp4955 = temp4954 ^ temp4954;
    assign temp4956 = temp4955 ^ temp4955;
    assign temp4957 = temp4956 ^ temp4956;
    assign temp4958 = temp4957 ^ temp4957;
    assign temp4959 = temp4958 ^ temp4958;
    assign temp4960 = temp4959 ^ temp4959;
    assign temp4961 = temp4960 ^ temp4960;
    assign temp4962 = temp4961 ^ temp4961;
    assign temp4963 = temp4962 ^ temp4962;
    assign temp4964 = temp4963 ^ temp4963;
    assign temp4965 = temp4964 ^ temp4964;
    assign temp4966 = temp4965 ^ temp4965;
    assign temp4967 = temp4966 ^ temp4966;
    assign temp4968 = temp4967 ^ temp4967;
    assign temp4969 = temp4968 ^ temp4968;
    assign temp4970 = temp4969 ^ temp4969;
    assign temp4971 = temp4970 ^ temp4970;
    assign temp4972 = temp4971 ^ temp4971;
    assign temp4973 = temp4972 ^ temp4972;
    assign temp4974 = temp4973 ^ temp4973;
    assign temp4975 = temp4974 ^ temp4974;
    assign temp4976 = temp4975 ^ temp4975;
    assign temp4977 = temp4976 ^ temp4976;
    assign temp4978 = temp4977 ^ temp4977;
    assign temp4979 = temp4978 ^ temp4978;
    assign temp4980 = temp4979 ^ temp4979;
    assign temp4981 = temp4980 ^ temp4980;
    assign temp4982 = temp4981 ^ temp4981;
    assign temp4983 = temp4982 ^ temp4982;
    assign temp4984 = temp4983 ^ temp4983;
    assign temp4985 = temp4984 ^ temp4984;
    assign temp4986 = temp4985 ^ temp4985;
    assign temp4987 = temp4986 ^ temp4986;
    assign temp4988 = temp4987 ^ temp4987;
    assign temp4989 = temp4988 ^ temp4988;
    assign temp4990 = temp4989 ^ temp4989;
    assign temp4991 = temp4990 ^ temp4990;
    assign temp4992 = temp4991 ^ temp4991;
    assign temp4993 = temp4992 ^ temp4992;
    assign temp4994 = temp4993 ^ temp4993;
    assign temp4995 = temp4994 ^ temp4994;
    assign temp4996 = temp4995 ^ temp4995;
    assign temp4997 = temp4996 ^ temp4996;
    assign temp4998 = temp4997 ^ temp4997;
    assign temp4999 = temp4998 ^ temp4998;
    assign temp5000 = temp4999 ^ temp4999;
    assign temp5001 = temp5000 ^ temp5000;
    assign temp5002 = temp5001 ^ temp5001;
    assign temp5003 = temp5002 ^ temp5002;
    assign temp5004 = temp5003 ^ temp5003;
    assign temp5005 = temp5004 ^ temp5004;
    assign temp5006 = temp5005 ^ temp5005;
    assign temp5007 = temp5006 ^ temp5006;
    assign temp5008 = temp5007 ^ temp5007;
    assign temp5009 = temp5008 ^ temp5008;
    assign temp5010 = temp5009 ^ temp5009;
    assign temp5011 = temp5010 ^ temp5010;
    assign temp5012 = temp5011 ^ temp5011;
    assign temp5013 = temp5012 ^ temp5012;
    assign temp5014 = temp5013 ^ temp5013;
    assign temp5015 = temp5014 ^ temp5014;
    assign temp5016 = temp5015 ^ temp5015;
    assign temp5017 = temp5016 ^ temp5016;
    assign temp5018 = temp5017 ^ temp5017;
    assign temp5019 = temp5018 ^ temp5018;
    assign temp5020 = temp5019 ^ temp5019;
    assign temp5021 = temp5020 ^ temp5020;
    assign temp5022 = temp5021 ^ temp5021;
    assign temp5023 = temp5022 ^ temp5022;
    assign temp5024 = temp5023 ^ temp5023;
    assign temp5025 = temp5024 ^ temp5024;
    assign temp5026 = temp5025 ^ temp5025;
    assign temp5027 = temp5026 ^ temp5026;
    assign temp5028 = temp5027 ^ temp5027;
    assign temp5029 = temp5028 ^ temp5028;
    assign temp5030 = temp5029 ^ temp5029;
    assign temp5031 = temp5030 ^ temp5030;
    assign temp5032 = temp5031 ^ temp5031;
    assign temp5033 = temp5032 ^ temp5032;
    assign temp5034 = temp5033 ^ temp5033;
    assign temp5035 = temp5034 ^ temp5034;
    assign temp5036 = temp5035 ^ temp5035;
    assign temp5037 = temp5036 ^ temp5036;
    assign temp5038 = temp5037 ^ temp5037;
    assign temp5039 = temp5038 ^ temp5038;
    assign temp5040 = temp5039 ^ temp5039;
    assign temp5041 = temp5040 ^ temp5040;
    assign temp5042 = temp5041 ^ temp5041;
    assign temp5043 = temp5042 ^ temp5042;
    assign temp5044 = temp5043 ^ temp5043;
    assign temp5045 = temp5044 ^ temp5044;
    assign temp5046 = temp5045 ^ temp5045;
    assign temp5047 = temp5046 ^ temp5046;
    assign temp5048 = temp5047 ^ temp5047;
    assign temp5049 = temp5048 ^ temp5048;
    assign temp5050 = temp5049 ^ temp5049;
    assign temp5051 = temp5050 ^ temp5050;
    assign temp5052 = temp5051 ^ temp5051;
    assign temp5053 = temp5052 ^ temp5052;
    assign temp5054 = temp5053 ^ temp5053;
    assign temp5055 = temp5054 ^ temp5054;
    assign temp5056 = temp5055 ^ temp5055;
    assign temp5057 = temp5056 ^ temp5056;
    assign temp5058 = temp5057 ^ temp5057;
    assign temp5059 = temp5058 ^ temp5058;
    assign temp5060 = temp5059 ^ temp5059;
    assign temp5061 = temp5060 ^ temp5060;
    assign temp5062 = temp5061 ^ temp5061;
    assign temp5063 = temp5062 ^ temp5062;
    assign temp5064 = temp5063 ^ temp5063;
    assign temp5065 = temp5064 ^ temp5064;
    assign temp5066 = temp5065 ^ temp5065;
    assign temp5067 = temp5066 ^ temp5066;
    assign temp5068 = temp5067 ^ temp5067;
    assign temp5069 = temp5068 ^ temp5068;
    assign temp5070 = temp5069 ^ temp5069;
    assign temp5071 = temp5070 ^ temp5070;
    assign temp5072 = temp5071 ^ temp5071;
    assign temp5073 = temp5072 ^ temp5072;
    assign temp5074 = temp5073 ^ temp5073;
    assign temp5075 = temp5074 ^ temp5074;
    assign temp5076 = temp5075 ^ temp5075;
    assign temp5077 = temp5076 ^ temp5076;
    assign temp5078 = temp5077 ^ temp5077;
    assign temp5079 = temp5078 ^ temp5078;
    assign temp5080 = temp5079 ^ temp5079;
    assign temp5081 = temp5080 ^ temp5080;
    assign temp5082 = temp5081 ^ temp5081;
    assign temp5083 = temp5082 ^ temp5082;
    assign temp5084 = temp5083 ^ temp5083;
    assign temp5085 = temp5084 ^ temp5084;
    assign temp5086 = temp5085 ^ temp5085;
    assign temp5087 = temp5086 ^ temp5086;
    assign temp5088 = temp5087 ^ temp5087;
    assign temp5089 = temp5088 ^ temp5088;
    assign temp5090 = temp5089 ^ temp5089;
    assign temp5091 = temp5090 ^ temp5090;
    assign temp5092 = temp5091 ^ temp5091;
    assign temp5093 = temp5092 ^ temp5092;
    assign temp5094 = temp5093 ^ temp5093;
    assign temp5095 = temp5094 ^ temp5094;
    assign temp5096 = temp5095 ^ temp5095;
    assign temp5097 = temp5096 ^ temp5096;
    assign temp5098 = temp5097 ^ temp5097;
    assign temp5099 = temp5098 ^ temp5098;
    assign temp5100 = temp5099 ^ temp5099;
    assign temp5101 = temp5100 ^ temp5100;
    assign temp5102 = temp5101 ^ temp5101;
    assign temp5103 = temp5102 ^ temp5102;
    assign temp5104 = temp5103 ^ temp5103;
    assign temp5105 = temp5104 ^ temp5104;
    assign temp5106 = temp5105 ^ temp5105;
    assign temp5107 = temp5106 ^ temp5106;
    assign temp5108 = temp5107 ^ temp5107;
    assign temp5109 = temp5108 ^ temp5108;
    assign temp5110 = temp5109 ^ temp5109;
    assign temp5111 = temp5110 ^ temp5110;
    assign temp5112 = temp5111 ^ temp5111;
    assign temp5113 = temp5112 ^ temp5112;
    assign temp5114 = temp5113 ^ temp5113;
    assign temp5115 = temp5114 ^ temp5114;
    assign temp5116 = temp5115 ^ temp5115;
    assign temp5117 = temp5116 ^ temp5116;
    assign temp5118 = temp5117 ^ temp5117;
    assign temp5119 = temp5118 ^ temp5118;
    assign temp5120 = temp5119 ^ temp5119;
    assign temp5121 = temp5120 ^ temp5120;
    assign temp5122 = temp5121 ^ temp5121;
    assign temp5123 = temp5122 ^ temp5122;
    assign temp5124 = temp5123 ^ temp5123;
    assign temp5125 = temp5124 ^ temp5124;
    assign temp5126 = temp5125 ^ temp5125;
    assign temp5127 = temp5126 ^ temp5126;
    assign temp5128 = temp5127 ^ temp5127;
    assign temp5129 = temp5128 ^ temp5128;
    assign temp5130 = temp5129 ^ temp5129;
    assign temp5131 = temp5130 ^ temp5130;
    assign temp5132 = temp5131 ^ temp5131;
    assign temp5133 = temp5132 ^ temp5132;
    assign temp5134 = temp5133 ^ temp5133;
    assign temp5135 = temp5134 ^ temp5134;
    assign temp5136 = temp5135 ^ temp5135;
    assign temp5137 = temp5136 ^ temp5136;
    assign temp5138 = temp5137 ^ temp5137;
    assign temp5139 = temp5138 ^ temp5138;
    assign temp5140 = temp5139 ^ temp5139;
    assign temp5141 = temp5140 ^ temp5140;
    assign temp5142 = temp5141 ^ temp5141;
    assign temp5143 = temp5142 ^ temp5142;
    assign temp5144 = temp5143 ^ temp5143;
    assign temp5145 = temp5144 ^ temp5144;
    assign temp5146 = temp5145 ^ temp5145;
    assign temp5147 = temp5146 ^ temp5146;
    assign temp5148 = temp5147 ^ temp5147;
    assign temp5149 = temp5148 ^ temp5148;
    assign temp5150 = temp5149 ^ temp5149;
    assign temp5151 = temp5150 ^ temp5150;
    assign temp5152 = temp5151 ^ temp5151;
    assign temp5153 = temp5152 ^ temp5152;
    assign temp5154 = temp5153 ^ temp5153;
    assign temp5155 = temp5154 ^ temp5154;
    assign temp5156 = temp5155 ^ temp5155;
    assign temp5157 = temp5156 ^ temp5156;
    assign temp5158 = temp5157 ^ temp5157;
    assign temp5159 = temp5158 ^ temp5158;
    assign temp5160 = temp5159 ^ temp5159;
    assign temp5161 = temp5160 ^ temp5160;
    assign temp5162 = temp5161 ^ temp5161;
    assign temp5163 = temp5162 ^ temp5162;
    assign temp5164 = temp5163 ^ temp5163;
    assign temp5165 = temp5164 ^ temp5164;
    assign temp5166 = temp5165 ^ temp5165;
    assign temp5167 = temp5166 ^ temp5166;
    assign temp5168 = temp5167 ^ temp5167;
    assign temp5169 = temp5168 ^ temp5168;
    assign temp5170 = temp5169 ^ temp5169;
    assign temp5171 = temp5170 ^ temp5170;
    assign temp5172 = temp5171 ^ temp5171;
    assign temp5173 = temp5172 ^ temp5172;
    assign temp5174 = temp5173 ^ temp5173;
    assign temp5175 = temp5174 ^ temp5174;
    assign temp5176 = temp5175 ^ temp5175;
    assign temp5177 = temp5176 ^ temp5176;
    assign temp5178 = temp5177 ^ temp5177;
    assign temp5179 = temp5178 ^ temp5178;
    assign temp5180 = temp5179 ^ temp5179;
    assign temp5181 = temp5180 ^ temp5180;
    assign temp5182 = temp5181 ^ temp5181;
    assign temp5183 = temp5182 ^ temp5182;
    assign temp5184 = temp5183 ^ temp5183;
    assign temp5185 = temp5184 ^ temp5184;
    assign temp5186 = temp5185 ^ temp5185;
    assign temp5187 = temp5186 ^ temp5186;
    assign temp5188 = temp5187 ^ temp5187;
    assign temp5189 = temp5188 ^ temp5188;
    assign temp5190 = temp5189 ^ temp5189;
    assign temp5191 = temp5190 ^ temp5190;
    assign temp5192 = temp5191 ^ temp5191;
    assign temp5193 = temp5192 ^ temp5192;
    assign temp5194 = temp5193 ^ temp5193;
    assign temp5195 = temp5194 ^ temp5194;
    assign temp5196 = temp5195 ^ temp5195;
    assign temp5197 = temp5196 ^ temp5196;
    assign temp5198 = temp5197 ^ temp5197;
    assign temp5199 = temp5198 ^ temp5198;
    assign temp5200 = temp5199 ^ temp5199;
    assign temp5201 = temp5200 ^ temp5200;
    assign temp5202 = temp5201 ^ temp5201;
    assign temp5203 = temp5202 ^ temp5202;
    assign temp5204 = temp5203 ^ temp5203;
    assign temp5205 = temp5204 ^ temp5204;
    assign temp5206 = temp5205 ^ temp5205;
    assign temp5207 = temp5206 ^ temp5206;
    assign temp5208 = temp5207 ^ temp5207;
    assign temp5209 = temp5208 ^ temp5208;
    assign temp5210 = temp5209 ^ temp5209;
    assign temp5211 = temp5210 ^ temp5210;
    assign temp5212 = temp5211 ^ temp5211;
    assign temp5213 = temp5212 ^ temp5212;
    assign temp5214 = temp5213 ^ temp5213;
    assign temp5215 = temp5214 ^ temp5214;
    assign temp5216 = temp5215 ^ temp5215;
    assign temp5217 = temp5216 ^ temp5216;
    assign temp5218 = temp5217 ^ temp5217;
    assign temp5219 = temp5218 ^ temp5218;
    assign temp5220 = temp5219 ^ temp5219;
    assign temp5221 = temp5220 ^ temp5220;
    assign temp5222 = temp5221 ^ temp5221;
    assign temp5223 = temp5222 ^ temp5222;
    assign temp5224 = temp5223 ^ temp5223;
    assign temp5225 = temp5224 ^ temp5224;
    assign temp5226 = temp5225 ^ temp5225;
    assign temp5227 = temp5226 ^ temp5226;
    assign temp5228 = temp5227 ^ temp5227;
    assign temp5229 = temp5228 ^ temp5228;
    assign temp5230 = temp5229 ^ temp5229;
    assign temp5231 = temp5230 ^ temp5230;
    assign temp5232 = temp5231 ^ temp5231;
    assign temp5233 = temp5232 ^ temp5232;
    assign temp5234 = temp5233 ^ temp5233;
    assign temp5235 = temp5234 ^ temp5234;
    assign temp5236 = temp5235 ^ temp5235;
    assign temp5237 = temp5236 ^ temp5236;
    assign temp5238 = temp5237 ^ temp5237;
    assign temp5239 = temp5238 ^ temp5238;
    assign temp5240 = temp5239 ^ temp5239;
    assign temp5241 = temp5240 ^ temp5240;
    assign temp5242 = temp5241 ^ temp5241;
    assign temp5243 = temp5242 ^ temp5242;
    assign temp5244 = temp5243 ^ temp5243;
    assign temp5245 = temp5244 ^ temp5244;
    assign temp5246 = temp5245 ^ temp5245;
    assign temp5247 = temp5246 ^ temp5246;
    assign temp5248 = temp5247 ^ temp5247;
    assign temp5249 = temp5248 ^ temp5248;
    assign temp5250 = temp5249 ^ temp5249;
    assign temp5251 = temp5250 ^ temp5250;
    assign temp5252 = temp5251 ^ temp5251;
    assign temp5253 = temp5252 ^ temp5252;
    assign temp5254 = temp5253 ^ temp5253;
    assign temp5255 = temp5254 ^ temp5254;
    assign temp5256 = temp5255 ^ temp5255;
    assign temp5257 = temp5256 ^ temp5256;
    assign temp5258 = temp5257 ^ temp5257;
    assign temp5259 = temp5258 ^ temp5258;
    assign temp5260 = temp5259 ^ temp5259;
    assign temp5261 = temp5260 ^ temp5260;
    assign temp5262 = temp5261 ^ temp5261;
    assign temp5263 = temp5262 ^ temp5262;
    assign temp5264 = temp5263 ^ temp5263;
    assign temp5265 = temp5264 ^ temp5264;
    assign temp5266 = temp5265 ^ temp5265;
    assign temp5267 = temp5266 ^ temp5266;
    assign temp5268 = temp5267 ^ temp5267;
    assign temp5269 = temp5268 ^ temp5268;
    assign temp5270 = temp5269 ^ temp5269;
    assign temp5271 = temp5270 ^ temp5270;
    assign temp5272 = temp5271 ^ temp5271;
    assign temp5273 = temp5272 ^ temp5272;
    assign temp5274 = temp5273 ^ temp5273;
    assign temp5275 = temp5274 ^ temp5274;
    assign temp5276 = temp5275 ^ temp5275;
    assign temp5277 = temp5276 ^ temp5276;
    assign temp5278 = temp5277 ^ temp5277;
    assign temp5279 = temp5278 ^ temp5278;
    assign temp5280 = temp5279 ^ temp5279;
    assign temp5281 = temp5280 ^ temp5280;
    assign temp5282 = temp5281 ^ temp5281;
    assign temp5283 = temp5282 ^ temp5282;
    assign temp5284 = temp5283 ^ temp5283;
    assign temp5285 = temp5284 ^ temp5284;
    assign temp5286 = temp5285 ^ temp5285;
    assign temp5287 = temp5286 ^ temp5286;
    assign temp5288 = temp5287 ^ temp5287;
    assign temp5289 = temp5288 ^ temp5288;
    assign temp5290 = temp5289 ^ temp5289;
    assign temp5291 = temp5290 ^ temp5290;
    assign temp5292 = temp5291 ^ temp5291;
    assign temp5293 = temp5292 ^ temp5292;
    assign temp5294 = temp5293 ^ temp5293;
    assign temp5295 = temp5294 ^ temp5294;
    assign temp5296 = temp5295 ^ temp5295;
    assign temp5297 = temp5296 ^ temp5296;
    assign temp5298 = temp5297 ^ temp5297;
    assign temp5299 = temp5298 ^ temp5298;
    assign temp5300 = temp5299 ^ temp5299;
    assign temp5301 = temp5300 ^ temp5300;
    assign temp5302 = temp5301 ^ temp5301;
    assign temp5303 = temp5302 ^ temp5302;
    assign temp5304 = temp5303 ^ temp5303;
    assign temp5305 = temp5304 ^ temp5304;
    assign temp5306 = temp5305 ^ temp5305;
    assign temp5307 = temp5306 ^ temp5306;
    assign temp5308 = temp5307 ^ temp5307;
    assign temp5309 = temp5308 ^ temp5308;
    assign temp5310 = temp5309 ^ temp5309;
    assign temp5311 = temp5310 ^ temp5310;
    assign temp5312 = temp5311 ^ temp5311;
    assign temp5313 = temp5312 ^ temp5312;
    assign temp5314 = temp5313 ^ temp5313;
    assign temp5315 = temp5314 ^ temp5314;
    assign temp5316 = temp5315 ^ temp5315;
    assign temp5317 = temp5316 ^ temp5316;
    assign temp5318 = temp5317 ^ temp5317;
    assign temp5319 = temp5318 ^ temp5318;
    assign temp5320 = temp5319 ^ temp5319;
    assign temp5321 = temp5320 ^ temp5320;
    assign temp5322 = temp5321 ^ temp5321;
    assign temp5323 = temp5322 ^ temp5322;
    assign temp5324 = temp5323 ^ temp5323;
    assign temp5325 = temp5324 ^ temp5324;
    assign temp5326 = temp5325 ^ temp5325;
    assign temp5327 = temp5326 ^ temp5326;
    assign temp5328 = temp5327 ^ temp5327;
    assign temp5329 = temp5328 ^ temp5328;
    assign temp5330 = temp5329 ^ temp5329;
    assign temp5331 = temp5330 ^ temp5330;
    assign temp5332 = temp5331 ^ temp5331;
    assign temp5333 = temp5332 ^ temp5332;
    assign temp5334 = temp5333 ^ temp5333;
    assign temp5335 = temp5334 ^ temp5334;
    assign temp5336 = temp5335 ^ temp5335;
    assign temp5337 = temp5336 ^ temp5336;
    assign temp5338 = temp5337 ^ temp5337;
    assign temp5339 = temp5338 ^ temp5338;
    assign temp5340 = temp5339 ^ temp5339;
    assign temp5341 = temp5340 ^ temp5340;
    assign temp5342 = temp5341 ^ temp5341;
    assign temp5343 = temp5342 ^ temp5342;
    assign temp5344 = temp5343 ^ temp5343;
    assign temp5345 = temp5344 ^ temp5344;
    assign temp5346 = temp5345 ^ temp5345;
    assign temp5347 = temp5346 ^ temp5346;
    assign temp5348 = temp5347 ^ temp5347;
    assign temp5349 = temp5348 ^ temp5348;
    assign temp5350 = temp5349 ^ temp5349;
    assign temp5351 = temp5350 ^ temp5350;
    assign temp5352 = temp5351 ^ temp5351;
    assign temp5353 = temp5352 ^ temp5352;
    assign temp5354 = temp5353 ^ temp5353;
    assign temp5355 = temp5354 ^ temp5354;
    assign temp5356 = temp5355 ^ temp5355;
    assign temp5357 = temp5356 ^ temp5356;
    assign temp5358 = temp5357 ^ temp5357;
    assign temp5359 = temp5358 ^ temp5358;
    assign temp5360 = temp5359 ^ temp5359;
    assign temp5361 = temp5360 ^ temp5360;
    assign temp5362 = temp5361 ^ temp5361;
    assign temp5363 = temp5362 ^ temp5362;
    assign temp5364 = temp5363 ^ temp5363;
    assign temp5365 = temp5364 ^ temp5364;
    assign temp5366 = temp5365 ^ temp5365;
    assign temp5367 = temp5366 ^ temp5366;
    assign temp5368 = temp5367 ^ temp5367;
    assign temp5369 = temp5368 ^ temp5368;
    assign temp5370 = temp5369 ^ temp5369;
    assign temp5371 = temp5370 ^ temp5370;
    assign temp5372 = temp5371 ^ temp5371;
    assign temp5373 = temp5372 ^ temp5372;
    assign temp5374 = temp5373 ^ temp5373;
    assign temp5375 = temp5374 ^ temp5374;
    assign temp5376 = temp5375 ^ temp5375;
    assign temp5377 = temp5376 ^ temp5376;
    assign temp5378 = temp5377 ^ temp5377;
    assign temp5379 = temp5378 ^ temp5378;
    assign temp5380 = temp5379 ^ temp5379;
    assign temp5381 = temp5380 ^ temp5380;
    assign temp5382 = temp5381 ^ temp5381;
    assign temp5383 = temp5382 ^ temp5382;
    assign temp5384 = temp5383 ^ temp5383;
    assign temp5385 = temp5384 ^ temp5384;
    assign temp5386 = temp5385 ^ temp5385;
    assign temp5387 = temp5386 ^ temp5386;
    assign temp5388 = temp5387 ^ temp5387;
    assign temp5389 = temp5388 ^ temp5388;
    assign temp5390 = temp5389 ^ temp5389;
    assign temp5391 = temp5390 ^ temp5390;
    assign temp5392 = temp5391 ^ temp5391;
    assign temp5393 = temp5392 ^ temp5392;
    assign temp5394 = temp5393 ^ temp5393;
    assign temp5395 = temp5394 ^ temp5394;
    assign temp5396 = temp5395 ^ temp5395;
    assign temp5397 = temp5396 ^ temp5396;
    assign temp5398 = temp5397 ^ temp5397;
    assign temp5399 = temp5398 ^ temp5398;
    assign temp5400 = temp5399 ^ temp5399;
    assign temp5401 = temp5400 ^ temp5400;
    assign temp5402 = temp5401 ^ temp5401;
    assign temp5403 = temp5402 ^ temp5402;
    assign temp5404 = temp5403 ^ temp5403;
    assign temp5405 = temp5404 ^ temp5404;
    assign temp5406 = temp5405 ^ temp5405;
    assign temp5407 = temp5406 ^ temp5406;
    assign temp5408 = temp5407 ^ temp5407;
    assign temp5409 = temp5408 ^ temp5408;
    assign temp5410 = temp5409 ^ temp5409;
    assign temp5411 = temp5410 ^ temp5410;
    assign temp5412 = temp5411 ^ temp5411;
    assign temp5413 = temp5412 ^ temp5412;
    assign temp5414 = temp5413 ^ temp5413;
    assign temp5415 = temp5414 ^ temp5414;
    assign temp5416 = temp5415 ^ temp5415;
    assign temp5417 = temp5416 ^ temp5416;
    assign temp5418 = temp5417 ^ temp5417;
    assign temp5419 = temp5418 ^ temp5418;
    assign temp5420 = temp5419 ^ temp5419;
    assign temp5421 = temp5420 ^ temp5420;
    assign temp5422 = temp5421 ^ temp5421;
    assign temp5423 = temp5422 ^ temp5422;
    assign temp5424 = temp5423 ^ temp5423;
    assign temp5425 = temp5424 ^ temp5424;
    assign temp5426 = temp5425 ^ temp5425;
    assign temp5427 = temp5426 ^ temp5426;
    assign temp5428 = temp5427 ^ temp5427;
    assign temp5429 = temp5428 ^ temp5428;
    assign temp5430 = temp5429 ^ temp5429;
    assign temp5431 = temp5430 ^ temp5430;
    assign temp5432 = temp5431 ^ temp5431;
    assign temp5433 = temp5432 ^ temp5432;
    assign temp5434 = temp5433 ^ temp5433;
    assign temp5435 = temp5434 ^ temp5434;
    assign temp5436 = temp5435 ^ temp5435;
    assign temp5437 = temp5436 ^ temp5436;
    assign temp5438 = temp5437 ^ temp5437;
    assign temp5439 = temp5438 ^ temp5438;
    assign temp5440 = temp5439 ^ temp5439;
    assign temp5441 = temp5440 ^ temp5440;
    assign temp5442 = temp5441 ^ temp5441;
    assign temp5443 = temp5442 ^ temp5442;
    assign temp5444 = temp5443 ^ temp5443;
    assign temp5445 = temp5444 ^ temp5444;
    assign temp5446 = temp5445 ^ temp5445;
    assign temp5447 = temp5446 ^ temp5446;
    assign temp5448 = temp5447 ^ temp5447;
    assign temp5449 = temp5448 ^ temp5448;
    assign temp5450 = temp5449 ^ temp5449;
    assign temp5451 = temp5450 ^ temp5450;
    assign temp5452 = temp5451 ^ temp5451;
    assign temp5453 = temp5452 ^ temp5452;
    assign temp5454 = temp5453 ^ temp5453;
    assign temp5455 = temp5454 ^ temp5454;
    assign temp5456 = temp5455 ^ temp5455;
    assign temp5457 = temp5456 ^ temp5456;
    assign temp5458 = temp5457 ^ temp5457;
    assign temp5459 = temp5458 ^ temp5458;
    assign temp5460 = temp5459 ^ temp5459;
    assign temp5461 = temp5460 ^ temp5460;
    assign temp5462 = temp5461 ^ temp5461;
    assign temp5463 = temp5462 ^ temp5462;
    assign temp5464 = temp5463 ^ temp5463;
    assign temp5465 = temp5464 ^ temp5464;
    assign temp5466 = temp5465 ^ temp5465;
    assign temp5467 = temp5466 ^ temp5466;
    assign temp5468 = temp5467 ^ temp5467;
    assign temp5469 = temp5468 ^ temp5468;
    assign temp5470 = temp5469 ^ temp5469;
    assign temp5471 = temp5470 ^ temp5470;
    assign temp5472 = temp5471 ^ temp5471;
    assign temp5473 = temp5472 ^ temp5472;
    assign temp5474 = temp5473 ^ temp5473;
    assign temp5475 = temp5474 ^ temp5474;
    assign temp5476 = temp5475 ^ temp5475;
    assign temp5477 = temp5476 ^ temp5476;
    assign temp5478 = temp5477 ^ temp5477;
    assign temp5479 = temp5478 ^ temp5478;
    assign temp5480 = temp5479 ^ temp5479;
    assign temp5481 = temp5480 ^ temp5480;
    assign temp5482 = temp5481 ^ temp5481;
    assign temp5483 = temp5482 ^ temp5482;
    assign temp5484 = temp5483 ^ temp5483;
    assign temp5485 = temp5484 ^ temp5484;
    assign temp5486 = temp5485 ^ temp5485;
    assign temp5487 = temp5486 ^ temp5486;
    assign temp5488 = temp5487 ^ temp5487;
    assign temp5489 = temp5488 ^ temp5488;
    assign temp5490 = temp5489 ^ temp5489;
    assign temp5491 = temp5490 ^ temp5490;
    assign temp5492 = temp5491 ^ temp5491;
    assign temp5493 = temp5492 ^ temp5492;
    assign temp5494 = temp5493 ^ temp5493;
    assign temp5495 = temp5494 ^ temp5494;
    assign temp5496 = temp5495 ^ temp5495;
    assign temp5497 = temp5496 ^ temp5496;
    assign temp5498 = temp5497 ^ temp5497;
    assign temp5499 = temp5498 ^ temp5498;
    assign temp5500 = temp5499 ^ temp5499;
    assign temp5501 = temp5500 ^ temp5500;
    assign temp5502 = temp5501 ^ temp5501;
    assign temp5503 = temp5502 ^ temp5502;
    assign temp5504 = temp5503 ^ temp5503;
    assign temp5505 = temp5504 ^ temp5504;
    assign temp5506 = temp5505 ^ temp5505;
    assign temp5507 = temp5506 ^ temp5506;
    assign temp5508 = temp5507 ^ temp5507;
    assign temp5509 = temp5508 ^ temp5508;
    assign temp5510 = temp5509 ^ temp5509;
    assign temp5511 = temp5510 ^ temp5510;
    assign temp5512 = temp5511 ^ temp5511;
    assign temp5513 = temp5512 ^ temp5512;
    assign temp5514 = temp5513 ^ temp5513;
    assign temp5515 = temp5514 ^ temp5514;
    assign temp5516 = temp5515 ^ temp5515;
    assign temp5517 = temp5516 ^ temp5516;
    assign temp5518 = temp5517 ^ temp5517;
    assign temp5519 = temp5518 ^ temp5518;
    assign temp5520 = temp5519 ^ temp5519;
    assign temp5521 = temp5520 ^ temp5520;
    assign temp5522 = temp5521 ^ temp5521;
    assign temp5523 = temp5522 ^ temp5522;
    assign temp5524 = temp5523 ^ temp5523;
    assign temp5525 = temp5524 ^ temp5524;
    assign temp5526 = temp5525 ^ temp5525;
    assign temp5527 = temp5526 ^ temp5526;
    assign temp5528 = temp5527 ^ temp5527;
    assign temp5529 = temp5528 ^ temp5528;
    assign temp5530 = temp5529 ^ temp5529;
    assign temp5531 = temp5530 ^ temp5530;
    assign temp5532 = temp5531 ^ temp5531;
    assign temp5533 = temp5532 ^ temp5532;
    assign temp5534 = temp5533 ^ temp5533;
    assign temp5535 = temp5534 ^ temp5534;
    assign temp5536 = temp5535 ^ temp5535;
    assign temp5537 = temp5536 ^ temp5536;
    assign temp5538 = temp5537 ^ temp5537;
    assign temp5539 = temp5538 ^ temp5538;
    assign temp5540 = temp5539 ^ temp5539;
    assign temp5541 = temp5540 ^ temp5540;
    assign temp5542 = temp5541 ^ temp5541;
    assign temp5543 = temp5542 ^ temp5542;
    assign temp5544 = temp5543 ^ temp5543;
    assign temp5545 = temp5544 ^ temp5544;
    assign temp5546 = temp5545 ^ temp5545;
    assign temp5547 = temp5546 ^ temp5546;
    assign temp5548 = temp5547 ^ temp5547;
    assign temp5549 = temp5548 ^ temp5548;
    assign temp5550 = temp5549 ^ temp5549;
    assign temp5551 = temp5550 ^ temp5550;
    assign temp5552 = temp5551 ^ temp5551;
    assign temp5553 = temp5552 ^ temp5552;
    assign temp5554 = temp5553 ^ temp5553;
    assign temp5555 = temp5554 ^ temp5554;
    assign temp5556 = temp5555 ^ temp5555;
    assign temp5557 = temp5556 ^ temp5556;
    assign temp5558 = temp5557 ^ temp5557;
    assign temp5559 = temp5558 ^ temp5558;
    assign temp5560 = temp5559 ^ temp5559;
    assign temp5561 = temp5560 ^ temp5560;
    assign temp5562 = temp5561 ^ temp5561;
    assign temp5563 = temp5562 ^ temp5562;
    assign temp5564 = temp5563 ^ temp5563;
    assign temp5565 = temp5564 ^ temp5564;
    assign temp5566 = temp5565 ^ temp5565;
    assign temp5567 = temp5566 ^ temp5566;
    assign temp5568 = temp5567 ^ temp5567;
    assign temp5569 = temp5568 ^ temp5568;
    assign temp5570 = temp5569 ^ temp5569;
    assign temp5571 = temp5570 ^ temp5570;
    assign temp5572 = temp5571 ^ temp5571;
    assign temp5573 = temp5572 ^ temp5572;
    assign temp5574 = temp5573 ^ temp5573;
    assign temp5575 = temp5574 ^ temp5574;
    assign temp5576 = temp5575 ^ temp5575;
    assign temp5577 = temp5576 ^ temp5576;
    assign temp5578 = temp5577 ^ temp5577;
    assign temp5579 = temp5578 ^ temp5578;
    assign temp5580 = temp5579 ^ temp5579;
    assign temp5581 = temp5580 ^ temp5580;
    assign temp5582 = temp5581 ^ temp5581;
    assign temp5583 = temp5582 ^ temp5582;
    assign temp5584 = temp5583 ^ temp5583;
    assign temp5585 = temp5584 ^ temp5584;
    assign temp5586 = temp5585 ^ temp5585;
    assign temp5587 = temp5586 ^ temp5586;
    assign temp5588 = temp5587 ^ temp5587;
    assign temp5589 = temp5588 ^ temp5588;
    assign temp5590 = temp5589 ^ temp5589;
    assign temp5591 = temp5590 ^ temp5590;
    assign temp5592 = temp5591 ^ temp5591;
    assign temp5593 = temp5592 ^ temp5592;
    assign temp5594 = temp5593 ^ temp5593;
    assign temp5595 = temp5594 ^ temp5594;
    assign temp5596 = temp5595 ^ temp5595;
    assign temp5597 = temp5596 ^ temp5596;
    assign temp5598 = temp5597 ^ temp5597;
    assign temp5599 = temp5598 ^ temp5598;
    assign temp5600 = temp5599 ^ temp5599;
    assign temp5601 = temp5600 ^ temp5600;
    assign temp5602 = temp5601 ^ temp5601;
    assign temp5603 = temp5602 ^ temp5602;
    assign temp5604 = temp5603 ^ temp5603;
    assign temp5605 = temp5604 ^ temp5604;
    assign temp5606 = temp5605 ^ temp5605;
    assign temp5607 = temp5606 ^ temp5606;
    assign temp5608 = temp5607 ^ temp5607;
    assign temp5609 = temp5608 ^ temp5608;
    assign temp5610 = temp5609 ^ temp5609;
    assign temp5611 = temp5610 ^ temp5610;
    assign temp5612 = temp5611 ^ temp5611;
    assign temp5613 = temp5612 ^ temp5612;
    assign temp5614 = temp5613 ^ temp5613;
    assign temp5615 = temp5614 ^ temp5614;
    assign temp5616 = temp5615 ^ temp5615;
    assign temp5617 = temp5616 ^ temp5616;
    assign temp5618 = temp5617 ^ temp5617;
    assign temp5619 = temp5618 ^ temp5618;
    assign temp5620 = temp5619 ^ temp5619;
    assign temp5621 = temp5620 ^ temp5620;
    assign temp5622 = temp5621 ^ temp5621;
    assign temp5623 = temp5622 ^ temp5622;
    assign temp5624 = temp5623 ^ temp5623;
    assign temp5625 = temp5624 ^ temp5624;
    assign temp5626 = temp5625 ^ temp5625;
    assign temp5627 = temp5626 ^ temp5626;
    assign temp5628 = temp5627 ^ temp5627;
    assign temp5629 = temp5628 ^ temp5628;
    assign temp5630 = temp5629 ^ temp5629;
    assign temp5631 = temp5630 ^ temp5630;
    assign temp5632 = temp5631 ^ temp5631;
    assign temp5633 = temp5632 ^ temp5632;
    assign temp5634 = temp5633 ^ temp5633;
    assign temp5635 = temp5634 ^ temp5634;
    assign temp5636 = temp5635 ^ temp5635;
    assign temp5637 = temp5636 ^ temp5636;
    assign temp5638 = temp5637 ^ temp5637;
    assign temp5639 = temp5638 ^ temp5638;
    assign temp5640 = temp5639 ^ temp5639;
    assign temp5641 = temp5640 ^ temp5640;
    assign temp5642 = temp5641 ^ temp5641;
    assign temp5643 = temp5642 ^ temp5642;
    assign temp5644 = temp5643 ^ temp5643;
    assign temp5645 = temp5644 ^ temp5644;
    assign temp5646 = temp5645 ^ temp5645;
    assign temp5647 = temp5646 ^ temp5646;
    assign temp5648 = temp5647 ^ temp5647;
    assign temp5649 = temp5648 ^ temp5648;
    assign temp5650 = temp5649 ^ temp5649;
    assign temp5651 = temp5650 ^ temp5650;
    assign temp5652 = temp5651 ^ temp5651;
    assign temp5653 = temp5652 ^ temp5652;
    assign temp5654 = temp5653 ^ temp5653;
    assign temp5655 = temp5654 ^ temp5654;
    assign temp5656 = temp5655 ^ temp5655;
    assign temp5657 = temp5656 ^ temp5656;
    assign temp5658 = temp5657 ^ temp5657;
    assign temp5659 = temp5658 ^ temp5658;
    assign temp5660 = temp5659 ^ temp5659;
    assign temp5661 = temp5660 ^ temp5660;
    assign temp5662 = temp5661 ^ temp5661;
    assign temp5663 = temp5662 ^ temp5662;
    assign temp5664 = temp5663 ^ temp5663;
    assign temp5665 = temp5664 ^ temp5664;
    assign temp5666 = temp5665 ^ temp5665;
    assign temp5667 = temp5666 ^ temp5666;
    assign temp5668 = temp5667 ^ temp5667;
    assign temp5669 = temp5668 ^ temp5668;
    assign temp5670 = temp5669 ^ temp5669;
    assign temp5671 = temp5670 ^ temp5670;
    assign temp5672 = temp5671 ^ temp5671;
    assign temp5673 = temp5672 ^ temp5672;
    assign temp5674 = temp5673 ^ temp5673;
    assign temp5675 = temp5674 ^ temp5674;
    assign temp5676 = temp5675 ^ temp5675;
    assign temp5677 = temp5676 ^ temp5676;
    assign temp5678 = temp5677 ^ temp5677;
    assign temp5679 = temp5678 ^ temp5678;
    assign temp5680 = temp5679 ^ temp5679;
    assign temp5681 = temp5680 ^ temp5680;
    assign temp5682 = temp5681 ^ temp5681;
    assign temp5683 = temp5682 ^ temp5682;
    assign temp5684 = temp5683 ^ temp5683;
    assign temp5685 = temp5684 ^ temp5684;
    assign temp5686 = temp5685 ^ temp5685;
    assign temp5687 = temp5686 ^ temp5686;
    assign temp5688 = temp5687 ^ temp5687;
    assign temp5689 = temp5688 ^ temp5688;
    assign temp5690 = temp5689 ^ temp5689;
    assign temp5691 = temp5690 ^ temp5690;
    assign temp5692 = temp5691 ^ temp5691;
    assign temp5693 = temp5692 ^ temp5692;
    assign temp5694 = temp5693 ^ temp5693;
    assign temp5695 = temp5694 ^ temp5694;
    assign temp5696 = temp5695 ^ temp5695;
    assign temp5697 = temp5696 ^ temp5696;
    assign temp5698 = temp5697 ^ temp5697;
    assign temp5699 = temp5698 ^ temp5698;
    assign temp5700 = temp5699 ^ temp5699;
    assign temp5701 = temp5700 ^ temp5700;
    assign temp5702 = temp5701 ^ temp5701;
    assign temp5703 = temp5702 ^ temp5702;
    assign temp5704 = temp5703 ^ temp5703;
    assign temp5705 = temp5704 ^ temp5704;
    assign temp5706 = temp5705 ^ temp5705;
    assign temp5707 = temp5706 ^ temp5706;
    assign temp5708 = temp5707 ^ temp5707;
    assign temp5709 = temp5708 ^ temp5708;
    assign temp5710 = temp5709 ^ temp5709;
    assign temp5711 = temp5710 ^ temp5710;
    assign temp5712 = temp5711 ^ temp5711;
    assign temp5713 = temp5712 ^ temp5712;
    assign temp5714 = temp5713 ^ temp5713;
    assign temp5715 = temp5714 ^ temp5714;
    assign temp5716 = temp5715 ^ temp5715;
    assign temp5717 = temp5716 ^ temp5716;
    assign temp5718 = temp5717 ^ temp5717;
    assign temp5719 = temp5718 ^ temp5718;
    assign temp5720 = temp5719 ^ temp5719;
    assign temp5721 = temp5720 ^ temp5720;
    assign temp5722 = temp5721 ^ temp5721;
    assign temp5723 = temp5722 ^ temp5722;
    assign temp5724 = temp5723 ^ temp5723;
    assign temp5725 = temp5724 ^ temp5724;
    assign temp5726 = temp5725 ^ temp5725;
    assign temp5727 = temp5726 ^ temp5726;
    assign temp5728 = temp5727 ^ temp5727;
    assign temp5729 = temp5728 ^ temp5728;
    assign temp5730 = temp5729 ^ temp5729;
    assign temp5731 = temp5730 ^ temp5730;
    assign temp5732 = temp5731 ^ temp5731;
    assign temp5733 = temp5732 ^ temp5732;
    assign temp5734 = temp5733 ^ temp5733;
    assign temp5735 = temp5734 ^ temp5734;
    assign temp5736 = temp5735 ^ temp5735;
    assign temp5737 = temp5736 ^ temp5736;
    assign temp5738 = temp5737 ^ temp5737;
    assign temp5739 = temp5738 ^ temp5738;
    assign temp5740 = temp5739 ^ temp5739;
    assign temp5741 = temp5740 ^ temp5740;
    assign temp5742 = temp5741 ^ temp5741;
    assign temp5743 = temp5742 ^ temp5742;
    assign temp5744 = temp5743 ^ temp5743;
    assign temp5745 = temp5744 ^ temp5744;
    assign temp5746 = temp5745 ^ temp5745;
    assign temp5747 = temp5746 ^ temp5746;
    assign temp5748 = temp5747 ^ temp5747;
    assign temp5749 = temp5748 ^ temp5748;
    assign temp5750 = temp5749 ^ temp5749;
    assign temp5751 = temp5750 ^ temp5750;
    assign temp5752 = temp5751 ^ temp5751;
    assign temp5753 = temp5752 ^ temp5752;
    assign temp5754 = temp5753 ^ temp5753;
    assign temp5755 = temp5754 ^ temp5754;
    assign temp5756 = temp5755 ^ temp5755;
    assign temp5757 = temp5756 ^ temp5756;
    assign temp5758 = temp5757 ^ temp5757;
    assign temp5759 = temp5758 ^ temp5758;
    assign temp5760 = temp5759 ^ temp5759;
    assign temp5761 = temp5760 ^ temp5760;
    assign temp5762 = temp5761 ^ temp5761;
    assign temp5763 = temp5762 ^ temp5762;
    assign temp5764 = temp5763 ^ temp5763;
    assign temp5765 = temp5764 ^ temp5764;
    assign temp5766 = temp5765 ^ temp5765;
    assign temp5767 = temp5766 ^ temp5766;
    assign temp5768 = temp5767 ^ temp5767;
    assign temp5769 = temp5768 ^ temp5768;
    assign temp5770 = temp5769 ^ temp5769;
    assign temp5771 = temp5770 ^ temp5770;
    assign temp5772 = temp5771 ^ temp5771;
    assign temp5773 = temp5772 ^ temp5772;
    assign temp5774 = temp5773 ^ temp5773;
    assign temp5775 = temp5774 ^ temp5774;
    assign temp5776 = temp5775 ^ temp5775;
    assign temp5777 = temp5776 ^ temp5776;
    assign temp5778 = temp5777 ^ temp5777;
    assign temp5779 = temp5778 ^ temp5778;
    assign temp5780 = temp5779 ^ temp5779;
    assign temp5781 = temp5780 ^ temp5780;
    assign temp5782 = temp5781 ^ temp5781;
    assign temp5783 = temp5782 ^ temp5782;
    assign temp5784 = temp5783 ^ temp5783;
    assign temp5785 = temp5784 ^ temp5784;
    assign temp5786 = temp5785 ^ temp5785;
    assign temp5787 = temp5786 ^ temp5786;
    assign temp5788 = temp5787 ^ temp5787;
    assign temp5789 = temp5788 ^ temp5788;
    assign temp5790 = temp5789 ^ temp5789;
    assign temp5791 = temp5790 ^ temp5790;
    assign temp5792 = temp5791 ^ temp5791;
    assign temp5793 = temp5792 ^ temp5792;
    assign temp5794 = temp5793 ^ temp5793;
    assign temp5795 = temp5794 ^ temp5794;
    assign temp5796 = temp5795 ^ temp5795;
    assign temp5797 = temp5796 ^ temp5796;
    assign temp5798 = temp5797 ^ temp5797;
    assign temp5799 = temp5798 ^ temp5798;
    assign temp5800 = temp5799 ^ temp5799;
    assign temp5801 = temp5800 ^ temp5800;
    assign temp5802 = temp5801 ^ temp5801;
    assign temp5803 = temp5802 ^ temp5802;
    assign temp5804 = temp5803 ^ temp5803;
    assign temp5805 = temp5804 ^ temp5804;
    assign temp5806 = temp5805 ^ temp5805;
    assign temp5807 = temp5806 ^ temp5806;
    assign temp5808 = temp5807 ^ temp5807;
    assign temp5809 = temp5808 ^ temp5808;
    assign temp5810 = temp5809 ^ temp5809;
    assign temp5811 = temp5810 ^ temp5810;
    assign temp5812 = temp5811 ^ temp5811;
    assign temp5813 = temp5812 ^ temp5812;
    assign temp5814 = temp5813 ^ temp5813;
    assign temp5815 = temp5814 ^ temp5814;
    assign temp5816 = temp5815 ^ temp5815;
    assign temp5817 = temp5816 ^ temp5816;
    assign temp5818 = temp5817 ^ temp5817;
    assign temp5819 = temp5818 ^ temp5818;
    assign temp5820 = temp5819 ^ temp5819;
    assign temp5821 = temp5820 ^ temp5820;
    assign temp5822 = temp5821 ^ temp5821;
    assign temp5823 = temp5822 ^ temp5822;
    assign temp5824 = temp5823 ^ temp5823;
    assign temp5825 = temp5824 ^ temp5824;
    assign temp5826 = temp5825 ^ temp5825;
    assign temp5827 = temp5826 ^ temp5826;
    assign temp5828 = temp5827 ^ temp5827;
    assign temp5829 = temp5828 ^ temp5828;
    assign temp5830 = temp5829 ^ temp5829;
    assign temp5831 = temp5830 ^ temp5830;
    assign temp5832 = temp5831 ^ temp5831;
    assign temp5833 = temp5832 ^ temp5832;
    assign temp5834 = temp5833 ^ temp5833;
    assign temp5835 = temp5834 ^ temp5834;
    assign temp5836 = temp5835 ^ temp5835;
    assign temp5837 = temp5836 ^ temp5836;
    assign temp5838 = temp5837 ^ temp5837;
    assign temp5839 = temp5838 ^ temp5838;
    assign temp5840 = temp5839 ^ temp5839;
    assign temp5841 = temp5840 ^ temp5840;
    assign temp5842 = temp5841 ^ temp5841;
    assign temp5843 = temp5842 ^ temp5842;
    assign temp5844 = temp5843 ^ temp5843;
    assign temp5845 = temp5844 ^ temp5844;
    assign temp5846 = temp5845 ^ temp5845;
    assign temp5847 = temp5846 ^ temp5846;
    assign temp5848 = temp5847 ^ temp5847;
    assign temp5849 = temp5848 ^ temp5848;
    assign temp5850 = temp5849 ^ temp5849;
    assign temp5851 = temp5850 ^ temp5850;
    assign temp5852 = temp5851 ^ temp5851;
    assign temp5853 = temp5852 ^ temp5852;
    assign temp5854 = temp5853 ^ temp5853;
    assign temp5855 = temp5854 ^ temp5854;
    assign temp5856 = temp5855 ^ temp5855;
    assign temp5857 = temp5856 ^ temp5856;
    assign temp5858 = temp5857 ^ temp5857;
    assign temp5859 = temp5858 ^ temp5858;
    assign temp5860 = temp5859 ^ temp5859;
    assign temp5861 = temp5860 ^ temp5860;
    assign temp5862 = temp5861 ^ temp5861;
    assign temp5863 = temp5862 ^ temp5862;
    assign temp5864 = temp5863 ^ temp5863;
    assign temp5865 = temp5864 ^ temp5864;
    assign temp5866 = temp5865 ^ temp5865;
    assign temp5867 = temp5866 ^ temp5866;
    assign temp5868 = temp5867 ^ temp5867;
    assign temp5869 = temp5868 ^ temp5868;
    assign temp5870 = temp5869 ^ temp5869;
    assign temp5871 = temp5870 ^ temp5870;
    assign temp5872 = temp5871 ^ temp5871;
    assign temp5873 = temp5872 ^ temp5872;
    assign temp5874 = temp5873 ^ temp5873;
    assign temp5875 = temp5874 ^ temp5874;
    assign temp5876 = temp5875 ^ temp5875;
    assign temp5877 = temp5876 ^ temp5876;
    assign temp5878 = temp5877 ^ temp5877;
    assign temp5879 = temp5878 ^ temp5878;
    assign temp5880 = temp5879 ^ temp5879;
    assign temp5881 = temp5880 ^ temp5880;
    assign temp5882 = temp5881 ^ temp5881;
    assign temp5883 = temp5882 ^ temp5882;
    assign temp5884 = temp5883 ^ temp5883;
    assign temp5885 = temp5884 ^ temp5884;
    assign temp5886 = temp5885 ^ temp5885;
    assign temp5887 = temp5886 ^ temp5886;
    assign temp5888 = temp5887 ^ temp5887;
    assign temp5889 = temp5888 ^ temp5888;
    assign temp5890 = temp5889 ^ temp5889;
    assign temp5891 = temp5890 ^ temp5890;
    assign temp5892 = temp5891 ^ temp5891;
    assign temp5893 = temp5892 ^ temp5892;
    assign temp5894 = temp5893 ^ temp5893;
    assign temp5895 = temp5894 ^ temp5894;
    assign temp5896 = temp5895 ^ temp5895;
    assign temp5897 = temp5896 ^ temp5896;
    assign temp5898 = temp5897 ^ temp5897;
    assign temp5899 = temp5898 ^ temp5898;
    assign temp5900 = temp5899 ^ temp5899;
    assign temp5901 = temp5900 ^ temp5900;
    assign temp5902 = temp5901 ^ temp5901;
    assign temp5903 = temp5902 ^ temp5902;
    assign temp5904 = temp5903 ^ temp5903;
    assign temp5905 = temp5904 ^ temp5904;
    assign temp5906 = temp5905 ^ temp5905;
    assign temp5907 = temp5906 ^ temp5906;
    assign temp5908 = temp5907 ^ temp5907;
    assign temp5909 = temp5908 ^ temp5908;
    assign temp5910 = temp5909 ^ temp5909;
    assign temp5911 = temp5910 ^ temp5910;
    assign temp5912 = temp5911 ^ temp5911;
    assign temp5913 = temp5912 ^ temp5912;
    assign temp5914 = temp5913 ^ temp5913;
    assign temp5915 = temp5914 ^ temp5914;
    assign temp5916 = temp5915 ^ temp5915;
    assign temp5917 = temp5916 ^ temp5916;
    assign temp5918 = temp5917 ^ temp5917;
    assign temp5919 = temp5918 ^ temp5918;
    assign temp5920 = temp5919 ^ temp5919;
    assign temp5921 = temp5920 ^ temp5920;
    assign temp5922 = temp5921 ^ temp5921;
    assign temp5923 = temp5922 ^ temp5922;
    assign temp5924 = temp5923 ^ temp5923;
    assign temp5925 = temp5924 ^ temp5924;
    assign temp5926 = temp5925 ^ temp5925;
    assign temp5927 = temp5926 ^ temp5926;
    assign temp5928 = temp5927 ^ temp5927;
    assign temp5929 = temp5928 ^ temp5928;
    assign temp5930 = temp5929 ^ temp5929;
    assign temp5931 = temp5930 ^ temp5930;
    assign temp5932 = temp5931 ^ temp5931;
    assign temp5933 = temp5932 ^ temp5932;
    assign temp5934 = temp5933 ^ temp5933;
    assign temp5935 = temp5934 ^ temp5934;
    assign temp5936 = temp5935 ^ temp5935;
    assign temp5937 = temp5936 ^ temp5936;
    assign temp5938 = temp5937 ^ temp5937;
    assign temp5939 = temp5938 ^ temp5938;
    assign temp5940 = temp5939 ^ temp5939;
    assign temp5941 = temp5940 ^ temp5940;
    assign temp5942 = temp5941 ^ temp5941;
    assign temp5943 = temp5942 ^ temp5942;
    assign temp5944 = temp5943 ^ temp5943;
    assign temp5945 = temp5944 ^ temp5944;
    assign temp5946 = temp5945 ^ temp5945;
    assign temp5947 = temp5946 ^ temp5946;
    assign temp5948 = temp5947 ^ temp5947;
    assign temp5949 = temp5948 ^ temp5948;
    assign temp5950 = temp5949 ^ temp5949;
    assign temp5951 = temp5950 ^ temp5950;
    assign temp5952 = temp5951 ^ temp5951;
    assign temp5953 = temp5952 ^ temp5952;
    assign temp5954 = temp5953 ^ temp5953;
    assign temp5955 = temp5954 ^ temp5954;
    assign temp5956 = temp5955 ^ temp5955;
    assign temp5957 = temp5956 ^ temp5956;
    assign temp5958 = temp5957 ^ temp5957;
    assign temp5959 = temp5958 ^ temp5958;
    assign temp5960 = temp5959 ^ temp5959;
    assign temp5961 = temp5960 ^ temp5960;
    assign temp5962 = temp5961 ^ temp5961;
    assign temp5963 = temp5962 ^ temp5962;
    assign temp5964 = temp5963 ^ temp5963;
    assign temp5965 = temp5964 ^ temp5964;
    assign temp5966 = temp5965 ^ temp5965;
    assign temp5967 = temp5966 ^ temp5966;
    assign temp5968 = temp5967 ^ temp5967;
    assign temp5969 = temp5968 ^ temp5968;
    assign temp5970 = temp5969 ^ temp5969;
    assign temp5971 = temp5970 ^ temp5970;
    assign temp5972 = temp5971 ^ temp5971;
    assign temp5973 = temp5972 ^ temp5972;
    assign temp5974 = temp5973 ^ temp5973;
    assign temp5975 = temp5974 ^ temp5974;
    assign temp5976 = temp5975 ^ temp5975;
    assign temp5977 = temp5976 ^ temp5976;
    assign temp5978 = temp5977 ^ temp5977;
    assign temp5979 = temp5978 ^ temp5978;
    assign temp5980 = temp5979 ^ temp5979;
    assign temp5981 = temp5980 ^ temp5980;
    assign temp5982 = temp5981 ^ temp5981;
    assign temp5983 = temp5982 ^ temp5982;
    assign temp5984 = temp5983 ^ temp5983;
    assign temp5985 = temp5984 ^ temp5984;
    assign temp5986 = temp5985 ^ temp5985;
    assign temp5987 = temp5986 ^ temp5986;
    assign temp5988 = temp5987 ^ temp5987;
    assign temp5989 = temp5988 ^ temp5988;
    assign temp5990 = temp5989 ^ temp5989;
    assign temp5991 = temp5990 ^ temp5990;
    assign temp5992 = temp5991 ^ temp5991;
    assign temp5993 = temp5992 ^ temp5992;
    assign temp5994 = temp5993 ^ temp5993;
    assign temp5995 = temp5994 ^ temp5994;
    assign temp5996 = temp5995 ^ temp5995;
    assign temp5997 = temp5996 ^ temp5996;
    assign temp5998 = temp5997 ^ temp5997;
    assign temp5999 = temp5998 ^ temp5998;
    assign temp6000 = temp5999 ^ temp5999;
    assign temp6001 = temp6000 ^ temp6000;
    assign temp6002 = temp6001 ^ temp6001;
    assign temp6003 = temp6002 ^ temp6002;
    assign temp6004 = temp6003 ^ temp6003;
    assign temp6005 = temp6004 ^ temp6004;
    assign temp6006 = temp6005 ^ temp6005;
    assign temp6007 = temp6006 ^ temp6006;
    assign temp6008 = temp6007 ^ temp6007;
    assign temp6009 = temp6008 ^ temp6008;
    assign temp6010 = temp6009 ^ temp6009;
    assign temp6011 = temp6010 ^ temp6010;
    assign temp6012 = temp6011 ^ temp6011;
    assign temp6013 = temp6012 ^ temp6012;
    assign temp6014 = temp6013 ^ temp6013;
    assign temp6015 = temp6014 ^ temp6014;
    assign temp6016 = temp6015 ^ temp6015;
    assign temp6017 = temp6016 ^ temp6016;
    assign temp6018 = temp6017 ^ temp6017;
    assign temp6019 = temp6018 ^ temp6018;
    assign temp6020 = temp6019 ^ temp6019;
    assign temp6021 = temp6020 ^ temp6020;
    assign temp6022 = temp6021 ^ temp6021;
    assign temp6023 = temp6022 ^ temp6022;
    assign temp6024 = temp6023 ^ temp6023;
    assign temp6025 = temp6024 ^ temp6024;
    assign temp6026 = temp6025 ^ temp6025;
    assign temp6027 = temp6026 ^ temp6026;
    assign temp6028 = temp6027 ^ temp6027;
    assign temp6029 = temp6028 ^ temp6028;
    assign temp6030 = temp6029 ^ temp6029;
    assign temp6031 = temp6030 ^ temp6030;
    assign temp6032 = temp6031 ^ temp6031;
    assign temp6033 = temp6032 ^ temp6032;
    assign temp6034 = temp6033 ^ temp6033;
    assign temp6035 = temp6034 ^ temp6034;
    assign temp6036 = temp6035 ^ temp6035;
    assign temp6037 = temp6036 ^ temp6036;
    assign temp6038 = temp6037 ^ temp6037;
    assign temp6039 = temp6038 ^ temp6038;
    assign temp6040 = temp6039 ^ temp6039;
    assign temp6041 = temp6040 ^ temp6040;
    assign temp6042 = temp6041 ^ temp6041;
    assign temp6043 = temp6042 ^ temp6042;
    assign temp6044 = temp6043 ^ temp6043;
    assign temp6045 = temp6044 ^ temp6044;
    assign temp6046 = temp6045 ^ temp6045;
    assign temp6047 = temp6046 ^ temp6046;
    assign temp6048 = temp6047 ^ temp6047;
    assign temp6049 = temp6048 ^ temp6048;
    assign temp6050 = temp6049 ^ temp6049;
    assign temp6051 = temp6050 ^ temp6050;
    assign temp6052 = temp6051 ^ temp6051;
    assign temp6053 = temp6052 ^ temp6052;
    assign temp6054 = temp6053 ^ temp6053;
    assign temp6055 = temp6054 ^ temp6054;
    assign temp6056 = temp6055 ^ temp6055;
    assign temp6057 = temp6056 ^ temp6056;
    assign temp6058 = temp6057 ^ temp6057;
    assign temp6059 = temp6058 ^ temp6058;
    assign temp6060 = temp6059 ^ temp6059;
    assign temp6061 = temp6060 ^ temp6060;
    assign temp6062 = temp6061 ^ temp6061;
    assign temp6063 = temp6062 ^ temp6062;
    assign temp6064 = temp6063 ^ temp6063;
    assign temp6065 = temp6064 ^ temp6064;
    assign temp6066 = temp6065 ^ temp6065;
    assign temp6067 = temp6066 ^ temp6066;
    assign temp6068 = temp6067 ^ temp6067;
    assign temp6069 = temp6068 ^ temp6068;
    assign temp6070 = temp6069 ^ temp6069;
    assign temp6071 = temp6070 ^ temp6070;
    assign temp6072 = temp6071 ^ temp6071;
    assign temp6073 = temp6072 ^ temp6072;
    assign temp6074 = temp6073 ^ temp6073;
    assign temp6075 = temp6074 ^ temp6074;
    assign temp6076 = temp6075 ^ temp6075;
    assign temp6077 = temp6076 ^ temp6076;
    assign temp6078 = temp6077 ^ temp6077;
    assign temp6079 = temp6078 ^ temp6078;
    assign temp6080 = temp6079 ^ temp6079;
    assign temp6081 = temp6080 ^ temp6080;
    assign temp6082 = temp6081 ^ temp6081;
    assign temp6083 = temp6082 ^ temp6082;
    assign temp6084 = temp6083 ^ temp6083;
    assign temp6085 = temp6084 ^ temp6084;
    assign temp6086 = temp6085 ^ temp6085;
    assign temp6087 = temp6086 ^ temp6086;
    assign temp6088 = temp6087 ^ temp6087;
    assign temp6089 = temp6088 ^ temp6088;
    assign temp6090 = temp6089 ^ temp6089;
    assign temp6091 = temp6090 ^ temp6090;
    assign temp6092 = temp6091 ^ temp6091;
    assign temp6093 = temp6092 ^ temp6092;
    assign temp6094 = temp6093 ^ temp6093;
    assign temp6095 = temp6094 ^ temp6094;
    assign temp6096 = temp6095 ^ temp6095;
    assign temp6097 = temp6096 ^ temp6096;
    assign temp6098 = temp6097 ^ temp6097;
    assign temp6099 = temp6098 ^ temp6098;
    assign temp6100 = temp6099 ^ temp6099;
    assign temp6101 = temp6100 ^ temp6100;
    assign temp6102 = temp6101 ^ temp6101;
    assign temp6103 = temp6102 ^ temp6102;
    assign temp6104 = temp6103 ^ temp6103;
    assign temp6105 = temp6104 ^ temp6104;
    assign temp6106 = temp6105 ^ temp6105;
    assign temp6107 = temp6106 ^ temp6106;
    assign temp6108 = temp6107 ^ temp6107;
    assign temp6109 = temp6108 ^ temp6108;
    assign temp6110 = temp6109 ^ temp6109;
    assign temp6111 = temp6110 ^ temp6110;
    assign temp6112 = temp6111 ^ temp6111;
    assign temp6113 = temp6112 ^ temp6112;
    assign temp6114 = temp6113 ^ temp6113;
    assign temp6115 = temp6114 ^ temp6114;
    assign temp6116 = temp6115 ^ temp6115;
    assign temp6117 = temp6116 ^ temp6116;
    assign temp6118 = temp6117 ^ temp6117;
    assign temp6119 = temp6118 ^ temp6118;
    assign temp6120 = temp6119 ^ temp6119;
    assign temp6121 = temp6120 ^ temp6120;
    assign temp6122 = temp6121 ^ temp6121;
    assign temp6123 = temp6122 ^ temp6122;
    assign temp6124 = temp6123 ^ temp6123;
    assign temp6125 = temp6124 ^ temp6124;
    assign temp6126 = temp6125 ^ temp6125;
    assign temp6127 = temp6126 ^ temp6126;
    assign temp6128 = temp6127 ^ temp6127;
    assign temp6129 = temp6128 ^ temp6128;
    assign temp6130 = temp6129 ^ temp6129;
    assign temp6131 = temp6130 ^ temp6130;
    assign temp6132 = temp6131 ^ temp6131;
    assign temp6133 = temp6132 ^ temp6132;
    assign temp6134 = temp6133 ^ temp6133;
    assign temp6135 = temp6134 ^ temp6134;
    assign temp6136 = temp6135 ^ temp6135;
    assign temp6137 = temp6136 ^ temp6136;
    assign temp6138 = temp6137 ^ temp6137;
    assign temp6139 = temp6138 ^ temp6138;
    assign temp6140 = temp6139 ^ temp6139;
    assign temp6141 = temp6140 ^ temp6140;
    assign temp6142 = temp6141 ^ temp6141;
    assign temp6143 = temp6142 ^ temp6142;
    assign temp6144 = temp6143 ^ temp6143;
    assign temp6145 = temp6144 ^ temp6144;
    assign temp6146 = temp6145 ^ temp6145;
    assign temp6147 = temp6146 ^ temp6146;
    assign temp6148 = temp6147 ^ temp6147;
    assign temp6149 = temp6148 ^ temp6148;
    assign temp6150 = temp6149 ^ temp6149;
    assign temp6151 = temp6150 ^ temp6150;
    assign temp6152 = temp6151 ^ temp6151;
    assign temp6153 = temp6152 ^ temp6152;
    assign temp6154 = temp6153 ^ temp6153;
    assign temp6155 = temp6154 ^ temp6154;
    assign temp6156 = temp6155 ^ temp6155;
    assign temp6157 = temp6156 ^ temp6156;
    assign temp6158 = temp6157 ^ temp6157;
    assign temp6159 = temp6158 ^ temp6158;
    assign temp6160 = temp6159 ^ temp6159;
    assign temp6161 = temp6160 ^ temp6160;
    assign temp6162 = temp6161 ^ temp6161;
    assign temp6163 = temp6162 ^ temp6162;
    assign temp6164 = temp6163 ^ temp6163;
    assign temp6165 = temp6164 ^ temp6164;
    assign temp6166 = temp6165 ^ temp6165;
    assign temp6167 = temp6166 ^ temp6166;
    assign temp6168 = temp6167 ^ temp6167;
    assign temp6169 = temp6168 ^ temp6168;
    assign temp6170 = temp6169 ^ temp6169;
    assign temp6171 = temp6170 ^ temp6170;
    assign temp6172 = temp6171 ^ temp6171;
    assign temp6173 = temp6172 ^ temp6172;
    assign temp6174 = temp6173 ^ temp6173;
    assign temp6175 = temp6174 ^ temp6174;
    assign temp6176 = temp6175 ^ temp6175;
    assign temp6177 = temp6176 ^ temp6176;
    assign temp6178 = temp6177 ^ temp6177;
    assign temp6179 = temp6178 ^ temp6178;
    assign temp6180 = temp6179 ^ temp6179;
    assign temp6181 = temp6180 ^ temp6180;
    assign temp6182 = temp6181 ^ temp6181;
    assign temp6183 = temp6182 ^ temp6182;
    assign temp6184 = temp6183 ^ temp6183;
    assign temp6185 = temp6184 ^ temp6184;
    assign temp6186 = temp6185 ^ temp6185;
    assign temp6187 = temp6186 ^ temp6186;
    assign temp6188 = temp6187 ^ temp6187;
    assign temp6189 = temp6188 ^ temp6188;
    assign temp6190 = temp6189 ^ temp6189;
    assign temp6191 = temp6190 ^ temp6190;
    assign temp6192 = temp6191 ^ temp6191;
    assign temp6193 = temp6192 ^ temp6192;
    assign temp6194 = temp6193 ^ temp6193;
    assign temp6195 = temp6194 ^ temp6194;
    assign temp6196 = temp6195 ^ temp6195;
    assign temp6197 = temp6196 ^ temp6196;
    assign temp6198 = temp6197 ^ temp6197;
    assign temp6199 = temp6198 ^ temp6198;
    assign temp6200 = temp6199 ^ temp6199;
    assign temp6201 = temp6200 ^ temp6200;
    assign temp6202 = temp6201 ^ temp6201;
    assign temp6203 = temp6202 ^ temp6202;
    assign temp6204 = temp6203 ^ temp6203;
    assign temp6205 = temp6204 ^ temp6204;
    assign temp6206 = temp6205 ^ temp6205;
    assign temp6207 = temp6206 ^ temp6206;
    assign temp6208 = temp6207 ^ temp6207;
    assign temp6209 = temp6208 ^ temp6208;
    assign temp6210 = temp6209 ^ temp6209;
    assign temp6211 = temp6210 ^ temp6210;
    assign temp6212 = temp6211 ^ temp6211;
    assign temp6213 = temp6212 ^ temp6212;
    assign temp6214 = temp6213 ^ temp6213;
    assign temp6215 = temp6214 ^ temp6214;
    assign temp6216 = temp6215 ^ temp6215;
    assign temp6217 = temp6216 ^ temp6216;
    assign temp6218 = temp6217 ^ temp6217;
    assign temp6219 = temp6218 ^ temp6218;
    assign temp6220 = temp6219 ^ temp6219;
    assign temp6221 = temp6220 ^ temp6220;
    assign temp6222 = temp6221 ^ temp6221;
    assign temp6223 = temp6222 ^ temp6222;
    assign temp6224 = temp6223 ^ temp6223;
    assign temp6225 = temp6224 ^ temp6224;
    assign temp6226 = temp6225 ^ temp6225;
    assign temp6227 = temp6226 ^ temp6226;
    assign temp6228 = temp6227 ^ temp6227;
    assign temp6229 = temp6228 ^ temp6228;
    assign temp6230 = temp6229 ^ temp6229;
    assign temp6231 = temp6230 ^ temp6230;
    assign temp6232 = temp6231 ^ temp6231;
    assign temp6233 = temp6232 ^ temp6232;
    assign temp6234 = temp6233 ^ temp6233;
    assign temp6235 = temp6234 ^ temp6234;
    assign temp6236 = temp6235 ^ temp6235;
    assign temp6237 = temp6236 ^ temp6236;
    assign temp6238 = temp6237 ^ temp6237;
    assign temp6239 = temp6238 ^ temp6238;
    assign temp6240 = temp6239 ^ temp6239;
    assign temp6241 = temp6240 ^ temp6240;
    assign temp6242 = temp6241 ^ temp6241;
    assign temp6243 = temp6242 ^ temp6242;
    assign temp6244 = temp6243 ^ temp6243;
    assign temp6245 = temp6244 ^ temp6244;
    assign temp6246 = temp6245 ^ temp6245;
    assign temp6247 = temp6246 ^ temp6246;
    assign temp6248 = temp6247 ^ temp6247;
    assign temp6249 = temp6248 ^ temp6248;
    assign temp6250 = temp6249 ^ temp6249;
    assign temp6251 = temp6250 ^ temp6250;
    assign temp6252 = temp6251 ^ temp6251;
    assign temp6253 = temp6252 ^ temp6252;
    assign temp6254 = temp6253 ^ temp6253;
    assign temp6255 = temp6254 ^ temp6254;
    assign temp6256 = temp6255 ^ temp6255;
    assign temp6257 = temp6256 ^ temp6256;
    assign temp6258 = temp6257 ^ temp6257;
    assign temp6259 = temp6258 ^ temp6258;
    assign temp6260 = temp6259 ^ temp6259;
    assign temp6261 = temp6260 ^ temp6260;
    assign temp6262 = temp6261 ^ temp6261;
    assign temp6263 = temp6262 ^ temp6262;
    assign temp6264 = temp6263 ^ temp6263;
    assign temp6265 = temp6264 ^ temp6264;
    assign temp6266 = temp6265 ^ temp6265;
    assign temp6267 = temp6266 ^ temp6266;
    assign temp6268 = temp6267 ^ temp6267;
    assign temp6269 = temp6268 ^ temp6268;
    assign temp6270 = temp6269 ^ temp6269;
    assign temp6271 = temp6270 ^ temp6270;
    assign temp6272 = temp6271 ^ temp6271;
    assign temp6273 = temp6272 ^ temp6272;
    assign temp6274 = temp6273 ^ temp6273;
    assign temp6275 = temp6274 ^ temp6274;
    assign temp6276 = temp6275 ^ temp6275;
    assign temp6277 = temp6276 ^ temp6276;
    assign temp6278 = temp6277 ^ temp6277;
    assign temp6279 = temp6278 ^ temp6278;
    assign temp6280 = temp6279 ^ temp6279;
    assign temp6281 = temp6280 ^ temp6280;
    assign temp6282 = temp6281 ^ temp6281;
    assign temp6283 = temp6282 ^ temp6282;
    assign temp6284 = temp6283 ^ temp6283;
    assign temp6285 = temp6284 ^ temp6284;
    assign temp6286 = temp6285 ^ temp6285;
    assign temp6287 = temp6286 ^ temp6286;
    assign temp6288 = temp6287 ^ temp6287;
    assign temp6289 = temp6288 ^ temp6288;
    assign temp6290 = temp6289 ^ temp6289;
    assign temp6291 = temp6290 ^ temp6290;
    assign temp6292 = temp6291 ^ temp6291;
    assign temp6293 = temp6292 ^ temp6292;
    assign temp6294 = temp6293 ^ temp6293;
    assign temp6295 = temp6294 ^ temp6294;
    assign temp6296 = temp6295 ^ temp6295;
    assign temp6297 = temp6296 ^ temp6296;
    assign temp6298 = temp6297 ^ temp6297;
    assign temp6299 = temp6298 ^ temp6298;
    assign temp6300 = temp6299 ^ temp6299;
    assign temp6301 = temp6300 ^ temp6300;
    assign temp6302 = temp6301 ^ temp6301;
    assign temp6303 = temp6302 ^ temp6302;
    assign temp6304 = temp6303 ^ temp6303;
    assign temp6305 = temp6304 ^ temp6304;
    assign temp6306 = temp6305 ^ temp6305;
    assign temp6307 = temp6306 ^ temp6306;
    assign temp6308 = temp6307 ^ temp6307;
    assign temp6309 = temp6308 ^ temp6308;
    assign temp6310 = temp6309 ^ temp6309;
    assign temp6311 = temp6310 ^ temp6310;
    assign temp6312 = temp6311 ^ temp6311;
    assign temp6313 = temp6312 ^ temp6312;
    assign temp6314 = temp6313 ^ temp6313;
    assign temp6315 = temp6314 ^ temp6314;
    assign temp6316 = temp6315 ^ temp6315;
    assign temp6317 = temp6316 ^ temp6316;
    assign temp6318 = temp6317 ^ temp6317;
    assign temp6319 = temp6318 ^ temp6318;
    assign temp6320 = temp6319 ^ temp6319;
    assign temp6321 = temp6320 ^ temp6320;
    assign temp6322 = temp6321 ^ temp6321;
    assign temp6323 = temp6322 ^ temp6322;
    assign temp6324 = temp6323 ^ temp6323;
    assign temp6325 = temp6324 ^ temp6324;
    assign temp6326 = temp6325 ^ temp6325;
    assign temp6327 = temp6326 ^ temp6326;
    assign temp6328 = temp6327 ^ temp6327;
    assign temp6329 = temp6328 ^ temp6328;
    assign temp6330 = temp6329 ^ temp6329;
    assign temp6331 = temp6330 ^ temp6330;
    assign temp6332 = temp6331 ^ temp6331;
    assign temp6333 = temp6332 ^ temp6332;
    assign temp6334 = temp6333 ^ temp6333;
    assign temp6335 = temp6334 ^ temp6334;
    assign temp6336 = temp6335 ^ temp6335;
    assign temp6337 = temp6336 ^ temp6336;
    assign temp6338 = temp6337 ^ temp6337;
    assign temp6339 = temp6338 ^ temp6338;
    assign temp6340 = temp6339 ^ temp6339;
    assign temp6341 = temp6340 ^ temp6340;
    assign temp6342 = temp6341 ^ temp6341;
    assign temp6343 = temp6342 ^ temp6342;
    assign temp6344 = temp6343 ^ temp6343;
    assign temp6345 = temp6344 ^ temp6344;
    assign temp6346 = temp6345 ^ temp6345;
    assign temp6347 = temp6346 ^ temp6346;
    assign temp6348 = temp6347 ^ temp6347;
    assign temp6349 = temp6348 ^ temp6348;
    assign temp6350 = temp6349 ^ temp6349;
    assign temp6351 = temp6350 ^ temp6350;
    assign temp6352 = temp6351 ^ temp6351;
    assign temp6353 = temp6352 ^ temp6352;
    assign temp6354 = temp6353 ^ temp6353;
    assign temp6355 = temp6354 ^ temp6354;
    assign temp6356 = temp6355 ^ temp6355;
    assign temp6357 = temp6356 ^ temp6356;
    assign temp6358 = temp6357 ^ temp6357;
    assign temp6359 = temp6358 ^ temp6358;
    assign temp6360 = temp6359 ^ temp6359;
    assign temp6361 = temp6360 ^ temp6360;
    assign temp6362 = temp6361 ^ temp6361;
    assign temp6363 = temp6362 ^ temp6362;
    assign temp6364 = temp6363 ^ temp6363;
    assign temp6365 = temp6364 ^ temp6364;
    assign temp6366 = temp6365 ^ temp6365;
    assign temp6367 = temp6366 ^ temp6366;
    assign temp6368 = temp6367 ^ temp6367;
    assign temp6369 = temp6368 ^ temp6368;
    assign temp6370 = temp6369 ^ temp6369;
    assign temp6371 = temp6370 ^ temp6370;
    assign temp6372 = temp6371 ^ temp6371;
    assign temp6373 = temp6372 ^ temp6372;
    assign temp6374 = temp6373 ^ temp6373;
    assign temp6375 = temp6374 ^ temp6374;
    assign temp6376 = temp6375 ^ temp6375;
    assign temp6377 = temp6376 ^ temp6376;
    assign temp6378 = temp6377 ^ temp6377;
    assign temp6379 = temp6378 ^ temp6378;
    assign temp6380 = temp6379 ^ temp6379;
    assign temp6381 = temp6380 ^ temp6380;
    assign temp6382 = temp6381 ^ temp6381;
    assign temp6383 = temp6382 ^ temp6382;
    assign temp6384 = temp6383 ^ temp6383;
    assign temp6385 = temp6384 ^ temp6384;
    assign temp6386 = temp6385 ^ temp6385;
    assign temp6387 = temp6386 ^ temp6386;
    assign temp6388 = temp6387 ^ temp6387;
    assign temp6389 = temp6388 ^ temp6388;
    assign temp6390 = temp6389 ^ temp6389;
    assign temp6391 = temp6390 ^ temp6390;
    assign temp6392 = temp6391 ^ temp6391;
    assign temp6393 = temp6392 ^ temp6392;
    assign temp6394 = temp6393 ^ temp6393;
    assign temp6395 = temp6394 ^ temp6394;
    assign temp6396 = temp6395 ^ temp6395;
    assign temp6397 = temp6396 ^ temp6396;
    assign temp6398 = temp6397 ^ temp6397;
    assign temp6399 = temp6398 ^ temp6398;
    assign temp6400 = temp6399 ^ temp6399;
    assign temp6401 = temp6400 ^ temp6400;
    assign temp6402 = temp6401 ^ temp6401;
    assign temp6403 = temp6402 ^ temp6402;
    assign temp6404 = temp6403 ^ temp6403;
    assign temp6405 = temp6404 ^ temp6404;
    assign temp6406 = temp6405 ^ temp6405;
    assign temp6407 = temp6406 ^ temp6406;
    assign temp6408 = temp6407 ^ temp6407;
    assign temp6409 = temp6408 ^ temp6408;
    assign temp6410 = temp6409 ^ temp6409;
    assign temp6411 = temp6410 ^ temp6410;
    assign temp6412 = temp6411 ^ temp6411;
    assign temp6413 = temp6412 ^ temp6412;
    assign temp6414 = temp6413 ^ temp6413;
    assign temp6415 = temp6414 ^ temp6414;
    assign temp6416 = temp6415 ^ temp6415;
    assign temp6417 = temp6416 ^ temp6416;
    assign temp6418 = temp6417 ^ temp6417;
    assign temp6419 = temp6418 ^ temp6418;
    assign temp6420 = temp6419 ^ temp6419;
    assign temp6421 = temp6420 ^ temp6420;
    assign temp6422 = temp6421 ^ temp6421;
    assign temp6423 = temp6422 ^ temp6422;
    assign temp6424 = temp6423 ^ temp6423;
    assign temp6425 = temp6424 ^ temp6424;
    assign temp6426 = temp6425 ^ temp6425;
    assign temp6427 = temp6426 ^ temp6426;
    assign temp6428 = temp6427 ^ temp6427;
    assign temp6429 = temp6428 ^ temp6428;
    assign temp6430 = temp6429 ^ temp6429;
    assign temp6431 = temp6430 ^ temp6430;
    assign temp6432 = temp6431 ^ temp6431;
    assign temp6433 = temp6432 ^ temp6432;
    assign temp6434 = temp6433 ^ temp6433;
    assign temp6435 = temp6434 ^ temp6434;
    assign temp6436 = temp6435 ^ temp6435;
    assign temp6437 = temp6436 ^ temp6436;
    assign temp6438 = temp6437 ^ temp6437;
    assign temp6439 = temp6438 ^ temp6438;
    assign temp6440 = temp6439 ^ temp6439;
    assign temp6441 = temp6440 ^ temp6440;
    assign temp6442 = temp6441 ^ temp6441;
    assign temp6443 = temp6442 ^ temp6442;
    assign temp6444 = temp6443 ^ temp6443;
    assign temp6445 = temp6444 ^ temp6444;
    assign temp6446 = temp6445 ^ temp6445;
    assign temp6447 = temp6446 ^ temp6446;
    assign temp6448 = temp6447 ^ temp6447;
    assign temp6449 = temp6448 ^ temp6448;
    assign temp6450 = temp6449 ^ temp6449;
    assign temp6451 = temp6450 ^ temp6450;
    assign temp6452 = temp6451 ^ temp6451;
    assign temp6453 = temp6452 ^ temp6452;
    assign temp6454 = temp6453 ^ temp6453;
    assign temp6455 = temp6454 ^ temp6454;
    assign temp6456 = temp6455 ^ temp6455;
    assign temp6457 = temp6456 ^ temp6456;
    assign temp6458 = temp6457 ^ temp6457;
    assign temp6459 = temp6458 ^ temp6458;
    assign temp6460 = temp6459 ^ temp6459;
    assign temp6461 = temp6460 ^ temp6460;
    assign temp6462 = temp6461 ^ temp6461;
    assign temp6463 = temp6462 ^ temp6462;
    assign temp6464 = temp6463 ^ temp6463;
    assign temp6465 = temp6464 ^ temp6464;
    assign temp6466 = temp6465 ^ temp6465;
    assign temp6467 = temp6466 ^ temp6466;
    assign temp6468 = temp6467 ^ temp6467;
    assign temp6469 = temp6468 ^ temp6468;
    assign temp6470 = temp6469 ^ temp6469;
    assign temp6471 = temp6470 ^ temp6470;
    assign temp6472 = temp6471 ^ temp6471;
    assign temp6473 = temp6472 ^ temp6472;
    assign temp6474 = temp6473 ^ temp6473;
    assign temp6475 = temp6474 ^ temp6474;
    assign temp6476 = temp6475 ^ temp6475;
    assign temp6477 = temp6476 ^ temp6476;
    assign temp6478 = temp6477 ^ temp6477;
    assign temp6479 = temp6478 ^ temp6478;
    assign temp6480 = temp6479 ^ temp6479;
    assign temp6481 = temp6480 ^ temp6480;
    assign temp6482 = temp6481 ^ temp6481;
    assign temp6483 = temp6482 ^ temp6482;
    assign temp6484 = temp6483 ^ temp6483;
    assign temp6485 = temp6484 ^ temp6484;
    assign temp6486 = temp6485 ^ temp6485;
    assign temp6487 = temp6486 ^ temp6486;
    assign temp6488 = temp6487 ^ temp6487;
    assign temp6489 = temp6488 ^ temp6488;
    assign temp6490 = temp6489 ^ temp6489;
    assign temp6491 = temp6490 ^ temp6490;
    assign temp6492 = temp6491 ^ temp6491;
    assign temp6493 = temp6492 ^ temp6492;
    assign temp6494 = temp6493 ^ temp6493;
    assign temp6495 = temp6494 ^ temp6494;
    assign temp6496 = temp6495 ^ temp6495;
    assign temp6497 = temp6496 ^ temp6496;
    assign temp6498 = temp6497 ^ temp6497;
    assign temp6499 = temp6498 ^ temp6498;
    assign temp6500 = temp6499 ^ temp6499;
    assign temp6501 = temp6500 ^ temp6500;
    assign temp6502 = temp6501 ^ temp6501;
    assign temp6503 = temp6502 ^ temp6502;
    assign temp6504 = temp6503 ^ temp6503;
    assign temp6505 = temp6504 ^ temp6504;
    assign temp6506 = temp6505 ^ temp6505;
    assign temp6507 = temp6506 ^ temp6506;
    assign temp6508 = temp6507 ^ temp6507;
    assign temp6509 = temp6508 ^ temp6508;
    assign temp6510 = temp6509 ^ temp6509;
    assign temp6511 = temp6510 ^ temp6510;
    assign temp6512 = temp6511 ^ temp6511;
    assign temp6513 = temp6512 ^ temp6512;
    assign temp6514 = temp6513 ^ temp6513;
    assign temp6515 = temp6514 ^ temp6514;
    assign temp6516 = temp6515 ^ temp6515;
    assign temp6517 = temp6516 ^ temp6516;
    assign temp6518 = temp6517 ^ temp6517;
    assign temp6519 = temp6518 ^ temp6518;
    assign temp6520 = temp6519 ^ temp6519;
    assign temp6521 = temp6520 ^ temp6520;
    assign temp6522 = temp6521 ^ temp6521;
    assign temp6523 = temp6522 ^ temp6522;
    assign temp6524 = temp6523 ^ temp6523;
    assign temp6525 = temp6524 ^ temp6524;
    assign temp6526 = temp6525 ^ temp6525;
    assign temp6527 = temp6526 ^ temp6526;
    assign temp6528 = temp6527 ^ temp6527;
    assign temp6529 = temp6528 ^ temp6528;
    assign temp6530 = temp6529 ^ temp6529;
    assign temp6531 = temp6530 ^ temp6530;
    assign temp6532 = temp6531 ^ temp6531;
    assign temp6533 = temp6532 ^ temp6532;
    assign temp6534 = temp6533 ^ temp6533;
    assign temp6535 = temp6534 ^ temp6534;
    assign temp6536 = temp6535 ^ temp6535;
    assign temp6537 = temp6536 ^ temp6536;
    assign temp6538 = temp6537 ^ temp6537;
    assign temp6539 = temp6538 ^ temp6538;
    assign temp6540 = temp6539 ^ temp6539;
    assign temp6541 = temp6540 ^ temp6540;
    assign temp6542 = temp6541 ^ temp6541;
    assign temp6543 = temp6542 ^ temp6542;
    assign temp6544 = temp6543 ^ temp6543;
    assign temp6545 = temp6544 ^ temp6544;
    assign temp6546 = temp6545 ^ temp6545;
    assign temp6547 = temp6546 ^ temp6546;
    assign temp6548 = temp6547 ^ temp6547;
    assign temp6549 = temp6548 ^ temp6548;
    assign temp6550 = temp6549 ^ temp6549;
    assign temp6551 = temp6550 ^ temp6550;
    assign temp6552 = temp6551 ^ temp6551;
    assign temp6553 = temp6552 ^ temp6552;
    assign temp6554 = temp6553 ^ temp6553;
    assign temp6555 = temp6554 ^ temp6554;
    assign temp6556 = temp6555 ^ temp6555;
    assign temp6557 = temp6556 ^ temp6556;
    assign temp6558 = temp6557 ^ temp6557;
    assign temp6559 = temp6558 ^ temp6558;
    assign temp6560 = temp6559 ^ temp6559;
    assign temp6561 = temp6560 ^ temp6560;
    assign temp6562 = temp6561 ^ temp6561;
    assign temp6563 = temp6562 ^ temp6562;
    assign temp6564 = temp6563 ^ temp6563;
    assign temp6565 = temp6564 ^ temp6564;
    assign temp6566 = temp6565 ^ temp6565;
    assign temp6567 = temp6566 ^ temp6566;
    assign temp6568 = temp6567 ^ temp6567;
    assign temp6569 = temp6568 ^ temp6568;
    assign temp6570 = temp6569 ^ temp6569;
    assign temp6571 = temp6570 ^ temp6570;
    assign temp6572 = temp6571 ^ temp6571;
    assign temp6573 = temp6572 ^ temp6572;
    assign temp6574 = temp6573 ^ temp6573;
    assign temp6575 = temp6574 ^ temp6574;
    assign temp6576 = temp6575 ^ temp6575;
    assign temp6577 = temp6576 ^ temp6576;
    assign temp6578 = temp6577 ^ temp6577;
    assign temp6579 = temp6578 ^ temp6578;
    assign temp6580 = temp6579 ^ temp6579;
    assign temp6581 = temp6580 ^ temp6580;
    assign temp6582 = temp6581 ^ temp6581;
    assign temp6583 = temp6582 ^ temp6582;
    assign temp6584 = temp6583 ^ temp6583;
    assign temp6585 = temp6584 ^ temp6584;
    assign temp6586 = temp6585 ^ temp6585;
    assign temp6587 = temp6586 ^ temp6586;
    assign temp6588 = temp6587 ^ temp6587;
    assign temp6589 = temp6588 ^ temp6588;
    assign temp6590 = temp6589 ^ temp6589;
    assign temp6591 = temp6590 ^ temp6590;
    assign temp6592 = temp6591 ^ temp6591;
    assign temp6593 = temp6592 ^ temp6592;
    assign temp6594 = temp6593 ^ temp6593;
    assign temp6595 = temp6594 ^ temp6594;
    assign temp6596 = temp6595 ^ temp6595;
    assign temp6597 = temp6596 ^ temp6596;
    assign temp6598 = temp6597 ^ temp6597;
    assign temp6599 = temp6598 ^ temp6598;
    assign temp6600 = temp6599 ^ temp6599;
    assign temp6601 = temp6600 ^ temp6600;
    assign temp6602 = temp6601 ^ temp6601;
    assign temp6603 = temp6602 ^ temp6602;
    assign temp6604 = temp6603 ^ temp6603;
    assign temp6605 = temp6604 ^ temp6604;
    assign temp6606 = temp6605 ^ temp6605;
    assign temp6607 = temp6606 ^ temp6606;
    assign temp6608 = temp6607 ^ temp6607;
    assign temp6609 = temp6608 ^ temp6608;
    assign temp6610 = temp6609 ^ temp6609;
    assign temp6611 = temp6610 ^ temp6610;
    assign temp6612 = temp6611 ^ temp6611;
    assign temp6613 = temp6612 ^ temp6612;
    assign temp6614 = temp6613 ^ temp6613;
    assign temp6615 = temp6614 ^ temp6614;
    assign temp6616 = temp6615 ^ temp6615;
    assign temp6617 = temp6616 ^ temp6616;
    assign temp6618 = temp6617 ^ temp6617;
    assign temp6619 = temp6618 ^ temp6618;
    assign temp6620 = temp6619 ^ temp6619;
    assign temp6621 = temp6620 ^ temp6620;
    assign temp6622 = temp6621 ^ temp6621;
    assign temp6623 = temp6622 ^ temp6622;
    assign temp6624 = temp6623 ^ temp6623;
    assign temp6625 = temp6624 ^ temp6624;
    assign temp6626 = temp6625 ^ temp6625;
    assign temp6627 = temp6626 ^ temp6626;
    assign temp6628 = temp6627 ^ temp6627;
    assign temp6629 = temp6628 ^ temp6628;
    assign temp6630 = temp6629 ^ temp6629;
    assign temp6631 = temp6630 ^ temp6630;
    assign temp6632 = temp6631 ^ temp6631;
    assign temp6633 = temp6632 ^ temp6632;
    assign temp6634 = temp6633 ^ temp6633;
    assign temp6635 = temp6634 ^ temp6634;
    assign temp6636 = temp6635 ^ temp6635;
    assign temp6637 = temp6636 ^ temp6636;
    assign temp6638 = temp6637 ^ temp6637;
    assign temp6639 = temp6638 ^ temp6638;
    assign temp6640 = temp6639 ^ temp6639;
    assign temp6641 = temp6640 ^ temp6640;
    assign temp6642 = temp6641 ^ temp6641;
    assign temp6643 = temp6642 ^ temp6642;
    assign temp6644 = temp6643 ^ temp6643;
    assign temp6645 = temp6644 ^ temp6644;
    assign temp6646 = temp6645 ^ temp6645;
    assign temp6647 = temp6646 ^ temp6646;
    assign temp6648 = temp6647 ^ temp6647;
    assign temp6649 = temp6648 ^ temp6648;
    assign temp6650 = temp6649 ^ temp6649;
    assign temp6651 = temp6650 ^ temp6650;
    assign temp6652 = temp6651 ^ temp6651;
    assign temp6653 = temp6652 ^ temp6652;
    assign temp6654 = temp6653 ^ temp6653;
    assign temp6655 = temp6654 ^ temp6654;
    assign temp6656 = temp6655 ^ temp6655;
    assign temp6657 = temp6656 ^ temp6656;
    assign temp6658 = temp6657 ^ temp6657;
    assign temp6659 = temp6658 ^ temp6658;
    assign temp6660 = temp6659 ^ temp6659;
    assign temp6661 = temp6660 ^ temp6660;
    assign temp6662 = temp6661 ^ temp6661;
    assign temp6663 = temp6662 ^ temp6662;
    assign temp6664 = temp6663 ^ temp6663;
    assign temp6665 = temp6664 ^ temp6664;
    assign temp6666 = temp6665 ^ temp6665;
    assign temp6667 = temp6666 ^ temp6666;
    assign temp6668 = temp6667 ^ temp6667;
    assign temp6669 = temp6668 ^ temp6668;
    assign temp6670 = temp6669 ^ temp6669;
    assign temp6671 = temp6670 ^ temp6670;
    assign temp6672 = temp6671 ^ temp6671;
    assign temp6673 = temp6672 ^ temp6672;
    assign temp6674 = temp6673 ^ temp6673;
    assign temp6675 = temp6674 ^ temp6674;
    assign temp6676 = temp6675 ^ temp6675;
    assign temp6677 = temp6676 ^ temp6676;
    assign temp6678 = temp6677 ^ temp6677;
    assign temp6679 = temp6678 ^ temp6678;
    assign temp6680 = temp6679 ^ temp6679;
    assign temp6681 = temp6680 ^ temp6680;
    assign temp6682 = temp6681 ^ temp6681;
    assign temp6683 = temp6682 ^ temp6682;
    assign temp6684 = temp6683 ^ temp6683;
    assign temp6685 = temp6684 ^ temp6684;
    assign temp6686 = temp6685 ^ temp6685;
    assign temp6687 = temp6686 ^ temp6686;
    assign temp6688 = temp6687 ^ temp6687;
    assign temp6689 = temp6688 ^ temp6688;
    assign temp6690 = temp6689 ^ temp6689;
    assign temp6691 = temp6690 ^ temp6690;
    assign temp6692 = temp6691 ^ temp6691;
    assign temp6693 = temp6692 ^ temp6692;
    assign temp6694 = temp6693 ^ temp6693;
    assign temp6695 = temp6694 ^ temp6694;
    assign temp6696 = temp6695 ^ temp6695;
    assign temp6697 = temp6696 ^ temp6696;
    assign temp6698 = temp6697 ^ temp6697;
    assign temp6699 = temp6698 ^ temp6698;
    assign temp6700 = temp6699 ^ temp6699;
    assign temp6701 = temp6700 ^ temp6700;
    assign temp6702 = temp6701 ^ temp6701;
    assign temp6703 = temp6702 ^ temp6702;
    assign temp6704 = temp6703 ^ temp6703;
    assign temp6705 = temp6704 ^ temp6704;
    assign temp6706 = temp6705 ^ temp6705;
    assign temp6707 = temp6706 ^ temp6706;
    assign temp6708 = temp6707 ^ temp6707;
    assign temp6709 = temp6708 ^ temp6708;
    assign temp6710 = temp6709 ^ temp6709;
    assign temp6711 = temp6710 ^ temp6710;
    assign temp6712 = temp6711 ^ temp6711;
    assign temp6713 = temp6712 ^ temp6712;
    assign temp6714 = temp6713 ^ temp6713;
    assign temp6715 = temp6714 ^ temp6714;
    assign temp6716 = temp6715 ^ temp6715;
    assign temp6717 = temp6716 ^ temp6716;
    assign temp6718 = temp6717 ^ temp6717;
    assign temp6719 = temp6718 ^ temp6718;
    assign temp6720 = temp6719 ^ temp6719;
    assign temp6721 = temp6720 ^ temp6720;
    assign temp6722 = temp6721 ^ temp6721;
    assign temp6723 = temp6722 ^ temp6722;
    assign temp6724 = temp6723 ^ temp6723;
    assign temp6725 = temp6724 ^ temp6724;
    assign temp6726 = temp6725 ^ temp6725;
    assign temp6727 = temp6726 ^ temp6726;
    assign temp6728 = temp6727 ^ temp6727;
    assign temp6729 = temp6728 ^ temp6728;
    assign temp6730 = temp6729 ^ temp6729;
    assign temp6731 = temp6730 ^ temp6730;
    assign temp6732 = temp6731 ^ temp6731;
    assign temp6733 = temp6732 ^ temp6732;
    assign temp6734 = temp6733 ^ temp6733;
    assign temp6735 = temp6734 ^ temp6734;
    assign temp6736 = temp6735 ^ temp6735;
    assign temp6737 = temp6736 ^ temp6736;
    assign temp6738 = temp6737 ^ temp6737;
    assign temp6739 = temp6738 ^ temp6738;
    assign temp6740 = temp6739 ^ temp6739;
    assign temp6741 = temp6740 ^ temp6740;
    assign temp6742 = temp6741 ^ temp6741;
    assign temp6743 = temp6742 ^ temp6742;
    assign temp6744 = temp6743 ^ temp6743;
    assign temp6745 = temp6744 ^ temp6744;
    assign temp6746 = temp6745 ^ temp6745;
    assign temp6747 = temp6746 ^ temp6746;
    assign temp6748 = temp6747 ^ temp6747;
    assign temp6749 = temp6748 ^ temp6748;
    assign temp6750 = temp6749 ^ temp6749;
    assign temp6751 = temp6750 ^ temp6750;
    assign temp6752 = temp6751 ^ temp6751;
    assign temp6753 = temp6752 ^ temp6752;
    assign temp6754 = temp6753 ^ temp6753;
    assign temp6755 = temp6754 ^ temp6754;
    assign temp6756 = temp6755 ^ temp6755;
    assign temp6757 = temp6756 ^ temp6756;
    assign temp6758 = temp6757 ^ temp6757;
    assign temp6759 = temp6758 ^ temp6758;
    assign temp6760 = temp6759 ^ temp6759;
    assign temp6761 = temp6760 ^ temp6760;
    assign temp6762 = temp6761 ^ temp6761;
    assign temp6763 = temp6762 ^ temp6762;
    assign temp6764 = temp6763 ^ temp6763;
    assign temp6765 = temp6764 ^ temp6764;
    assign temp6766 = temp6765 ^ temp6765;
    assign temp6767 = temp6766 ^ temp6766;
    assign temp6768 = temp6767 ^ temp6767;
    assign temp6769 = temp6768 ^ temp6768;
    assign temp6770 = temp6769 ^ temp6769;
    assign temp6771 = temp6770 ^ temp6770;
    assign temp6772 = temp6771 ^ temp6771;
    assign temp6773 = temp6772 ^ temp6772;
    assign temp6774 = temp6773 ^ temp6773;
    assign temp6775 = temp6774 ^ temp6774;
    assign temp6776 = temp6775 ^ temp6775;
    assign temp6777 = temp6776 ^ temp6776;
    assign temp6778 = temp6777 ^ temp6777;
    assign temp6779 = temp6778 ^ temp6778;
    assign temp6780 = temp6779 ^ temp6779;
    assign temp6781 = temp6780 ^ temp6780;
    assign temp6782 = temp6781 ^ temp6781;
    assign temp6783 = temp6782 ^ temp6782;
    assign temp6784 = temp6783 ^ temp6783;
    assign temp6785 = temp6784 ^ temp6784;
    assign temp6786 = temp6785 ^ temp6785;
    assign temp6787 = temp6786 ^ temp6786;
    assign temp6788 = temp6787 ^ temp6787;
    assign temp6789 = temp6788 ^ temp6788;
    assign temp6790 = temp6789 ^ temp6789;
    assign temp6791 = temp6790 ^ temp6790;
    assign temp6792 = temp6791 ^ temp6791;
    assign temp6793 = temp6792 ^ temp6792;
    assign temp6794 = temp6793 ^ temp6793;
    assign temp6795 = temp6794 ^ temp6794;
    assign temp6796 = temp6795 ^ temp6795;
    assign temp6797 = temp6796 ^ temp6796;
    assign temp6798 = temp6797 ^ temp6797;
    assign temp6799 = temp6798 ^ temp6798;
    assign temp6800 = temp6799 ^ temp6799;
    assign temp6801 = temp6800 ^ temp6800;
    assign temp6802 = temp6801 ^ temp6801;
    assign temp6803 = temp6802 ^ temp6802;
    assign temp6804 = temp6803 ^ temp6803;
    assign temp6805 = temp6804 ^ temp6804;
    assign temp6806 = temp6805 ^ temp6805;
    assign temp6807 = temp6806 ^ temp6806;
    assign temp6808 = temp6807 ^ temp6807;
    assign temp6809 = temp6808 ^ temp6808;
    assign temp6810 = temp6809 ^ temp6809;
    assign temp6811 = temp6810 ^ temp6810;
    assign temp6812 = temp6811 ^ temp6811;
    assign temp6813 = temp6812 ^ temp6812;
    assign temp6814 = temp6813 ^ temp6813;
    assign temp6815 = temp6814 ^ temp6814;
    assign temp6816 = temp6815 ^ temp6815;
    assign temp6817 = temp6816 ^ temp6816;
    assign temp6818 = temp6817 ^ temp6817;
    assign temp6819 = temp6818 ^ temp6818;
    assign temp6820 = temp6819 ^ temp6819;
    assign temp6821 = temp6820 ^ temp6820;
    assign temp6822 = temp6821 ^ temp6821;
    assign temp6823 = temp6822 ^ temp6822;
    assign temp6824 = temp6823 ^ temp6823;
    assign temp6825 = temp6824 ^ temp6824;
    assign temp6826 = temp6825 ^ temp6825;
    assign temp6827 = temp6826 ^ temp6826;
    assign temp6828 = temp6827 ^ temp6827;
    assign temp6829 = temp6828 ^ temp6828;
    assign temp6830 = temp6829 ^ temp6829;
    assign temp6831 = temp6830 ^ temp6830;
    assign temp6832 = temp6831 ^ temp6831;
    assign temp6833 = temp6832 ^ temp6832;
    assign temp6834 = temp6833 ^ temp6833;
    assign temp6835 = temp6834 ^ temp6834;
    assign temp6836 = temp6835 ^ temp6835;
    assign temp6837 = temp6836 ^ temp6836;
    assign temp6838 = temp6837 ^ temp6837;
    assign temp6839 = temp6838 ^ temp6838;
    assign temp6840 = temp6839 ^ temp6839;
    assign temp6841 = temp6840 ^ temp6840;
    assign temp6842 = temp6841 ^ temp6841;
    assign temp6843 = temp6842 ^ temp6842;
    assign temp6844 = temp6843 ^ temp6843;
    assign temp6845 = temp6844 ^ temp6844;
    assign temp6846 = temp6845 ^ temp6845;
    assign temp6847 = temp6846 ^ temp6846;
    assign temp6848 = temp6847 ^ temp6847;
    assign temp6849 = temp6848 ^ temp6848;
    assign temp6850 = temp6849 ^ temp6849;
    assign temp6851 = temp6850 ^ temp6850;
    assign temp6852 = temp6851 ^ temp6851;
    assign temp6853 = temp6852 ^ temp6852;
    assign temp6854 = temp6853 ^ temp6853;
    assign temp6855 = temp6854 ^ temp6854;
    assign temp6856 = temp6855 ^ temp6855;
    assign temp6857 = temp6856 ^ temp6856;
    assign temp6858 = temp6857 ^ temp6857;
    assign temp6859 = temp6858 ^ temp6858;
    assign temp6860 = temp6859 ^ temp6859;
    assign temp6861 = temp6860 ^ temp6860;
    assign temp6862 = temp6861 ^ temp6861;
    assign temp6863 = temp6862 ^ temp6862;
    assign temp6864 = temp6863 ^ temp6863;
    assign temp6865 = temp6864 ^ temp6864;
    assign temp6866 = temp6865 ^ temp6865;
    assign temp6867 = temp6866 ^ temp6866;
    assign temp6868 = temp6867 ^ temp6867;
    assign temp6869 = temp6868 ^ temp6868;
    assign temp6870 = temp6869 ^ temp6869;
    assign temp6871 = temp6870 ^ temp6870;
    assign temp6872 = temp6871 ^ temp6871;
    assign temp6873 = temp6872 ^ temp6872;
    assign temp6874 = temp6873 ^ temp6873;
    assign temp6875 = temp6874 ^ temp6874;
    assign temp6876 = temp6875 ^ temp6875;
    assign temp6877 = temp6876 ^ temp6876;
    assign temp6878 = temp6877 ^ temp6877;
    assign temp6879 = temp6878 ^ temp6878;
    assign temp6880 = temp6879 ^ temp6879;
    assign temp6881 = temp6880 ^ temp6880;
    assign temp6882 = temp6881 ^ temp6881;
    assign temp6883 = temp6882 ^ temp6882;
    assign temp6884 = temp6883 ^ temp6883;
    assign temp6885 = temp6884 ^ temp6884;
    assign temp6886 = temp6885 ^ temp6885;
    assign temp6887 = temp6886 ^ temp6886;
    assign temp6888 = temp6887 ^ temp6887;
    assign temp6889 = temp6888 ^ temp6888;
    assign temp6890 = temp6889 ^ temp6889;
    assign temp6891 = temp6890 ^ temp6890;
    assign temp6892 = temp6891 ^ temp6891;
    assign temp6893 = temp6892 ^ temp6892;
    assign temp6894 = temp6893 ^ temp6893;
    assign temp6895 = temp6894 ^ temp6894;
    assign temp6896 = temp6895 ^ temp6895;
    assign temp6897 = temp6896 ^ temp6896;
    assign temp6898 = temp6897 ^ temp6897;
    assign temp6899 = temp6898 ^ temp6898;
    assign temp6900 = temp6899 ^ temp6899;
    assign temp6901 = temp6900 ^ temp6900;
    assign temp6902 = temp6901 ^ temp6901;
    assign temp6903 = temp6902 ^ temp6902;
    assign temp6904 = temp6903 ^ temp6903;
    assign temp6905 = temp6904 ^ temp6904;
    assign temp6906 = temp6905 ^ temp6905;
    assign temp6907 = temp6906 ^ temp6906;
    assign temp6908 = temp6907 ^ temp6907;
    assign temp6909 = temp6908 ^ temp6908;
    assign temp6910 = temp6909 ^ temp6909;
    assign temp6911 = temp6910 ^ temp6910;
    assign temp6912 = temp6911 ^ temp6911;
    assign temp6913 = temp6912 ^ temp6912;
    assign temp6914 = temp6913 ^ temp6913;
    assign temp6915 = temp6914 ^ temp6914;
    assign temp6916 = temp6915 ^ temp6915;
    assign temp6917 = temp6916 ^ temp6916;
    assign temp6918 = temp6917 ^ temp6917;
    assign temp6919 = temp6918 ^ temp6918;
    assign temp6920 = temp6919 ^ temp6919;
    assign temp6921 = temp6920 ^ temp6920;
    assign temp6922 = temp6921 ^ temp6921;
    assign temp6923 = temp6922 ^ temp6922;
    assign temp6924 = temp6923 ^ temp6923;
    assign temp6925 = temp6924 ^ temp6924;
    assign temp6926 = temp6925 ^ temp6925;
    assign temp6927 = temp6926 ^ temp6926;
    assign temp6928 = temp6927 ^ temp6927;
    assign temp6929 = temp6928 ^ temp6928;
    assign temp6930 = temp6929 ^ temp6929;
    assign temp6931 = temp6930 ^ temp6930;
    assign temp6932 = temp6931 ^ temp6931;
    assign temp6933 = temp6932 ^ temp6932;
    assign temp6934 = temp6933 ^ temp6933;
    assign temp6935 = temp6934 ^ temp6934;
    assign temp6936 = temp6935 ^ temp6935;
    assign temp6937 = temp6936 ^ temp6936;
    assign temp6938 = temp6937 ^ temp6937;
    assign temp6939 = temp6938 ^ temp6938;
    assign temp6940 = temp6939 ^ temp6939;
    assign temp6941 = temp6940 ^ temp6940;
    assign temp6942 = temp6941 ^ temp6941;
    assign temp6943 = temp6942 ^ temp6942;
    assign temp6944 = temp6943 ^ temp6943;
    assign temp6945 = temp6944 ^ temp6944;
    assign temp6946 = temp6945 ^ temp6945;
    assign temp6947 = temp6946 ^ temp6946;
    assign temp6948 = temp6947 ^ temp6947;
    assign temp6949 = temp6948 ^ temp6948;
    assign temp6950 = temp6949 ^ temp6949;
    assign temp6951 = temp6950 ^ temp6950;
    assign temp6952 = temp6951 ^ temp6951;
    assign temp6953 = temp6952 ^ temp6952;
    assign temp6954 = temp6953 ^ temp6953;
    assign temp6955 = temp6954 ^ temp6954;
    assign temp6956 = temp6955 ^ temp6955;
    assign temp6957 = temp6956 ^ temp6956;
    assign temp6958 = temp6957 ^ temp6957;
    assign temp6959 = temp6958 ^ temp6958;
    assign temp6960 = temp6959 ^ temp6959;
    assign temp6961 = temp6960 ^ temp6960;
    assign temp6962 = temp6961 ^ temp6961;
    assign temp6963 = temp6962 ^ temp6962;
    assign temp6964 = temp6963 ^ temp6963;
    assign temp6965 = temp6964 ^ temp6964;
    assign temp6966 = temp6965 ^ temp6965;
    assign temp6967 = temp6966 ^ temp6966;
    assign temp6968 = temp6967 ^ temp6967;
    assign temp6969 = temp6968 ^ temp6968;
    assign temp6970 = temp6969 ^ temp6969;
    assign temp6971 = temp6970 ^ temp6970;
    assign temp6972 = temp6971 ^ temp6971;
    assign temp6973 = temp6972 ^ temp6972;
    assign temp6974 = temp6973 ^ temp6973;
    assign temp6975 = temp6974 ^ temp6974;
    assign temp6976 = temp6975 ^ temp6975;
    assign temp6977 = temp6976 ^ temp6976;
    assign temp6978 = temp6977 ^ temp6977;
    assign temp6979 = temp6978 ^ temp6978;
    assign temp6980 = temp6979 ^ temp6979;
    assign temp6981 = temp6980 ^ temp6980;
    assign temp6982 = temp6981 ^ temp6981;
    assign temp6983 = temp6982 ^ temp6982;
    assign temp6984 = temp6983 ^ temp6983;
    assign temp6985 = temp6984 ^ temp6984;
    assign temp6986 = temp6985 ^ temp6985;
    assign temp6987 = temp6986 ^ temp6986;
    assign temp6988 = temp6987 ^ temp6987;
    assign temp6989 = temp6988 ^ temp6988;
    assign temp6990 = temp6989 ^ temp6989;
    assign temp6991 = temp6990 ^ temp6990;
    assign temp6992 = temp6991 ^ temp6991;
    assign temp6993 = temp6992 ^ temp6992;
    assign temp6994 = temp6993 ^ temp6993;
    assign temp6995 = temp6994 ^ temp6994;
    assign temp6996 = temp6995 ^ temp6995;
    assign temp6997 = temp6996 ^ temp6996;
    assign temp6998 = temp6997 ^ temp6997;
    assign temp6999 = temp6998 ^ temp6998;
    assign temp7000 = temp6999 ^ temp6999;
    assign temp7001 = temp7000 ^ temp7000;
    assign temp7002 = temp7001 ^ temp7001;
    assign temp7003 = temp7002 ^ temp7002;
    assign temp7004 = temp7003 ^ temp7003;
    assign temp7005 = temp7004 ^ temp7004;
    assign temp7006 = temp7005 ^ temp7005;
    assign temp7007 = temp7006 ^ temp7006;
    assign temp7008 = temp7007 ^ temp7007;
    assign temp7009 = temp7008 ^ temp7008;
    assign temp7010 = temp7009 ^ temp7009;
    assign temp7011 = temp7010 ^ temp7010;
    assign temp7012 = temp7011 ^ temp7011;
    assign temp7013 = temp7012 ^ temp7012;
    assign temp7014 = temp7013 ^ temp7013;
    assign temp7015 = temp7014 ^ temp7014;
    assign temp7016 = temp7015 ^ temp7015;
    assign temp7017 = temp7016 ^ temp7016;
    assign temp7018 = temp7017 ^ temp7017;
    assign temp7019 = temp7018 ^ temp7018;
    assign temp7020 = temp7019 ^ temp7019;
    assign temp7021 = temp7020 ^ temp7020;
    assign temp7022 = temp7021 ^ temp7021;
    assign temp7023 = temp7022 ^ temp7022;
    assign temp7024 = temp7023 ^ temp7023;
    assign temp7025 = temp7024 ^ temp7024;
    assign temp7026 = temp7025 ^ temp7025;
    assign temp7027 = temp7026 ^ temp7026;
    assign temp7028 = temp7027 ^ temp7027;
    assign temp7029 = temp7028 ^ temp7028;
    assign temp7030 = temp7029 ^ temp7029;
    assign temp7031 = temp7030 ^ temp7030;
    assign temp7032 = temp7031 ^ temp7031;
    assign temp7033 = temp7032 ^ temp7032;
    assign temp7034 = temp7033 ^ temp7033;
    assign temp7035 = temp7034 ^ temp7034;
    assign temp7036 = temp7035 ^ temp7035;
    assign temp7037 = temp7036 ^ temp7036;
    assign temp7038 = temp7037 ^ temp7037;
    assign temp7039 = temp7038 ^ temp7038;
    assign temp7040 = temp7039 ^ temp7039;
    assign temp7041 = temp7040 ^ temp7040;
    assign temp7042 = temp7041 ^ temp7041;
    assign temp7043 = temp7042 ^ temp7042;
    assign temp7044 = temp7043 ^ temp7043;
    assign temp7045 = temp7044 ^ temp7044;
    assign temp7046 = temp7045 ^ temp7045;
    assign temp7047 = temp7046 ^ temp7046;
    assign temp7048 = temp7047 ^ temp7047;
    assign temp7049 = temp7048 ^ temp7048;
    assign temp7050 = temp7049 ^ temp7049;
    assign temp7051 = temp7050 ^ temp7050;
    assign temp7052 = temp7051 ^ temp7051;
    assign temp7053 = temp7052 ^ temp7052;
    assign temp7054 = temp7053 ^ temp7053;
    assign temp7055 = temp7054 ^ temp7054;
    assign temp7056 = temp7055 ^ temp7055;
    assign temp7057 = temp7056 ^ temp7056;
    assign temp7058 = temp7057 ^ temp7057;
    assign temp7059 = temp7058 ^ temp7058;
    assign temp7060 = temp7059 ^ temp7059;
    assign temp7061 = temp7060 ^ temp7060;
    assign temp7062 = temp7061 ^ temp7061;
    assign temp7063 = temp7062 ^ temp7062;
    assign temp7064 = temp7063 ^ temp7063;
    assign temp7065 = temp7064 ^ temp7064;
    assign temp7066 = temp7065 ^ temp7065;
    assign temp7067 = temp7066 ^ temp7066;
    assign temp7068 = temp7067 ^ temp7067;
    assign temp7069 = temp7068 ^ temp7068;
    assign temp7070 = temp7069 ^ temp7069;
    assign temp7071 = temp7070 ^ temp7070;
    assign temp7072 = temp7071 ^ temp7071;
    assign temp7073 = temp7072 ^ temp7072;
    assign temp7074 = temp7073 ^ temp7073;
    assign temp7075 = temp7074 ^ temp7074;
    assign temp7076 = temp7075 ^ temp7075;
    assign temp7077 = temp7076 ^ temp7076;
    assign temp7078 = temp7077 ^ temp7077;
    assign temp7079 = temp7078 ^ temp7078;
    assign temp7080 = temp7079 ^ temp7079;
    assign temp7081 = temp7080 ^ temp7080;
    assign temp7082 = temp7081 ^ temp7081;
    assign temp7083 = temp7082 ^ temp7082;
    assign temp7084 = temp7083 ^ temp7083;
    assign temp7085 = temp7084 ^ temp7084;
    assign temp7086 = temp7085 ^ temp7085;
    assign temp7087 = temp7086 ^ temp7086;
    assign temp7088 = temp7087 ^ temp7087;
    assign temp7089 = temp7088 ^ temp7088;
    assign temp7090 = temp7089 ^ temp7089;
    assign temp7091 = temp7090 ^ temp7090;
    assign temp7092 = temp7091 ^ temp7091;
    assign temp7093 = temp7092 ^ temp7092;
    assign temp7094 = temp7093 ^ temp7093;
    assign temp7095 = temp7094 ^ temp7094;
    assign temp7096 = temp7095 ^ temp7095;
    assign temp7097 = temp7096 ^ temp7096;
    assign temp7098 = temp7097 ^ temp7097;
    assign temp7099 = temp7098 ^ temp7098;
    assign temp7100 = temp7099 ^ temp7099;
    assign temp7101 = temp7100 ^ temp7100;
    assign temp7102 = temp7101 ^ temp7101;
    assign temp7103 = temp7102 ^ temp7102;
    assign temp7104 = temp7103 ^ temp7103;
    assign temp7105 = temp7104 ^ temp7104;
    assign temp7106 = temp7105 ^ temp7105;
    assign temp7107 = temp7106 ^ temp7106;
    assign temp7108 = temp7107 ^ temp7107;
    assign temp7109 = temp7108 ^ temp7108;
    assign temp7110 = temp7109 ^ temp7109;
    assign temp7111 = temp7110 ^ temp7110;
    assign temp7112 = temp7111 ^ temp7111;
    assign temp7113 = temp7112 ^ temp7112;
    assign temp7114 = temp7113 ^ temp7113;
    assign temp7115 = temp7114 ^ temp7114;
    assign temp7116 = temp7115 ^ temp7115;
    assign temp7117 = temp7116 ^ temp7116;
    assign temp7118 = temp7117 ^ temp7117;
    assign temp7119 = temp7118 ^ temp7118;
    assign temp7120 = temp7119 ^ temp7119;
    assign temp7121 = temp7120 ^ temp7120;
    assign temp7122 = temp7121 ^ temp7121;
    assign temp7123 = temp7122 ^ temp7122;
    assign temp7124 = temp7123 ^ temp7123;
    assign temp7125 = temp7124 ^ temp7124;
    assign temp7126 = temp7125 ^ temp7125;
    assign temp7127 = temp7126 ^ temp7126;
    assign temp7128 = temp7127 ^ temp7127;
    assign temp7129 = temp7128 ^ temp7128;
    assign temp7130 = temp7129 ^ temp7129;
    assign temp7131 = temp7130 ^ temp7130;
    assign temp7132 = temp7131 ^ temp7131;
    assign temp7133 = temp7132 ^ temp7132;
    assign temp7134 = temp7133 ^ temp7133;
    assign temp7135 = temp7134 ^ temp7134;
    assign temp7136 = temp7135 ^ temp7135;
    assign temp7137 = temp7136 ^ temp7136;
    assign temp7138 = temp7137 ^ temp7137;
    assign temp7139 = temp7138 ^ temp7138;
    assign temp7140 = temp7139 ^ temp7139;
    assign temp7141 = temp7140 ^ temp7140;
    assign temp7142 = temp7141 ^ temp7141;
    assign temp7143 = temp7142 ^ temp7142;
    assign temp7144 = temp7143 ^ temp7143;
    assign temp7145 = temp7144 ^ temp7144;
    assign temp7146 = temp7145 ^ temp7145;
    assign temp7147 = temp7146 ^ temp7146;
    assign temp7148 = temp7147 ^ temp7147;
    assign temp7149 = temp7148 ^ temp7148;
    assign temp7150 = temp7149 ^ temp7149;
    assign temp7151 = temp7150 ^ temp7150;
    assign temp7152 = temp7151 ^ temp7151;
    assign temp7153 = temp7152 ^ temp7152;
    assign temp7154 = temp7153 ^ temp7153;
    assign temp7155 = temp7154 ^ temp7154;
    assign temp7156 = temp7155 ^ temp7155;
    assign temp7157 = temp7156 ^ temp7156;
    assign temp7158 = temp7157 ^ temp7157;
    assign temp7159 = temp7158 ^ temp7158;
    assign temp7160 = temp7159 ^ temp7159;
    assign temp7161 = temp7160 ^ temp7160;
    assign temp7162 = temp7161 ^ temp7161;
    assign temp7163 = temp7162 ^ temp7162;
    assign temp7164 = temp7163 ^ temp7163;
    assign temp7165 = temp7164 ^ temp7164;
    assign temp7166 = temp7165 ^ temp7165;
    assign temp7167 = temp7166 ^ temp7166;
    assign temp7168 = temp7167 ^ temp7167;
    assign temp7169 = temp7168 ^ temp7168;
    assign temp7170 = temp7169 ^ temp7169;
    assign temp7171 = temp7170 ^ temp7170;
    assign temp7172 = temp7171 ^ temp7171;
    assign temp7173 = temp7172 ^ temp7172;
    assign temp7174 = temp7173 ^ temp7173;
    assign temp7175 = temp7174 ^ temp7174;
    assign temp7176 = temp7175 ^ temp7175;
    assign temp7177 = temp7176 ^ temp7176;
    assign temp7178 = temp7177 ^ temp7177;
    assign temp7179 = temp7178 ^ temp7178;
    assign temp7180 = temp7179 ^ temp7179;
    assign temp7181 = temp7180 ^ temp7180;
    assign temp7182 = temp7181 ^ temp7181;
    assign temp7183 = temp7182 ^ temp7182;
    assign temp7184 = temp7183 ^ temp7183;
    assign temp7185 = temp7184 ^ temp7184;
    assign temp7186 = temp7185 ^ temp7185;
    assign temp7187 = temp7186 ^ temp7186;
    assign temp7188 = temp7187 ^ temp7187;
    assign temp7189 = temp7188 ^ temp7188;
    assign temp7190 = temp7189 ^ temp7189;
    assign temp7191 = temp7190 ^ temp7190;
    assign temp7192 = temp7191 ^ temp7191;
    assign temp7193 = temp7192 ^ temp7192;
    assign temp7194 = temp7193 ^ temp7193;
    assign temp7195 = temp7194 ^ temp7194;
    assign temp7196 = temp7195 ^ temp7195;
    assign temp7197 = temp7196 ^ temp7196;
    assign temp7198 = temp7197 ^ temp7197;
    assign temp7199 = temp7198 ^ temp7198;
    assign temp7200 = temp7199 ^ temp7199;
    assign temp7201 = temp7200 ^ temp7200;
    assign temp7202 = temp7201 ^ temp7201;
    assign temp7203 = temp7202 ^ temp7202;
    assign temp7204 = temp7203 ^ temp7203;
    assign temp7205 = temp7204 ^ temp7204;
    assign temp7206 = temp7205 ^ temp7205;
    assign temp7207 = temp7206 ^ temp7206;
    assign temp7208 = temp7207 ^ temp7207;
    assign temp7209 = temp7208 ^ temp7208;
    assign temp7210 = temp7209 ^ temp7209;
    assign temp7211 = temp7210 ^ temp7210;
    assign temp7212 = temp7211 ^ temp7211;
    assign temp7213 = temp7212 ^ temp7212;
    assign temp7214 = temp7213 ^ temp7213;
    assign temp7215 = temp7214 ^ temp7214;
    assign temp7216 = temp7215 ^ temp7215;
    assign temp7217 = temp7216 ^ temp7216;
    assign temp7218 = temp7217 ^ temp7217;
    assign temp7219 = temp7218 ^ temp7218;
    assign temp7220 = temp7219 ^ temp7219;
    assign temp7221 = temp7220 ^ temp7220;
    assign temp7222 = temp7221 ^ temp7221;
    assign temp7223 = temp7222 ^ temp7222;
    assign temp7224 = temp7223 ^ temp7223;
    assign temp7225 = temp7224 ^ temp7224;
    assign temp7226 = temp7225 ^ temp7225;
    assign temp7227 = temp7226 ^ temp7226;
    assign temp7228 = temp7227 ^ temp7227;
    assign temp7229 = temp7228 ^ temp7228;
    assign temp7230 = temp7229 ^ temp7229;
    assign temp7231 = temp7230 ^ temp7230;
    assign temp7232 = temp7231 ^ temp7231;
    assign temp7233 = temp7232 ^ temp7232;
    assign temp7234 = temp7233 ^ temp7233;
    assign temp7235 = temp7234 ^ temp7234;
    assign temp7236 = temp7235 ^ temp7235;
    assign temp7237 = temp7236 ^ temp7236;
    assign temp7238 = temp7237 ^ temp7237;
    assign temp7239 = temp7238 ^ temp7238;
    assign temp7240 = temp7239 ^ temp7239;
    assign temp7241 = temp7240 ^ temp7240;
    assign temp7242 = temp7241 ^ temp7241;
    assign temp7243 = temp7242 ^ temp7242;
    assign temp7244 = temp7243 ^ temp7243;
    assign temp7245 = temp7244 ^ temp7244;
    assign temp7246 = temp7245 ^ temp7245;
    assign temp7247 = temp7246 ^ temp7246;
    assign temp7248 = temp7247 ^ temp7247;
    assign temp7249 = temp7248 ^ temp7248;
    assign temp7250 = temp7249 ^ temp7249;
    assign temp7251 = temp7250 ^ temp7250;
    assign temp7252 = temp7251 ^ temp7251;
    assign temp7253 = temp7252 ^ temp7252;
    assign temp7254 = temp7253 ^ temp7253;
    assign temp7255 = temp7254 ^ temp7254;
    assign temp7256 = temp7255 ^ temp7255;
    assign temp7257 = temp7256 ^ temp7256;
    assign temp7258 = temp7257 ^ temp7257;
    assign temp7259 = temp7258 ^ temp7258;
    assign temp7260 = temp7259 ^ temp7259;
    assign temp7261 = temp7260 ^ temp7260;
    assign temp7262 = temp7261 ^ temp7261;
    assign temp7263 = temp7262 ^ temp7262;
    assign temp7264 = temp7263 ^ temp7263;
    assign temp7265 = temp7264 ^ temp7264;
    assign temp7266 = temp7265 ^ temp7265;
    assign temp7267 = temp7266 ^ temp7266;
    assign temp7268 = temp7267 ^ temp7267;
    assign temp7269 = temp7268 ^ temp7268;
    assign temp7270 = temp7269 ^ temp7269;
    assign temp7271 = temp7270 ^ temp7270;
    assign temp7272 = temp7271 ^ temp7271;
    assign temp7273 = temp7272 ^ temp7272;
    assign temp7274 = temp7273 ^ temp7273;
    assign temp7275 = temp7274 ^ temp7274;
    assign temp7276 = temp7275 ^ temp7275;
    assign temp7277 = temp7276 ^ temp7276;
    assign temp7278 = temp7277 ^ temp7277;
    assign temp7279 = temp7278 ^ temp7278;
    assign temp7280 = temp7279 ^ temp7279;
    assign temp7281 = temp7280 ^ temp7280;
    assign temp7282 = temp7281 ^ temp7281;
    assign temp7283 = temp7282 ^ temp7282;
    assign temp7284 = temp7283 ^ temp7283;
    assign temp7285 = temp7284 ^ temp7284;
    assign temp7286 = temp7285 ^ temp7285;
    assign temp7287 = temp7286 ^ temp7286;
    assign temp7288 = temp7287 ^ temp7287;
    assign temp7289 = temp7288 ^ temp7288;
    assign temp7290 = temp7289 ^ temp7289;
    assign temp7291 = temp7290 ^ temp7290;
    assign temp7292 = temp7291 ^ temp7291;
    assign temp7293 = temp7292 ^ temp7292;
    assign temp7294 = temp7293 ^ temp7293;
    assign temp7295 = temp7294 ^ temp7294;
    assign temp7296 = temp7295 ^ temp7295;
    assign temp7297 = temp7296 ^ temp7296;
    assign temp7298 = temp7297 ^ temp7297;
    assign temp7299 = temp7298 ^ temp7298;
    assign temp7300 = temp7299 ^ temp7299;
    assign temp7301 = temp7300 ^ temp7300;
    assign temp7302 = temp7301 ^ temp7301;
    assign temp7303 = temp7302 ^ temp7302;
    assign temp7304 = temp7303 ^ temp7303;
    assign temp7305 = temp7304 ^ temp7304;
    assign temp7306 = temp7305 ^ temp7305;
    assign temp7307 = temp7306 ^ temp7306;
    assign temp7308 = temp7307 ^ temp7307;
    assign temp7309 = temp7308 ^ temp7308;
    assign temp7310 = temp7309 ^ temp7309;
    assign temp7311 = temp7310 ^ temp7310;
    assign temp7312 = temp7311 ^ temp7311;
    assign temp7313 = temp7312 ^ temp7312;
    assign temp7314 = temp7313 ^ temp7313;
    assign temp7315 = temp7314 ^ temp7314;
    assign temp7316 = temp7315 ^ temp7315;
    assign temp7317 = temp7316 ^ temp7316;
    assign temp7318 = temp7317 ^ temp7317;
    assign temp7319 = temp7318 ^ temp7318;
    assign temp7320 = temp7319 ^ temp7319;
    assign temp7321 = temp7320 ^ temp7320;
    assign temp7322 = temp7321 ^ temp7321;
    assign temp7323 = temp7322 ^ temp7322;
    assign temp7324 = temp7323 ^ temp7323;
    assign temp7325 = temp7324 ^ temp7324;
    assign temp7326 = temp7325 ^ temp7325;
    assign temp7327 = temp7326 ^ temp7326;
    assign temp7328 = temp7327 ^ temp7327;
    assign temp7329 = temp7328 ^ temp7328;
    assign temp7330 = temp7329 ^ temp7329;
    assign temp7331 = temp7330 ^ temp7330;
    assign temp7332 = temp7331 ^ temp7331;
    assign temp7333 = temp7332 ^ temp7332;
    assign temp7334 = temp7333 ^ temp7333;
    assign temp7335 = temp7334 ^ temp7334;
    assign temp7336 = temp7335 ^ temp7335;
    assign temp7337 = temp7336 ^ temp7336;
    assign temp7338 = temp7337 ^ temp7337;
    assign temp7339 = temp7338 ^ temp7338;
    assign temp7340 = temp7339 ^ temp7339;
    assign temp7341 = temp7340 ^ temp7340;
    assign temp7342 = temp7341 ^ temp7341;
    assign temp7343 = temp7342 ^ temp7342;
    assign temp7344 = temp7343 ^ temp7343;
    assign temp7345 = temp7344 ^ temp7344;
    assign temp7346 = temp7345 ^ temp7345;
    assign temp7347 = temp7346 ^ temp7346;
    assign temp7348 = temp7347 ^ temp7347;
    assign temp7349 = temp7348 ^ temp7348;
    assign temp7350 = temp7349 ^ temp7349;
    assign temp7351 = temp7350 ^ temp7350;
    assign temp7352 = temp7351 ^ temp7351;
    assign temp7353 = temp7352 ^ temp7352;
    assign temp7354 = temp7353 ^ temp7353;
    assign temp7355 = temp7354 ^ temp7354;
    assign temp7356 = temp7355 ^ temp7355;
    assign temp7357 = temp7356 ^ temp7356;
    assign temp7358 = temp7357 ^ temp7357;
    assign temp7359 = temp7358 ^ temp7358;
    assign temp7360 = temp7359 ^ temp7359;
    assign temp7361 = temp7360 ^ temp7360;
    assign temp7362 = temp7361 ^ temp7361;
    assign temp7363 = temp7362 ^ temp7362;
    assign temp7364 = temp7363 ^ temp7363;
    assign temp7365 = temp7364 ^ temp7364;
    assign temp7366 = temp7365 ^ temp7365;
    assign temp7367 = temp7366 ^ temp7366;
    assign temp7368 = temp7367 ^ temp7367;
    assign temp7369 = temp7368 ^ temp7368;
    assign temp7370 = temp7369 ^ temp7369;
    assign temp7371 = temp7370 ^ temp7370;
    assign temp7372 = temp7371 ^ temp7371;
    assign temp7373 = temp7372 ^ temp7372;
    assign temp7374 = temp7373 ^ temp7373;
    assign temp7375 = temp7374 ^ temp7374;
    assign temp7376 = temp7375 ^ temp7375;
    assign temp7377 = temp7376 ^ temp7376;
    assign temp7378 = temp7377 ^ temp7377;
    assign temp7379 = temp7378 ^ temp7378;
    assign temp7380 = temp7379 ^ temp7379;
    assign temp7381 = temp7380 ^ temp7380;
    assign temp7382 = temp7381 ^ temp7381;
    assign temp7383 = temp7382 ^ temp7382;
    assign temp7384 = temp7383 ^ temp7383;
    assign temp7385 = temp7384 ^ temp7384;
    assign temp7386 = temp7385 ^ temp7385;
    assign temp7387 = temp7386 ^ temp7386;
    assign temp7388 = temp7387 ^ temp7387;
    assign temp7389 = temp7388 ^ temp7388;
    assign temp7390 = temp7389 ^ temp7389;
    assign temp7391 = temp7390 ^ temp7390;
    assign temp7392 = temp7391 ^ temp7391;
    assign temp7393 = temp7392 ^ temp7392;
    assign temp7394 = temp7393 ^ temp7393;
    assign temp7395 = temp7394 ^ temp7394;
    assign temp7396 = temp7395 ^ temp7395;
    assign temp7397 = temp7396 ^ temp7396;
    assign temp7398 = temp7397 ^ temp7397;
    assign temp7399 = temp7398 ^ temp7398;
    assign temp7400 = temp7399 ^ temp7399;
    assign temp7401 = temp7400 ^ temp7400;
    assign temp7402 = temp7401 ^ temp7401;
    assign temp7403 = temp7402 ^ temp7402;
    assign temp7404 = temp7403 ^ temp7403;
    assign temp7405 = temp7404 ^ temp7404;
    assign temp7406 = temp7405 ^ temp7405;
    assign temp7407 = temp7406 ^ temp7406;
    assign temp7408 = temp7407 ^ temp7407;
    assign temp7409 = temp7408 ^ temp7408;
    assign temp7410 = temp7409 ^ temp7409;
    assign temp7411 = temp7410 ^ temp7410;
    assign temp7412 = temp7411 ^ temp7411;
    assign temp7413 = temp7412 ^ temp7412;
    assign temp7414 = temp7413 ^ temp7413;
    assign temp7415 = temp7414 ^ temp7414;
    assign temp7416 = temp7415 ^ temp7415;
    assign temp7417 = temp7416 ^ temp7416;
    assign temp7418 = temp7417 ^ temp7417;
    assign temp7419 = temp7418 ^ temp7418;
    assign temp7420 = temp7419 ^ temp7419;
    assign temp7421 = temp7420 ^ temp7420;
    assign temp7422 = temp7421 ^ temp7421;
    assign temp7423 = temp7422 ^ temp7422;
    assign temp7424 = temp7423 ^ temp7423;
    assign temp7425 = temp7424 ^ temp7424;
    assign temp7426 = temp7425 ^ temp7425;
    assign temp7427 = temp7426 ^ temp7426;
    assign temp7428 = temp7427 ^ temp7427;
    assign temp7429 = temp7428 ^ temp7428;
    assign temp7430 = temp7429 ^ temp7429;
    assign temp7431 = temp7430 ^ temp7430;
    assign temp7432 = temp7431 ^ temp7431;
    assign temp7433 = temp7432 ^ temp7432;
    assign temp7434 = temp7433 ^ temp7433;
    assign temp7435 = temp7434 ^ temp7434;
    assign temp7436 = temp7435 ^ temp7435;
    assign temp7437 = temp7436 ^ temp7436;
    assign temp7438 = temp7437 ^ temp7437;
    assign temp7439 = temp7438 ^ temp7438;
    assign temp7440 = temp7439 ^ temp7439;
    assign temp7441 = temp7440 ^ temp7440;
    assign temp7442 = temp7441 ^ temp7441;
    assign temp7443 = temp7442 ^ temp7442;
    assign temp7444 = temp7443 ^ temp7443;
    assign temp7445 = temp7444 ^ temp7444;
    assign temp7446 = temp7445 ^ temp7445;
    assign temp7447 = temp7446 ^ temp7446;
    assign temp7448 = temp7447 ^ temp7447;
    assign temp7449 = temp7448 ^ temp7448;
    assign temp7450 = temp7449 ^ temp7449;
    assign temp7451 = temp7450 ^ temp7450;
    assign temp7452 = temp7451 ^ temp7451;
    assign temp7453 = temp7452 ^ temp7452;
    assign temp7454 = temp7453 ^ temp7453;
    assign temp7455 = temp7454 ^ temp7454;
    assign temp7456 = temp7455 ^ temp7455;
    assign temp7457 = temp7456 ^ temp7456;
    assign temp7458 = temp7457 ^ temp7457;
    assign temp7459 = temp7458 ^ temp7458;
    assign temp7460 = temp7459 ^ temp7459;
    assign temp7461 = temp7460 ^ temp7460;
    assign temp7462 = temp7461 ^ temp7461;
    assign temp7463 = temp7462 ^ temp7462;
    assign temp7464 = temp7463 ^ temp7463;
    assign temp7465 = temp7464 ^ temp7464;
    assign temp7466 = temp7465 ^ temp7465;
    assign temp7467 = temp7466 ^ temp7466;
    assign temp7468 = temp7467 ^ temp7467;
    assign temp7469 = temp7468 ^ temp7468;
    assign temp7470 = temp7469 ^ temp7469;
    assign temp7471 = temp7470 ^ temp7470;
    assign temp7472 = temp7471 ^ temp7471;
    assign temp7473 = temp7472 ^ temp7472;
    assign temp7474 = temp7473 ^ temp7473;
    assign temp7475 = temp7474 ^ temp7474;
    assign temp7476 = temp7475 ^ temp7475;
    assign temp7477 = temp7476 ^ temp7476;
    assign temp7478 = temp7477 ^ temp7477;
    assign temp7479 = temp7478 ^ temp7478;
    assign temp7480 = temp7479 ^ temp7479;
    assign temp7481 = temp7480 ^ temp7480;
    assign temp7482 = temp7481 ^ temp7481;
    assign temp7483 = temp7482 ^ temp7482;
    assign temp7484 = temp7483 ^ temp7483;
    assign temp7485 = temp7484 ^ temp7484;
    assign temp7486 = temp7485 ^ temp7485;
    assign temp7487 = temp7486 ^ temp7486;
    assign temp7488 = temp7487 ^ temp7487;
    assign temp7489 = temp7488 ^ temp7488;
    assign temp7490 = temp7489 ^ temp7489;
    assign temp7491 = temp7490 ^ temp7490;
    assign temp7492 = temp7491 ^ temp7491;
    assign temp7493 = temp7492 ^ temp7492;
    assign temp7494 = temp7493 ^ temp7493;
    assign temp7495 = temp7494 ^ temp7494;
    assign temp7496 = temp7495 ^ temp7495;
    assign temp7497 = temp7496 ^ temp7496;
    assign temp7498 = temp7497 ^ temp7497;
    assign temp7499 = temp7498 ^ temp7498;
    assign temp7500 = temp7499 ^ temp7499;
    assign temp7501 = temp7500 ^ temp7500;
    assign temp7502 = temp7501 ^ temp7501;
    assign temp7503 = temp7502 ^ temp7502;
    assign temp7504 = temp7503 ^ temp7503;
    assign temp7505 = temp7504 ^ temp7504;
    assign temp7506 = temp7505 ^ temp7505;
    assign temp7507 = temp7506 ^ temp7506;
    assign temp7508 = temp7507 ^ temp7507;
    assign temp7509 = temp7508 ^ temp7508;
    assign temp7510 = temp7509 ^ temp7509;
    assign temp7511 = temp7510 ^ temp7510;
    assign temp7512 = temp7511 ^ temp7511;
    assign temp7513 = temp7512 ^ temp7512;
    assign temp7514 = temp7513 ^ temp7513;
    assign temp7515 = temp7514 ^ temp7514;
    assign temp7516 = temp7515 ^ temp7515;
    assign temp7517 = temp7516 ^ temp7516;
    assign temp7518 = temp7517 ^ temp7517;
    assign temp7519 = temp7518 ^ temp7518;
    assign temp7520 = temp7519 ^ temp7519;
    assign temp7521 = temp7520 ^ temp7520;
    assign temp7522 = temp7521 ^ temp7521;
    assign temp7523 = temp7522 ^ temp7522;
    assign temp7524 = temp7523 ^ temp7523;
    assign temp7525 = temp7524 ^ temp7524;
    assign temp7526 = temp7525 ^ temp7525;
    assign temp7527 = temp7526 ^ temp7526;
    assign temp7528 = temp7527 ^ temp7527;
    assign temp7529 = temp7528 ^ temp7528;
    assign temp7530 = temp7529 ^ temp7529;
    assign temp7531 = temp7530 ^ temp7530;
    assign temp7532 = temp7531 ^ temp7531;
    assign temp7533 = temp7532 ^ temp7532;
    assign temp7534 = temp7533 ^ temp7533;
    assign temp7535 = temp7534 ^ temp7534;
    assign temp7536 = temp7535 ^ temp7535;
    assign temp7537 = temp7536 ^ temp7536;
    assign temp7538 = temp7537 ^ temp7537;
    assign temp7539 = temp7538 ^ temp7538;
    assign temp7540 = temp7539 ^ temp7539;
    assign temp7541 = temp7540 ^ temp7540;
    assign temp7542 = temp7541 ^ temp7541;
    assign temp7543 = temp7542 ^ temp7542;
    assign temp7544 = temp7543 ^ temp7543;
    assign temp7545 = temp7544 ^ temp7544;
    assign temp7546 = temp7545 ^ temp7545;
    assign temp7547 = temp7546 ^ temp7546;
    assign temp7548 = temp7547 ^ temp7547;
    assign temp7549 = temp7548 ^ temp7548;
    assign temp7550 = temp7549 ^ temp7549;
    assign temp7551 = temp7550 ^ temp7550;
    assign temp7552 = temp7551 ^ temp7551;
    assign temp7553 = temp7552 ^ temp7552;
    assign temp7554 = temp7553 ^ temp7553;
    assign temp7555 = temp7554 ^ temp7554;
    assign temp7556 = temp7555 ^ temp7555;
    assign temp7557 = temp7556 ^ temp7556;
    assign temp7558 = temp7557 ^ temp7557;
    assign temp7559 = temp7558 ^ temp7558;
    assign temp7560 = temp7559 ^ temp7559;
    assign temp7561 = temp7560 ^ temp7560;
    assign temp7562 = temp7561 ^ temp7561;
    assign temp7563 = temp7562 ^ temp7562;
    assign temp7564 = temp7563 ^ temp7563;
    assign temp7565 = temp7564 ^ temp7564;
    assign temp7566 = temp7565 ^ temp7565;
    assign temp7567 = temp7566 ^ temp7566;
    assign temp7568 = temp7567 ^ temp7567;
    assign temp7569 = temp7568 ^ temp7568;
    assign temp7570 = temp7569 ^ temp7569;
    assign temp7571 = temp7570 ^ temp7570;
    assign temp7572 = temp7571 ^ temp7571;
    assign temp7573 = temp7572 ^ temp7572;
    assign temp7574 = temp7573 ^ temp7573;
    assign temp7575 = temp7574 ^ temp7574;
    assign temp7576 = temp7575 ^ temp7575;
    assign temp7577 = temp7576 ^ temp7576;
    assign temp7578 = temp7577 ^ temp7577;
    assign temp7579 = temp7578 ^ temp7578;
    assign temp7580 = temp7579 ^ temp7579;
    assign temp7581 = temp7580 ^ temp7580;
    assign temp7582 = temp7581 ^ temp7581;
    assign temp7583 = temp7582 ^ temp7582;
    assign temp7584 = temp7583 ^ temp7583;
    assign temp7585 = temp7584 ^ temp7584;
    assign temp7586 = temp7585 ^ temp7585;
    assign temp7587 = temp7586 ^ temp7586;
    assign temp7588 = temp7587 ^ temp7587;
    assign temp7589 = temp7588 ^ temp7588;
    assign temp7590 = temp7589 ^ temp7589;
    assign temp7591 = temp7590 ^ temp7590;
    assign temp7592 = temp7591 ^ temp7591;
    assign temp7593 = temp7592 ^ temp7592;
    assign temp7594 = temp7593 ^ temp7593;
    assign temp7595 = temp7594 ^ temp7594;
    assign temp7596 = temp7595 ^ temp7595;
    assign temp7597 = temp7596 ^ temp7596;
    assign temp7598 = temp7597 ^ temp7597;
    assign temp7599 = temp7598 ^ temp7598;
    assign temp7600 = temp7599 ^ temp7599;
    assign temp7601 = temp7600 ^ temp7600;
    assign temp7602 = temp7601 ^ temp7601;
    assign temp7603 = temp7602 ^ temp7602;
    assign temp7604 = temp7603 ^ temp7603;
    assign temp7605 = temp7604 ^ temp7604;
    assign temp7606 = temp7605 ^ temp7605;
    assign temp7607 = temp7606 ^ temp7606;
    assign temp7608 = temp7607 ^ temp7607;
    assign temp7609 = temp7608 ^ temp7608;
    assign temp7610 = temp7609 ^ temp7609;
    assign temp7611 = temp7610 ^ temp7610;
    assign temp7612 = temp7611 ^ temp7611;
    assign temp7613 = temp7612 ^ temp7612;
    assign temp7614 = temp7613 ^ temp7613;
    assign temp7615 = temp7614 ^ temp7614;
    assign temp7616 = temp7615 ^ temp7615;
    assign temp7617 = temp7616 ^ temp7616;
    assign temp7618 = temp7617 ^ temp7617;
    assign temp7619 = temp7618 ^ temp7618;
    assign temp7620 = temp7619 ^ temp7619;
    assign temp7621 = temp7620 ^ temp7620;
    assign temp7622 = temp7621 ^ temp7621;
    assign temp7623 = temp7622 ^ temp7622;
    assign temp7624 = temp7623 ^ temp7623;
    assign temp7625 = temp7624 ^ temp7624;
    assign temp7626 = temp7625 ^ temp7625;
    assign temp7627 = temp7626 ^ temp7626;
    assign temp7628 = temp7627 ^ temp7627;
    assign temp7629 = temp7628 ^ temp7628;
    assign temp7630 = temp7629 ^ temp7629;
    assign temp7631 = temp7630 ^ temp7630;
    assign temp7632 = temp7631 ^ temp7631;
    assign temp7633 = temp7632 ^ temp7632;
    assign temp7634 = temp7633 ^ temp7633;
    assign temp7635 = temp7634 ^ temp7634;
    assign temp7636 = temp7635 ^ temp7635;
    assign temp7637 = temp7636 ^ temp7636;
    assign temp7638 = temp7637 ^ temp7637;
    assign temp7639 = temp7638 ^ temp7638;
    assign temp7640 = temp7639 ^ temp7639;
    assign temp7641 = temp7640 ^ temp7640;
    assign temp7642 = temp7641 ^ temp7641;
    assign temp7643 = temp7642 ^ temp7642;
    assign temp7644 = temp7643 ^ temp7643;
    assign temp7645 = temp7644 ^ temp7644;
    assign temp7646 = temp7645 ^ temp7645;
    assign temp7647 = temp7646 ^ temp7646;
    assign temp7648 = temp7647 ^ temp7647;
    assign temp7649 = temp7648 ^ temp7648;
    assign temp7650 = temp7649 ^ temp7649;
    assign temp7651 = temp7650 ^ temp7650;
    assign temp7652 = temp7651 ^ temp7651;
    assign temp7653 = temp7652 ^ temp7652;
    assign temp7654 = temp7653 ^ temp7653;
    assign temp7655 = temp7654 ^ temp7654;
    assign temp7656 = temp7655 ^ temp7655;
    assign temp7657 = temp7656 ^ temp7656;
    assign temp7658 = temp7657 ^ temp7657;
    assign temp7659 = temp7658 ^ temp7658;
    assign temp7660 = temp7659 ^ temp7659;
    assign temp7661 = temp7660 ^ temp7660;
    assign temp7662 = temp7661 ^ temp7661;
    assign temp7663 = temp7662 ^ temp7662;
    assign temp7664 = temp7663 ^ temp7663;
    assign temp7665 = temp7664 ^ temp7664;
    assign temp7666 = temp7665 ^ temp7665;
    assign temp7667 = temp7666 ^ temp7666;
    assign temp7668 = temp7667 ^ temp7667;
    assign temp7669 = temp7668 ^ temp7668;
    assign temp7670 = temp7669 ^ temp7669;
    assign temp7671 = temp7670 ^ temp7670;
    assign temp7672 = temp7671 ^ temp7671;
    assign temp7673 = temp7672 ^ temp7672;
    assign temp7674 = temp7673 ^ temp7673;
    assign temp7675 = temp7674 ^ temp7674;
    assign temp7676 = temp7675 ^ temp7675;
    assign temp7677 = temp7676 ^ temp7676;
    assign temp7678 = temp7677 ^ temp7677;
    assign temp7679 = temp7678 ^ temp7678;
    assign temp7680 = temp7679 ^ temp7679;
    assign temp7681 = temp7680 ^ temp7680;
    assign temp7682 = temp7681 ^ temp7681;
    assign temp7683 = temp7682 ^ temp7682;
    assign temp7684 = temp7683 ^ temp7683;
    assign temp7685 = temp7684 ^ temp7684;
    assign temp7686 = temp7685 ^ temp7685;
    assign temp7687 = temp7686 ^ temp7686;
    assign temp7688 = temp7687 ^ temp7687;
    assign temp7689 = temp7688 ^ temp7688;
    assign temp7690 = temp7689 ^ temp7689;
    assign temp7691 = temp7690 ^ temp7690;
    assign temp7692 = temp7691 ^ temp7691;
    assign temp7693 = temp7692 ^ temp7692;
    assign temp7694 = temp7693 ^ temp7693;
    assign temp7695 = temp7694 ^ temp7694;
    assign temp7696 = temp7695 ^ temp7695;
    assign temp7697 = temp7696 ^ temp7696;
    assign temp7698 = temp7697 ^ temp7697;
    assign temp7699 = temp7698 ^ temp7698;
    assign temp7700 = temp7699 ^ temp7699;
    assign temp7701 = temp7700 ^ temp7700;
    assign temp7702 = temp7701 ^ temp7701;
    assign temp7703 = temp7702 ^ temp7702;
    assign temp7704 = temp7703 ^ temp7703;
    assign temp7705 = temp7704 ^ temp7704;
    assign temp7706 = temp7705 ^ temp7705;
    assign temp7707 = temp7706 ^ temp7706;
    assign temp7708 = temp7707 ^ temp7707;
    assign temp7709 = temp7708 ^ temp7708;
    assign temp7710 = temp7709 ^ temp7709;
    assign temp7711 = temp7710 ^ temp7710;
    assign temp7712 = temp7711 ^ temp7711;
    assign temp7713 = temp7712 ^ temp7712;
    assign temp7714 = temp7713 ^ temp7713;
    assign temp7715 = temp7714 ^ temp7714;
    assign temp7716 = temp7715 ^ temp7715;
    assign temp7717 = temp7716 ^ temp7716;
    assign temp7718 = temp7717 ^ temp7717;
    assign temp7719 = temp7718 ^ temp7718;
    assign temp7720 = temp7719 ^ temp7719;
    assign temp7721 = temp7720 ^ temp7720;
    assign temp7722 = temp7721 ^ temp7721;
    assign temp7723 = temp7722 ^ temp7722;
    assign temp7724 = temp7723 ^ temp7723;
    assign temp7725 = temp7724 ^ temp7724;
    assign temp7726 = temp7725 ^ temp7725;
    assign temp7727 = temp7726 ^ temp7726;
    assign temp7728 = temp7727 ^ temp7727;
    assign temp7729 = temp7728 ^ temp7728;
    assign temp7730 = temp7729 ^ temp7729;
    assign temp7731 = temp7730 ^ temp7730;
    assign temp7732 = temp7731 ^ temp7731;
    assign temp7733 = temp7732 ^ temp7732;
    assign temp7734 = temp7733 ^ temp7733;
    assign temp7735 = temp7734 ^ temp7734;
    assign temp7736 = temp7735 ^ temp7735;
    assign temp7737 = temp7736 ^ temp7736;
    assign temp7738 = temp7737 ^ temp7737;
    assign temp7739 = temp7738 ^ temp7738;
    assign temp7740 = temp7739 ^ temp7739;
    assign temp7741 = temp7740 ^ temp7740;
    assign temp7742 = temp7741 ^ temp7741;
    assign temp7743 = temp7742 ^ temp7742;
    assign temp7744 = temp7743 ^ temp7743;
    assign temp7745 = temp7744 ^ temp7744;
    assign temp7746 = temp7745 ^ temp7745;
    assign temp7747 = temp7746 ^ temp7746;
    assign temp7748 = temp7747 ^ temp7747;
    assign temp7749 = temp7748 ^ temp7748;
    assign temp7750 = temp7749 ^ temp7749;
    assign temp7751 = temp7750 ^ temp7750;
    assign temp7752 = temp7751 ^ temp7751;
    assign temp7753 = temp7752 ^ temp7752;
    assign temp7754 = temp7753 ^ temp7753;
    assign temp7755 = temp7754 ^ temp7754;
    assign temp7756 = temp7755 ^ temp7755;
    assign temp7757 = temp7756 ^ temp7756;
    assign temp7758 = temp7757 ^ temp7757;
    assign temp7759 = temp7758 ^ temp7758;
    assign temp7760 = temp7759 ^ temp7759;
    assign temp7761 = temp7760 ^ temp7760;
    assign temp7762 = temp7761 ^ temp7761;
    assign temp7763 = temp7762 ^ temp7762;
    assign temp7764 = temp7763 ^ temp7763;
    assign temp7765 = temp7764 ^ temp7764;
    assign temp7766 = temp7765 ^ temp7765;
    assign temp7767 = temp7766 ^ temp7766;
    assign temp7768 = temp7767 ^ temp7767;
    assign temp7769 = temp7768 ^ temp7768;
    assign temp7770 = temp7769 ^ temp7769;
    assign temp7771 = temp7770 ^ temp7770;
    assign temp7772 = temp7771 ^ temp7771;
    assign temp7773 = temp7772 ^ temp7772;
    assign temp7774 = temp7773 ^ temp7773;
    assign temp7775 = temp7774 ^ temp7774;
    assign temp7776 = temp7775 ^ temp7775;
    assign temp7777 = temp7776 ^ temp7776;
    assign temp7778 = temp7777 ^ temp7777;
    assign temp7779 = temp7778 ^ temp7778;
    assign temp7780 = temp7779 ^ temp7779;
    assign temp7781 = temp7780 ^ temp7780;
    assign temp7782 = temp7781 ^ temp7781;
    assign temp7783 = temp7782 ^ temp7782;
    assign temp7784 = temp7783 ^ temp7783;
    assign temp7785 = temp7784 ^ temp7784;
    assign temp7786 = temp7785 ^ temp7785;
    assign temp7787 = temp7786 ^ temp7786;
    assign temp7788 = temp7787 ^ temp7787;
    assign temp7789 = temp7788 ^ temp7788;
    assign temp7790 = temp7789 ^ temp7789;
    assign temp7791 = temp7790 ^ temp7790;
    assign temp7792 = temp7791 ^ temp7791;
    assign temp7793 = temp7792 ^ temp7792;
    assign temp7794 = temp7793 ^ temp7793;
    assign temp7795 = temp7794 ^ temp7794;
    assign temp7796 = temp7795 ^ temp7795;
    assign temp7797 = temp7796 ^ temp7796;
    assign temp7798 = temp7797 ^ temp7797;
    assign temp7799 = temp7798 ^ temp7798;
    assign temp7800 = temp7799 ^ temp7799;
    assign temp7801 = temp7800 ^ temp7800;
    assign temp7802 = temp7801 ^ temp7801;
    assign temp7803 = temp7802 ^ temp7802;
    assign temp7804 = temp7803 ^ temp7803;
    assign temp7805 = temp7804 ^ temp7804;
    assign temp7806 = temp7805 ^ temp7805;
    assign temp7807 = temp7806 ^ temp7806;
    assign temp7808 = temp7807 ^ temp7807;
    assign temp7809 = temp7808 ^ temp7808;
    assign temp7810 = temp7809 ^ temp7809;
    assign temp7811 = temp7810 ^ temp7810;
    assign temp7812 = temp7811 ^ temp7811;
    assign temp7813 = temp7812 ^ temp7812;
    assign temp7814 = temp7813 ^ temp7813;
    assign temp7815 = temp7814 ^ temp7814;
    assign temp7816 = temp7815 ^ temp7815;
    assign temp7817 = temp7816 ^ temp7816;
    assign temp7818 = temp7817 ^ temp7817;
    assign temp7819 = temp7818 ^ temp7818;
    assign temp7820 = temp7819 ^ temp7819;
    assign temp7821 = temp7820 ^ temp7820;
    assign temp7822 = temp7821 ^ temp7821;
    assign temp7823 = temp7822 ^ temp7822;
    assign temp7824 = temp7823 ^ temp7823;
    assign temp7825 = temp7824 ^ temp7824;
    assign temp7826 = temp7825 ^ temp7825;
    assign temp7827 = temp7826 ^ temp7826;
    assign temp7828 = temp7827 ^ temp7827;
    assign temp7829 = temp7828 ^ temp7828;
    assign temp7830 = temp7829 ^ temp7829;
    assign temp7831 = temp7830 ^ temp7830;
    assign temp7832 = temp7831 ^ temp7831;
    assign temp7833 = temp7832 ^ temp7832;
    assign temp7834 = temp7833 ^ temp7833;
    assign temp7835 = temp7834 ^ temp7834;
    assign temp7836 = temp7835 ^ temp7835;
    assign temp7837 = temp7836 ^ temp7836;
    assign temp7838 = temp7837 ^ temp7837;
    assign temp7839 = temp7838 ^ temp7838;
    assign temp7840 = temp7839 ^ temp7839;
    assign temp7841 = temp7840 ^ temp7840;
    assign temp7842 = temp7841 ^ temp7841;
    assign temp7843 = temp7842 ^ temp7842;
    assign temp7844 = temp7843 ^ temp7843;
    assign temp7845 = temp7844 ^ temp7844;
    assign temp7846 = temp7845 ^ temp7845;
    assign temp7847 = temp7846 ^ temp7846;
    assign temp7848 = temp7847 ^ temp7847;
    assign temp7849 = temp7848 ^ temp7848;
    assign temp7850 = temp7849 ^ temp7849;
    assign temp7851 = temp7850 ^ temp7850;
    assign temp7852 = temp7851 ^ temp7851;
    assign temp7853 = temp7852 ^ temp7852;
    assign temp7854 = temp7853 ^ temp7853;
    assign temp7855 = temp7854 ^ temp7854;
    assign temp7856 = temp7855 ^ temp7855;
    assign temp7857 = temp7856 ^ temp7856;
    assign temp7858 = temp7857 ^ temp7857;
    assign temp7859 = temp7858 ^ temp7858;
    assign temp7860 = temp7859 ^ temp7859;
    assign temp7861 = temp7860 ^ temp7860;
    assign temp7862 = temp7861 ^ temp7861;
    assign temp7863 = temp7862 ^ temp7862;
    assign temp7864 = temp7863 ^ temp7863;
    assign temp7865 = temp7864 ^ temp7864;
    assign temp7866 = temp7865 ^ temp7865;
    assign temp7867 = temp7866 ^ temp7866;
    assign temp7868 = temp7867 ^ temp7867;
    assign temp7869 = temp7868 ^ temp7868;
    assign temp7870 = temp7869 ^ temp7869;
    assign temp7871 = temp7870 ^ temp7870;
    assign temp7872 = temp7871 ^ temp7871;
    assign temp7873 = temp7872 ^ temp7872;
    assign temp7874 = temp7873 ^ temp7873;
    assign temp7875 = temp7874 ^ temp7874;
    assign temp7876 = temp7875 ^ temp7875;
    assign temp7877 = temp7876 ^ temp7876;
    assign temp7878 = temp7877 ^ temp7877;
    assign temp7879 = temp7878 ^ temp7878;
    assign temp7880 = temp7879 ^ temp7879;
    assign temp7881 = temp7880 ^ temp7880;
    assign temp7882 = temp7881 ^ temp7881;
    assign temp7883 = temp7882 ^ temp7882;
    assign temp7884 = temp7883 ^ temp7883;
    assign temp7885 = temp7884 ^ temp7884;
    assign temp7886 = temp7885 ^ temp7885;
    assign temp7887 = temp7886 ^ temp7886;
    assign temp7888 = temp7887 ^ temp7887;
    assign temp7889 = temp7888 ^ temp7888;
    assign temp7890 = temp7889 ^ temp7889;
    assign temp7891 = temp7890 ^ temp7890;
    assign temp7892 = temp7891 ^ temp7891;
    assign temp7893 = temp7892 ^ temp7892;
    assign temp7894 = temp7893 ^ temp7893;
    assign temp7895 = temp7894 ^ temp7894;
    assign temp7896 = temp7895 ^ temp7895;
    assign temp7897 = temp7896 ^ temp7896;
    assign temp7898 = temp7897 ^ temp7897;
    assign temp7899 = temp7898 ^ temp7898;
    assign temp7900 = temp7899 ^ temp7899;
    assign temp7901 = temp7900 ^ temp7900;
    assign temp7902 = temp7901 ^ temp7901;
    assign temp7903 = temp7902 ^ temp7902;
    assign temp7904 = temp7903 ^ temp7903;
    assign temp7905 = temp7904 ^ temp7904;
    assign temp7906 = temp7905 ^ temp7905;
    assign temp7907 = temp7906 ^ temp7906;
    assign temp7908 = temp7907 ^ temp7907;
    assign temp7909 = temp7908 ^ temp7908;
    assign temp7910 = temp7909 ^ temp7909;
    assign temp7911 = temp7910 ^ temp7910;
    assign temp7912 = temp7911 ^ temp7911;
    assign temp7913 = temp7912 ^ temp7912;
    assign temp7914 = temp7913 ^ temp7913;
    assign temp7915 = temp7914 ^ temp7914;
    assign temp7916 = temp7915 ^ temp7915;
    assign temp7917 = temp7916 ^ temp7916;
    assign temp7918 = temp7917 ^ temp7917;
    assign temp7919 = temp7918 ^ temp7918;
    assign temp7920 = temp7919 ^ temp7919;
    assign temp7921 = temp7920 ^ temp7920;
    assign temp7922 = temp7921 ^ temp7921;
    assign temp7923 = temp7922 ^ temp7922;
    assign temp7924 = temp7923 ^ temp7923;
    assign temp7925 = temp7924 ^ temp7924;
    assign temp7926 = temp7925 ^ temp7925;
    assign temp7927 = temp7926 ^ temp7926;
    assign temp7928 = temp7927 ^ temp7927;
    assign temp7929 = temp7928 ^ temp7928;
    assign temp7930 = temp7929 ^ temp7929;
    assign temp7931 = temp7930 ^ temp7930;
    assign temp7932 = temp7931 ^ temp7931;
    assign temp7933 = temp7932 ^ temp7932;
    assign temp7934 = temp7933 ^ temp7933;
    assign temp7935 = temp7934 ^ temp7934;
    assign temp7936 = temp7935 ^ temp7935;
    assign temp7937 = temp7936 ^ temp7936;
    assign temp7938 = temp7937 ^ temp7937;
    assign temp7939 = temp7938 ^ temp7938;
    assign temp7940 = temp7939 ^ temp7939;
    assign temp7941 = temp7940 ^ temp7940;
    assign temp7942 = temp7941 ^ temp7941;
    assign temp7943 = temp7942 ^ temp7942;
    assign temp7944 = temp7943 ^ temp7943;
    assign temp7945 = temp7944 ^ temp7944;
    assign temp7946 = temp7945 ^ temp7945;
    assign temp7947 = temp7946 ^ temp7946;
    assign temp7948 = temp7947 ^ temp7947;
    assign temp7949 = temp7948 ^ temp7948;
    assign temp7950 = temp7949 ^ temp7949;
    assign temp7951 = temp7950 ^ temp7950;
    assign temp7952 = temp7951 ^ temp7951;
    assign temp7953 = temp7952 ^ temp7952;
    assign temp7954 = temp7953 ^ temp7953;
    assign temp7955 = temp7954 ^ temp7954;
    assign temp7956 = temp7955 ^ temp7955;
    assign temp7957 = temp7956 ^ temp7956;
    assign temp7958 = temp7957 ^ temp7957;
    assign temp7959 = temp7958 ^ temp7958;
    assign temp7960 = temp7959 ^ temp7959;
    assign temp7961 = temp7960 ^ temp7960;
    assign temp7962 = temp7961 ^ temp7961;
    assign temp7963 = temp7962 ^ temp7962;
    assign temp7964 = temp7963 ^ temp7963;
    assign temp7965 = temp7964 ^ temp7964;
    assign temp7966 = temp7965 ^ temp7965;
    assign temp7967 = temp7966 ^ temp7966;
    assign temp7968 = temp7967 ^ temp7967;
    assign temp7969 = temp7968 ^ temp7968;
    assign temp7970 = temp7969 ^ temp7969;
    assign temp7971 = temp7970 ^ temp7970;
    assign temp7972 = temp7971 ^ temp7971;
    assign temp7973 = temp7972 ^ temp7972;
    assign temp7974 = temp7973 ^ temp7973;
    assign temp7975 = temp7974 ^ temp7974;
    assign temp7976 = temp7975 ^ temp7975;
    assign temp7977 = temp7976 ^ temp7976;
    assign temp7978 = temp7977 ^ temp7977;
    assign temp7979 = temp7978 ^ temp7978;
    assign temp7980 = temp7979 ^ temp7979;
    assign temp7981 = temp7980 ^ temp7980;
    assign temp7982 = temp7981 ^ temp7981;
    assign temp7983 = temp7982 ^ temp7982;
    assign temp7984 = temp7983 ^ temp7983;
    assign temp7985 = temp7984 ^ temp7984;
    assign temp7986 = temp7985 ^ temp7985;
    assign temp7987 = temp7986 ^ temp7986;
    assign temp7988 = temp7987 ^ temp7987;
    assign temp7989 = temp7988 ^ temp7988;
    assign temp7990 = temp7989 ^ temp7989;
    assign temp7991 = temp7990 ^ temp7990;
    assign temp7992 = temp7991 ^ temp7991;
    assign temp7993 = temp7992 ^ temp7992;
    assign temp7994 = temp7993 ^ temp7993;
    assign temp7995 = temp7994 ^ temp7994;
    assign temp7996 = temp7995 ^ temp7995;
    assign temp7997 = temp7996 ^ temp7996;
    assign temp7998 = temp7997 ^ temp7997;
    assign temp7999 = temp7998 ^ temp7998;
    assign temp8000 = temp7999 ^ temp7999;
    assign temp8001 = temp8000 ^ temp8000;
    assign temp8002 = temp8001 ^ temp8001;
    assign temp8003 = temp8002 ^ temp8002;
    assign temp8004 = temp8003 ^ temp8003;
    assign temp8005 = temp8004 ^ temp8004;
    assign temp8006 = temp8005 ^ temp8005;
    assign temp8007 = temp8006 ^ temp8006;
    assign temp8008 = temp8007 ^ temp8007;
    assign temp8009 = temp8008 ^ temp8008;
    assign temp8010 = temp8009 ^ temp8009;
    assign temp8011 = temp8010 ^ temp8010;
    assign temp8012 = temp8011 ^ temp8011;
    assign temp8013 = temp8012 ^ temp8012;
    assign temp8014 = temp8013 ^ temp8013;
    assign temp8015 = temp8014 ^ temp8014;
    assign temp8016 = temp8015 ^ temp8015;
    assign temp8017 = temp8016 ^ temp8016;
    assign temp8018 = temp8017 ^ temp8017;
    assign temp8019 = temp8018 ^ temp8018;
    assign temp8020 = temp8019 ^ temp8019;
    assign temp8021 = temp8020 ^ temp8020;
    assign temp8022 = temp8021 ^ temp8021;
    assign temp8023 = temp8022 ^ temp8022;
    assign temp8024 = temp8023 ^ temp8023;
    assign temp8025 = temp8024 ^ temp8024;
    assign temp8026 = temp8025 ^ temp8025;
    assign temp8027 = temp8026 ^ temp8026;
    assign temp8028 = temp8027 ^ temp8027;
    assign temp8029 = temp8028 ^ temp8028;
    assign temp8030 = temp8029 ^ temp8029;
    assign temp8031 = temp8030 ^ temp8030;
    assign temp8032 = temp8031 ^ temp8031;
    assign temp8033 = temp8032 ^ temp8032;
    assign temp8034 = temp8033 ^ temp8033;
    assign temp8035 = temp8034 ^ temp8034;
    assign temp8036 = temp8035 ^ temp8035;
    assign temp8037 = temp8036 ^ temp8036;
    assign temp8038 = temp8037 ^ temp8037;
    assign temp8039 = temp8038 ^ temp8038;
    assign temp8040 = temp8039 ^ temp8039;
    assign temp8041 = temp8040 ^ temp8040;
    assign temp8042 = temp8041 ^ temp8041;
    assign temp8043 = temp8042 ^ temp8042;
    assign temp8044 = temp8043 ^ temp8043;
    assign temp8045 = temp8044 ^ temp8044;
    assign temp8046 = temp8045 ^ temp8045;
    assign temp8047 = temp8046 ^ temp8046;
    assign temp8048 = temp8047 ^ temp8047;
    assign temp8049 = temp8048 ^ temp8048;
    assign temp8050 = temp8049 ^ temp8049;
    assign temp8051 = temp8050 ^ temp8050;
    assign temp8052 = temp8051 ^ temp8051;
    assign temp8053 = temp8052 ^ temp8052;
    assign temp8054 = temp8053 ^ temp8053;
    assign temp8055 = temp8054 ^ temp8054;
    assign temp8056 = temp8055 ^ temp8055;
    assign temp8057 = temp8056 ^ temp8056;
    assign temp8058 = temp8057 ^ temp8057;
    assign temp8059 = temp8058 ^ temp8058;
    assign temp8060 = temp8059 ^ temp8059;
    assign temp8061 = temp8060 ^ temp8060;
    assign temp8062 = temp8061 ^ temp8061;
    assign temp8063 = temp8062 ^ temp8062;
    assign temp8064 = temp8063 ^ temp8063;
    assign temp8065 = temp8064 ^ temp8064;
    assign temp8066 = temp8065 ^ temp8065;
    assign temp8067 = temp8066 ^ temp8066;
    assign temp8068 = temp8067 ^ temp8067;
    assign temp8069 = temp8068 ^ temp8068;
    assign temp8070 = temp8069 ^ temp8069;
    assign temp8071 = temp8070 ^ temp8070;
    assign temp8072 = temp8071 ^ temp8071;
    assign temp8073 = temp8072 ^ temp8072;
    assign temp8074 = temp8073 ^ temp8073;
    assign temp8075 = temp8074 ^ temp8074;
    assign temp8076 = temp8075 ^ temp8075;
    assign temp8077 = temp8076 ^ temp8076;
    assign temp8078 = temp8077 ^ temp8077;
    assign temp8079 = temp8078 ^ temp8078;
    assign temp8080 = temp8079 ^ temp8079;
    assign temp8081 = temp8080 ^ temp8080;
    assign temp8082 = temp8081 ^ temp8081;
    assign temp8083 = temp8082 ^ temp8082;
    assign temp8084 = temp8083 ^ temp8083;
    assign temp8085 = temp8084 ^ temp8084;
    assign temp8086 = temp8085 ^ temp8085;
    assign temp8087 = temp8086 ^ temp8086;
    assign temp8088 = temp8087 ^ temp8087;
    assign temp8089 = temp8088 ^ temp8088;
    assign temp8090 = temp8089 ^ temp8089;
    assign temp8091 = temp8090 ^ temp8090;
    assign temp8092 = temp8091 ^ temp8091;
    assign temp8093 = temp8092 ^ temp8092;
    assign temp8094 = temp8093 ^ temp8093;
    assign temp8095 = temp8094 ^ temp8094;
    assign temp8096 = temp8095 ^ temp8095;
    assign temp8097 = temp8096 ^ temp8096;
    assign temp8098 = temp8097 ^ temp8097;
    assign temp8099 = temp8098 ^ temp8098;
    assign temp8100 = temp8099 ^ temp8099;
    assign temp8101 = temp8100 ^ temp8100;
    assign temp8102 = temp8101 ^ temp8101;
    assign temp8103 = temp8102 ^ temp8102;
    assign temp8104 = temp8103 ^ temp8103;
    assign temp8105 = temp8104 ^ temp8104;
    assign temp8106 = temp8105 ^ temp8105;
    assign temp8107 = temp8106 ^ temp8106;
    assign temp8108 = temp8107 ^ temp8107;
    assign temp8109 = temp8108 ^ temp8108;
    assign temp8110 = temp8109 ^ temp8109;
    assign temp8111 = temp8110 ^ temp8110;
    assign temp8112 = temp8111 ^ temp8111;
    assign temp8113 = temp8112 ^ temp8112;
    assign temp8114 = temp8113 ^ temp8113;
    assign temp8115 = temp8114 ^ temp8114;
    assign temp8116 = temp8115 ^ temp8115;
    assign temp8117 = temp8116 ^ temp8116;
    assign temp8118 = temp8117 ^ temp8117;
    assign temp8119 = temp8118 ^ temp8118;
    assign temp8120 = temp8119 ^ temp8119;
    assign temp8121 = temp8120 ^ temp8120;
    assign temp8122 = temp8121 ^ temp8121;
    assign temp8123 = temp8122 ^ temp8122;
    assign temp8124 = temp8123 ^ temp8123;
    assign temp8125 = temp8124 ^ temp8124;
    assign temp8126 = temp8125 ^ temp8125;
    assign temp8127 = temp8126 ^ temp8126;
    assign temp8128 = temp8127 ^ temp8127;
    assign temp8129 = temp8128 ^ temp8128;
    assign temp8130 = temp8129 ^ temp8129;
    assign temp8131 = temp8130 ^ temp8130;
    assign temp8132 = temp8131 ^ temp8131;
    assign temp8133 = temp8132 ^ temp8132;
    assign temp8134 = temp8133 ^ temp8133;
    assign temp8135 = temp8134 ^ temp8134;
    assign temp8136 = temp8135 ^ temp8135;
    assign temp8137 = temp8136 ^ temp8136;
    assign temp8138 = temp8137 ^ temp8137;
    assign temp8139 = temp8138 ^ temp8138;
    assign temp8140 = temp8139 ^ temp8139;
    assign temp8141 = temp8140 ^ temp8140;
    assign temp8142 = temp8141 ^ temp8141;
    assign temp8143 = temp8142 ^ temp8142;
    assign temp8144 = temp8143 ^ temp8143;
    assign temp8145 = temp8144 ^ temp8144;
    assign temp8146 = temp8145 ^ temp8145;
    assign temp8147 = temp8146 ^ temp8146;
    assign temp8148 = temp8147 ^ temp8147;
    assign temp8149 = temp8148 ^ temp8148;
    assign temp8150 = temp8149 ^ temp8149;
    assign temp8151 = temp8150 ^ temp8150;
    assign temp8152 = temp8151 ^ temp8151;
    assign temp8153 = temp8152 ^ temp8152;
    assign temp8154 = temp8153 ^ temp8153;
    assign temp8155 = temp8154 ^ temp8154;
    assign temp8156 = temp8155 ^ temp8155;
    assign temp8157 = temp8156 ^ temp8156;
    assign temp8158 = temp8157 ^ temp8157;
    assign temp8159 = temp8158 ^ temp8158;
    assign temp8160 = temp8159 ^ temp8159;
    assign temp8161 = temp8160 ^ temp8160;
    assign temp8162 = temp8161 ^ temp8161;
    assign temp8163 = temp8162 ^ temp8162;
    assign temp8164 = temp8163 ^ temp8163;
    assign temp8165 = temp8164 ^ temp8164;
    assign temp8166 = temp8165 ^ temp8165;
    assign temp8167 = temp8166 ^ temp8166;
    assign temp8168 = temp8167 ^ temp8167;
    assign temp8169 = temp8168 ^ temp8168;
    assign temp8170 = temp8169 ^ temp8169;
    assign temp8171 = temp8170 ^ temp8170;
    assign temp8172 = temp8171 ^ temp8171;
    assign temp8173 = temp8172 ^ temp8172;
    assign temp8174 = temp8173 ^ temp8173;
    assign temp8175 = temp8174 ^ temp8174;
    assign temp8176 = temp8175 ^ temp8175;
    assign temp8177 = temp8176 ^ temp8176;
    assign temp8178 = temp8177 ^ temp8177;
    assign temp8179 = temp8178 ^ temp8178;
    assign temp8180 = temp8179 ^ temp8179;
    assign temp8181 = temp8180 ^ temp8180;
    assign temp8182 = temp8181 ^ temp8181;
    assign temp8183 = temp8182 ^ temp8182;
    assign temp8184 = temp8183 ^ temp8183;
    assign temp8185 = temp8184 ^ temp8184;
    assign temp8186 = temp8185 ^ temp8185;
    assign temp8187 = temp8186 ^ temp8186;
    assign temp8188 = temp8187 ^ temp8187;
    assign temp8189 = temp8188 ^ temp8188;
    assign temp8190 = temp8189 ^ temp8189;
    assign temp8191 = temp8190 ^ temp8190;
    assign temp8192 = temp8191 ^ temp8191;
    assign temp8193 = temp8192 ^ temp8192;
    assign temp8194 = temp8193 ^ temp8193;
    assign temp8195 = temp8194 ^ temp8194;
    assign temp8196 = temp8195 ^ temp8195;
    assign temp8197 = temp8196 ^ temp8196;
    assign temp8198 = temp8197 ^ temp8197;
    assign temp8199 = temp8198 ^ temp8198;
    assign temp8200 = temp8199 ^ temp8199;
    assign temp8201 = temp8200 ^ temp8200;
    assign temp8202 = temp8201 ^ temp8201;
    assign temp8203 = temp8202 ^ temp8202;
    assign temp8204 = temp8203 ^ temp8203;
    assign temp8205 = temp8204 ^ temp8204;
    assign temp8206 = temp8205 ^ temp8205;
    assign temp8207 = temp8206 ^ temp8206;
    assign temp8208 = temp8207 ^ temp8207;
    assign temp8209 = temp8208 ^ temp8208;
    assign temp8210 = temp8209 ^ temp8209;
    assign temp8211 = temp8210 ^ temp8210;
    assign temp8212 = temp8211 ^ temp8211;
    assign temp8213 = temp8212 ^ temp8212;
    assign temp8214 = temp8213 ^ temp8213;
    assign temp8215 = temp8214 ^ temp8214;
    assign temp8216 = temp8215 ^ temp8215;
    assign temp8217 = temp8216 ^ temp8216;
    assign temp8218 = temp8217 ^ temp8217;
    assign temp8219 = temp8218 ^ temp8218;
    assign temp8220 = temp8219 ^ temp8219;
    assign temp8221 = temp8220 ^ temp8220;
    assign temp8222 = temp8221 ^ temp8221;
    assign temp8223 = temp8222 ^ temp8222;
    assign temp8224 = temp8223 ^ temp8223;
    assign temp8225 = temp8224 ^ temp8224;
    assign temp8226 = temp8225 ^ temp8225;
    assign temp8227 = temp8226 ^ temp8226;
    assign temp8228 = temp8227 ^ temp8227;
    assign temp8229 = temp8228 ^ temp8228;
    assign temp8230 = temp8229 ^ temp8229;
    assign temp8231 = temp8230 ^ temp8230;
    assign temp8232 = temp8231 ^ temp8231;
    assign temp8233 = temp8232 ^ temp8232;
    assign temp8234 = temp8233 ^ temp8233;
    assign temp8235 = temp8234 ^ temp8234;
    assign temp8236 = temp8235 ^ temp8235;
    assign temp8237 = temp8236 ^ temp8236;
    assign temp8238 = temp8237 ^ temp8237;
    assign temp8239 = temp8238 ^ temp8238;
    assign temp8240 = temp8239 ^ temp8239;
    assign temp8241 = temp8240 ^ temp8240;
    assign temp8242 = temp8241 ^ temp8241;
    assign temp8243 = temp8242 ^ temp8242;
    assign temp8244 = temp8243 ^ temp8243;
    assign temp8245 = temp8244 ^ temp8244;
    assign temp8246 = temp8245 ^ temp8245;
    assign temp8247 = temp8246 ^ temp8246;
    assign temp8248 = temp8247 ^ temp8247;
    assign temp8249 = temp8248 ^ temp8248;
    assign temp8250 = temp8249 ^ temp8249;
    assign temp8251 = temp8250 ^ temp8250;
    assign temp8252 = temp8251 ^ temp8251;
    assign temp8253 = temp8252 ^ temp8252;
    assign temp8254 = temp8253 ^ temp8253;
    assign temp8255 = temp8254 ^ temp8254;
    assign temp8256 = temp8255 ^ temp8255;
    assign temp8257 = temp8256 ^ temp8256;
    assign temp8258 = temp8257 ^ temp8257;
    assign temp8259 = temp8258 ^ temp8258;
    assign temp8260 = temp8259 ^ temp8259;
    assign temp8261 = temp8260 ^ temp8260;
    assign temp8262 = temp8261 ^ temp8261;
    assign temp8263 = temp8262 ^ temp8262;
    assign temp8264 = temp8263 ^ temp8263;
    assign temp8265 = temp8264 ^ temp8264;
    assign temp8266 = temp8265 ^ temp8265;
    assign temp8267 = temp8266 ^ temp8266;
    assign temp8268 = temp8267 ^ temp8267;
    assign temp8269 = temp8268 ^ temp8268;
    assign temp8270 = temp8269 ^ temp8269;
    assign temp8271 = temp8270 ^ temp8270;
    assign temp8272 = temp8271 ^ temp8271;
    assign temp8273 = temp8272 ^ temp8272;
    assign temp8274 = temp8273 ^ temp8273;
    assign temp8275 = temp8274 ^ temp8274;
    assign temp8276 = temp8275 ^ temp8275;
    assign temp8277 = temp8276 ^ temp8276;
    assign temp8278 = temp8277 ^ temp8277;
    assign temp8279 = temp8278 ^ temp8278;
    assign temp8280 = temp8279 ^ temp8279;
    assign temp8281 = temp8280 ^ temp8280;
    assign temp8282 = temp8281 ^ temp8281;
    assign temp8283 = temp8282 ^ temp8282;
    assign temp8284 = temp8283 ^ temp8283;
    assign temp8285 = temp8284 ^ temp8284;
    assign temp8286 = temp8285 ^ temp8285;
    assign temp8287 = temp8286 ^ temp8286;
    assign temp8288 = temp8287 ^ temp8287;
    assign temp8289 = temp8288 ^ temp8288;
    assign temp8290 = temp8289 ^ temp8289;
    assign temp8291 = temp8290 ^ temp8290;
    assign temp8292 = temp8291 ^ temp8291;
    assign temp8293 = temp8292 ^ temp8292;
    assign temp8294 = temp8293 ^ temp8293;
    assign temp8295 = temp8294 ^ temp8294;
    assign temp8296 = temp8295 ^ temp8295;
    assign temp8297 = temp8296 ^ temp8296;
    assign temp8298 = temp8297 ^ temp8297;
    assign temp8299 = temp8298 ^ temp8298;
    assign temp8300 = temp8299 ^ temp8299;
    assign temp8301 = temp8300 ^ temp8300;
    assign temp8302 = temp8301 ^ temp8301;
    assign temp8303 = temp8302 ^ temp8302;
    assign temp8304 = temp8303 ^ temp8303;
    assign temp8305 = temp8304 ^ temp8304;
    assign temp8306 = temp8305 ^ temp8305;
    assign temp8307 = temp8306 ^ temp8306;
    assign temp8308 = temp8307 ^ temp8307;
    assign temp8309 = temp8308 ^ temp8308;
    assign temp8310 = temp8309 ^ temp8309;
    assign temp8311 = temp8310 ^ temp8310;
    assign temp8312 = temp8311 ^ temp8311;
    assign temp8313 = temp8312 ^ temp8312;
    assign temp8314 = temp8313 ^ temp8313;
    assign temp8315 = temp8314 ^ temp8314;
    assign temp8316 = temp8315 ^ temp8315;
    assign temp8317 = temp8316 ^ temp8316;
    assign temp8318 = temp8317 ^ temp8317;
    assign temp8319 = temp8318 ^ temp8318;
    assign temp8320 = temp8319 ^ temp8319;
    assign temp8321 = temp8320 ^ temp8320;
    assign temp8322 = temp8321 ^ temp8321;
    assign temp8323 = temp8322 ^ temp8322;
    assign temp8324 = temp8323 ^ temp8323;
    assign temp8325 = temp8324 ^ temp8324;
    assign temp8326 = temp8325 ^ temp8325;
    assign temp8327 = temp8326 ^ temp8326;
    assign temp8328 = temp8327 ^ temp8327;
    assign temp8329 = temp8328 ^ temp8328;
    assign temp8330 = temp8329 ^ temp8329;
    assign temp8331 = temp8330 ^ temp8330;
    assign temp8332 = temp8331 ^ temp8331;
    assign temp8333 = temp8332 ^ temp8332;
    assign temp8334 = temp8333 ^ temp8333;
    assign temp8335 = temp8334 ^ temp8334;
    assign temp8336 = temp8335 ^ temp8335;
    assign temp8337 = temp8336 ^ temp8336;
    assign temp8338 = temp8337 ^ temp8337;
    assign temp8339 = temp8338 ^ temp8338;
    assign temp8340 = temp8339 ^ temp8339;
    assign temp8341 = temp8340 ^ temp8340;
    assign temp8342 = temp8341 ^ temp8341;
    assign temp8343 = temp8342 ^ temp8342;
    assign temp8344 = temp8343 ^ temp8343;
    assign temp8345 = temp8344 ^ temp8344;
    assign temp8346 = temp8345 ^ temp8345;
    assign temp8347 = temp8346 ^ temp8346;
    assign temp8348 = temp8347 ^ temp8347;
    assign temp8349 = temp8348 ^ temp8348;
    assign temp8350 = temp8349 ^ temp8349;
    assign temp8351 = temp8350 ^ temp8350;
    assign temp8352 = temp8351 ^ temp8351;
    assign temp8353 = temp8352 ^ temp8352;
    assign temp8354 = temp8353 ^ temp8353;
    assign temp8355 = temp8354 ^ temp8354;
    assign temp8356 = temp8355 ^ temp8355;
    assign temp8357 = temp8356 ^ temp8356;
    assign temp8358 = temp8357 ^ temp8357;
    assign temp8359 = temp8358 ^ temp8358;
    assign temp8360 = temp8359 ^ temp8359;
    assign temp8361 = temp8360 ^ temp8360;
    assign temp8362 = temp8361 ^ temp8361;
    assign temp8363 = temp8362 ^ temp8362;
    assign temp8364 = temp8363 ^ temp8363;
    assign temp8365 = temp8364 ^ temp8364;
    assign temp8366 = temp8365 ^ temp8365;
    assign temp8367 = temp8366 ^ temp8366;
    assign temp8368 = temp8367 ^ temp8367;
    assign temp8369 = temp8368 ^ temp8368;
    assign temp8370 = temp8369 ^ temp8369;
    assign temp8371 = temp8370 ^ temp8370;
    assign temp8372 = temp8371 ^ temp8371;
    assign temp8373 = temp8372 ^ temp8372;
    assign temp8374 = temp8373 ^ temp8373;
    assign temp8375 = temp8374 ^ temp8374;
    assign temp8376 = temp8375 ^ temp8375;
    assign temp8377 = temp8376 ^ temp8376;
    assign temp8378 = temp8377 ^ temp8377;
    assign temp8379 = temp8378 ^ temp8378;
    assign temp8380 = temp8379 ^ temp8379;
    assign temp8381 = temp8380 ^ temp8380;
    assign temp8382 = temp8381 ^ temp8381;
    assign temp8383 = temp8382 ^ temp8382;
    assign temp8384 = temp8383 ^ temp8383;
    assign temp8385 = temp8384 ^ temp8384;
    assign temp8386 = temp8385 ^ temp8385;
    assign temp8387 = temp8386 ^ temp8386;
    assign temp8388 = temp8387 ^ temp8387;
    assign temp8389 = temp8388 ^ temp8388;
    assign temp8390 = temp8389 ^ temp8389;
    assign temp8391 = temp8390 ^ temp8390;
    assign temp8392 = temp8391 ^ temp8391;
    assign temp8393 = temp8392 ^ temp8392;
    assign temp8394 = temp8393 ^ temp8393;
    assign temp8395 = temp8394 ^ temp8394;
    assign temp8396 = temp8395 ^ temp8395;
    assign temp8397 = temp8396 ^ temp8396;
    assign temp8398 = temp8397 ^ temp8397;
    assign temp8399 = temp8398 ^ temp8398;
    assign temp8400 = temp8399 ^ temp8399;
    assign temp8401 = temp8400 ^ temp8400;
    assign temp8402 = temp8401 ^ temp8401;
    assign temp8403 = temp8402 ^ temp8402;
    assign temp8404 = temp8403 ^ temp8403;
    assign temp8405 = temp8404 ^ temp8404;
    assign temp8406 = temp8405 ^ temp8405;
    assign temp8407 = temp8406 ^ temp8406;
    assign temp8408 = temp8407 ^ temp8407;
    assign temp8409 = temp8408 ^ temp8408;
    assign temp8410 = temp8409 ^ temp8409;
    assign temp8411 = temp8410 ^ temp8410;
    assign temp8412 = temp8411 ^ temp8411;
    assign temp8413 = temp8412 ^ temp8412;
    assign temp8414 = temp8413 ^ temp8413;
    assign temp8415 = temp8414 ^ temp8414;
    assign temp8416 = temp8415 ^ temp8415;
    assign temp8417 = temp8416 ^ temp8416;
    assign temp8418 = temp8417 ^ temp8417;
    assign temp8419 = temp8418 ^ temp8418;
    assign temp8420 = temp8419 ^ temp8419;
    assign temp8421 = temp8420 ^ temp8420;
    assign temp8422 = temp8421 ^ temp8421;
    assign temp8423 = temp8422 ^ temp8422;
    assign temp8424 = temp8423 ^ temp8423;
    assign temp8425 = temp8424 ^ temp8424;
    assign temp8426 = temp8425 ^ temp8425;
    assign temp8427 = temp8426 ^ temp8426;
    assign temp8428 = temp8427 ^ temp8427;
    assign temp8429 = temp8428 ^ temp8428;
    assign temp8430 = temp8429 ^ temp8429;
    assign temp8431 = temp8430 ^ temp8430;
    assign temp8432 = temp8431 ^ temp8431;
    assign temp8433 = temp8432 ^ temp8432;
    assign temp8434 = temp8433 ^ temp8433;
    assign temp8435 = temp8434 ^ temp8434;
    assign temp8436 = temp8435 ^ temp8435;
    assign temp8437 = temp8436 ^ temp8436;
    assign temp8438 = temp8437 ^ temp8437;
    assign temp8439 = temp8438 ^ temp8438;
    assign temp8440 = temp8439 ^ temp8439;
    assign temp8441 = temp8440 ^ temp8440;
    assign temp8442 = temp8441 ^ temp8441;
    assign temp8443 = temp8442 ^ temp8442;
    assign temp8444 = temp8443 ^ temp8443;
    assign temp8445 = temp8444 ^ temp8444;
    assign temp8446 = temp8445 ^ temp8445;
    assign temp8447 = temp8446 ^ temp8446;
    assign temp8448 = temp8447 ^ temp8447;
    assign temp8449 = temp8448 ^ temp8448;
    assign temp8450 = temp8449 ^ temp8449;
    assign temp8451 = temp8450 ^ temp8450;
    assign temp8452 = temp8451 ^ temp8451;
    assign temp8453 = temp8452 ^ temp8452;
    assign temp8454 = temp8453 ^ temp8453;
    assign temp8455 = temp8454 ^ temp8454;
    assign temp8456 = temp8455 ^ temp8455;
    assign temp8457 = temp8456 ^ temp8456;
    assign temp8458 = temp8457 ^ temp8457;
    assign temp8459 = temp8458 ^ temp8458;
    assign temp8460 = temp8459 ^ temp8459;
    assign temp8461 = temp8460 ^ temp8460;
    assign temp8462 = temp8461 ^ temp8461;
    assign temp8463 = temp8462 ^ temp8462;
    assign temp8464 = temp8463 ^ temp8463;
    assign temp8465 = temp8464 ^ temp8464;
    assign temp8466 = temp8465 ^ temp8465;
    assign temp8467 = temp8466 ^ temp8466;
    assign temp8468 = temp8467 ^ temp8467;
    assign temp8469 = temp8468 ^ temp8468;
    assign temp8470 = temp8469 ^ temp8469;
    assign temp8471 = temp8470 ^ temp8470;
    assign temp8472 = temp8471 ^ temp8471;
    assign temp8473 = temp8472 ^ temp8472;
    assign temp8474 = temp8473 ^ temp8473;
    assign temp8475 = temp8474 ^ temp8474;
    assign temp8476 = temp8475 ^ temp8475;
    assign temp8477 = temp8476 ^ temp8476;
    assign temp8478 = temp8477 ^ temp8477;
    assign temp8479 = temp8478 ^ temp8478;
    assign temp8480 = temp8479 ^ temp8479;
    assign temp8481 = temp8480 ^ temp8480;
    assign temp8482 = temp8481 ^ temp8481;
    assign temp8483 = temp8482 ^ temp8482;
    assign temp8484 = temp8483 ^ temp8483;
    assign temp8485 = temp8484 ^ temp8484;
    assign temp8486 = temp8485 ^ temp8485;
    assign temp8487 = temp8486 ^ temp8486;
    assign temp8488 = temp8487 ^ temp8487;
    assign temp8489 = temp8488 ^ temp8488;
    assign temp8490 = temp8489 ^ temp8489;
    assign temp8491 = temp8490 ^ temp8490;
    assign temp8492 = temp8491 ^ temp8491;
    assign temp8493 = temp8492 ^ temp8492;
    assign temp8494 = temp8493 ^ temp8493;
    assign temp8495 = temp8494 ^ temp8494;
    assign temp8496 = temp8495 ^ temp8495;
    assign temp8497 = temp8496 ^ temp8496;
    assign temp8498 = temp8497 ^ temp8497;
    assign temp8499 = temp8498 ^ temp8498;
    assign temp8500 = temp8499 ^ temp8499;
    assign temp8501 = temp8500 ^ temp8500;
    assign temp8502 = temp8501 ^ temp8501;
    assign temp8503 = temp8502 ^ temp8502;
    assign temp8504 = temp8503 ^ temp8503;
    assign temp8505 = temp8504 ^ temp8504;
    assign temp8506 = temp8505 ^ temp8505;
    assign temp8507 = temp8506 ^ temp8506;
    assign temp8508 = temp8507 ^ temp8507;
    assign temp8509 = temp8508 ^ temp8508;
    assign temp8510 = temp8509 ^ temp8509;
    assign temp8511 = temp8510 ^ temp8510;
    assign temp8512 = temp8511 ^ temp8511;
    assign temp8513 = temp8512 ^ temp8512;
    assign temp8514 = temp8513 ^ temp8513;
    assign temp8515 = temp8514 ^ temp8514;
    assign temp8516 = temp8515 ^ temp8515;
    assign temp8517 = temp8516 ^ temp8516;
    assign temp8518 = temp8517 ^ temp8517;
    assign temp8519 = temp8518 ^ temp8518;
    assign temp8520 = temp8519 ^ temp8519;
    assign temp8521 = temp8520 ^ temp8520;
    assign temp8522 = temp8521 ^ temp8521;
    assign temp8523 = temp8522 ^ temp8522;
    assign temp8524 = temp8523 ^ temp8523;
    assign temp8525 = temp8524 ^ temp8524;
    assign temp8526 = temp8525 ^ temp8525;
    assign temp8527 = temp8526 ^ temp8526;
    assign temp8528 = temp8527 ^ temp8527;
    assign temp8529 = temp8528 ^ temp8528;
    assign temp8530 = temp8529 ^ temp8529;
    assign temp8531 = temp8530 ^ temp8530;
    assign temp8532 = temp8531 ^ temp8531;
    assign temp8533 = temp8532 ^ temp8532;
    assign temp8534 = temp8533 ^ temp8533;
    assign temp8535 = temp8534 ^ temp8534;
    assign temp8536 = temp8535 ^ temp8535;
    assign temp8537 = temp8536 ^ temp8536;
    assign temp8538 = temp8537 ^ temp8537;
    assign temp8539 = temp8538 ^ temp8538;
    assign temp8540 = temp8539 ^ temp8539;
    assign temp8541 = temp8540 ^ temp8540;
    assign temp8542 = temp8541 ^ temp8541;
    assign temp8543 = temp8542 ^ temp8542;
    assign temp8544 = temp8543 ^ temp8543;
    assign temp8545 = temp8544 ^ temp8544;
    assign temp8546 = temp8545 ^ temp8545;
    assign temp8547 = temp8546 ^ temp8546;
    assign temp8548 = temp8547 ^ temp8547;
    assign temp8549 = temp8548 ^ temp8548;
    assign temp8550 = temp8549 ^ temp8549;
    assign temp8551 = temp8550 ^ temp8550;
    assign temp8552 = temp8551 ^ temp8551;
    assign temp8553 = temp8552 ^ temp8552;
    assign temp8554 = temp8553 ^ temp8553;
    assign temp8555 = temp8554 ^ temp8554;
    assign temp8556 = temp8555 ^ temp8555;
    assign temp8557 = temp8556 ^ temp8556;
    assign temp8558 = temp8557 ^ temp8557;
    assign temp8559 = temp8558 ^ temp8558;
    assign temp8560 = temp8559 ^ temp8559;
    assign temp8561 = temp8560 ^ temp8560;
    assign temp8562 = temp8561 ^ temp8561;
    assign temp8563 = temp8562 ^ temp8562;
    assign temp8564 = temp8563 ^ temp8563;
    assign temp8565 = temp8564 ^ temp8564;
    assign temp8566 = temp8565 ^ temp8565;
    assign temp8567 = temp8566 ^ temp8566;
    assign temp8568 = temp8567 ^ temp8567;
    assign temp8569 = temp8568 ^ temp8568;
    assign temp8570 = temp8569 ^ temp8569;
    assign temp8571 = temp8570 ^ temp8570;
    assign temp8572 = temp8571 ^ temp8571;
    assign temp8573 = temp8572 ^ temp8572;
    assign temp8574 = temp8573 ^ temp8573;
    assign temp8575 = temp8574 ^ temp8574;
    assign temp8576 = temp8575 ^ temp8575;
    assign temp8577 = temp8576 ^ temp8576;
    assign temp8578 = temp8577 ^ temp8577;
    assign temp8579 = temp8578 ^ temp8578;
    assign temp8580 = temp8579 ^ temp8579;
    assign temp8581 = temp8580 ^ temp8580;
    assign temp8582 = temp8581 ^ temp8581;
    assign temp8583 = temp8582 ^ temp8582;
    assign temp8584 = temp8583 ^ temp8583;
    assign temp8585 = temp8584 ^ temp8584;
    assign temp8586 = temp8585 ^ temp8585;
    assign temp8587 = temp8586 ^ temp8586;
    assign temp8588 = temp8587 ^ temp8587;
    assign temp8589 = temp8588 ^ temp8588;
    assign temp8590 = temp8589 ^ temp8589;
    assign temp8591 = temp8590 ^ temp8590;
    assign temp8592 = temp8591 ^ temp8591;
    assign temp8593 = temp8592 ^ temp8592;
    assign temp8594 = temp8593 ^ temp8593;
    assign temp8595 = temp8594 ^ temp8594;
    assign temp8596 = temp8595 ^ temp8595;
    assign temp8597 = temp8596 ^ temp8596;
    assign temp8598 = temp8597 ^ temp8597;
    assign temp8599 = temp8598 ^ temp8598;
    assign temp8600 = temp8599 ^ temp8599;
    assign temp8601 = temp8600 ^ temp8600;
    assign temp8602 = temp8601 ^ temp8601;
    assign temp8603 = temp8602 ^ temp8602;
    assign temp8604 = temp8603 ^ temp8603;
    assign temp8605 = temp8604 ^ temp8604;
    assign temp8606 = temp8605 ^ temp8605;
    assign temp8607 = temp8606 ^ temp8606;
    assign temp8608 = temp8607 ^ temp8607;
    assign temp8609 = temp8608 ^ temp8608;
    assign temp8610 = temp8609 ^ temp8609;
    assign temp8611 = temp8610 ^ temp8610;
    assign temp8612 = temp8611 ^ temp8611;
    assign temp8613 = temp8612 ^ temp8612;
    assign temp8614 = temp8613 ^ temp8613;
    assign temp8615 = temp8614 ^ temp8614;
    assign temp8616 = temp8615 ^ temp8615;
    assign temp8617 = temp8616 ^ temp8616;
    assign temp8618 = temp8617 ^ temp8617;
    assign temp8619 = temp8618 ^ temp8618;
    assign temp8620 = temp8619 ^ temp8619;
    assign temp8621 = temp8620 ^ temp8620;
    assign temp8622 = temp8621 ^ temp8621;
    assign temp8623 = temp8622 ^ temp8622;
    assign temp8624 = temp8623 ^ temp8623;
    assign temp8625 = temp8624 ^ temp8624;
    assign temp8626 = temp8625 ^ temp8625;
    assign temp8627 = temp8626 ^ temp8626;
    assign temp8628 = temp8627 ^ temp8627;
    assign temp8629 = temp8628 ^ temp8628;
    assign temp8630 = temp8629 ^ temp8629;
    assign temp8631 = temp8630 ^ temp8630;
    assign temp8632 = temp8631 ^ temp8631;
    assign temp8633 = temp8632 ^ temp8632;
    assign temp8634 = temp8633 ^ temp8633;
    assign temp8635 = temp8634 ^ temp8634;
    assign temp8636 = temp8635 ^ temp8635;
    assign temp8637 = temp8636 ^ temp8636;
    assign temp8638 = temp8637 ^ temp8637;
    assign temp8639 = temp8638 ^ temp8638;
    assign temp8640 = temp8639 ^ temp8639;
    assign temp8641 = temp8640 ^ temp8640;
    assign temp8642 = temp8641 ^ temp8641;
    assign temp8643 = temp8642 ^ temp8642;
    assign temp8644 = temp8643 ^ temp8643;
    assign temp8645 = temp8644 ^ temp8644;
    assign temp8646 = temp8645 ^ temp8645;
    assign temp8647 = temp8646 ^ temp8646;
    assign temp8648 = temp8647 ^ temp8647;
    assign temp8649 = temp8648 ^ temp8648;
    assign temp8650 = temp8649 ^ temp8649;
    assign temp8651 = temp8650 ^ temp8650;
    assign temp8652 = temp8651 ^ temp8651;
    assign temp8653 = temp8652 ^ temp8652;
    assign temp8654 = temp8653 ^ temp8653;
    assign temp8655 = temp8654 ^ temp8654;
    assign temp8656 = temp8655 ^ temp8655;
    assign temp8657 = temp8656 ^ temp8656;
    assign temp8658 = temp8657 ^ temp8657;
    assign temp8659 = temp8658 ^ temp8658;
    assign temp8660 = temp8659 ^ temp8659;
    assign temp8661 = temp8660 ^ temp8660;
    assign temp8662 = temp8661 ^ temp8661;
    assign temp8663 = temp8662 ^ temp8662;
    assign temp8664 = temp8663 ^ temp8663;
    assign temp8665 = temp8664 ^ temp8664;
    assign temp8666 = temp8665 ^ temp8665;
    assign temp8667 = temp8666 ^ temp8666;
    assign temp8668 = temp8667 ^ temp8667;
    assign temp8669 = temp8668 ^ temp8668;
    assign temp8670 = temp8669 ^ temp8669;
    assign temp8671 = temp8670 ^ temp8670;
    assign temp8672 = temp8671 ^ temp8671;
    assign temp8673 = temp8672 ^ temp8672;
    assign temp8674 = temp8673 ^ temp8673;
    assign temp8675 = temp8674 ^ temp8674;
    assign temp8676 = temp8675 ^ temp8675;
    assign temp8677 = temp8676 ^ temp8676;
    assign temp8678 = temp8677 ^ temp8677;
    assign temp8679 = temp8678 ^ temp8678;
    assign temp8680 = temp8679 ^ temp8679;
    assign temp8681 = temp8680 ^ temp8680;
    assign temp8682 = temp8681 ^ temp8681;
    assign temp8683 = temp8682 ^ temp8682;
    assign temp8684 = temp8683 ^ temp8683;
    assign temp8685 = temp8684 ^ temp8684;
    assign temp8686 = temp8685 ^ temp8685;
    assign temp8687 = temp8686 ^ temp8686;
    assign temp8688 = temp8687 ^ temp8687;
    assign temp8689 = temp8688 ^ temp8688;
    assign temp8690 = temp8689 ^ temp8689;
    assign temp8691 = temp8690 ^ temp8690;
    assign temp8692 = temp8691 ^ temp8691;
    assign temp8693 = temp8692 ^ temp8692;
    assign temp8694 = temp8693 ^ temp8693;
    assign temp8695 = temp8694 ^ temp8694;
    assign temp8696 = temp8695 ^ temp8695;
    assign temp8697 = temp8696 ^ temp8696;
    assign temp8698 = temp8697 ^ temp8697;
    assign temp8699 = temp8698 ^ temp8698;
    assign temp8700 = temp8699 ^ temp8699;
    assign temp8701 = temp8700 ^ temp8700;
    assign temp8702 = temp8701 ^ temp8701;
    assign temp8703 = temp8702 ^ temp8702;
    assign temp8704 = temp8703 ^ temp8703;
    assign temp8705 = temp8704 ^ temp8704;
    assign temp8706 = temp8705 ^ temp8705;
    assign temp8707 = temp8706 ^ temp8706;
    assign temp8708 = temp8707 ^ temp8707;
    assign temp8709 = temp8708 ^ temp8708;
    assign temp8710 = temp8709 ^ temp8709;
    assign temp8711 = temp8710 ^ temp8710;
    assign temp8712 = temp8711 ^ temp8711;
    assign temp8713 = temp8712 ^ temp8712;
    assign temp8714 = temp8713 ^ temp8713;
    assign temp8715 = temp8714 ^ temp8714;
    assign temp8716 = temp8715 ^ temp8715;
    assign temp8717 = temp8716 ^ temp8716;
    assign temp8718 = temp8717 ^ temp8717;
    assign temp8719 = temp8718 ^ temp8718;
    assign temp8720 = temp8719 ^ temp8719;
    assign temp8721 = temp8720 ^ temp8720;
    assign temp8722 = temp8721 ^ temp8721;
    assign temp8723 = temp8722 ^ temp8722;
    assign temp8724 = temp8723 ^ temp8723;
    assign temp8725 = temp8724 ^ temp8724;
    assign temp8726 = temp8725 ^ temp8725;
    assign temp8727 = temp8726 ^ temp8726;
    assign temp8728 = temp8727 ^ temp8727;
    assign temp8729 = temp8728 ^ temp8728;
    assign temp8730 = temp8729 ^ temp8729;
    assign temp8731 = temp8730 ^ temp8730;
    assign temp8732 = temp8731 ^ temp8731;
    assign temp8733 = temp8732 ^ temp8732;
    assign temp8734 = temp8733 ^ temp8733;
    assign temp8735 = temp8734 ^ temp8734;
    assign temp8736 = temp8735 ^ temp8735;
    assign temp8737 = temp8736 ^ temp8736;
    assign temp8738 = temp8737 ^ temp8737;
    assign temp8739 = temp8738 ^ temp8738;
    assign temp8740 = temp8739 ^ temp8739;
    assign temp8741 = temp8740 ^ temp8740;
    assign temp8742 = temp8741 ^ temp8741;
    assign temp8743 = temp8742 ^ temp8742;
    assign temp8744 = temp8743 ^ temp8743;
    assign temp8745 = temp8744 ^ temp8744;
    assign temp8746 = temp8745 ^ temp8745;
    assign temp8747 = temp8746 ^ temp8746;
    assign temp8748 = temp8747 ^ temp8747;
    assign temp8749 = temp8748 ^ temp8748;
    assign temp8750 = temp8749 ^ temp8749;
    assign temp8751 = temp8750 ^ temp8750;
    assign temp8752 = temp8751 ^ temp8751;
    assign temp8753 = temp8752 ^ temp8752;
    assign temp8754 = temp8753 ^ temp8753;
    assign temp8755 = temp8754 ^ temp8754;
    assign temp8756 = temp8755 ^ temp8755;
    assign temp8757 = temp8756 ^ temp8756;
    assign temp8758 = temp8757 ^ temp8757;
    assign temp8759 = temp8758 ^ temp8758;
    assign temp8760 = temp8759 ^ temp8759;
    assign temp8761 = temp8760 ^ temp8760;
    assign temp8762 = temp8761 ^ temp8761;
    assign temp8763 = temp8762 ^ temp8762;
    assign temp8764 = temp8763 ^ temp8763;
    assign temp8765 = temp8764 ^ temp8764;
    assign temp8766 = temp8765 ^ temp8765;
    assign temp8767 = temp8766 ^ temp8766;
    assign temp8768 = temp8767 ^ temp8767;
    assign temp8769 = temp8768 ^ temp8768;
    assign temp8770 = temp8769 ^ temp8769;
    assign temp8771 = temp8770 ^ temp8770;
    assign temp8772 = temp8771 ^ temp8771;
    assign temp8773 = temp8772 ^ temp8772;
    assign temp8774 = temp8773 ^ temp8773;
    assign temp8775 = temp8774 ^ temp8774;
    assign temp8776 = temp8775 ^ temp8775;
    assign temp8777 = temp8776 ^ temp8776;
    assign temp8778 = temp8777 ^ temp8777;
    assign temp8779 = temp8778 ^ temp8778;
    assign temp8780 = temp8779 ^ temp8779;
    assign temp8781 = temp8780 ^ temp8780;
    assign temp8782 = temp8781 ^ temp8781;
    assign temp8783 = temp8782 ^ temp8782;
    assign temp8784 = temp8783 ^ temp8783;
    assign temp8785 = temp8784 ^ temp8784;
    assign temp8786 = temp8785 ^ temp8785;
    assign temp8787 = temp8786 ^ temp8786;
    assign temp8788 = temp8787 ^ temp8787;
    assign temp8789 = temp8788 ^ temp8788;
    assign temp8790 = temp8789 ^ temp8789;
    assign temp8791 = temp8790 ^ temp8790;
    assign temp8792 = temp8791 ^ temp8791;
    assign temp8793 = temp8792 ^ temp8792;
    assign temp8794 = temp8793 ^ temp8793;
    assign temp8795 = temp8794 ^ temp8794;
    assign temp8796 = temp8795 ^ temp8795;
    assign temp8797 = temp8796 ^ temp8796;
    assign temp8798 = temp8797 ^ temp8797;
    assign temp8799 = temp8798 ^ temp8798;
    assign temp8800 = temp8799 ^ temp8799;
    assign temp8801 = temp8800 ^ temp8800;
    assign temp8802 = temp8801 ^ temp8801;
    assign temp8803 = temp8802 ^ temp8802;
    assign temp8804 = temp8803 ^ temp8803;
    assign temp8805 = temp8804 ^ temp8804;
    assign temp8806 = temp8805 ^ temp8805;
    assign temp8807 = temp8806 ^ temp8806;
    assign temp8808 = temp8807 ^ temp8807;
    assign temp8809 = temp8808 ^ temp8808;
    assign temp8810 = temp8809 ^ temp8809;
    assign temp8811 = temp8810 ^ temp8810;
    assign temp8812 = temp8811 ^ temp8811;
    assign temp8813 = temp8812 ^ temp8812;
    assign temp8814 = temp8813 ^ temp8813;
    assign temp8815 = temp8814 ^ temp8814;
    assign temp8816 = temp8815 ^ temp8815;
    assign temp8817 = temp8816 ^ temp8816;
    assign temp8818 = temp8817 ^ temp8817;
    assign temp8819 = temp8818 ^ temp8818;
    assign temp8820 = temp8819 ^ temp8819;
    assign temp8821 = temp8820 ^ temp8820;
    assign temp8822 = temp8821 ^ temp8821;
    assign temp8823 = temp8822 ^ temp8822;
    assign temp8824 = temp8823 ^ temp8823;
    assign temp8825 = temp8824 ^ temp8824;
    assign temp8826 = temp8825 ^ temp8825;
    assign temp8827 = temp8826 ^ temp8826;
    assign temp8828 = temp8827 ^ temp8827;
    assign temp8829 = temp8828 ^ temp8828;
    assign temp8830 = temp8829 ^ temp8829;
    assign temp8831 = temp8830 ^ temp8830;
    assign temp8832 = temp8831 ^ temp8831;
    assign temp8833 = temp8832 ^ temp8832;
    assign temp8834 = temp8833 ^ temp8833;
    assign temp8835 = temp8834 ^ temp8834;
    assign temp8836 = temp8835 ^ temp8835;
    assign temp8837 = temp8836 ^ temp8836;
    assign temp8838 = temp8837 ^ temp8837;
    assign temp8839 = temp8838 ^ temp8838;
    assign temp8840 = temp8839 ^ temp8839;
    assign temp8841 = temp8840 ^ temp8840;
    assign temp8842 = temp8841 ^ temp8841;
    assign temp8843 = temp8842 ^ temp8842;
    assign temp8844 = temp8843 ^ temp8843;
    assign temp8845 = temp8844 ^ temp8844;
    assign temp8846 = temp8845 ^ temp8845;
    assign temp8847 = temp8846 ^ temp8846;
    assign temp8848 = temp8847 ^ temp8847;
    assign temp8849 = temp8848 ^ temp8848;
    assign temp8850 = temp8849 ^ temp8849;
    assign temp8851 = temp8850 ^ temp8850;
    assign temp8852 = temp8851 ^ temp8851;
    assign temp8853 = temp8852 ^ temp8852;
    assign temp8854 = temp8853 ^ temp8853;
    assign temp8855 = temp8854 ^ temp8854;
    assign temp8856 = temp8855 ^ temp8855;
    assign temp8857 = temp8856 ^ temp8856;
    assign temp8858 = temp8857 ^ temp8857;
    assign temp8859 = temp8858 ^ temp8858;
    assign temp8860 = temp8859 ^ temp8859;
    assign temp8861 = temp8860 ^ temp8860;
    assign temp8862 = temp8861 ^ temp8861;
    assign temp8863 = temp8862 ^ temp8862;
    assign temp8864 = temp8863 ^ temp8863;
    assign temp8865 = temp8864 ^ temp8864;
    assign temp8866 = temp8865 ^ temp8865;
    assign temp8867 = temp8866 ^ temp8866;
    assign temp8868 = temp8867 ^ temp8867;
    assign temp8869 = temp8868 ^ temp8868;
    assign temp8870 = temp8869 ^ temp8869;
    assign temp8871 = temp8870 ^ temp8870;
    assign temp8872 = temp8871 ^ temp8871;
    assign temp8873 = temp8872 ^ temp8872;
    assign temp8874 = temp8873 ^ temp8873;
    assign temp8875 = temp8874 ^ temp8874;
    assign temp8876 = temp8875 ^ temp8875;
    assign temp8877 = temp8876 ^ temp8876;
    assign temp8878 = temp8877 ^ temp8877;
    assign temp8879 = temp8878 ^ temp8878;
    assign temp8880 = temp8879 ^ temp8879;
    assign temp8881 = temp8880 ^ temp8880;
    assign temp8882 = temp8881 ^ temp8881;
    assign temp8883 = temp8882 ^ temp8882;
    assign temp8884 = temp8883 ^ temp8883;
    assign temp8885 = temp8884 ^ temp8884;
    assign temp8886 = temp8885 ^ temp8885;
    assign temp8887 = temp8886 ^ temp8886;
    assign temp8888 = temp8887 ^ temp8887;
    assign temp8889 = temp8888 ^ temp8888;
    assign temp8890 = temp8889 ^ temp8889;
    assign temp8891 = temp8890 ^ temp8890;
    assign temp8892 = temp8891 ^ temp8891;
    assign temp8893 = temp8892 ^ temp8892;
    assign temp8894 = temp8893 ^ temp8893;
    assign temp8895 = temp8894 ^ temp8894;
    assign temp8896 = temp8895 ^ temp8895;
    assign temp8897 = temp8896 ^ temp8896;
    assign temp8898 = temp8897 ^ temp8897;
    assign temp8899 = temp8898 ^ temp8898;
    assign temp8900 = temp8899 ^ temp8899;
    assign temp8901 = temp8900 ^ temp8900;
    assign temp8902 = temp8901 ^ temp8901;
    assign temp8903 = temp8902 ^ temp8902;
    assign temp8904 = temp8903 ^ temp8903;
    assign temp8905 = temp8904 ^ temp8904;
    assign temp8906 = temp8905 ^ temp8905;
    assign temp8907 = temp8906 ^ temp8906;
    assign temp8908 = temp8907 ^ temp8907;
    assign temp8909 = temp8908 ^ temp8908;
    assign temp8910 = temp8909 ^ temp8909;
    assign temp8911 = temp8910 ^ temp8910;
    assign temp8912 = temp8911 ^ temp8911;
    assign temp8913 = temp8912 ^ temp8912;
    assign temp8914 = temp8913 ^ temp8913;
    assign temp8915 = temp8914 ^ temp8914;
    assign temp8916 = temp8915 ^ temp8915;
    assign temp8917 = temp8916 ^ temp8916;
    assign temp8918 = temp8917 ^ temp8917;
    assign temp8919 = temp8918 ^ temp8918;
    assign temp8920 = temp8919 ^ temp8919;
    assign temp8921 = temp8920 ^ temp8920;
    assign temp8922 = temp8921 ^ temp8921;
    assign temp8923 = temp8922 ^ temp8922;
    assign temp8924 = temp8923 ^ temp8923;
    assign temp8925 = temp8924 ^ temp8924;
    assign temp8926 = temp8925 ^ temp8925;
    assign temp8927 = temp8926 ^ temp8926;
    assign temp8928 = temp8927 ^ temp8927;
    assign temp8929 = temp8928 ^ temp8928;
    assign temp8930 = temp8929 ^ temp8929;
    assign temp8931 = temp8930 ^ temp8930;
    assign temp8932 = temp8931 ^ temp8931;
    assign temp8933 = temp8932 ^ temp8932;
    assign temp8934 = temp8933 ^ temp8933;
    assign temp8935 = temp8934 ^ temp8934;
    assign temp8936 = temp8935 ^ temp8935;
    assign temp8937 = temp8936 ^ temp8936;
    assign temp8938 = temp8937 ^ temp8937;
    assign temp8939 = temp8938 ^ temp8938;
    assign temp8940 = temp8939 ^ temp8939;
    assign temp8941 = temp8940 ^ temp8940;
    assign temp8942 = temp8941 ^ temp8941;
    assign temp8943 = temp8942 ^ temp8942;
    assign temp8944 = temp8943 ^ temp8943;
    assign temp8945 = temp8944 ^ temp8944;
    assign temp8946 = temp8945 ^ temp8945;
    assign temp8947 = temp8946 ^ temp8946;
    assign temp8948 = temp8947 ^ temp8947;
    assign temp8949 = temp8948 ^ temp8948;
    assign temp8950 = temp8949 ^ temp8949;
    assign temp8951 = temp8950 ^ temp8950;
    assign temp8952 = temp8951 ^ temp8951;
    assign temp8953 = temp8952 ^ temp8952;
    assign temp8954 = temp8953 ^ temp8953;
    assign temp8955 = temp8954 ^ temp8954;
    assign temp8956 = temp8955 ^ temp8955;
    assign temp8957 = temp8956 ^ temp8956;
    assign temp8958 = temp8957 ^ temp8957;
    assign temp8959 = temp8958 ^ temp8958;
    assign temp8960 = temp8959 ^ temp8959;
    assign temp8961 = temp8960 ^ temp8960;
    assign temp8962 = temp8961 ^ temp8961;
    assign temp8963 = temp8962 ^ temp8962;
    assign temp8964 = temp8963 ^ temp8963;
    assign temp8965 = temp8964 ^ temp8964;
    assign temp8966 = temp8965 ^ temp8965;
    assign temp8967 = temp8966 ^ temp8966;
    assign temp8968 = temp8967 ^ temp8967;
    assign temp8969 = temp8968 ^ temp8968;
    assign temp8970 = temp8969 ^ temp8969;
    assign temp8971 = temp8970 ^ temp8970;
    assign temp8972 = temp8971 ^ temp8971;
    assign temp8973 = temp8972 ^ temp8972;
    assign temp8974 = temp8973 ^ temp8973;
    assign temp8975 = temp8974 ^ temp8974;
    assign temp8976 = temp8975 ^ temp8975;
    assign temp8977 = temp8976 ^ temp8976;
    assign temp8978 = temp8977 ^ temp8977;
    assign temp8979 = temp8978 ^ temp8978;
    assign temp8980 = temp8979 ^ temp8979;
    assign temp8981 = temp8980 ^ temp8980;
    assign temp8982 = temp8981 ^ temp8981;
    assign temp8983 = temp8982 ^ temp8982;
    assign temp8984 = temp8983 ^ temp8983;
    assign temp8985 = temp8984 ^ temp8984;
    assign temp8986 = temp8985 ^ temp8985;
    assign temp8987 = temp8986 ^ temp8986;
    assign temp8988 = temp8987 ^ temp8987;
    assign temp8989 = temp8988 ^ temp8988;
    assign temp8990 = temp8989 ^ temp8989;
    assign temp8991 = temp8990 ^ temp8990;
    assign temp8992 = temp8991 ^ temp8991;
    assign temp8993 = temp8992 ^ temp8992;
    assign temp8994 = temp8993 ^ temp8993;
    assign temp8995 = temp8994 ^ temp8994;
    assign temp8996 = temp8995 ^ temp8995;
    assign temp8997 = temp8996 ^ temp8996;
    assign temp8998 = temp8997 ^ temp8997;
    assign temp8999 = temp8998 ^ temp8998;
    assign temp9000 = temp8999 ^ temp8999;
    assign temp9001 = temp9000 ^ temp9000;
    assign temp9002 = temp9001 ^ temp9001;
    assign temp9003 = temp9002 ^ temp9002;
    assign temp9004 = temp9003 ^ temp9003;
    assign temp9005 = temp9004 ^ temp9004;
    assign temp9006 = temp9005 ^ temp9005;
    assign temp9007 = temp9006 ^ temp9006;
    assign temp9008 = temp9007 ^ temp9007;
    assign temp9009 = temp9008 ^ temp9008;
    assign temp9010 = temp9009 ^ temp9009;
    assign temp9011 = temp9010 ^ temp9010;
    assign temp9012 = temp9011 ^ temp9011;
    assign temp9013 = temp9012 ^ temp9012;
    assign temp9014 = temp9013 ^ temp9013;
    assign temp9015 = temp9014 ^ temp9014;
    assign temp9016 = temp9015 ^ temp9015;
    assign temp9017 = temp9016 ^ temp9016;
    assign temp9018 = temp9017 ^ temp9017;
    assign temp9019 = temp9018 ^ temp9018;
    assign temp9020 = temp9019 ^ temp9019;
    assign temp9021 = temp9020 ^ temp9020;
    assign temp9022 = temp9021 ^ temp9021;
    assign temp9023 = temp9022 ^ temp9022;
    assign temp9024 = temp9023 ^ temp9023;
    assign temp9025 = temp9024 ^ temp9024;
    assign temp9026 = temp9025 ^ temp9025;
    assign temp9027 = temp9026 ^ temp9026;
    assign temp9028 = temp9027 ^ temp9027;
    assign temp9029 = temp9028 ^ temp9028;
    assign temp9030 = temp9029 ^ temp9029;
    assign temp9031 = temp9030 ^ temp9030;
    assign temp9032 = temp9031 ^ temp9031;
    assign temp9033 = temp9032 ^ temp9032;
    assign temp9034 = temp9033 ^ temp9033;
    assign temp9035 = temp9034 ^ temp9034;
    assign temp9036 = temp9035 ^ temp9035;
    assign temp9037 = temp9036 ^ temp9036;
    assign temp9038 = temp9037 ^ temp9037;
    assign temp9039 = temp9038 ^ temp9038;
    assign temp9040 = temp9039 ^ temp9039;
    assign temp9041 = temp9040 ^ temp9040;
    assign temp9042 = temp9041 ^ temp9041;
    assign temp9043 = temp9042 ^ temp9042;
    assign temp9044 = temp9043 ^ temp9043;
    assign temp9045 = temp9044 ^ temp9044;
    assign temp9046 = temp9045 ^ temp9045;
    assign temp9047 = temp9046 ^ temp9046;
    assign temp9048 = temp9047 ^ temp9047;
    assign temp9049 = temp9048 ^ temp9048;
    assign temp9050 = temp9049 ^ temp9049;
    assign temp9051 = temp9050 ^ temp9050;
    assign temp9052 = temp9051 ^ temp9051;
    assign temp9053 = temp9052 ^ temp9052;
    assign temp9054 = temp9053 ^ temp9053;
    assign temp9055 = temp9054 ^ temp9054;
    assign temp9056 = temp9055 ^ temp9055;
    assign temp9057 = temp9056 ^ temp9056;
    assign temp9058 = temp9057 ^ temp9057;
    assign temp9059 = temp9058 ^ temp9058;
    assign temp9060 = temp9059 ^ temp9059;
    assign temp9061 = temp9060 ^ temp9060;
    assign temp9062 = temp9061 ^ temp9061;
    assign temp9063 = temp9062 ^ temp9062;
    assign temp9064 = temp9063 ^ temp9063;
    assign temp9065 = temp9064 ^ temp9064;
    assign temp9066 = temp9065 ^ temp9065;
    assign temp9067 = temp9066 ^ temp9066;
    assign temp9068 = temp9067 ^ temp9067;
    assign temp9069 = temp9068 ^ temp9068;
    assign temp9070 = temp9069 ^ temp9069;
    assign temp9071 = temp9070 ^ temp9070;
    assign temp9072 = temp9071 ^ temp9071;
    assign temp9073 = temp9072 ^ temp9072;
    assign temp9074 = temp9073 ^ temp9073;
    assign temp9075 = temp9074 ^ temp9074;
    assign temp9076 = temp9075 ^ temp9075;
    assign temp9077 = temp9076 ^ temp9076;
    assign temp9078 = temp9077 ^ temp9077;
    assign temp9079 = temp9078 ^ temp9078;
    assign temp9080 = temp9079 ^ temp9079;
    assign temp9081 = temp9080 ^ temp9080;
    assign temp9082 = temp9081 ^ temp9081;
    assign temp9083 = temp9082 ^ temp9082;
    assign temp9084 = temp9083 ^ temp9083;
    assign temp9085 = temp9084 ^ temp9084;
    assign temp9086 = temp9085 ^ temp9085;
    assign temp9087 = temp9086 ^ temp9086;
    assign temp9088 = temp9087 ^ temp9087;
    assign temp9089 = temp9088 ^ temp9088;
    assign temp9090 = temp9089 ^ temp9089;
    assign temp9091 = temp9090 ^ temp9090;
    assign temp9092 = temp9091 ^ temp9091;
    assign temp9093 = temp9092 ^ temp9092;
    assign temp9094 = temp9093 ^ temp9093;
    assign temp9095 = temp9094 ^ temp9094;
    assign temp9096 = temp9095 ^ temp9095;
    assign temp9097 = temp9096 ^ temp9096;
    assign temp9098 = temp9097 ^ temp9097;
    assign temp9099 = temp9098 ^ temp9098;
    assign temp9100 = temp9099 ^ temp9099;
    assign temp9101 = temp9100 ^ temp9100;
    assign temp9102 = temp9101 ^ temp9101;
    assign temp9103 = temp9102 ^ temp9102;
    assign temp9104 = temp9103 ^ temp9103;
    assign temp9105 = temp9104 ^ temp9104;
    assign temp9106 = temp9105 ^ temp9105;
    assign temp9107 = temp9106 ^ temp9106;
    assign temp9108 = temp9107 ^ temp9107;
    assign temp9109 = temp9108 ^ temp9108;
    assign temp9110 = temp9109 ^ temp9109;
    assign temp9111 = temp9110 ^ temp9110;
    assign temp9112 = temp9111 ^ temp9111;
    assign temp9113 = temp9112 ^ temp9112;
    assign temp9114 = temp9113 ^ temp9113;
    assign temp9115 = temp9114 ^ temp9114;
    assign temp9116 = temp9115 ^ temp9115;
    assign temp9117 = temp9116 ^ temp9116;
    assign temp9118 = temp9117 ^ temp9117;
    assign temp9119 = temp9118 ^ temp9118;
    assign temp9120 = temp9119 ^ temp9119;
    assign temp9121 = temp9120 ^ temp9120;
    assign temp9122 = temp9121 ^ temp9121;
    assign temp9123 = temp9122 ^ temp9122;
    assign temp9124 = temp9123 ^ temp9123;
    assign temp9125 = temp9124 ^ temp9124;
    assign temp9126 = temp9125 ^ temp9125;
    assign temp9127 = temp9126 ^ temp9126;
    assign temp9128 = temp9127 ^ temp9127;
    assign temp9129 = temp9128 ^ temp9128;
    assign temp9130 = temp9129 ^ temp9129;
    assign temp9131 = temp9130 ^ temp9130;
    assign temp9132 = temp9131 ^ temp9131;
    assign temp9133 = temp9132 ^ temp9132;
    assign temp9134 = temp9133 ^ temp9133;
    assign temp9135 = temp9134 ^ temp9134;
    assign temp9136 = temp9135 ^ temp9135;
    assign temp9137 = temp9136 ^ temp9136;
    assign temp9138 = temp9137 ^ temp9137;
    assign temp9139 = temp9138 ^ temp9138;
    assign temp9140 = temp9139 ^ temp9139;
    assign temp9141 = temp9140 ^ temp9140;
    assign temp9142 = temp9141 ^ temp9141;
    assign temp9143 = temp9142 ^ temp9142;
    assign temp9144 = temp9143 ^ temp9143;
    assign temp9145 = temp9144 ^ temp9144;
    assign temp9146 = temp9145 ^ temp9145;
    assign temp9147 = temp9146 ^ temp9146;
    assign temp9148 = temp9147 ^ temp9147;
    assign temp9149 = temp9148 ^ temp9148;
    assign temp9150 = temp9149 ^ temp9149;
    assign temp9151 = temp9150 ^ temp9150;
    assign temp9152 = temp9151 ^ temp9151;
    assign temp9153 = temp9152 ^ temp9152;
    assign temp9154 = temp9153 ^ temp9153;
    assign temp9155 = temp9154 ^ temp9154;
    assign temp9156 = temp9155 ^ temp9155;
    assign temp9157 = temp9156 ^ temp9156;
    assign temp9158 = temp9157 ^ temp9157;
    assign temp9159 = temp9158 ^ temp9158;
    assign temp9160 = temp9159 ^ temp9159;
    assign temp9161 = temp9160 ^ temp9160;
    assign temp9162 = temp9161 ^ temp9161;
    assign temp9163 = temp9162 ^ temp9162;
    assign temp9164 = temp9163 ^ temp9163;
    assign temp9165 = temp9164 ^ temp9164;
    assign temp9166 = temp9165 ^ temp9165;
    assign temp9167 = temp9166 ^ temp9166;
    assign temp9168 = temp9167 ^ temp9167;
    assign temp9169 = temp9168 ^ temp9168;
    assign temp9170 = temp9169 ^ temp9169;
    assign temp9171 = temp9170 ^ temp9170;
    assign temp9172 = temp9171 ^ temp9171;
    assign temp9173 = temp9172 ^ temp9172;
    assign temp9174 = temp9173 ^ temp9173;
    assign temp9175 = temp9174 ^ temp9174;
    assign temp9176 = temp9175 ^ temp9175;
    assign temp9177 = temp9176 ^ temp9176;
    assign temp9178 = temp9177 ^ temp9177;
    assign temp9179 = temp9178 ^ temp9178;
    assign temp9180 = temp9179 ^ temp9179;
    assign temp9181 = temp9180 ^ temp9180;
    assign temp9182 = temp9181 ^ temp9181;
    assign temp9183 = temp9182 ^ temp9182;
    assign temp9184 = temp9183 ^ temp9183;
    assign temp9185 = temp9184 ^ temp9184;
    assign temp9186 = temp9185 ^ temp9185;
    assign temp9187 = temp9186 ^ temp9186;
    assign temp9188 = temp9187 ^ temp9187;
    assign temp9189 = temp9188 ^ temp9188;
    assign temp9190 = temp9189 ^ temp9189;
    assign temp9191 = temp9190 ^ temp9190;
    assign temp9192 = temp9191 ^ temp9191;
    assign temp9193 = temp9192 ^ temp9192;
    assign temp9194 = temp9193 ^ temp9193;
    assign temp9195 = temp9194 ^ temp9194;
    assign temp9196 = temp9195 ^ temp9195;
    assign temp9197 = temp9196 ^ temp9196;
    assign temp9198 = temp9197 ^ temp9197;
    assign temp9199 = temp9198 ^ temp9198;
    assign temp9200 = temp9199 ^ temp9199;
    assign temp9201 = temp9200 ^ temp9200;
    assign temp9202 = temp9201 ^ temp9201;
    assign temp9203 = temp9202 ^ temp9202;
    assign temp9204 = temp9203 ^ temp9203;
    assign temp9205 = temp9204 ^ temp9204;
    assign temp9206 = temp9205 ^ temp9205;
    assign temp9207 = temp9206 ^ temp9206;
    assign temp9208 = temp9207 ^ temp9207;
    assign temp9209 = temp9208 ^ temp9208;
    assign temp9210 = temp9209 ^ temp9209;
    assign temp9211 = temp9210 ^ temp9210;
    assign temp9212 = temp9211 ^ temp9211;
    assign temp9213 = temp9212 ^ temp9212;
    assign temp9214 = temp9213 ^ temp9213;
    assign temp9215 = temp9214 ^ temp9214;
    assign temp9216 = temp9215 ^ temp9215;
    assign temp9217 = temp9216 ^ temp9216;
    assign temp9218 = temp9217 ^ temp9217;
    assign temp9219 = temp9218 ^ temp9218;
    assign temp9220 = temp9219 ^ temp9219;
    assign temp9221 = temp9220 ^ temp9220;
    assign temp9222 = temp9221 ^ temp9221;
    assign temp9223 = temp9222 ^ temp9222;
    assign temp9224 = temp9223 ^ temp9223;
    assign temp9225 = temp9224 ^ temp9224;
    assign temp9226 = temp9225 ^ temp9225;
    assign temp9227 = temp9226 ^ temp9226;
    assign temp9228 = temp9227 ^ temp9227;
    assign temp9229 = temp9228 ^ temp9228;
    assign temp9230 = temp9229 ^ temp9229;
    assign temp9231 = temp9230 ^ temp9230;
    assign temp9232 = temp9231 ^ temp9231;
    assign temp9233 = temp9232 ^ temp9232;
    assign temp9234 = temp9233 ^ temp9233;
    assign temp9235 = temp9234 ^ temp9234;
    assign temp9236 = temp9235 ^ temp9235;
    assign temp9237 = temp9236 ^ temp9236;
    assign temp9238 = temp9237 ^ temp9237;
    assign temp9239 = temp9238 ^ temp9238;
    assign temp9240 = temp9239 ^ temp9239;
    assign temp9241 = temp9240 ^ temp9240;
    assign temp9242 = temp9241 ^ temp9241;
    assign temp9243 = temp9242 ^ temp9242;
    assign temp9244 = temp9243 ^ temp9243;
    assign temp9245 = temp9244 ^ temp9244;
    assign temp9246 = temp9245 ^ temp9245;
    assign temp9247 = temp9246 ^ temp9246;
    assign temp9248 = temp9247 ^ temp9247;
    assign temp9249 = temp9248 ^ temp9248;
    assign temp9250 = temp9249 ^ temp9249;
    assign temp9251 = temp9250 ^ temp9250;
    assign temp9252 = temp9251 ^ temp9251;
    assign temp9253 = temp9252 ^ temp9252;
    assign temp9254 = temp9253 ^ temp9253;
    assign temp9255 = temp9254 ^ temp9254;
    assign temp9256 = temp9255 ^ temp9255;
    assign temp9257 = temp9256 ^ temp9256;
    assign temp9258 = temp9257 ^ temp9257;
    assign temp9259 = temp9258 ^ temp9258;
    assign temp9260 = temp9259 ^ temp9259;
    assign temp9261 = temp9260 ^ temp9260;
    assign temp9262 = temp9261 ^ temp9261;
    assign temp9263 = temp9262 ^ temp9262;
    assign temp9264 = temp9263 ^ temp9263;
    assign temp9265 = temp9264 ^ temp9264;
    assign temp9266 = temp9265 ^ temp9265;
    assign temp9267 = temp9266 ^ temp9266;
    assign temp9268 = temp9267 ^ temp9267;
    assign temp9269 = temp9268 ^ temp9268;
    assign temp9270 = temp9269 ^ temp9269;
    assign temp9271 = temp9270 ^ temp9270;
    assign temp9272 = temp9271 ^ temp9271;
    assign temp9273 = temp9272 ^ temp9272;
    assign temp9274 = temp9273 ^ temp9273;
    assign temp9275 = temp9274 ^ temp9274;
    assign temp9276 = temp9275 ^ temp9275;
    assign temp9277 = temp9276 ^ temp9276;
    assign temp9278 = temp9277 ^ temp9277;
    assign temp9279 = temp9278 ^ temp9278;
    assign temp9280 = temp9279 ^ temp9279;
    assign temp9281 = temp9280 ^ temp9280;
    assign temp9282 = temp9281 ^ temp9281;
    assign temp9283 = temp9282 ^ temp9282;
    assign temp9284 = temp9283 ^ temp9283;
    assign temp9285 = temp9284 ^ temp9284;
    assign temp9286 = temp9285 ^ temp9285;
    assign temp9287 = temp9286 ^ temp9286;
    assign temp9288 = temp9287 ^ temp9287;
    assign temp9289 = temp9288 ^ temp9288;
    assign temp9290 = temp9289 ^ temp9289;
    assign temp9291 = temp9290 ^ temp9290;
    assign temp9292 = temp9291 ^ temp9291;
    assign temp9293 = temp9292 ^ temp9292;
    assign temp9294 = temp9293 ^ temp9293;
    assign temp9295 = temp9294 ^ temp9294;
    assign temp9296 = temp9295 ^ temp9295;
    assign temp9297 = temp9296 ^ temp9296;
    assign temp9298 = temp9297 ^ temp9297;
    assign temp9299 = temp9298 ^ temp9298;
    assign temp9300 = temp9299 ^ temp9299;
    assign temp9301 = temp9300 ^ temp9300;
    assign temp9302 = temp9301 ^ temp9301;
    assign temp9303 = temp9302 ^ temp9302;
    assign temp9304 = temp9303 ^ temp9303;
    assign temp9305 = temp9304 ^ temp9304;
    assign temp9306 = temp9305 ^ temp9305;
    assign temp9307 = temp9306 ^ temp9306;
    assign temp9308 = temp9307 ^ temp9307;
    assign temp9309 = temp9308 ^ temp9308;
    assign temp9310 = temp9309 ^ temp9309;
    assign temp9311 = temp9310 ^ temp9310;
    assign temp9312 = temp9311 ^ temp9311;
    assign temp9313 = temp9312 ^ temp9312;
    assign temp9314 = temp9313 ^ temp9313;
    assign temp9315 = temp9314 ^ temp9314;
    assign temp9316 = temp9315 ^ temp9315;
    assign temp9317 = temp9316 ^ temp9316;
    assign temp9318 = temp9317 ^ temp9317;
    assign temp9319 = temp9318 ^ temp9318;
    assign temp9320 = temp9319 ^ temp9319;
    assign temp9321 = temp9320 ^ temp9320;
    assign temp9322 = temp9321 ^ temp9321;
    assign temp9323 = temp9322 ^ temp9322;
    assign temp9324 = temp9323 ^ temp9323;
    assign temp9325 = temp9324 ^ temp9324;
    assign temp9326 = temp9325 ^ temp9325;
    assign temp9327 = temp9326 ^ temp9326;
    assign temp9328 = temp9327 ^ temp9327;
    assign temp9329 = temp9328 ^ temp9328;
    assign temp9330 = temp9329 ^ temp9329;
    assign temp9331 = temp9330 ^ temp9330;
    assign temp9332 = temp9331 ^ temp9331;
    assign temp9333 = temp9332 ^ temp9332;
    assign temp9334 = temp9333 ^ temp9333;
    assign temp9335 = temp9334 ^ temp9334;
    assign temp9336 = temp9335 ^ temp9335;
    assign temp9337 = temp9336 ^ temp9336;
    assign temp9338 = temp9337 ^ temp9337;
    assign temp9339 = temp9338 ^ temp9338;
    assign temp9340 = temp9339 ^ temp9339;
    assign temp9341 = temp9340 ^ temp9340;
    assign temp9342 = temp9341 ^ temp9341;
    assign temp9343 = temp9342 ^ temp9342;
    assign temp9344 = temp9343 ^ temp9343;
    assign temp9345 = temp9344 ^ temp9344;
    assign temp9346 = temp9345 ^ temp9345;
    assign temp9347 = temp9346 ^ temp9346;
    assign temp9348 = temp9347 ^ temp9347;
    assign temp9349 = temp9348 ^ temp9348;
    assign temp9350 = temp9349 ^ temp9349;
    assign temp9351 = temp9350 ^ temp9350;
    assign temp9352 = temp9351 ^ temp9351;
    assign temp9353 = temp9352 ^ temp9352;
    assign temp9354 = temp9353 ^ temp9353;
    assign temp9355 = temp9354 ^ temp9354;
    assign temp9356 = temp9355 ^ temp9355;
    assign temp9357 = temp9356 ^ temp9356;
    assign temp9358 = temp9357 ^ temp9357;
    assign temp9359 = temp9358 ^ temp9358;
    assign temp9360 = temp9359 ^ temp9359;
    assign temp9361 = temp9360 ^ temp9360;
    assign temp9362 = temp9361 ^ temp9361;
    assign temp9363 = temp9362 ^ temp9362;
    assign temp9364 = temp9363 ^ temp9363;
    assign temp9365 = temp9364 ^ temp9364;
    assign temp9366 = temp9365 ^ temp9365;
    assign temp9367 = temp9366 ^ temp9366;
    assign temp9368 = temp9367 ^ temp9367;
    assign temp9369 = temp9368 ^ temp9368;
    assign temp9370 = temp9369 ^ temp9369;
    assign temp9371 = temp9370 ^ temp9370;
    assign temp9372 = temp9371 ^ temp9371;
    assign temp9373 = temp9372 ^ temp9372;
    assign temp9374 = temp9373 ^ temp9373;
    assign temp9375 = temp9374 ^ temp9374;
    assign temp9376 = temp9375 ^ temp9375;
    assign temp9377 = temp9376 ^ temp9376;
    assign temp9378 = temp9377 ^ temp9377;
    assign temp9379 = temp9378 ^ temp9378;
    assign temp9380 = temp9379 ^ temp9379;
    assign temp9381 = temp9380 ^ temp9380;
    assign temp9382 = temp9381 ^ temp9381;
    assign temp9383 = temp9382 ^ temp9382;
    assign temp9384 = temp9383 ^ temp9383;
    assign temp9385 = temp9384 ^ temp9384;
    assign temp9386 = temp9385 ^ temp9385;
    assign temp9387 = temp9386 ^ temp9386;
    assign temp9388 = temp9387 ^ temp9387;
    assign temp9389 = temp9388 ^ temp9388;
    assign temp9390 = temp9389 ^ temp9389;
    assign temp9391 = temp9390 ^ temp9390;
    assign temp9392 = temp9391 ^ temp9391;
    assign temp9393 = temp9392 ^ temp9392;
    assign temp9394 = temp9393 ^ temp9393;
    assign temp9395 = temp9394 ^ temp9394;
    assign temp9396 = temp9395 ^ temp9395;
    assign temp9397 = temp9396 ^ temp9396;
    assign temp9398 = temp9397 ^ temp9397;
    assign temp9399 = temp9398 ^ temp9398;
    assign temp9400 = temp9399 ^ temp9399;
    assign temp9401 = temp9400 ^ temp9400;
    assign temp9402 = temp9401 ^ temp9401;
    assign temp9403 = temp9402 ^ temp9402;
    assign temp9404 = temp9403 ^ temp9403;
    assign temp9405 = temp9404 ^ temp9404;
    assign temp9406 = temp9405 ^ temp9405;
    assign temp9407 = temp9406 ^ temp9406;
    assign temp9408 = temp9407 ^ temp9407;
    assign temp9409 = temp9408 ^ temp9408;
    assign temp9410 = temp9409 ^ temp9409;
    assign temp9411 = temp9410 ^ temp9410;
    assign temp9412 = temp9411 ^ temp9411;
    assign temp9413 = temp9412 ^ temp9412;
    assign temp9414 = temp9413 ^ temp9413;
    assign temp9415 = temp9414 ^ temp9414;
    assign temp9416 = temp9415 ^ temp9415;
    assign temp9417 = temp9416 ^ temp9416;
    assign temp9418 = temp9417 ^ temp9417;
    assign temp9419 = temp9418 ^ temp9418;
    assign temp9420 = temp9419 ^ temp9419;
    assign temp9421 = temp9420 ^ temp9420;
    assign temp9422 = temp9421 ^ temp9421;
    assign temp9423 = temp9422 ^ temp9422;
    assign temp9424 = temp9423 ^ temp9423;
    assign temp9425 = temp9424 ^ temp9424;
    assign temp9426 = temp9425 ^ temp9425;
    assign temp9427 = temp9426 ^ temp9426;
    assign temp9428 = temp9427 ^ temp9427;
    assign temp9429 = temp9428 ^ temp9428;
    assign temp9430 = temp9429 ^ temp9429;
    assign temp9431 = temp9430 ^ temp9430;
    assign temp9432 = temp9431 ^ temp9431;
    assign temp9433 = temp9432 ^ temp9432;
    assign temp9434 = temp9433 ^ temp9433;
    assign temp9435 = temp9434 ^ temp9434;
    assign temp9436 = temp9435 ^ temp9435;
    assign temp9437 = temp9436 ^ temp9436;
    assign temp9438 = temp9437 ^ temp9437;
    assign temp9439 = temp9438 ^ temp9438;
    assign temp9440 = temp9439 ^ temp9439;
    assign temp9441 = temp9440 ^ temp9440;
    assign temp9442 = temp9441 ^ temp9441;
    assign temp9443 = temp9442 ^ temp9442;
    assign temp9444 = temp9443 ^ temp9443;
    assign temp9445 = temp9444 ^ temp9444;
    assign temp9446 = temp9445 ^ temp9445;
    assign temp9447 = temp9446 ^ temp9446;
    assign temp9448 = temp9447 ^ temp9447;
    assign temp9449 = temp9448 ^ temp9448;
    assign temp9450 = temp9449 ^ temp9449;
    assign temp9451 = temp9450 ^ temp9450;
    assign temp9452 = temp9451 ^ temp9451;
    assign temp9453 = temp9452 ^ temp9452;
    assign temp9454 = temp9453 ^ temp9453;
    assign temp9455 = temp9454 ^ temp9454;
    assign temp9456 = temp9455 ^ temp9455;
    assign temp9457 = temp9456 ^ temp9456;
    assign temp9458 = temp9457 ^ temp9457;
    assign temp9459 = temp9458 ^ temp9458;
    assign temp9460 = temp9459 ^ temp9459;
    assign temp9461 = temp9460 ^ temp9460;
    assign temp9462 = temp9461 ^ temp9461;
    assign temp9463 = temp9462 ^ temp9462;
    assign temp9464 = temp9463 ^ temp9463;
    assign temp9465 = temp9464 ^ temp9464;
    assign temp9466 = temp9465 ^ temp9465;
    assign temp9467 = temp9466 ^ temp9466;
    assign temp9468 = temp9467 ^ temp9467;
    assign temp9469 = temp9468 ^ temp9468;
    assign temp9470 = temp9469 ^ temp9469;
    assign temp9471 = temp9470 ^ temp9470;
    assign temp9472 = temp9471 ^ temp9471;
    assign temp9473 = temp9472 ^ temp9472;
    assign temp9474 = temp9473 ^ temp9473;
    assign temp9475 = temp9474 ^ temp9474;
    assign temp9476 = temp9475 ^ temp9475;
    assign temp9477 = temp9476 ^ temp9476;
    assign temp9478 = temp9477 ^ temp9477;
    assign temp9479 = temp9478 ^ temp9478;
    assign temp9480 = temp9479 ^ temp9479;
    assign temp9481 = temp9480 ^ temp9480;
    assign temp9482 = temp9481 ^ temp9481;
    assign temp9483 = temp9482 ^ temp9482;
    assign temp9484 = temp9483 ^ temp9483;
    assign temp9485 = temp9484 ^ temp9484;
    assign temp9486 = temp9485 ^ temp9485;
    assign temp9487 = temp9486 ^ temp9486;
    assign temp9488 = temp9487 ^ temp9487;
    assign temp9489 = temp9488 ^ temp9488;
    assign temp9490 = temp9489 ^ temp9489;
    assign temp9491 = temp9490 ^ temp9490;
    assign temp9492 = temp9491 ^ temp9491;
    assign temp9493 = temp9492 ^ temp9492;
    assign temp9494 = temp9493 ^ temp9493;
    assign temp9495 = temp9494 ^ temp9494;
    assign temp9496 = temp9495 ^ temp9495;
    assign temp9497 = temp9496 ^ temp9496;
    assign temp9498 = temp9497 ^ temp9497;
    assign temp9499 = temp9498 ^ temp9498;
    assign temp9500 = temp9499 ^ temp9499;
    assign temp9501 = temp9500 ^ temp9500;
    assign temp9502 = temp9501 ^ temp9501;
    assign temp9503 = temp9502 ^ temp9502;
    assign temp9504 = temp9503 ^ temp9503;
    assign temp9505 = temp9504 ^ temp9504;
    assign temp9506 = temp9505 ^ temp9505;
    assign temp9507 = temp9506 ^ temp9506;
    assign temp9508 = temp9507 ^ temp9507;
    assign temp9509 = temp9508 ^ temp9508;
    assign temp9510 = temp9509 ^ temp9509;
    assign temp9511 = temp9510 ^ temp9510;
    assign temp9512 = temp9511 ^ temp9511;
    assign temp9513 = temp9512 ^ temp9512;
    assign temp9514 = temp9513 ^ temp9513;
    assign temp9515 = temp9514 ^ temp9514;
    assign temp9516 = temp9515 ^ temp9515;
    assign temp9517 = temp9516 ^ temp9516;
    assign temp9518 = temp9517 ^ temp9517;
    assign temp9519 = temp9518 ^ temp9518;
    assign temp9520 = temp9519 ^ temp9519;
    assign temp9521 = temp9520 ^ temp9520;
    assign temp9522 = temp9521 ^ temp9521;
    assign temp9523 = temp9522 ^ temp9522;
    assign temp9524 = temp9523 ^ temp9523;
    assign temp9525 = temp9524 ^ temp9524;
    assign temp9526 = temp9525 ^ temp9525;
    assign temp9527 = temp9526 ^ temp9526;
    assign temp9528 = temp9527 ^ temp9527;
    assign temp9529 = temp9528 ^ temp9528;
    assign temp9530 = temp9529 ^ temp9529;
    assign temp9531 = temp9530 ^ temp9530;
    assign temp9532 = temp9531 ^ temp9531;
    assign temp9533 = temp9532 ^ temp9532;
    assign temp9534 = temp9533 ^ temp9533;
    assign temp9535 = temp9534 ^ temp9534;
    assign temp9536 = temp9535 ^ temp9535;
    assign temp9537 = temp9536 ^ temp9536;
    assign temp9538 = temp9537 ^ temp9537;
    assign temp9539 = temp9538 ^ temp9538;
    assign temp9540 = temp9539 ^ temp9539;
    assign temp9541 = temp9540 ^ temp9540;
    assign temp9542 = temp9541 ^ temp9541;
    assign temp9543 = temp9542 ^ temp9542;
    assign temp9544 = temp9543 ^ temp9543;
    assign temp9545 = temp9544 ^ temp9544;
    assign temp9546 = temp9545 ^ temp9545;
    assign temp9547 = temp9546 ^ temp9546;
    assign temp9548 = temp9547 ^ temp9547;
    assign temp9549 = temp9548 ^ temp9548;
    assign temp9550 = temp9549 ^ temp9549;
    assign temp9551 = temp9550 ^ temp9550;
    assign temp9552 = temp9551 ^ temp9551;
    assign temp9553 = temp9552 ^ temp9552;
    assign temp9554 = temp9553 ^ temp9553;
    assign temp9555 = temp9554 ^ temp9554;
    assign temp9556 = temp9555 ^ temp9555;
    assign temp9557 = temp9556 ^ temp9556;
    assign temp9558 = temp9557 ^ temp9557;
    assign temp9559 = temp9558 ^ temp9558;
    assign temp9560 = temp9559 ^ temp9559;
    assign temp9561 = temp9560 ^ temp9560;
    assign temp9562 = temp9561 ^ temp9561;
    assign temp9563 = temp9562 ^ temp9562;
    assign temp9564 = temp9563 ^ temp9563;
    assign temp9565 = temp9564 ^ temp9564;
    assign temp9566 = temp9565 ^ temp9565;
    assign temp9567 = temp9566 ^ temp9566;
    assign temp9568 = temp9567 ^ temp9567;
    assign temp9569 = temp9568 ^ temp9568;
    assign temp9570 = temp9569 ^ temp9569;
    assign temp9571 = temp9570 ^ temp9570;
    assign temp9572 = temp9571 ^ temp9571;
    assign temp9573 = temp9572 ^ temp9572;
    assign temp9574 = temp9573 ^ temp9573;
    assign temp9575 = temp9574 ^ temp9574;
    assign temp9576 = temp9575 ^ temp9575;
    assign temp9577 = temp9576 ^ temp9576;
    assign temp9578 = temp9577 ^ temp9577;
    assign temp9579 = temp9578 ^ temp9578;
    assign temp9580 = temp9579 ^ temp9579;
    assign temp9581 = temp9580 ^ temp9580;
    assign temp9582 = temp9581 ^ temp9581;
    assign temp9583 = temp9582 ^ temp9582;
    assign temp9584 = temp9583 ^ temp9583;
    assign temp9585 = temp9584 ^ temp9584;
    assign temp9586 = temp9585 ^ temp9585;
    assign temp9587 = temp9586 ^ temp9586;
    assign temp9588 = temp9587 ^ temp9587;
    assign temp9589 = temp9588 ^ temp9588;
    assign temp9590 = temp9589 ^ temp9589;
    assign temp9591 = temp9590 ^ temp9590;
    assign temp9592 = temp9591 ^ temp9591;
    assign temp9593 = temp9592 ^ temp9592;
    assign temp9594 = temp9593 ^ temp9593;
    assign temp9595 = temp9594 ^ temp9594;
    assign temp9596 = temp9595 ^ temp9595;
    assign temp9597 = temp9596 ^ temp9596;
    assign temp9598 = temp9597 ^ temp9597;
    assign temp9599 = temp9598 ^ temp9598;
    assign temp9600 = temp9599 ^ temp9599;
    assign temp9601 = temp9600 ^ temp9600;
    assign temp9602 = temp9601 ^ temp9601;
    assign temp9603 = temp9602 ^ temp9602;
    assign temp9604 = temp9603 ^ temp9603;
    assign temp9605 = temp9604 ^ temp9604;
    assign temp9606 = temp9605 ^ temp9605;
    assign temp9607 = temp9606 ^ temp9606;
    assign temp9608 = temp9607 ^ temp9607;
    assign temp9609 = temp9608 ^ temp9608;
    assign temp9610 = temp9609 ^ temp9609;
    assign temp9611 = temp9610 ^ temp9610;
    assign temp9612 = temp9611 ^ temp9611;
    assign temp9613 = temp9612 ^ temp9612;
    assign temp9614 = temp9613 ^ temp9613;
    assign temp9615 = temp9614 ^ temp9614;
    assign temp9616 = temp9615 ^ temp9615;
    assign temp9617 = temp9616 ^ temp9616;
    assign temp9618 = temp9617 ^ temp9617;
    assign temp9619 = temp9618 ^ temp9618;
    assign temp9620 = temp9619 ^ temp9619;
    assign temp9621 = temp9620 ^ temp9620;
    assign temp9622 = temp9621 ^ temp9621;
    assign temp9623 = temp9622 ^ temp9622;
    assign temp9624 = temp9623 ^ temp9623;
    assign temp9625 = temp9624 ^ temp9624;
    assign temp9626 = temp9625 ^ temp9625;
    assign temp9627 = temp9626 ^ temp9626;
    assign temp9628 = temp9627 ^ temp9627;
    assign temp9629 = temp9628 ^ temp9628;
    assign temp9630 = temp9629 ^ temp9629;
    assign temp9631 = temp9630 ^ temp9630;
    assign temp9632 = temp9631 ^ temp9631;
    assign temp9633 = temp9632 ^ temp9632;
    assign temp9634 = temp9633 ^ temp9633;
    assign temp9635 = temp9634 ^ temp9634;
    assign temp9636 = temp9635 ^ temp9635;
    assign temp9637 = temp9636 ^ temp9636;
    assign temp9638 = temp9637 ^ temp9637;
    assign temp9639 = temp9638 ^ temp9638;
    assign temp9640 = temp9639 ^ temp9639;
    assign temp9641 = temp9640 ^ temp9640;
    assign temp9642 = temp9641 ^ temp9641;
    assign temp9643 = temp9642 ^ temp9642;
    assign temp9644 = temp9643 ^ temp9643;
    assign temp9645 = temp9644 ^ temp9644;
    assign temp9646 = temp9645 ^ temp9645;
    assign temp9647 = temp9646 ^ temp9646;
    assign temp9648 = temp9647 ^ temp9647;
    assign temp9649 = temp9648 ^ temp9648;
    assign temp9650 = temp9649 ^ temp9649;
    assign temp9651 = temp9650 ^ temp9650;
    assign temp9652 = temp9651 ^ temp9651;
    assign temp9653 = temp9652 ^ temp9652;
    assign temp9654 = temp9653 ^ temp9653;
    assign temp9655 = temp9654 ^ temp9654;
    assign temp9656 = temp9655 ^ temp9655;
    assign temp9657 = temp9656 ^ temp9656;
    assign temp9658 = temp9657 ^ temp9657;
    assign temp9659 = temp9658 ^ temp9658;
    assign temp9660 = temp9659 ^ temp9659;
    assign temp9661 = temp9660 ^ temp9660;
    assign temp9662 = temp9661 ^ temp9661;
    assign temp9663 = temp9662 ^ temp9662;
    assign temp9664 = temp9663 ^ temp9663;
    assign temp9665 = temp9664 ^ temp9664;
    assign temp9666 = temp9665 ^ temp9665;
    assign temp9667 = temp9666 ^ temp9666;
    assign temp9668 = temp9667 ^ temp9667;
    assign temp9669 = temp9668 ^ temp9668;
    assign temp9670 = temp9669 ^ temp9669;
    assign temp9671 = temp9670 ^ temp9670;
    assign temp9672 = temp9671 ^ temp9671;
    assign temp9673 = temp9672 ^ temp9672;
    assign temp9674 = temp9673 ^ temp9673;
    assign temp9675 = temp9674 ^ temp9674;
    assign temp9676 = temp9675 ^ temp9675;
    assign temp9677 = temp9676 ^ temp9676;
    assign temp9678 = temp9677 ^ temp9677;
    assign temp9679 = temp9678 ^ temp9678;
    assign temp9680 = temp9679 ^ temp9679;
    assign temp9681 = temp9680 ^ temp9680;
    assign temp9682 = temp9681 ^ temp9681;
    assign temp9683 = temp9682 ^ temp9682;
    assign temp9684 = temp9683 ^ temp9683;
    assign temp9685 = temp9684 ^ temp9684;
    assign temp9686 = temp9685 ^ temp9685;
    assign temp9687 = temp9686 ^ temp9686;
    assign temp9688 = temp9687 ^ temp9687;
    assign temp9689 = temp9688 ^ temp9688;
    assign temp9690 = temp9689 ^ temp9689;
    assign temp9691 = temp9690 ^ temp9690;
    assign temp9692 = temp9691 ^ temp9691;
    assign temp9693 = temp9692 ^ temp9692;
    assign temp9694 = temp9693 ^ temp9693;
    assign temp9695 = temp9694 ^ temp9694;
    assign temp9696 = temp9695 ^ temp9695;
    assign temp9697 = temp9696 ^ temp9696;
    assign temp9698 = temp9697 ^ temp9697;
    assign temp9699 = temp9698 ^ temp9698;
    assign temp9700 = temp9699 ^ temp9699;
    assign temp9701 = temp9700 ^ temp9700;
    assign temp9702 = temp9701 ^ temp9701;
    assign temp9703 = temp9702 ^ temp9702;
    assign temp9704 = temp9703 ^ temp9703;
    assign temp9705 = temp9704 ^ temp9704;
    assign temp9706 = temp9705 ^ temp9705;
    assign temp9707 = temp9706 ^ temp9706;
    assign temp9708 = temp9707 ^ temp9707;
    assign temp9709 = temp9708 ^ temp9708;
    assign temp9710 = temp9709 ^ temp9709;
    assign temp9711 = temp9710 ^ temp9710;
    assign temp9712 = temp9711 ^ temp9711;
    assign temp9713 = temp9712 ^ temp9712;
    assign temp9714 = temp9713 ^ temp9713;
    assign temp9715 = temp9714 ^ temp9714;
    assign temp9716 = temp9715 ^ temp9715;
    assign temp9717 = temp9716 ^ temp9716;
    assign temp9718 = temp9717 ^ temp9717;
    assign temp9719 = temp9718 ^ temp9718;
    assign temp9720 = temp9719 ^ temp9719;
    assign temp9721 = temp9720 ^ temp9720;
    assign temp9722 = temp9721 ^ temp9721;
    assign temp9723 = temp9722 ^ temp9722;
    assign temp9724 = temp9723 ^ temp9723;
    assign temp9725 = temp9724 ^ temp9724;
    assign temp9726 = temp9725 ^ temp9725;
    assign temp9727 = temp9726 ^ temp9726;
    assign temp9728 = temp9727 ^ temp9727;
    assign temp9729 = temp9728 ^ temp9728;
    assign temp9730 = temp9729 ^ temp9729;
    assign temp9731 = temp9730 ^ temp9730;
    assign temp9732 = temp9731 ^ temp9731;
    assign temp9733 = temp9732 ^ temp9732;
    assign temp9734 = temp9733 ^ temp9733;
    assign temp9735 = temp9734 ^ temp9734;
    assign temp9736 = temp9735 ^ temp9735;
    assign temp9737 = temp9736 ^ temp9736;
    assign temp9738 = temp9737 ^ temp9737;
    assign temp9739 = temp9738 ^ temp9738;
    assign temp9740 = temp9739 ^ temp9739;
    assign temp9741 = temp9740 ^ temp9740;
    assign temp9742 = temp9741 ^ temp9741;
    assign temp9743 = temp9742 ^ temp9742;
    assign temp9744 = temp9743 ^ temp9743;
    assign temp9745 = temp9744 ^ temp9744;
    assign temp9746 = temp9745 ^ temp9745;
    assign temp9747 = temp9746 ^ temp9746;
    assign temp9748 = temp9747 ^ temp9747;
    assign temp9749 = temp9748 ^ temp9748;
    assign temp9750 = temp9749 ^ temp9749;
    assign temp9751 = temp9750 ^ temp9750;
    assign temp9752 = temp9751 ^ temp9751;
    assign temp9753 = temp9752 ^ temp9752;
    assign temp9754 = temp9753 ^ temp9753;
    assign temp9755 = temp9754 ^ temp9754;
    assign temp9756 = temp9755 ^ temp9755;
    assign temp9757 = temp9756 ^ temp9756;
    assign temp9758 = temp9757 ^ temp9757;
    assign temp9759 = temp9758 ^ temp9758;
    assign temp9760 = temp9759 ^ temp9759;
    assign temp9761 = temp9760 ^ temp9760;
    assign temp9762 = temp9761 ^ temp9761;
    assign temp9763 = temp9762 ^ temp9762;
    assign temp9764 = temp9763 ^ temp9763;
    assign temp9765 = temp9764 ^ temp9764;
    assign temp9766 = temp9765 ^ temp9765;
    assign temp9767 = temp9766 ^ temp9766;
    assign temp9768 = temp9767 ^ temp9767;
    assign temp9769 = temp9768 ^ temp9768;
    assign temp9770 = temp9769 ^ temp9769;
    assign temp9771 = temp9770 ^ temp9770;
    assign temp9772 = temp9771 ^ temp9771;
    assign temp9773 = temp9772 ^ temp9772;
    assign temp9774 = temp9773 ^ temp9773;
    assign temp9775 = temp9774 ^ temp9774;
    assign temp9776 = temp9775 ^ temp9775;
    assign temp9777 = temp9776 ^ temp9776;
    assign temp9778 = temp9777 ^ temp9777;
    assign temp9779 = temp9778 ^ temp9778;
    assign temp9780 = temp9779 ^ temp9779;
    assign temp9781 = temp9780 ^ temp9780;
    assign temp9782 = temp9781 ^ temp9781;
    assign temp9783 = temp9782 ^ temp9782;
    assign temp9784 = temp9783 ^ temp9783;
    assign temp9785 = temp9784 ^ temp9784;
    assign temp9786 = temp9785 ^ temp9785;
    assign temp9787 = temp9786 ^ temp9786;
    assign temp9788 = temp9787 ^ temp9787;
    assign temp9789 = temp9788 ^ temp9788;
    assign temp9790 = temp9789 ^ temp9789;
    assign temp9791 = temp9790 ^ temp9790;
    assign temp9792 = temp9791 ^ temp9791;
    assign temp9793 = temp9792 ^ temp9792;
    assign temp9794 = temp9793 ^ temp9793;
    assign temp9795 = temp9794 ^ temp9794;
    assign temp9796 = temp9795 ^ temp9795;
    assign temp9797 = temp9796 ^ temp9796;
    assign temp9798 = temp9797 ^ temp9797;
    assign temp9799 = temp9798 ^ temp9798;
    assign temp9800 = temp9799 ^ temp9799;
    assign temp9801 = temp9800 ^ temp9800;
    assign temp9802 = temp9801 ^ temp9801;
    assign temp9803 = temp9802 ^ temp9802;
    assign temp9804 = temp9803 ^ temp9803;
    assign temp9805 = temp9804 ^ temp9804;
    assign temp9806 = temp9805 ^ temp9805;
    assign temp9807 = temp9806 ^ temp9806;
    assign temp9808 = temp9807 ^ temp9807;
    assign temp9809 = temp9808 ^ temp9808;
    assign temp9810 = temp9809 ^ temp9809;
    assign temp9811 = temp9810 ^ temp9810;
    assign temp9812 = temp9811 ^ temp9811;
    assign temp9813 = temp9812 ^ temp9812;
    assign temp9814 = temp9813 ^ temp9813;
    assign temp9815 = temp9814 ^ temp9814;
    assign temp9816 = temp9815 ^ temp9815;
    assign temp9817 = temp9816 ^ temp9816;
    assign temp9818 = temp9817 ^ temp9817;
    assign temp9819 = temp9818 ^ temp9818;
    assign temp9820 = temp9819 ^ temp9819;
    assign temp9821 = temp9820 ^ temp9820;
    assign temp9822 = temp9821 ^ temp9821;
    assign temp9823 = temp9822 ^ temp9822;
    assign temp9824 = temp9823 ^ temp9823;
    assign temp9825 = temp9824 ^ temp9824;
    assign temp9826 = temp9825 ^ temp9825;
    assign temp9827 = temp9826 ^ temp9826;
    assign temp9828 = temp9827 ^ temp9827;
    assign temp9829 = temp9828 ^ temp9828;
    assign temp9830 = temp9829 ^ temp9829;
    assign temp9831 = temp9830 ^ temp9830;
    assign temp9832 = temp9831 ^ temp9831;
    assign temp9833 = temp9832 ^ temp9832;
    assign temp9834 = temp9833 ^ temp9833;
    assign temp9835 = temp9834 ^ temp9834;
    assign temp9836 = temp9835 ^ temp9835;
    assign temp9837 = temp9836 ^ temp9836;
    assign temp9838 = temp9837 ^ temp9837;
    assign temp9839 = temp9838 ^ temp9838;
    assign temp9840 = temp9839 ^ temp9839;
    assign temp9841 = temp9840 ^ temp9840;
    assign temp9842 = temp9841 ^ temp9841;
    assign temp9843 = temp9842 ^ temp9842;
    assign temp9844 = temp9843 ^ temp9843;
    assign temp9845 = temp9844 ^ temp9844;
    assign temp9846 = temp9845 ^ temp9845;
    assign temp9847 = temp9846 ^ temp9846;
    assign temp9848 = temp9847 ^ temp9847;
    assign temp9849 = temp9848 ^ temp9848;
    assign temp9850 = temp9849 ^ temp9849;
    assign temp9851 = temp9850 ^ temp9850;
    assign temp9852 = temp9851 ^ temp9851;
    assign temp9853 = temp9852 ^ temp9852;
    assign temp9854 = temp9853 ^ temp9853;
    assign temp9855 = temp9854 ^ temp9854;
    assign temp9856 = temp9855 ^ temp9855;
    assign temp9857 = temp9856 ^ temp9856;
    assign temp9858 = temp9857 ^ temp9857;
    assign temp9859 = temp9858 ^ temp9858;
    assign temp9860 = temp9859 ^ temp9859;
    assign temp9861 = temp9860 ^ temp9860;
    assign temp9862 = temp9861 ^ temp9861;
    assign temp9863 = temp9862 ^ temp9862;
    assign temp9864 = temp9863 ^ temp9863;
    assign temp9865 = temp9864 ^ temp9864;
    assign temp9866 = temp9865 ^ temp9865;
    assign temp9867 = temp9866 ^ temp9866;
    assign temp9868 = temp9867 ^ temp9867;
    assign temp9869 = temp9868 ^ temp9868;
    assign temp9870 = temp9869 ^ temp9869;
    assign temp9871 = temp9870 ^ temp9870;
    assign temp9872 = temp9871 ^ temp9871;
    assign temp9873 = temp9872 ^ temp9872;
    assign temp9874 = temp9873 ^ temp9873;
    assign temp9875 = temp9874 ^ temp9874;
    assign temp9876 = temp9875 ^ temp9875;
    assign temp9877 = temp9876 ^ temp9876;
    assign temp9878 = temp9877 ^ temp9877;
    assign temp9879 = temp9878 ^ temp9878;
    assign temp9880 = temp9879 ^ temp9879;
    assign temp9881 = temp9880 ^ temp9880;
    assign temp9882 = temp9881 ^ temp9881;
    assign temp9883 = temp9882 ^ temp9882;
    assign temp9884 = temp9883 ^ temp9883;
    assign temp9885 = temp9884 ^ temp9884;
    assign temp9886 = temp9885 ^ temp9885;
    assign temp9887 = temp9886 ^ temp9886;
    assign temp9888 = temp9887 ^ temp9887;
    assign temp9889 = temp9888 ^ temp9888;
    assign temp9890 = temp9889 ^ temp9889;
    assign temp9891 = temp9890 ^ temp9890;
    assign temp9892 = temp9891 ^ temp9891;
    assign temp9893 = temp9892 ^ temp9892;
    assign temp9894 = temp9893 ^ temp9893;
    assign temp9895 = temp9894 ^ temp9894;
    assign temp9896 = temp9895 ^ temp9895;
    assign temp9897 = temp9896 ^ temp9896;
    assign temp9898 = temp9897 ^ temp9897;
    assign temp9899 = temp9898 ^ temp9898;
    assign temp9900 = temp9899 ^ temp9899;
    assign temp9901 = temp9900 ^ temp9900;
    assign temp9902 = temp9901 ^ temp9901;
    assign temp9903 = temp9902 ^ temp9902;
    assign temp9904 = temp9903 ^ temp9903;
    assign temp9905 = temp9904 ^ temp9904;
    assign temp9906 = temp9905 ^ temp9905;
    assign temp9907 = temp9906 ^ temp9906;
    assign temp9908 = temp9907 ^ temp9907;
    assign temp9909 = temp9908 ^ temp9908;
    assign temp9910 = temp9909 ^ temp9909;
    assign temp9911 = temp9910 ^ temp9910;
    assign temp9912 = temp9911 ^ temp9911;
    assign temp9913 = temp9912 ^ temp9912;
    assign temp9914 = temp9913 ^ temp9913;
    assign temp9915 = temp9914 ^ temp9914;
    assign temp9916 = temp9915 ^ temp9915;
    assign temp9917 = temp9916 ^ temp9916;
    assign temp9918 = temp9917 ^ temp9917;
    assign temp9919 = temp9918 ^ temp9918;
    assign temp9920 = temp9919 ^ temp9919;
    assign temp9921 = temp9920 ^ temp9920;
    assign temp9922 = temp9921 ^ temp9921;
    assign temp9923 = temp9922 ^ temp9922;
    assign temp9924 = temp9923 ^ temp9923;
    assign temp9925 = temp9924 ^ temp9924;
    assign temp9926 = temp9925 ^ temp9925;
    assign temp9927 = temp9926 ^ temp9926;
    assign temp9928 = temp9927 ^ temp9927;
    assign temp9929 = temp9928 ^ temp9928;
    assign temp9930 = temp9929 ^ temp9929;
    assign temp9931 = temp9930 ^ temp9930;
    assign temp9932 = temp9931 ^ temp9931;
    assign temp9933 = temp9932 ^ temp9932;
    assign temp9934 = temp9933 ^ temp9933;
    assign temp9935 = temp9934 ^ temp9934;
    assign temp9936 = temp9935 ^ temp9935;
    assign temp9937 = temp9936 ^ temp9936;
    assign temp9938 = temp9937 ^ temp9937;
    assign temp9939 = temp9938 ^ temp9938;
    assign temp9940 = temp9939 ^ temp9939;
    assign temp9941 = temp9940 ^ temp9940;
    assign temp9942 = temp9941 ^ temp9941;
    assign temp9943 = temp9942 ^ temp9942;
    assign temp9944 = temp9943 ^ temp9943;
    assign temp9945 = temp9944 ^ temp9944;
    assign temp9946 = temp9945 ^ temp9945;
    assign temp9947 = temp9946 ^ temp9946;
    assign temp9948 = temp9947 ^ temp9947;
    assign temp9949 = temp9948 ^ temp9948;
    assign temp9950 = temp9949 ^ temp9949;
    assign temp9951 = temp9950 ^ temp9950;
    assign temp9952 = temp9951 ^ temp9951;
    assign temp9953 = temp9952 ^ temp9952;
    assign temp9954 = temp9953 ^ temp9953;
    assign temp9955 = temp9954 ^ temp9954;
    assign temp9956 = temp9955 ^ temp9955;
    assign temp9957 = temp9956 ^ temp9956;
    assign temp9958 = temp9957 ^ temp9957;
    assign temp9959 = temp9958 ^ temp9958;
    assign temp9960 = temp9959 ^ temp9959;
    assign temp9961 = temp9960 ^ temp9960;
    assign temp9962 = temp9961 ^ temp9961;
    assign temp9963 = temp9962 ^ temp9962;
    assign temp9964 = temp9963 ^ temp9963;
    assign temp9965 = temp9964 ^ temp9964;
    assign temp9966 = temp9965 ^ temp9965;
    assign temp9967 = temp9966 ^ temp9966;
    assign temp9968 = temp9967 ^ temp9967;
    assign temp9969 = temp9968 ^ temp9968;
    assign temp9970 = temp9969 ^ temp9969;
    assign temp9971 = temp9970 ^ temp9970;
    assign temp9972 = temp9971 ^ temp9971;
    assign temp9973 = temp9972 ^ temp9972;
    assign temp9974 = temp9973 ^ temp9973;
    assign temp9975 = temp9974 ^ temp9974;
    assign temp9976 = temp9975 ^ temp9975;
    assign temp9977 = temp9976 ^ temp9976;
    assign temp9978 = temp9977 ^ temp9977;
    assign temp9979 = temp9978 ^ temp9978;
    assign temp9980 = temp9979 ^ temp9979;
    assign temp9981 = temp9980 ^ temp9980;
    assign temp9982 = temp9981 ^ temp9981;
    assign temp9983 = temp9982 ^ temp9982;
    assign temp9984 = temp9983 ^ temp9983;
    assign temp9985 = temp9984 ^ temp9984;
    assign temp9986 = temp9985 ^ temp9985;
    assign temp9987 = temp9986 ^ temp9986;
    assign temp9988 = temp9987 ^ temp9987;
    assign temp9989 = temp9988 ^ temp9988;
    assign temp9990 = temp9989 ^ temp9989;
    assign temp9991 = temp9990 ^ temp9990;
    assign temp9992 = temp9991 ^ temp9991;
    assign temp9993 = temp9992 ^ temp9992;
    assign temp9994 = temp9993 ^ temp9993;
    assign temp9995 = temp9994 ^ temp9994;
    assign temp9996 = temp9995 ^ temp9995;
    assign temp9997 = temp9996 ^ temp9996;
    assign temp9998 = temp9997 ^ temp9997;
    assign z = temp9998 ^ temp9998;


endmodule