module sum_gld (
  input  [2:0] a,
  input  [2:0] b,
  output [3:0] o
);


assign o = a + b;

endmodule 
