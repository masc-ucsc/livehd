module Cell(
  input   clock,
  input   reset,
  input   io_neighbors_0,
  input   io_neighbors_1,
  input   io_neighbors_2,
  input   io_neighbors_3,
  input   io_neighbors_4,
  input   io_neighbors_5,
  input   io_neighbors_6,
  input   io_neighbors_7,
  output  io_out,
  input   io_running,
  input   io_writeEnable,
  input   io_writeValue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  isAlive; // @[Life.scala 16:24]
  wire [3:0] _T_1 = {{3'd0}, io_neighbors_7}; // @[Life.scala 26:81]
  wire [2:0] _GEN_6 = {{2'd0}, io_neighbors_6}; // @[Life.scala 26:81]
  wire [2:0] _T_4 = _GEN_6 + _T_1[2:0]; // @[Life.scala 26:81]
  wire [2:0] _GEN_7 = {{2'd0}, io_neighbors_5}; // @[Life.scala 26:81]
  wire [2:0] _T_6 = _GEN_7 + _T_4; // @[Life.scala 26:81]
  wire [2:0] _GEN_8 = {{2'd0}, io_neighbors_4}; // @[Life.scala 26:81]
  wire [2:0] _T_8 = _GEN_8 + _T_6; // @[Life.scala 26:81]
  wire [2:0] _GEN_9 = {{2'd0}, io_neighbors_3}; // @[Life.scala 26:81]
  wire [2:0] _T_10 = _GEN_9 + _T_8; // @[Life.scala 26:81]
  wire [2:0] _GEN_10 = {{2'd0}, io_neighbors_2}; // @[Life.scala 26:81]
  wire [2:0] _T_12 = _GEN_10 + _T_10; // @[Life.scala 26:81]
  wire [2:0] _GEN_11 = {{2'd0}, io_neighbors_1}; // @[Life.scala 26:81]
  wire [2:0] _T_14 = _GEN_11 + _T_12; // @[Life.scala 26:81]
  wire [2:0] _GEN_12 = {{2'd0}, io_neighbors_0}; // @[Life.scala 26:81]
  wire [2:0] _T_16 = _GEN_12 + _T_14; // @[Life.scala 26:81]
  wire  _T_18 = _T_16 < 3'h4; // @[Life.scala 31:24]
  wire  _T_21 = ~isAlive & _T_16 == 3'h3; // @[Life.scala 37:21]
  assign io_out = isAlive; // @[Life.scala 46:10]
  always @(posedge clock) begin
    if (reset) begin // @[Life.scala 16:24]
      isAlive <= 1'h0; // @[Life.scala 16:24]
    end else if (~io_running) begin // @[Life.scala 18:21]
      if (io_writeEnable) begin // @[Life.scala 19:26]
        isAlive <= io_writeValue; // @[Life.scala 20:15]
      end
    end else if (isAlive) begin // @[Life.scala 28:19]
      if (_T_16 < 3'h2) begin // @[Life.scala 29:25]
        isAlive <= 1'h0; // @[Life.scala 30:17]
      end else begin
        isAlive <= _T_18;
      end
    end else begin
      isAlive <= _T_21;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isAlive = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Life(
  input        clock,
  input        reset,
  output       io_state_0_0,
  output       io_state_0_1,
  output       io_state_0_2,
  output       io_state_0_3,
  output       io_state_0_4,
  output       io_state_0_5,
  output       io_state_0_6,
  output       io_state_0_7,
  output       io_state_0_8,
  output       io_state_0_9,
  output       io_state_0_10,
  output       io_state_0_11,
  output       io_state_1_0,
  output       io_state_1_1,
  output       io_state_1_2,
  output       io_state_1_3,
  output       io_state_1_4,
  output       io_state_1_5,
  output       io_state_1_6,
  output       io_state_1_7,
  output       io_state_1_8,
  output       io_state_1_9,
  output       io_state_1_10,
  output       io_state_1_11,
  output       io_state_2_0,
  output       io_state_2_1,
  output       io_state_2_2,
  output       io_state_2_3,
  output       io_state_2_4,
  output       io_state_2_5,
  output       io_state_2_6,
  output       io_state_2_7,
  output       io_state_2_8,
  output       io_state_2_9,
  output       io_state_2_10,
  output       io_state_2_11,
  output       io_state_3_0,
  output       io_state_3_1,
  output       io_state_3_2,
  output       io_state_3_3,
  output       io_state_3_4,
  output       io_state_3_5,
  output       io_state_3_6,
  output       io_state_3_7,
  output       io_state_3_8,
  output       io_state_3_9,
  output       io_state_3_10,
  output       io_state_3_11,
  output       io_state_4_0,
  output       io_state_4_1,
  output       io_state_4_2,
  output       io_state_4_3,
  output       io_state_4_4,
  output       io_state_4_5,
  output       io_state_4_6,
  output       io_state_4_7,
  output       io_state_4_8,
  output       io_state_4_9,
  output       io_state_4_10,
  output       io_state_4_11,
  output       io_state_5_0,
  output       io_state_5_1,
  output       io_state_5_2,
  output       io_state_5_3,
  output       io_state_5_4,
  output       io_state_5_5,
  output       io_state_5_6,
  output       io_state_5_7,
  output       io_state_5_8,
  output       io_state_5_9,
  output       io_state_5_10,
  output       io_state_5_11,
  output       io_state_6_0,
  output       io_state_6_1,
  output       io_state_6_2,
  output       io_state_6_3,
  output       io_state_6_4,
  output       io_state_6_5,
  output       io_state_6_6,
  output       io_state_6_7,
  output       io_state_6_8,
  output       io_state_6_9,
  output       io_state_6_10,
  output       io_state_6_11,
  output       io_state_7_0,
  output       io_state_7_1,
  output       io_state_7_2,
  output       io_state_7_3,
  output       io_state_7_4,
  output       io_state_7_5,
  output       io_state_7_6,
  output       io_state_7_7,
  output       io_state_7_8,
  output       io_state_7_9,
  output       io_state_7_10,
  output       io_state_7_11,
  output       io_state_8_0,
  output       io_state_8_1,
  output       io_state_8_2,
  output       io_state_8_3,
  output       io_state_8_4,
  output       io_state_8_5,
  output       io_state_8_6,
  output       io_state_8_7,
  output       io_state_8_8,
  output       io_state_8_9,
  output       io_state_8_10,
  output       io_state_8_11,
  output       io_state_9_0,
  output       io_state_9_1,
  output       io_state_9_2,
  output       io_state_9_3,
  output       io_state_9_4,
  output       io_state_9_5,
  output       io_state_9_6,
  output       io_state_9_7,
  output       io_state_9_8,
  output       io_state_9_9,
  output       io_state_9_10,
  output       io_state_9_11,
  output       io_state_10_0,
  output       io_state_10_1,
  output       io_state_10_2,
  output       io_state_10_3,
  output       io_state_10_4,
  output       io_state_10_5,
  output       io_state_10_6,
  output       io_state_10_7,
  output       io_state_10_8,
  output       io_state_10_9,
  output       io_state_10_10,
  output       io_state_10_11,
  output       io_state_11_0,
  output       io_state_11_1,
  output       io_state_11_2,
  output       io_state_11_3,
  output       io_state_11_4,
  output       io_state_11_5,
  output       io_state_11_6,
  output       io_state_11_7,
  output       io_state_11_8,
  output       io_state_11_9,
  output       io_state_11_10,
  output       io_state_11_11,
  input        io_running,
  input        io_writeValue,
  input  [3:0] io_writeRowAddress,
  input  [3:0] io_writeColAddress
);
  wire  Cell_clock; // @[Life.scala 59:52]
  wire  Cell_reset; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_io_out; // @[Life.scala 59:52]
  wire  Cell_io_running; // @[Life.scala 59:52]
  wire  Cell_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_1_clock; // @[Life.scala 59:52]
  wire  Cell_1_reset; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_1_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_1_io_out; // @[Life.scala 59:52]
  wire  Cell_1_io_running; // @[Life.scala 59:52]
  wire  Cell_1_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_1_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_2_clock; // @[Life.scala 59:52]
  wire  Cell_2_reset; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_2_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_2_io_out; // @[Life.scala 59:52]
  wire  Cell_2_io_running; // @[Life.scala 59:52]
  wire  Cell_2_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_2_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_3_clock; // @[Life.scala 59:52]
  wire  Cell_3_reset; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_3_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_3_io_out; // @[Life.scala 59:52]
  wire  Cell_3_io_running; // @[Life.scala 59:52]
  wire  Cell_3_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_3_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_4_clock; // @[Life.scala 59:52]
  wire  Cell_4_reset; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_4_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_4_io_out; // @[Life.scala 59:52]
  wire  Cell_4_io_running; // @[Life.scala 59:52]
  wire  Cell_4_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_4_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_5_clock; // @[Life.scala 59:52]
  wire  Cell_5_reset; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_5_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_5_io_out; // @[Life.scala 59:52]
  wire  Cell_5_io_running; // @[Life.scala 59:52]
  wire  Cell_5_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_5_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_6_clock; // @[Life.scala 59:52]
  wire  Cell_6_reset; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_6_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_6_io_out; // @[Life.scala 59:52]
  wire  Cell_6_io_running; // @[Life.scala 59:52]
  wire  Cell_6_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_6_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_7_clock; // @[Life.scala 59:52]
  wire  Cell_7_reset; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_7_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_7_io_out; // @[Life.scala 59:52]
  wire  Cell_7_io_running; // @[Life.scala 59:52]
  wire  Cell_7_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_7_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_8_clock; // @[Life.scala 59:52]
  wire  Cell_8_reset; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_8_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_8_io_out; // @[Life.scala 59:52]
  wire  Cell_8_io_running; // @[Life.scala 59:52]
  wire  Cell_8_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_8_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_9_clock; // @[Life.scala 59:52]
  wire  Cell_9_reset; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_9_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_9_io_out; // @[Life.scala 59:52]
  wire  Cell_9_io_running; // @[Life.scala 59:52]
  wire  Cell_9_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_9_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_10_clock; // @[Life.scala 59:52]
  wire  Cell_10_reset; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_10_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_10_io_out; // @[Life.scala 59:52]
  wire  Cell_10_io_running; // @[Life.scala 59:52]
  wire  Cell_10_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_10_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_11_clock; // @[Life.scala 59:52]
  wire  Cell_11_reset; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_11_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_11_io_out; // @[Life.scala 59:52]
  wire  Cell_11_io_running; // @[Life.scala 59:52]
  wire  Cell_11_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_11_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_12_clock; // @[Life.scala 59:52]
  wire  Cell_12_reset; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_12_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_12_io_out; // @[Life.scala 59:52]
  wire  Cell_12_io_running; // @[Life.scala 59:52]
  wire  Cell_12_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_12_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_13_clock; // @[Life.scala 59:52]
  wire  Cell_13_reset; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_13_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_13_io_out; // @[Life.scala 59:52]
  wire  Cell_13_io_running; // @[Life.scala 59:52]
  wire  Cell_13_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_13_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_14_clock; // @[Life.scala 59:52]
  wire  Cell_14_reset; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_14_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_14_io_out; // @[Life.scala 59:52]
  wire  Cell_14_io_running; // @[Life.scala 59:52]
  wire  Cell_14_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_14_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_15_clock; // @[Life.scala 59:52]
  wire  Cell_15_reset; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_15_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_15_io_out; // @[Life.scala 59:52]
  wire  Cell_15_io_running; // @[Life.scala 59:52]
  wire  Cell_15_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_15_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_16_clock; // @[Life.scala 59:52]
  wire  Cell_16_reset; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_16_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_16_io_out; // @[Life.scala 59:52]
  wire  Cell_16_io_running; // @[Life.scala 59:52]
  wire  Cell_16_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_16_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_17_clock; // @[Life.scala 59:52]
  wire  Cell_17_reset; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_17_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_17_io_out; // @[Life.scala 59:52]
  wire  Cell_17_io_running; // @[Life.scala 59:52]
  wire  Cell_17_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_17_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_18_clock; // @[Life.scala 59:52]
  wire  Cell_18_reset; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_18_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_18_io_out; // @[Life.scala 59:52]
  wire  Cell_18_io_running; // @[Life.scala 59:52]
  wire  Cell_18_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_18_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_19_clock; // @[Life.scala 59:52]
  wire  Cell_19_reset; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_19_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_19_io_out; // @[Life.scala 59:52]
  wire  Cell_19_io_running; // @[Life.scala 59:52]
  wire  Cell_19_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_19_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_20_clock; // @[Life.scala 59:52]
  wire  Cell_20_reset; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_20_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_20_io_out; // @[Life.scala 59:52]
  wire  Cell_20_io_running; // @[Life.scala 59:52]
  wire  Cell_20_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_20_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_21_clock; // @[Life.scala 59:52]
  wire  Cell_21_reset; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_21_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_21_io_out; // @[Life.scala 59:52]
  wire  Cell_21_io_running; // @[Life.scala 59:52]
  wire  Cell_21_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_21_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_22_clock; // @[Life.scala 59:52]
  wire  Cell_22_reset; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_22_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_22_io_out; // @[Life.scala 59:52]
  wire  Cell_22_io_running; // @[Life.scala 59:52]
  wire  Cell_22_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_22_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_23_clock; // @[Life.scala 59:52]
  wire  Cell_23_reset; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_23_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_23_io_out; // @[Life.scala 59:52]
  wire  Cell_23_io_running; // @[Life.scala 59:52]
  wire  Cell_23_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_23_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_24_clock; // @[Life.scala 59:52]
  wire  Cell_24_reset; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_24_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_24_io_out; // @[Life.scala 59:52]
  wire  Cell_24_io_running; // @[Life.scala 59:52]
  wire  Cell_24_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_24_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_25_clock; // @[Life.scala 59:52]
  wire  Cell_25_reset; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_25_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_25_io_out; // @[Life.scala 59:52]
  wire  Cell_25_io_running; // @[Life.scala 59:52]
  wire  Cell_25_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_25_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_26_clock; // @[Life.scala 59:52]
  wire  Cell_26_reset; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_26_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_26_io_out; // @[Life.scala 59:52]
  wire  Cell_26_io_running; // @[Life.scala 59:52]
  wire  Cell_26_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_26_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_27_clock; // @[Life.scala 59:52]
  wire  Cell_27_reset; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_27_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_27_io_out; // @[Life.scala 59:52]
  wire  Cell_27_io_running; // @[Life.scala 59:52]
  wire  Cell_27_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_27_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_28_clock; // @[Life.scala 59:52]
  wire  Cell_28_reset; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_28_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_28_io_out; // @[Life.scala 59:52]
  wire  Cell_28_io_running; // @[Life.scala 59:52]
  wire  Cell_28_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_28_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_29_clock; // @[Life.scala 59:52]
  wire  Cell_29_reset; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_29_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_29_io_out; // @[Life.scala 59:52]
  wire  Cell_29_io_running; // @[Life.scala 59:52]
  wire  Cell_29_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_29_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_30_clock; // @[Life.scala 59:52]
  wire  Cell_30_reset; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_30_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_30_io_out; // @[Life.scala 59:52]
  wire  Cell_30_io_running; // @[Life.scala 59:52]
  wire  Cell_30_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_30_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_31_clock; // @[Life.scala 59:52]
  wire  Cell_31_reset; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_31_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_31_io_out; // @[Life.scala 59:52]
  wire  Cell_31_io_running; // @[Life.scala 59:52]
  wire  Cell_31_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_31_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_32_clock; // @[Life.scala 59:52]
  wire  Cell_32_reset; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_32_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_32_io_out; // @[Life.scala 59:52]
  wire  Cell_32_io_running; // @[Life.scala 59:52]
  wire  Cell_32_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_32_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_33_clock; // @[Life.scala 59:52]
  wire  Cell_33_reset; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_33_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_33_io_out; // @[Life.scala 59:52]
  wire  Cell_33_io_running; // @[Life.scala 59:52]
  wire  Cell_33_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_33_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_34_clock; // @[Life.scala 59:52]
  wire  Cell_34_reset; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_34_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_34_io_out; // @[Life.scala 59:52]
  wire  Cell_34_io_running; // @[Life.scala 59:52]
  wire  Cell_34_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_34_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_35_clock; // @[Life.scala 59:52]
  wire  Cell_35_reset; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_35_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_35_io_out; // @[Life.scala 59:52]
  wire  Cell_35_io_running; // @[Life.scala 59:52]
  wire  Cell_35_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_35_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_36_clock; // @[Life.scala 59:52]
  wire  Cell_36_reset; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_36_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_36_io_out; // @[Life.scala 59:52]
  wire  Cell_36_io_running; // @[Life.scala 59:52]
  wire  Cell_36_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_36_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_37_clock; // @[Life.scala 59:52]
  wire  Cell_37_reset; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_37_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_37_io_out; // @[Life.scala 59:52]
  wire  Cell_37_io_running; // @[Life.scala 59:52]
  wire  Cell_37_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_37_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_38_clock; // @[Life.scala 59:52]
  wire  Cell_38_reset; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_38_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_38_io_out; // @[Life.scala 59:52]
  wire  Cell_38_io_running; // @[Life.scala 59:52]
  wire  Cell_38_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_38_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_39_clock; // @[Life.scala 59:52]
  wire  Cell_39_reset; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_39_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_39_io_out; // @[Life.scala 59:52]
  wire  Cell_39_io_running; // @[Life.scala 59:52]
  wire  Cell_39_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_39_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_40_clock; // @[Life.scala 59:52]
  wire  Cell_40_reset; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_40_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_40_io_out; // @[Life.scala 59:52]
  wire  Cell_40_io_running; // @[Life.scala 59:52]
  wire  Cell_40_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_40_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_41_clock; // @[Life.scala 59:52]
  wire  Cell_41_reset; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_41_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_41_io_out; // @[Life.scala 59:52]
  wire  Cell_41_io_running; // @[Life.scala 59:52]
  wire  Cell_41_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_41_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_42_clock; // @[Life.scala 59:52]
  wire  Cell_42_reset; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_42_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_42_io_out; // @[Life.scala 59:52]
  wire  Cell_42_io_running; // @[Life.scala 59:52]
  wire  Cell_42_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_42_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_43_clock; // @[Life.scala 59:52]
  wire  Cell_43_reset; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_43_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_43_io_out; // @[Life.scala 59:52]
  wire  Cell_43_io_running; // @[Life.scala 59:52]
  wire  Cell_43_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_43_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_44_clock; // @[Life.scala 59:52]
  wire  Cell_44_reset; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_44_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_44_io_out; // @[Life.scala 59:52]
  wire  Cell_44_io_running; // @[Life.scala 59:52]
  wire  Cell_44_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_44_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_45_clock; // @[Life.scala 59:52]
  wire  Cell_45_reset; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_45_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_45_io_out; // @[Life.scala 59:52]
  wire  Cell_45_io_running; // @[Life.scala 59:52]
  wire  Cell_45_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_45_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_46_clock; // @[Life.scala 59:52]
  wire  Cell_46_reset; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_46_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_46_io_out; // @[Life.scala 59:52]
  wire  Cell_46_io_running; // @[Life.scala 59:52]
  wire  Cell_46_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_46_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_47_clock; // @[Life.scala 59:52]
  wire  Cell_47_reset; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_47_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_47_io_out; // @[Life.scala 59:52]
  wire  Cell_47_io_running; // @[Life.scala 59:52]
  wire  Cell_47_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_47_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_48_clock; // @[Life.scala 59:52]
  wire  Cell_48_reset; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_48_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_48_io_out; // @[Life.scala 59:52]
  wire  Cell_48_io_running; // @[Life.scala 59:52]
  wire  Cell_48_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_48_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_49_clock; // @[Life.scala 59:52]
  wire  Cell_49_reset; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_49_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_49_io_out; // @[Life.scala 59:52]
  wire  Cell_49_io_running; // @[Life.scala 59:52]
  wire  Cell_49_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_49_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_50_clock; // @[Life.scala 59:52]
  wire  Cell_50_reset; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_50_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_50_io_out; // @[Life.scala 59:52]
  wire  Cell_50_io_running; // @[Life.scala 59:52]
  wire  Cell_50_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_50_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_51_clock; // @[Life.scala 59:52]
  wire  Cell_51_reset; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_51_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_51_io_out; // @[Life.scala 59:52]
  wire  Cell_51_io_running; // @[Life.scala 59:52]
  wire  Cell_51_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_51_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_52_clock; // @[Life.scala 59:52]
  wire  Cell_52_reset; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_52_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_52_io_out; // @[Life.scala 59:52]
  wire  Cell_52_io_running; // @[Life.scala 59:52]
  wire  Cell_52_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_52_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_53_clock; // @[Life.scala 59:52]
  wire  Cell_53_reset; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_53_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_53_io_out; // @[Life.scala 59:52]
  wire  Cell_53_io_running; // @[Life.scala 59:52]
  wire  Cell_53_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_53_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_54_clock; // @[Life.scala 59:52]
  wire  Cell_54_reset; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_54_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_54_io_out; // @[Life.scala 59:52]
  wire  Cell_54_io_running; // @[Life.scala 59:52]
  wire  Cell_54_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_54_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_55_clock; // @[Life.scala 59:52]
  wire  Cell_55_reset; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_55_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_55_io_out; // @[Life.scala 59:52]
  wire  Cell_55_io_running; // @[Life.scala 59:52]
  wire  Cell_55_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_55_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_56_clock; // @[Life.scala 59:52]
  wire  Cell_56_reset; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_56_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_56_io_out; // @[Life.scala 59:52]
  wire  Cell_56_io_running; // @[Life.scala 59:52]
  wire  Cell_56_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_56_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_57_clock; // @[Life.scala 59:52]
  wire  Cell_57_reset; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_57_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_57_io_out; // @[Life.scala 59:52]
  wire  Cell_57_io_running; // @[Life.scala 59:52]
  wire  Cell_57_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_57_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_58_clock; // @[Life.scala 59:52]
  wire  Cell_58_reset; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_58_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_58_io_out; // @[Life.scala 59:52]
  wire  Cell_58_io_running; // @[Life.scala 59:52]
  wire  Cell_58_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_58_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_59_clock; // @[Life.scala 59:52]
  wire  Cell_59_reset; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_59_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_59_io_out; // @[Life.scala 59:52]
  wire  Cell_59_io_running; // @[Life.scala 59:52]
  wire  Cell_59_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_59_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_60_clock; // @[Life.scala 59:52]
  wire  Cell_60_reset; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_60_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_60_io_out; // @[Life.scala 59:52]
  wire  Cell_60_io_running; // @[Life.scala 59:52]
  wire  Cell_60_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_60_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_61_clock; // @[Life.scala 59:52]
  wire  Cell_61_reset; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_61_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_61_io_out; // @[Life.scala 59:52]
  wire  Cell_61_io_running; // @[Life.scala 59:52]
  wire  Cell_61_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_61_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_62_clock; // @[Life.scala 59:52]
  wire  Cell_62_reset; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_62_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_62_io_out; // @[Life.scala 59:52]
  wire  Cell_62_io_running; // @[Life.scala 59:52]
  wire  Cell_62_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_62_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_63_clock; // @[Life.scala 59:52]
  wire  Cell_63_reset; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_63_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_63_io_out; // @[Life.scala 59:52]
  wire  Cell_63_io_running; // @[Life.scala 59:52]
  wire  Cell_63_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_63_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_64_clock; // @[Life.scala 59:52]
  wire  Cell_64_reset; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_64_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_64_io_out; // @[Life.scala 59:52]
  wire  Cell_64_io_running; // @[Life.scala 59:52]
  wire  Cell_64_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_64_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_65_clock; // @[Life.scala 59:52]
  wire  Cell_65_reset; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_65_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_65_io_out; // @[Life.scala 59:52]
  wire  Cell_65_io_running; // @[Life.scala 59:52]
  wire  Cell_65_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_65_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_66_clock; // @[Life.scala 59:52]
  wire  Cell_66_reset; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_66_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_66_io_out; // @[Life.scala 59:52]
  wire  Cell_66_io_running; // @[Life.scala 59:52]
  wire  Cell_66_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_66_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_67_clock; // @[Life.scala 59:52]
  wire  Cell_67_reset; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_67_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_67_io_out; // @[Life.scala 59:52]
  wire  Cell_67_io_running; // @[Life.scala 59:52]
  wire  Cell_67_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_67_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_68_clock; // @[Life.scala 59:52]
  wire  Cell_68_reset; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_68_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_68_io_out; // @[Life.scala 59:52]
  wire  Cell_68_io_running; // @[Life.scala 59:52]
  wire  Cell_68_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_68_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_69_clock; // @[Life.scala 59:52]
  wire  Cell_69_reset; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_69_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_69_io_out; // @[Life.scala 59:52]
  wire  Cell_69_io_running; // @[Life.scala 59:52]
  wire  Cell_69_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_69_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_70_clock; // @[Life.scala 59:52]
  wire  Cell_70_reset; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_70_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_70_io_out; // @[Life.scala 59:52]
  wire  Cell_70_io_running; // @[Life.scala 59:52]
  wire  Cell_70_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_70_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_71_clock; // @[Life.scala 59:52]
  wire  Cell_71_reset; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_71_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_71_io_out; // @[Life.scala 59:52]
  wire  Cell_71_io_running; // @[Life.scala 59:52]
  wire  Cell_71_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_71_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_72_clock; // @[Life.scala 59:52]
  wire  Cell_72_reset; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_72_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_72_io_out; // @[Life.scala 59:52]
  wire  Cell_72_io_running; // @[Life.scala 59:52]
  wire  Cell_72_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_72_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_73_clock; // @[Life.scala 59:52]
  wire  Cell_73_reset; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_73_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_73_io_out; // @[Life.scala 59:52]
  wire  Cell_73_io_running; // @[Life.scala 59:52]
  wire  Cell_73_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_73_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_74_clock; // @[Life.scala 59:52]
  wire  Cell_74_reset; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_74_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_74_io_out; // @[Life.scala 59:52]
  wire  Cell_74_io_running; // @[Life.scala 59:52]
  wire  Cell_74_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_74_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_75_clock; // @[Life.scala 59:52]
  wire  Cell_75_reset; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_75_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_75_io_out; // @[Life.scala 59:52]
  wire  Cell_75_io_running; // @[Life.scala 59:52]
  wire  Cell_75_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_75_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_76_clock; // @[Life.scala 59:52]
  wire  Cell_76_reset; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_76_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_76_io_out; // @[Life.scala 59:52]
  wire  Cell_76_io_running; // @[Life.scala 59:52]
  wire  Cell_76_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_76_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_77_clock; // @[Life.scala 59:52]
  wire  Cell_77_reset; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_77_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_77_io_out; // @[Life.scala 59:52]
  wire  Cell_77_io_running; // @[Life.scala 59:52]
  wire  Cell_77_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_77_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_78_clock; // @[Life.scala 59:52]
  wire  Cell_78_reset; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_78_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_78_io_out; // @[Life.scala 59:52]
  wire  Cell_78_io_running; // @[Life.scala 59:52]
  wire  Cell_78_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_78_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_79_clock; // @[Life.scala 59:52]
  wire  Cell_79_reset; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_79_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_79_io_out; // @[Life.scala 59:52]
  wire  Cell_79_io_running; // @[Life.scala 59:52]
  wire  Cell_79_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_79_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_80_clock; // @[Life.scala 59:52]
  wire  Cell_80_reset; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_80_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_80_io_out; // @[Life.scala 59:52]
  wire  Cell_80_io_running; // @[Life.scala 59:52]
  wire  Cell_80_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_80_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_81_clock; // @[Life.scala 59:52]
  wire  Cell_81_reset; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_81_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_81_io_out; // @[Life.scala 59:52]
  wire  Cell_81_io_running; // @[Life.scala 59:52]
  wire  Cell_81_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_81_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_82_clock; // @[Life.scala 59:52]
  wire  Cell_82_reset; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_82_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_82_io_out; // @[Life.scala 59:52]
  wire  Cell_82_io_running; // @[Life.scala 59:52]
  wire  Cell_82_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_82_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_83_clock; // @[Life.scala 59:52]
  wire  Cell_83_reset; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_83_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_83_io_out; // @[Life.scala 59:52]
  wire  Cell_83_io_running; // @[Life.scala 59:52]
  wire  Cell_83_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_83_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_84_clock; // @[Life.scala 59:52]
  wire  Cell_84_reset; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_84_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_84_io_out; // @[Life.scala 59:52]
  wire  Cell_84_io_running; // @[Life.scala 59:52]
  wire  Cell_84_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_84_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_85_clock; // @[Life.scala 59:52]
  wire  Cell_85_reset; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_85_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_85_io_out; // @[Life.scala 59:52]
  wire  Cell_85_io_running; // @[Life.scala 59:52]
  wire  Cell_85_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_85_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_86_clock; // @[Life.scala 59:52]
  wire  Cell_86_reset; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_86_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_86_io_out; // @[Life.scala 59:52]
  wire  Cell_86_io_running; // @[Life.scala 59:52]
  wire  Cell_86_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_86_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_87_clock; // @[Life.scala 59:52]
  wire  Cell_87_reset; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_87_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_87_io_out; // @[Life.scala 59:52]
  wire  Cell_87_io_running; // @[Life.scala 59:52]
  wire  Cell_87_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_87_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_88_clock; // @[Life.scala 59:52]
  wire  Cell_88_reset; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_88_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_88_io_out; // @[Life.scala 59:52]
  wire  Cell_88_io_running; // @[Life.scala 59:52]
  wire  Cell_88_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_88_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_89_clock; // @[Life.scala 59:52]
  wire  Cell_89_reset; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_89_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_89_io_out; // @[Life.scala 59:52]
  wire  Cell_89_io_running; // @[Life.scala 59:52]
  wire  Cell_89_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_89_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_90_clock; // @[Life.scala 59:52]
  wire  Cell_90_reset; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_90_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_90_io_out; // @[Life.scala 59:52]
  wire  Cell_90_io_running; // @[Life.scala 59:52]
  wire  Cell_90_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_90_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_91_clock; // @[Life.scala 59:52]
  wire  Cell_91_reset; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_91_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_91_io_out; // @[Life.scala 59:52]
  wire  Cell_91_io_running; // @[Life.scala 59:52]
  wire  Cell_91_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_91_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_92_clock; // @[Life.scala 59:52]
  wire  Cell_92_reset; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_92_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_92_io_out; // @[Life.scala 59:52]
  wire  Cell_92_io_running; // @[Life.scala 59:52]
  wire  Cell_92_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_92_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_93_clock; // @[Life.scala 59:52]
  wire  Cell_93_reset; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_93_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_93_io_out; // @[Life.scala 59:52]
  wire  Cell_93_io_running; // @[Life.scala 59:52]
  wire  Cell_93_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_93_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_94_clock; // @[Life.scala 59:52]
  wire  Cell_94_reset; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_94_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_94_io_out; // @[Life.scala 59:52]
  wire  Cell_94_io_running; // @[Life.scala 59:52]
  wire  Cell_94_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_94_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_95_clock; // @[Life.scala 59:52]
  wire  Cell_95_reset; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_95_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_95_io_out; // @[Life.scala 59:52]
  wire  Cell_95_io_running; // @[Life.scala 59:52]
  wire  Cell_95_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_95_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_96_clock; // @[Life.scala 59:52]
  wire  Cell_96_reset; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_96_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_96_io_out; // @[Life.scala 59:52]
  wire  Cell_96_io_running; // @[Life.scala 59:52]
  wire  Cell_96_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_96_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_97_clock; // @[Life.scala 59:52]
  wire  Cell_97_reset; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_97_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_97_io_out; // @[Life.scala 59:52]
  wire  Cell_97_io_running; // @[Life.scala 59:52]
  wire  Cell_97_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_97_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_98_clock; // @[Life.scala 59:52]
  wire  Cell_98_reset; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_98_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_98_io_out; // @[Life.scala 59:52]
  wire  Cell_98_io_running; // @[Life.scala 59:52]
  wire  Cell_98_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_98_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_99_clock; // @[Life.scala 59:52]
  wire  Cell_99_reset; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_99_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_99_io_out; // @[Life.scala 59:52]
  wire  Cell_99_io_running; // @[Life.scala 59:52]
  wire  Cell_99_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_99_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_100_clock; // @[Life.scala 59:52]
  wire  Cell_100_reset; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_100_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_100_io_out; // @[Life.scala 59:52]
  wire  Cell_100_io_running; // @[Life.scala 59:52]
  wire  Cell_100_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_100_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_101_clock; // @[Life.scala 59:52]
  wire  Cell_101_reset; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_101_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_101_io_out; // @[Life.scala 59:52]
  wire  Cell_101_io_running; // @[Life.scala 59:52]
  wire  Cell_101_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_101_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_102_clock; // @[Life.scala 59:52]
  wire  Cell_102_reset; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_102_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_102_io_out; // @[Life.scala 59:52]
  wire  Cell_102_io_running; // @[Life.scala 59:52]
  wire  Cell_102_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_102_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_103_clock; // @[Life.scala 59:52]
  wire  Cell_103_reset; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_103_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_103_io_out; // @[Life.scala 59:52]
  wire  Cell_103_io_running; // @[Life.scala 59:52]
  wire  Cell_103_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_103_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_104_clock; // @[Life.scala 59:52]
  wire  Cell_104_reset; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_104_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_104_io_out; // @[Life.scala 59:52]
  wire  Cell_104_io_running; // @[Life.scala 59:52]
  wire  Cell_104_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_104_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_105_clock; // @[Life.scala 59:52]
  wire  Cell_105_reset; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_105_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_105_io_out; // @[Life.scala 59:52]
  wire  Cell_105_io_running; // @[Life.scala 59:52]
  wire  Cell_105_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_105_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_106_clock; // @[Life.scala 59:52]
  wire  Cell_106_reset; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_106_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_106_io_out; // @[Life.scala 59:52]
  wire  Cell_106_io_running; // @[Life.scala 59:52]
  wire  Cell_106_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_106_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_107_clock; // @[Life.scala 59:52]
  wire  Cell_107_reset; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_107_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_107_io_out; // @[Life.scala 59:52]
  wire  Cell_107_io_running; // @[Life.scala 59:52]
  wire  Cell_107_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_107_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_108_clock; // @[Life.scala 59:52]
  wire  Cell_108_reset; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_108_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_108_io_out; // @[Life.scala 59:52]
  wire  Cell_108_io_running; // @[Life.scala 59:52]
  wire  Cell_108_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_108_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_109_clock; // @[Life.scala 59:52]
  wire  Cell_109_reset; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_109_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_109_io_out; // @[Life.scala 59:52]
  wire  Cell_109_io_running; // @[Life.scala 59:52]
  wire  Cell_109_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_109_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_110_clock; // @[Life.scala 59:52]
  wire  Cell_110_reset; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_110_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_110_io_out; // @[Life.scala 59:52]
  wire  Cell_110_io_running; // @[Life.scala 59:52]
  wire  Cell_110_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_110_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_111_clock; // @[Life.scala 59:52]
  wire  Cell_111_reset; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_111_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_111_io_out; // @[Life.scala 59:52]
  wire  Cell_111_io_running; // @[Life.scala 59:52]
  wire  Cell_111_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_111_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_112_clock; // @[Life.scala 59:52]
  wire  Cell_112_reset; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_112_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_112_io_out; // @[Life.scala 59:52]
  wire  Cell_112_io_running; // @[Life.scala 59:52]
  wire  Cell_112_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_112_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_113_clock; // @[Life.scala 59:52]
  wire  Cell_113_reset; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_113_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_113_io_out; // @[Life.scala 59:52]
  wire  Cell_113_io_running; // @[Life.scala 59:52]
  wire  Cell_113_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_113_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_114_clock; // @[Life.scala 59:52]
  wire  Cell_114_reset; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_114_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_114_io_out; // @[Life.scala 59:52]
  wire  Cell_114_io_running; // @[Life.scala 59:52]
  wire  Cell_114_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_114_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_115_clock; // @[Life.scala 59:52]
  wire  Cell_115_reset; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_115_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_115_io_out; // @[Life.scala 59:52]
  wire  Cell_115_io_running; // @[Life.scala 59:52]
  wire  Cell_115_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_115_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_116_clock; // @[Life.scala 59:52]
  wire  Cell_116_reset; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_116_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_116_io_out; // @[Life.scala 59:52]
  wire  Cell_116_io_running; // @[Life.scala 59:52]
  wire  Cell_116_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_116_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_117_clock; // @[Life.scala 59:52]
  wire  Cell_117_reset; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_117_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_117_io_out; // @[Life.scala 59:52]
  wire  Cell_117_io_running; // @[Life.scala 59:52]
  wire  Cell_117_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_117_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_118_clock; // @[Life.scala 59:52]
  wire  Cell_118_reset; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_118_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_118_io_out; // @[Life.scala 59:52]
  wire  Cell_118_io_running; // @[Life.scala 59:52]
  wire  Cell_118_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_118_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_119_clock; // @[Life.scala 59:52]
  wire  Cell_119_reset; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_119_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_119_io_out; // @[Life.scala 59:52]
  wire  Cell_119_io_running; // @[Life.scala 59:52]
  wire  Cell_119_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_119_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_120_clock; // @[Life.scala 59:52]
  wire  Cell_120_reset; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_120_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_120_io_out; // @[Life.scala 59:52]
  wire  Cell_120_io_running; // @[Life.scala 59:52]
  wire  Cell_120_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_120_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_121_clock; // @[Life.scala 59:52]
  wire  Cell_121_reset; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_121_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_121_io_out; // @[Life.scala 59:52]
  wire  Cell_121_io_running; // @[Life.scala 59:52]
  wire  Cell_121_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_121_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_122_clock; // @[Life.scala 59:52]
  wire  Cell_122_reset; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_122_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_122_io_out; // @[Life.scala 59:52]
  wire  Cell_122_io_running; // @[Life.scala 59:52]
  wire  Cell_122_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_122_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_123_clock; // @[Life.scala 59:52]
  wire  Cell_123_reset; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_123_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_123_io_out; // @[Life.scala 59:52]
  wire  Cell_123_io_running; // @[Life.scala 59:52]
  wire  Cell_123_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_123_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_124_clock; // @[Life.scala 59:52]
  wire  Cell_124_reset; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_124_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_124_io_out; // @[Life.scala 59:52]
  wire  Cell_124_io_running; // @[Life.scala 59:52]
  wire  Cell_124_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_124_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_125_clock; // @[Life.scala 59:52]
  wire  Cell_125_reset; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_125_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_125_io_out; // @[Life.scala 59:52]
  wire  Cell_125_io_running; // @[Life.scala 59:52]
  wire  Cell_125_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_125_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_126_clock; // @[Life.scala 59:52]
  wire  Cell_126_reset; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_126_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_126_io_out; // @[Life.scala 59:52]
  wire  Cell_126_io_running; // @[Life.scala 59:52]
  wire  Cell_126_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_126_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_127_clock; // @[Life.scala 59:52]
  wire  Cell_127_reset; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_127_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_127_io_out; // @[Life.scala 59:52]
  wire  Cell_127_io_running; // @[Life.scala 59:52]
  wire  Cell_127_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_127_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_128_clock; // @[Life.scala 59:52]
  wire  Cell_128_reset; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_128_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_128_io_out; // @[Life.scala 59:52]
  wire  Cell_128_io_running; // @[Life.scala 59:52]
  wire  Cell_128_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_128_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_129_clock; // @[Life.scala 59:52]
  wire  Cell_129_reset; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_129_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_129_io_out; // @[Life.scala 59:52]
  wire  Cell_129_io_running; // @[Life.scala 59:52]
  wire  Cell_129_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_129_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_130_clock; // @[Life.scala 59:52]
  wire  Cell_130_reset; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_130_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_130_io_out; // @[Life.scala 59:52]
  wire  Cell_130_io_running; // @[Life.scala 59:52]
  wire  Cell_130_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_130_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_131_clock; // @[Life.scala 59:52]
  wire  Cell_131_reset; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_131_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_131_io_out; // @[Life.scala 59:52]
  wire  Cell_131_io_running; // @[Life.scala 59:52]
  wire  Cell_131_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_131_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_132_clock; // @[Life.scala 59:52]
  wire  Cell_132_reset; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_132_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_132_io_out; // @[Life.scala 59:52]
  wire  Cell_132_io_running; // @[Life.scala 59:52]
  wire  Cell_132_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_132_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_133_clock; // @[Life.scala 59:52]
  wire  Cell_133_reset; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_133_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_133_io_out; // @[Life.scala 59:52]
  wire  Cell_133_io_running; // @[Life.scala 59:52]
  wire  Cell_133_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_133_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_134_clock; // @[Life.scala 59:52]
  wire  Cell_134_reset; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_134_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_134_io_out; // @[Life.scala 59:52]
  wire  Cell_134_io_running; // @[Life.scala 59:52]
  wire  Cell_134_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_134_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_135_clock; // @[Life.scala 59:52]
  wire  Cell_135_reset; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_135_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_135_io_out; // @[Life.scala 59:52]
  wire  Cell_135_io_running; // @[Life.scala 59:52]
  wire  Cell_135_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_135_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_136_clock; // @[Life.scala 59:52]
  wire  Cell_136_reset; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_136_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_136_io_out; // @[Life.scala 59:52]
  wire  Cell_136_io_running; // @[Life.scala 59:52]
  wire  Cell_136_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_136_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_137_clock; // @[Life.scala 59:52]
  wire  Cell_137_reset; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_137_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_137_io_out; // @[Life.scala 59:52]
  wire  Cell_137_io_running; // @[Life.scala 59:52]
  wire  Cell_137_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_137_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_138_clock; // @[Life.scala 59:52]
  wire  Cell_138_reset; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_138_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_138_io_out; // @[Life.scala 59:52]
  wire  Cell_138_io_running; // @[Life.scala 59:52]
  wire  Cell_138_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_138_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_139_clock; // @[Life.scala 59:52]
  wire  Cell_139_reset; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_139_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_139_io_out; // @[Life.scala 59:52]
  wire  Cell_139_io_running; // @[Life.scala 59:52]
  wire  Cell_139_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_139_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_140_clock; // @[Life.scala 59:52]
  wire  Cell_140_reset; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_140_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_140_io_out; // @[Life.scala 59:52]
  wire  Cell_140_io_running; // @[Life.scala 59:52]
  wire  Cell_140_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_140_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_141_clock; // @[Life.scala 59:52]
  wire  Cell_141_reset; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_141_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_141_io_out; // @[Life.scala 59:52]
  wire  Cell_141_io_running; // @[Life.scala 59:52]
  wire  Cell_141_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_141_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_142_clock; // @[Life.scala 59:52]
  wire  Cell_142_reset; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_142_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_142_io_out; // @[Life.scala 59:52]
  wire  Cell_142_io_running; // @[Life.scala 59:52]
  wire  Cell_142_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_142_io_writeValue; // @[Life.scala 59:52]
  wire  Cell_143_clock; // @[Life.scala 59:52]
  wire  Cell_143_reset; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_0; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_1; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_2; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_3; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_4; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_5; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_6; // @[Life.scala 59:52]
  wire  Cell_143_io_neighbors_7; // @[Life.scala 59:52]
  wire  Cell_143_io_out; // @[Life.scala 59:52]
  wire  Cell_143_io_running; // @[Life.scala 59:52]
  wire  Cell_143_io_writeEnable; // @[Life.scala 59:52]
  wire  Cell_143_io_writeValue; // @[Life.scala 59:52]
  Cell Cell ( // @[Life.scala 59:52]
    .clock(Cell_clock),
    .reset(Cell_reset),
    .io_neighbors_0(Cell_io_neighbors_0),
    .io_neighbors_1(Cell_io_neighbors_1),
    .io_neighbors_2(Cell_io_neighbors_2),
    .io_neighbors_3(Cell_io_neighbors_3),
    .io_neighbors_4(Cell_io_neighbors_4),
    .io_neighbors_5(Cell_io_neighbors_5),
    .io_neighbors_6(Cell_io_neighbors_6),
    .io_neighbors_7(Cell_io_neighbors_7),
    .io_out(Cell_io_out),
    .io_running(Cell_io_running),
    .io_writeEnable(Cell_io_writeEnable),
    .io_writeValue(Cell_io_writeValue)
  );
  Cell Cell_1 ( // @[Life.scala 59:52]
    .clock(Cell_1_clock),
    .reset(Cell_1_reset),
    .io_neighbors_0(Cell_1_io_neighbors_0),
    .io_neighbors_1(Cell_1_io_neighbors_1),
    .io_neighbors_2(Cell_1_io_neighbors_2),
    .io_neighbors_3(Cell_1_io_neighbors_3),
    .io_neighbors_4(Cell_1_io_neighbors_4),
    .io_neighbors_5(Cell_1_io_neighbors_5),
    .io_neighbors_6(Cell_1_io_neighbors_6),
    .io_neighbors_7(Cell_1_io_neighbors_7),
    .io_out(Cell_1_io_out),
    .io_running(Cell_1_io_running),
    .io_writeEnable(Cell_1_io_writeEnable),
    .io_writeValue(Cell_1_io_writeValue)
  );
  Cell Cell_2 ( // @[Life.scala 59:52]
    .clock(Cell_2_clock),
    .reset(Cell_2_reset),
    .io_neighbors_0(Cell_2_io_neighbors_0),
    .io_neighbors_1(Cell_2_io_neighbors_1),
    .io_neighbors_2(Cell_2_io_neighbors_2),
    .io_neighbors_3(Cell_2_io_neighbors_3),
    .io_neighbors_4(Cell_2_io_neighbors_4),
    .io_neighbors_5(Cell_2_io_neighbors_5),
    .io_neighbors_6(Cell_2_io_neighbors_6),
    .io_neighbors_7(Cell_2_io_neighbors_7),
    .io_out(Cell_2_io_out),
    .io_running(Cell_2_io_running),
    .io_writeEnable(Cell_2_io_writeEnable),
    .io_writeValue(Cell_2_io_writeValue)
  );
  Cell Cell_3 ( // @[Life.scala 59:52]
    .clock(Cell_3_clock),
    .reset(Cell_3_reset),
    .io_neighbors_0(Cell_3_io_neighbors_0),
    .io_neighbors_1(Cell_3_io_neighbors_1),
    .io_neighbors_2(Cell_3_io_neighbors_2),
    .io_neighbors_3(Cell_3_io_neighbors_3),
    .io_neighbors_4(Cell_3_io_neighbors_4),
    .io_neighbors_5(Cell_3_io_neighbors_5),
    .io_neighbors_6(Cell_3_io_neighbors_6),
    .io_neighbors_7(Cell_3_io_neighbors_7),
    .io_out(Cell_3_io_out),
    .io_running(Cell_3_io_running),
    .io_writeEnable(Cell_3_io_writeEnable),
    .io_writeValue(Cell_3_io_writeValue)
  );
  Cell Cell_4 ( // @[Life.scala 59:52]
    .clock(Cell_4_clock),
    .reset(Cell_4_reset),
    .io_neighbors_0(Cell_4_io_neighbors_0),
    .io_neighbors_1(Cell_4_io_neighbors_1),
    .io_neighbors_2(Cell_4_io_neighbors_2),
    .io_neighbors_3(Cell_4_io_neighbors_3),
    .io_neighbors_4(Cell_4_io_neighbors_4),
    .io_neighbors_5(Cell_4_io_neighbors_5),
    .io_neighbors_6(Cell_4_io_neighbors_6),
    .io_neighbors_7(Cell_4_io_neighbors_7),
    .io_out(Cell_4_io_out),
    .io_running(Cell_4_io_running),
    .io_writeEnable(Cell_4_io_writeEnable),
    .io_writeValue(Cell_4_io_writeValue)
  );
  Cell Cell_5 ( // @[Life.scala 59:52]
    .clock(Cell_5_clock),
    .reset(Cell_5_reset),
    .io_neighbors_0(Cell_5_io_neighbors_0),
    .io_neighbors_1(Cell_5_io_neighbors_1),
    .io_neighbors_2(Cell_5_io_neighbors_2),
    .io_neighbors_3(Cell_5_io_neighbors_3),
    .io_neighbors_4(Cell_5_io_neighbors_4),
    .io_neighbors_5(Cell_5_io_neighbors_5),
    .io_neighbors_6(Cell_5_io_neighbors_6),
    .io_neighbors_7(Cell_5_io_neighbors_7),
    .io_out(Cell_5_io_out),
    .io_running(Cell_5_io_running),
    .io_writeEnable(Cell_5_io_writeEnable),
    .io_writeValue(Cell_5_io_writeValue)
  );
  Cell Cell_6 ( // @[Life.scala 59:52]
    .clock(Cell_6_clock),
    .reset(Cell_6_reset),
    .io_neighbors_0(Cell_6_io_neighbors_0),
    .io_neighbors_1(Cell_6_io_neighbors_1),
    .io_neighbors_2(Cell_6_io_neighbors_2),
    .io_neighbors_3(Cell_6_io_neighbors_3),
    .io_neighbors_4(Cell_6_io_neighbors_4),
    .io_neighbors_5(Cell_6_io_neighbors_5),
    .io_neighbors_6(Cell_6_io_neighbors_6),
    .io_neighbors_7(Cell_6_io_neighbors_7),
    .io_out(Cell_6_io_out),
    .io_running(Cell_6_io_running),
    .io_writeEnable(Cell_6_io_writeEnable),
    .io_writeValue(Cell_6_io_writeValue)
  );
  Cell Cell_7 ( // @[Life.scala 59:52]
    .clock(Cell_7_clock),
    .reset(Cell_7_reset),
    .io_neighbors_0(Cell_7_io_neighbors_0),
    .io_neighbors_1(Cell_7_io_neighbors_1),
    .io_neighbors_2(Cell_7_io_neighbors_2),
    .io_neighbors_3(Cell_7_io_neighbors_3),
    .io_neighbors_4(Cell_7_io_neighbors_4),
    .io_neighbors_5(Cell_7_io_neighbors_5),
    .io_neighbors_6(Cell_7_io_neighbors_6),
    .io_neighbors_7(Cell_7_io_neighbors_7),
    .io_out(Cell_7_io_out),
    .io_running(Cell_7_io_running),
    .io_writeEnable(Cell_7_io_writeEnable),
    .io_writeValue(Cell_7_io_writeValue)
  );
  Cell Cell_8 ( // @[Life.scala 59:52]
    .clock(Cell_8_clock),
    .reset(Cell_8_reset),
    .io_neighbors_0(Cell_8_io_neighbors_0),
    .io_neighbors_1(Cell_8_io_neighbors_1),
    .io_neighbors_2(Cell_8_io_neighbors_2),
    .io_neighbors_3(Cell_8_io_neighbors_3),
    .io_neighbors_4(Cell_8_io_neighbors_4),
    .io_neighbors_5(Cell_8_io_neighbors_5),
    .io_neighbors_6(Cell_8_io_neighbors_6),
    .io_neighbors_7(Cell_8_io_neighbors_7),
    .io_out(Cell_8_io_out),
    .io_running(Cell_8_io_running),
    .io_writeEnable(Cell_8_io_writeEnable),
    .io_writeValue(Cell_8_io_writeValue)
  );
  Cell Cell_9 ( // @[Life.scala 59:52]
    .clock(Cell_9_clock),
    .reset(Cell_9_reset),
    .io_neighbors_0(Cell_9_io_neighbors_0),
    .io_neighbors_1(Cell_9_io_neighbors_1),
    .io_neighbors_2(Cell_9_io_neighbors_2),
    .io_neighbors_3(Cell_9_io_neighbors_3),
    .io_neighbors_4(Cell_9_io_neighbors_4),
    .io_neighbors_5(Cell_9_io_neighbors_5),
    .io_neighbors_6(Cell_9_io_neighbors_6),
    .io_neighbors_7(Cell_9_io_neighbors_7),
    .io_out(Cell_9_io_out),
    .io_running(Cell_9_io_running),
    .io_writeEnable(Cell_9_io_writeEnable),
    .io_writeValue(Cell_9_io_writeValue)
  );
  Cell Cell_10 ( // @[Life.scala 59:52]
    .clock(Cell_10_clock),
    .reset(Cell_10_reset),
    .io_neighbors_0(Cell_10_io_neighbors_0),
    .io_neighbors_1(Cell_10_io_neighbors_1),
    .io_neighbors_2(Cell_10_io_neighbors_2),
    .io_neighbors_3(Cell_10_io_neighbors_3),
    .io_neighbors_4(Cell_10_io_neighbors_4),
    .io_neighbors_5(Cell_10_io_neighbors_5),
    .io_neighbors_6(Cell_10_io_neighbors_6),
    .io_neighbors_7(Cell_10_io_neighbors_7),
    .io_out(Cell_10_io_out),
    .io_running(Cell_10_io_running),
    .io_writeEnable(Cell_10_io_writeEnable),
    .io_writeValue(Cell_10_io_writeValue)
  );
  Cell Cell_11 ( // @[Life.scala 59:52]
    .clock(Cell_11_clock),
    .reset(Cell_11_reset),
    .io_neighbors_0(Cell_11_io_neighbors_0),
    .io_neighbors_1(Cell_11_io_neighbors_1),
    .io_neighbors_2(Cell_11_io_neighbors_2),
    .io_neighbors_3(Cell_11_io_neighbors_3),
    .io_neighbors_4(Cell_11_io_neighbors_4),
    .io_neighbors_5(Cell_11_io_neighbors_5),
    .io_neighbors_6(Cell_11_io_neighbors_6),
    .io_neighbors_7(Cell_11_io_neighbors_7),
    .io_out(Cell_11_io_out),
    .io_running(Cell_11_io_running),
    .io_writeEnable(Cell_11_io_writeEnable),
    .io_writeValue(Cell_11_io_writeValue)
  );
  Cell Cell_12 ( // @[Life.scala 59:52]
    .clock(Cell_12_clock),
    .reset(Cell_12_reset),
    .io_neighbors_0(Cell_12_io_neighbors_0),
    .io_neighbors_1(Cell_12_io_neighbors_1),
    .io_neighbors_2(Cell_12_io_neighbors_2),
    .io_neighbors_3(Cell_12_io_neighbors_3),
    .io_neighbors_4(Cell_12_io_neighbors_4),
    .io_neighbors_5(Cell_12_io_neighbors_5),
    .io_neighbors_6(Cell_12_io_neighbors_6),
    .io_neighbors_7(Cell_12_io_neighbors_7),
    .io_out(Cell_12_io_out),
    .io_running(Cell_12_io_running),
    .io_writeEnable(Cell_12_io_writeEnable),
    .io_writeValue(Cell_12_io_writeValue)
  );
  Cell Cell_13 ( // @[Life.scala 59:52]
    .clock(Cell_13_clock),
    .reset(Cell_13_reset),
    .io_neighbors_0(Cell_13_io_neighbors_0),
    .io_neighbors_1(Cell_13_io_neighbors_1),
    .io_neighbors_2(Cell_13_io_neighbors_2),
    .io_neighbors_3(Cell_13_io_neighbors_3),
    .io_neighbors_4(Cell_13_io_neighbors_4),
    .io_neighbors_5(Cell_13_io_neighbors_5),
    .io_neighbors_6(Cell_13_io_neighbors_6),
    .io_neighbors_7(Cell_13_io_neighbors_7),
    .io_out(Cell_13_io_out),
    .io_running(Cell_13_io_running),
    .io_writeEnable(Cell_13_io_writeEnable),
    .io_writeValue(Cell_13_io_writeValue)
  );
  Cell Cell_14 ( // @[Life.scala 59:52]
    .clock(Cell_14_clock),
    .reset(Cell_14_reset),
    .io_neighbors_0(Cell_14_io_neighbors_0),
    .io_neighbors_1(Cell_14_io_neighbors_1),
    .io_neighbors_2(Cell_14_io_neighbors_2),
    .io_neighbors_3(Cell_14_io_neighbors_3),
    .io_neighbors_4(Cell_14_io_neighbors_4),
    .io_neighbors_5(Cell_14_io_neighbors_5),
    .io_neighbors_6(Cell_14_io_neighbors_6),
    .io_neighbors_7(Cell_14_io_neighbors_7),
    .io_out(Cell_14_io_out),
    .io_running(Cell_14_io_running),
    .io_writeEnable(Cell_14_io_writeEnable),
    .io_writeValue(Cell_14_io_writeValue)
  );
  Cell Cell_15 ( // @[Life.scala 59:52]
    .clock(Cell_15_clock),
    .reset(Cell_15_reset),
    .io_neighbors_0(Cell_15_io_neighbors_0),
    .io_neighbors_1(Cell_15_io_neighbors_1),
    .io_neighbors_2(Cell_15_io_neighbors_2),
    .io_neighbors_3(Cell_15_io_neighbors_3),
    .io_neighbors_4(Cell_15_io_neighbors_4),
    .io_neighbors_5(Cell_15_io_neighbors_5),
    .io_neighbors_6(Cell_15_io_neighbors_6),
    .io_neighbors_7(Cell_15_io_neighbors_7),
    .io_out(Cell_15_io_out),
    .io_running(Cell_15_io_running),
    .io_writeEnable(Cell_15_io_writeEnable),
    .io_writeValue(Cell_15_io_writeValue)
  );
  Cell Cell_16 ( // @[Life.scala 59:52]
    .clock(Cell_16_clock),
    .reset(Cell_16_reset),
    .io_neighbors_0(Cell_16_io_neighbors_0),
    .io_neighbors_1(Cell_16_io_neighbors_1),
    .io_neighbors_2(Cell_16_io_neighbors_2),
    .io_neighbors_3(Cell_16_io_neighbors_3),
    .io_neighbors_4(Cell_16_io_neighbors_4),
    .io_neighbors_5(Cell_16_io_neighbors_5),
    .io_neighbors_6(Cell_16_io_neighbors_6),
    .io_neighbors_7(Cell_16_io_neighbors_7),
    .io_out(Cell_16_io_out),
    .io_running(Cell_16_io_running),
    .io_writeEnable(Cell_16_io_writeEnable),
    .io_writeValue(Cell_16_io_writeValue)
  );
  Cell Cell_17 ( // @[Life.scala 59:52]
    .clock(Cell_17_clock),
    .reset(Cell_17_reset),
    .io_neighbors_0(Cell_17_io_neighbors_0),
    .io_neighbors_1(Cell_17_io_neighbors_1),
    .io_neighbors_2(Cell_17_io_neighbors_2),
    .io_neighbors_3(Cell_17_io_neighbors_3),
    .io_neighbors_4(Cell_17_io_neighbors_4),
    .io_neighbors_5(Cell_17_io_neighbors_5),
    .io_neighbors_6(Cell_17_io_neighbors_6),
    .io_neighbors_7(Cell_17_io_neighbors_7),
    .io_out(Cell_17_io_out),
    .io_running(Cell_17_io_running),
    .io_writeEnable(Cell_17_io_writeEnable),
    .io_writeValue(Cell_17_io_writeValue)
  );
  Cell Cell_18 ( // @[Life.scala 59:52]
    .clock(Cell_18_clock),
    .reset(Cell_18_reset),
    .io_neighbors_0(Cell_18_io_neighbors_0),
    .io_neighbors_1(Cell_18_io_neighbors_1),
    .io_neighbors_2(Cell_18_io_neighbors_2),
    .io_neighbors_3(Cell_18_io_neighbors_3),
    .io_neighbors_4(Cell_18_io_neighbors_4),
    .io_neighbors_5(Cell_18_io_neighbors_5),
    .io_neighbors_6(Cell_18_io_neighbors_6),
    .io_neighbors_7(Cell_18_io_neighbors_7),
    .io_out(Cell_18_io_out),
    .io_running(Cell_18_io_running),
    .io_writeEnable(Cell_18_io_writeEnable),
    .io_writeValue(Cell_18_io_writeValue)
  );
  Cell Cell_19 ( // @[Life.scala 59:52]
    .clock(Cell_19_clock),
    .reset(Cell_19_reset),
    .io_neighbors_0(Cell_19_io_neighbors_0),
    .io_neighbors_1(Cell_19_io_neighbors_1),
    .io_neighbors_2(Cell_19_io_neighbors_2),
    .io_neighbors_3(Cell_19_io_neighbors_3),
    .io_neighbors_4(Cell_19_io_neighbors_4),
    .io_neighbors_5(Cell_19_io_neighbors_5),
    .io_neighbors_6(Cell_19_io_neighbors_6),
    .io_neighbors_7(Cell_19_io_neighbors_7),
    .io_out(Cell_19_io_out),
    .io_running(Cell_19_io_running),
    .io_writeEnable(Cell_19_io_writeEnable),
    .io_writeValue(Cell_19_io_writeValue)
  );
  Cell Cell_20 ( // @[Life.scala 59:52]
    .clock(Cell_20_clock),
    .reset(Cell_20_reset),
    .io_neighbors_0(Cell_20_io_neighbors_0),
    .io_neighbors_1(Cell_20_io_neighbors_1),
    .io_neighbors_2(Cell_20_io_neighbors_2),
    .io_neighbors_3(Cell_20_io_neighbors_3),
    .io_neighbors_4(Cell_20_io_neighbors_4),
    .io_neighbors_5(Cell_20_io_neighbors_5),
    .io_neighbors_6(Cell_20_io_neighbors_6),
    .io_neighbors_7(Cell_20_io_neighbors_7),
    .io_out(Cell_20_io_out),
    .io_running(Cell_20_io_running),
    .io_writeEnable(Cell_20_io_writeEnable),
    .io_writeValue(Cell_20_io_writeValue)
  );
  Cell Cell_21 ( // @[Life.scala 59:52]
    .clock(Cell_21_clock),
    .reset(Cell_21_reset),
    .io_neighbors_0(Cell_21_io_neighbors_0),
    .io_neighbors_1(Cell_21_io_neighbors_1),
    .io_neighbors_2(Cell_21_io_neighbors_2),
    .io_neighbors_3(Cell_21_io_neighbors_3),
    .io_neighbors_4(Cell_21_io_neighbors_4),
    .io_neighbors_5(Cell_21_io_neighbors_5),
    .io_neighbors_6(Cell_21_io_neighbors_6),
    .io_neighbors_7(Cell_21_io_neighbors_7),
    .io_out(Cell_21_io_out),
    .io_running(Cell_21_io_running),
    .io_writeEnable(Cell_21_io_writeEnable),
    .io_writeValue(Cell_21_io_writeValue)
  );
  Cell Cell_22 ( // @[Life.scala 59:52]
    .clock(Cell_22_clock),
    .reset(Cell_22_reset),
    .io_neighbors_0(Cell_22_io_neighbors_0),
    .io_neighbors_1(Cell_22_io_neighbors_1),
    .io_neighbors_2(Cell_22_io_neighbors_2),
    .io_neighbors_3(Cell_22_io_neighbors_3),
    .io_neighbors_4(Cell_22_io_neighbors_4),
    .io_neighbors_5(Cell_22_io_neighbors_5),
    .io_neighbors_6(Cell_22_io_neighbors_6),
    .io_neighbors_7(Cell_22_io_neighbors_7),
    .io_out(Cell_22_io_out),
    .io_running(Cell_22_io_running),
    .io_writeEnable(Cell_22_io_writeEnable),
    .io_writeValue(Cell_22_io_writeValue)
  );
  Cell Cell_23 ( // @[Life.scala 59:52]
    .clock(Cell_23_clock),
    .reset(Cell_23_reset),
    .io_neighbors_0(Cell_23_io_neighbors_0),
    .io_neighbors_1(Cell_23_io_neighbors_1),
    .io_neighbors_2(Cell_23_io_neighbors_2),
    .io_neighbors_3(Cell_23_io_neighbors_3),
    .io_neighbors_4(Cell_23_io_neighbors_4),
    .io_neighbors_5(Cell_23_io_neighbors_5),
    .io_neighbors_6(Cell_23_io_neighbors_6),
    .io_neighbors_7(Cell_23_io_neighbors_7),
    .io_out(Cell_23_io_out),
    .io_running(Cell_23_io_running),
    .io_writeEnable(Cell_23_io_writeEnable),
    .io_writeValue(Cell_23_io_writeValue)
  );
  Cell Cell_24 ( // @[Life.scala 59:52]
    .clock(Cell_24_clock),
    .reset(Cell_24_reset),
    .io_neighbors_0(Cell_24_io_neighbors_0),
    .io_neighbors_1(Cell_24_io_neighbors_1),
    .io_neighbors_2(Cell_24_io_neighbors_2),
    .io_neighbors_3(Cell_24_io_neighbors_3),
    .io_neighbors_4(Cell_24_io_neighbors_4),
    .io_neighbors_5(Cell_24_io_neighbors_5),
    .io_neighbors_6(Cell_24_io_neighbors_6),
    .io_neighbors_7(Cell_24_io_neighbors_7),
    .io_out(Cell_24_io_out),
    .io_running(Cell_24_io_running),
    .io_writeEnable(Cell_24_io_writeEnable),
    .io_writeValue(Cell_24_io_writeValue)
  );
  Cell Cell_25 ( // @[Life.scala 59:52]
    .clock(Cell_25_clock),
    .reset(Cell_25_reset),
    .io_neighbors_0(Cell_25_io_neighbors_0),
    .io_neighbors_1(Cell_25_io_neighbors_1),
    .io_neighbors_2(Cell_25_io_neighbors_2),
    .io_neighbors_3(Cell_25_io_neighbors_3),
    .io_neighbors_4(Cell_25_io_neighbors_4),
    .io_neighbors_5(Cell_25_io_neighbors_5),
    .io_neighbors_6(Cell_25_io_neighbors_6),
    .io_neighbors_7(Cell_25_io_neighbors_7),
    .io_out(Cell_25_io_out),
    .io_running(Cell_25_io_running),
    .io_writeEnable(Cell_25_io_writeEnable),
    .io_writeValue(Cell_25_io_writeValue)
  );
  Cell Cell_26 ( // @[Life.scala 59:52]
    .clock(Cell_26_clock),
    .reset(Cell_26_reset),
    .io_neighbors_0(Cell_26_io_neighbors_0),
    .io_neighbors_1(Cell_26_io_neighbors_1),
    .io_neighbors_2(Cell_26_io_neighbors_2),
    .io_neighbors_3(Cell_26_io_neighbors_3),
    .io_neighbors_4(Cell_26_io_neighbors_4),
    .io_neighbors_5(Cell_26_io_neighbors_5),
    .io_neighbors_6(Cell_26_io_neighbors_6),
    .io_neighbors_7(Cell_26_io_neighbors_7),
    .io_out(Cell_26_io_out),
    .io_running(Cell_26_io_running),
    .io_writeEnable(Cell_26_io_writeEnable),
    .io_writeValue(Cell_26_io_writeValue)
  );
  Cell Cell_27 ( // @[Life.scala 59:52]
    .clock(Cell_27_clock),
    .reset(Cell_27_reset),
    .io_neighbors_0(Cell_27_io_neighbors_0),
    .io_neighbors_1(Cell_27_io_neighbors_1),
    .io_neighbors_2(Cell_27_io_neighbors_2),
    .io_neighbors_3(Cell_27_io_neighbors_3),
    .io_neighbors_4(Cell_27_io_neighbors_4),
    .io_neighbors_5(Cell_27_io_neighbors_5),
    .io_neighbors_6(Cell_27_io_neighbors_6),
    .io_neighbors_7(Cell_27_io_neighbors_7),
    .io_out(Cell_27_io_out),
    .io_running(Cell_27_io_running),
    .io_writeEnable(Cell_27_io_writeEnable),
    .io_writeValue(Cell_27_io_writeValue)
  );
  Cell Cell_28 ( // @[Life.scala 59:52]
    .clock(Cell_28_clock),
    .reset(Cell_28_reset),
    .io_neighbors_0(Cell_28_io_neighbors_0),
    .io_neighbors_1(Cell_28_io_neighbors_1),
    .io_neighbors_2(Cell_28_io_neighbors_2),
    .io_neighbors_3(Cell_28_io_neighbors_3),
    .io_neighbors_4(Cell_28_io_neighbors_4),
    .io_neighbors_5(Cell_28_io_neighbors_5),
    .io_neighbors_6(Cell_28_io_neighbors_6),
    .io_neighbors_7(Cell_28_io_neighbors_7),
    .io_out(Cell_28_io_out),
    .io_running(Cell_28_io_running),
    .io_writeEnable(Cell_28_io_writeEnable),
    .io_writeValue(Cell_28_io_writeValue)
  );
  Cell Cell_29 ( // @[Life.scala 59:52]
    .clock(Cell_29_clock),
    .reset(Cell_29_reset),
    .io_neighbors_0(Cell_29_io_neighbors_0),
    .io_neighbors_1(Cell_29_io_neighbors_1),
    .io_neighbors_2(Cell_29_io_neighbors_2),
    .io_neighbors_3(Cell_29_io_neighbors_3),
    .io_neighbors_4(Cell_29_io_neighbors_4),
    .io_neighbors_5(Cell_29_io_neighbors_5),
    .io_neighbors_6(Cell_29_io_neighbors_6),
    .io_neighbors_7(Cell_29_io_neighbors_7),
    .io_out(Cell_29_io_out),
    .io_running(Cell_29_io_running),
    .io_writeEnable(Cell_29_io_writeEnable),
    .io_writeValue(Cell_29_io_writeValue)
  );
  Cell Cell_30 ( // @[Life.scala 59:52]
    .clock(Cell_30_clock),
    .reset(Cell_30_reset),
    .io_neighbors_0(Cell_30_io_neighbors_0),
    .io_neighbors_1(Cell_30_io_neighbors_1),
    .io_neighbors_2(Cell_30_io_neighbors_2),
    .io_neighbors_3(Cell_30_io_neighbors_3),
    .io_neighbors_4(Cell_30_io_neighbors_4),
    .io_neighbors_5(Cell_30_io_neighbors_5),
    .io_neighbors_6(Cell_30_io_neighbors_6),
    .io_neighbors_7(Cell_30_io_neighbors_7),
    .io_out(Cell_30_io_out),
    .io_running(Cell_30_io_running),
    .io_writeEnable(Cell_30_io_writeEnable),
    .io_writeValue(Cell_30_io_writeValue)
  );
  Cell Cell_31 ( // @[Life.scala 59:52]
    .clock(Cell_31_clock),
    .reset(Cell_31_reset),
    .io_neighbors_0(Cell_31_io_neighbors_0),
    .io_neighbors_1(Cell_31_io_neighbors_1),
    .io_neighbors_2(Cell_31_io_neighbors_2),
    .io_neighbors_3(Cell_31_io_neighbors_3),
    .io_neighbors_4(Cell_31_io_neighbors_4),
    .io_neighbors_5(Cell_31_io_neighbors_5),
    .io_neighbors_6(Cell_31_io_neighbors_6),
    .io_neighbors_7(Cell_31_io_neighbors_7),
    .io_out(Cell_31_io_out),
    .io_running(Cell_31_io_running),
    .io_writeEnable(Cell_31_io_writeEnable),
    .io_writeValue(Cell_31_io_writeValue)
  );
  Cell Cell_32 ( // @[Life.scala 59:52]
    .clock(Cell_32_clock),
    .reset(Cell_32_reset),
    .io_neighbors_0(Cell_32_io_neighbors_0),
    .io_neighbors_1(Cell_32_io_neighbors_1),
    .io_neighbors_2(Cell_32_io_neighbors_2),
    .io_neighbors_3(Cell_32_io_neighbors_3),
    .io_neighbors_4(Cell_32_io_neighbors_4),
    .io_neighbors_5(Cell_32_io_neighbors_5),
    .io_neighbors_6(Cell_32_io_neighbors_6),
    .io_neighbors_7(Cell_32_io_neighbors_7),
    .io_out(Cell_32_io_out),
    .io_running(Cell_32_io_running),
    .io_writeEnable(Cell_32_io_writeEnable),
    .io_writeValue(Cell_32_io_writeValue)
  );
  Cell Cell_33 ( // @[Life.scala 59:52]
    .clock(Cell_33_clock),
    .reset(Cell_33_reset),
    .io_neighbors_0(Cell_33_io_neighbors_0),
    .io_neighbors_1(Cell_33_io_neighbors_1),
    .io_neighbors_2(Cell_33_io_neighbors_2),
    .io_neighbors_3(Cell_33_io_neighbors_3),
    .io_neighbors_4(Cell_33_io_neighbors_4),
    .io_neighbors_5(Cell_33_io_neighbors_5),
    .io_neighbors_6(Cell_33_io_neighbors_6),
    .io_neighbors_7(Cell_33_io_neighbors_7),
    .io_out(Cell_33_io_out),
    .io_running(Cell_33_io_running),
    .io_writeEnable(Cell_33_io_writeEnable),
    .io_writeValue(Cell_33_io_writeValue)
  );
  Cell Cell_34 ( // @[Life.scala 59:52]
    .clock(Cell_34_clock),
    .reset(Cell_34_reset),
    .io_neighbors_0(Cell_34_io_neighbors_0),
    .io_neighbors_1(Cell_34_io_neighbors_1),
    .io_neighbors_2(Cell_34_io_neighbors_2),
    .io_neighbors_3(Cell_34_io_neighbors_3),
    .io_neighbors_4(Cell_34_io_neighbors_4),
    .io_neighbors_5(Cell_34_io_neighbors_5),
    .io_neighbors_6(Cell_34_io_neighbors_6),
    .io_neighbors_7(Cell_34_io_neighbors_7),
    .io_out(Cell_34_io_out),
    .io_running(Cell_34_io_running),
    .io_writeEnable(Cell_34_io_writeEnable),
    .io_writeValue(Cell_34_io_writeValue)
  );
  Cell Cell_35 ( // @[Life.scala 59:52]
    .clock(Cell_35_clock),
    .reset(Cell_35_reset),
    .io_neighbors_0(Cell_35_io_neighbors_0),
    .io_neighbors_1(Cell_35_io_neighbors_1),
    .io_neighbors_2(Cell_35_io_neighbors_2),
    .io_neighbors_3(Cell_35_io_neighbors_3),
    .io_neighbors_4(Cell_35_io_neighbors_4),
    .io_neighbors_5(Cell_35_io_neighbors_5),
    .io_neighbors_6(Cell_35_io_neighbors_6),
    .io_neighbors_7(Cell_35_io_neighbors_7),
    .io_out(Cell_35_io_out),
    .io_running(Cell_35_io_running),
    .io_writeEnable(Cell_35_io_writeEnable),
    .io_writeValue(Cell_35_io_writeValue)
  );
  Cell Cell_36 ( // @[Life.scala 59:52]
    .clock(Cell_36_clock),
    .reset(Cell_36_reset),
    .io_neighbors_0(Cell_36_io_neighbors_0),
    .io_neighbors_1(Cell_36_io_neighbors_1),
    .io_neighbors_2(Cell_36_io_neighbors_2),
    .io_neighbors_3(Cell_36_io_neighbors_3),
    .io_neighbors_4(Cell_36_io_neighbors_4),
    .io_neighbors_5(Cell_36_io_neighbors_5),
    .io_neighbors_6(Cell_36_io_neighbors_6),
    .io_neighbors_7(Cell_36_io_neighbors_7),
    .io_out(Cell_36_io_out),
    .io_running(Cell_36_io_running),
    .io_writeEnable(Cell_36_io_writeEnable),
    .io_writeValue(Cell_36_io_writeValue)
  );
  Cell Cell_37 ( // @[Life.scala 59:52]
    .clock(Cell_37_clock),
    .reset(Cell_37_reset),
    .io_neighbors_0(Cell_37_io_neighbors_0),
    .io_neighbors_1(Cell_37_io_neighbors_1),
    .io_neighbors_2(Cell_37_io_neighbors_2),
    .io_neighbors_3(Cell_37_io_neighbors_3),
    .io_neighbors_4(Cell_37_io_neighbors_4),
    .io_neighbors_5(Cell_37_io_neighbors_5),
    .io_neighbors_6(Cell_37_io_neighbors_6),
    .io_neighbors_7(Cell_37_io_neighbors_7),
    .io_out(Cell_37_io_out),
    .io_running(Cell_37_io_running),
    .io_writeEnable(Cell_37_io_writeEnable),
    .io_writeValue(Cell_37_io_writeValue)
  );
  Cell Cell_38 ( // @[Life.scala 59:52]
    .clock(Cell_38_clock),
    .reset(Cell_38_reset),
    .io_neighbors_0(Cell_38_io_neighbors_0),
    .io_neighbors_1(Cell_38_io_neighbors_1),
    .io_neighbors_2(Cell_38_io_neighbors_2),
    .io_neighbors_3(Cell_38_io_neighbors_3),
    .io_neighbors_4(Cell_38_io_neighbors_4),
    .io_neighbors_5(Cell_38_io_neighbors_5),
    .io_neighbors_6(Cell_38_io_neighbors_6),
    .io_neighbors_7(Cell_38_io_neighbors_7),
    .io_out(Cell_38_io_out),
    .io_running(Cell_38_io_running),
    .io_writeEnable(Cell_38_io_writeEnable),
    .io_writeValue(Cell_38_io_writeValue)
  );
  Cell Cell_39 ( // @[Life.scala 59:52]
    .clock(Cell_39_clock),
    .reset(Cell_39_reset),
    .io_neighbors_0(Cell_39_io_neighbors_0),
    .io_neighbors_1(Cell_39_io_neighbors_1),
    .io_neighbors_2(Cell_39_io_neighbors_2),
    .io_neighbors_3(Cell_39_io_neighbors_3),
    .io_neighbors_4(Cell_39_io_neighbors_4),
    .io_neighbors_5(Cell_39_io_neighbors_5),
    .io_neighbors_6(Cell_39_io_neighbors_6),
    .io_neighbors_7(Cell_39_io_neighbors_7),
    .io_out(Cell_39_io_out),
    .io_running(Cell_39_io_running),
    .io_writeEnable(Cell_39_io_writeEnable),
    .io_writeValue(Cell_39_io_writeValue)
  );
  Cell Cell_40 ( // @[Life.scala 59:52]
    .clock(Cell_40_clock),
    .reset(Cell_40_reset),
    .io_neighbors_0(Cell_40_io_neighbors_0),
    .io_neighbors_1(Cell_40_io_neighbors_1),
    .io_neighbors_2(Cell_40_io_neighbors_2),
    .io_neighbors_3(Cell_40_io_neighbors_3),
    .io_neighbors_4(Cell_40_io_neighbors_4),
    .io_neighbors_5(Cell_40_io_neighbors_5),
    .io_neighbors_6(Cell_40_io_neighbors_6),
    .io_neighbors_7(Cell_40_io_neighbors_7),
    .io_out(Cell_40_io_out),
    .io_running(Cell_40_io_running),
    .io_writeEnable(Cell_40_io_writeEnable),
    .io_writeValue(Cell_40_io_writeValue)
  );
  Cell Cell_41 ( // @[Life.scala 59:52]
    .clock(Cell_41_clock),
    .reset(Cell_41_reset),
    .io_neighbors_0(Cell_41_io_neighbors_0),
    .io_neighbors_1(Cell_41_io_neighbors_1),
    .io_neighbors_2(Cell_41_io_neighbors_2),
    .io_neighbors_3(Cell_41_io_neighbors_3),
    .io_neighbors_4(Cell_41_io_neighbors_4),
    .io_neighbors_5(Cell_41_io_neighbors_5),
    .io_neighbors_6(Cell_41_io_neighbors_6),
    .io_neighbors_7(Cell_41_io_neighbors_7),
    .io_out(Cell_41_io_out),
    .io_running(Cell_41_io_running),
    .io_writeEnable(Cell_41_io_writeEnable),
    .io_writeValue(Cell_41_io_writeValue)
  );
  Cell Cell_42 ( // @[Life.scala 59:52]
    .clock(Cell_42_clock),
    .reset(Cell_42_reset),
    .io_neighbors_0(Cell_42_io_neighbors_0),
    .io_neighbors_1(Cell_42_io_neighbors_1),
    .io_neighbors_2(Cell_42_io_neighbors_2),
    .io_neighbors_3(Cell_42_io_neighbors_3),
    .io_neighbors_4(Cell_42_io_neighbors_4),
    .io_neighbors_5(Cell_42_io_neighbors_5),
    .io_neighbors_6(Cell_42_io_neighbors_6),
    .io_neighbors_7(Cell_42_io_neighbors_7),
    .io_out(Cell_42_io_out),
    .io_running(Cell_42_io_running),
    .io_writeEnable(Cell_42_io_writeEnable),
    .io_writeValue(Cell_42_io_writeValue)
  );
  Cell Cell_43 ( // @[Life.scala 59:52]
    .clock(Cell_43_clock),
    .reset(Cell_43_reset),
    .io_neighbors_0(Cell_43_io_neighbors_0),
    .io_neighbors_1(Cell_43_io_neighbors_1),
    .io_neighbors_2(Cell_43_io_neighbors_2),
    .io_neighbors_3(Cell_43_io_neighbors_3),
    .io_neighbors_4(Cell_43_io_neighbors_4),
    .io_neighbors_5(Cell_43_io_neighbors_5),
    .io_neighbors_6(Cell_43_io_neighbors_6),
    .io_neighbors_7(Cell_43_io_neighbors_7),
    .io_out(Cell_43_io_out),
    .io_running(Cell_43_io_running),
    .io_writeEnable(Cell_43_io_writeEnable),
    .io_writeValue(Cell_43_io_writeValue)
  );
  Cell Cell_44 ( // @[Life.scala 59:52]
    .clock(Cell_44_clock),
    .reset(Cell_44_reset),
    .io_neighbors_0(Cell_44_io_neighbors_0),
    .io_neighbors_1(Cell_44_io_neighbors_1),
    .io_neighbors_2(Cell_44_io_neighbors_2),
    .io_neighbors_3(Cell_44_io_neighbors_3),
    .io_neighbors_4(Cell_44_io_neighbors_4),
    .io_neighbors_5(Cell_44_io_neighbors_5),
    .io_neighbors_6(Cell_44_io_neighbors_6),
    .io_neighbors_7(Cell_44_io_neighbors_7),
    .io_out(Cell_44_io_out),
    .io_running(Cell_44_io_running),
    .io_writeEnable(Cell_44_io_writeEnable),
    .io_writeValue(Cell_44_io_writeValue)
  );
  Cell Cell_45 ( // @[Life.scala 59:52]
    .clock(Cell_45_clock),
    .reset(Cell_45_reset),
    .io_neighbors_0(Cell_45_io_neighbors_0),
    .io_neighbors_1(Cell_45_io_neighbors_1),
    .io_neighbors_2(Cell_45_io_neighbors_2),
    .io_neighbors_3(Cell_45_io_neighbors_3),
    .io_neighbors_4(Cell_45_io_neighbors_4),
    .io_neighbors_5(Cell_45_io_neighbors_5),
    .io_neighbors_6(Cell_45_io_neighbors_6),
    .io_neighbors_7(Cell_45_io_neighbors_7),
    .io_out(Cell_45_io_out),
    .io_running(Cell_45_io_running),
    .io_writeEnable(Cell_45_io_writeEnable),
    .io_writeValue(Cell_45_io_writeValue)
  );
  Cell Cell_46 ( // @[Life.scala 59:52]
    .clock(Cell_46_clock),
    .reset(Cell_46_reset),
    .io_neighbors_0(Cell_46_io_neighbors_0),
    .io_neighbors_1(Cell_46_io_neighbors_1),
    .io_neighbors_2(Cell_46_io_neighbors_2),
    .io_neighbors_3(Cell_46_io_neighbors_3),
    .io_neighbors_4(Cell_46_io_neighbors_4),
    .io_neighbors_5(Cell_46_io_neighbors_5),
    .io_neighbors_6(Cell_46_io_neighbors_6),
    .io_neighbors_7(Cell_46_io_neighbors_7),
    .io_out(Cell_46_io_out),
    .io_running(Cell_46_io_running),
    .io_writeEnable(Cell_46_io_writeEnable),
    .io_writeValue(Cell_46_io_writeValue)
  );
  Cell Cell_47 ( // @[Life.scala 59:52]
    .clock(Cell_47_clock),
    .reset(Cell_47_reset),
    .io_neighbors_0(Cell_47_io_neighbors_0),
    .io_neighbors_1(Cell_47_io_neighbors_1),
    .io_neighbors_2(Cell_47_io_neighbors_2),
    .io_neighbors_3(Cell_47_io_neighbors_3),
    .io_neighbors_4(Cell_47_io_neighbors_4),
    .io_neighbors_5(Cell_47_io_neighbors_5),
    .io_neighbors_6(Cell_47_io_neighbors_6),
    .io_neighbors_7(Cell_47_io_neighbors_7),
    .io_out(Cell_47_io_out),
    .io_running(Cell_47_io_running),
    .io_writeEnable(Cell_47_io_writeEnable),
    .io_writeValue(Cell_47_io_writeValue)
  );
  Cell Cell_48 ( // @[Life.scala 59:52]
    .clock(Cell_48_clock),
    .reset(Cell_48_reset),
    .io_neighbors_0(Cell_48_io_neighbors_0),
    .io_neighbors_1(Cell_48_io_neighbors_1),
    .io_neighbors_2(Cell_48_io_neighbors_2),
    .io_neighbors_3(Cell_48_io_neighbors_3),
    .io_neighbors_4(Cell_48_io_neighbors_4),
    .io_neighbors_5(Cell_48_io_neighbors_5),
    .io_neighbors_6(Cell_48_io_neighbors_6),
    .io_neighbors_7(Cell_48_io_neighbors_7),
    .io_out(Cell_48_io_out),
    .io_running(Cell_48_io_running),
    .io_writeEnable(Cell_48_io_writeEnable),
    .io_writeValue(Cell_48_io_writeValue)
  );
  Cell Cell_49 ( // @[Life.scala 59:52]
    .clock(Cell_49_clock),
    .reset(Cell_49_reset),
    .io_neighbors_0(Cell_49_io_neighbors_0),
    .io_neighbors_1(Cell_49_io_neighbors_1),
    .io_neighbors_2(Cell_49_io_neighbors_2),
    .io_neighbors_3(Cell_49_io_neighbors_3),
    .io_neighbors_4(Cell_49_io_neighbors_4),
    .io_neighbors_5(Cell_49_io_neighbors_5),
    .io_neighbors_6(Cell_49_io_neighbors_6),
    .io_neighbors_7(Cell_49_io_neighbors_7),
    .io_out(Cell_49_io_out),
    .io_running(Cell_49_io_running),
    .io_writeEnable(Cell_49_io_writeEnable),
    .io_writeValue(Cell_49_io_writeValue)
  );
  Cell Cell_50 ( // @[Life.scala 59:52]
    .clock(Cell_50_clock),
    .reset(Cell_50_reset),
    .io_neighbors_0(Cell_50_io_neighbors_0),
    .io_neighbors_1(Cell_50_io_neighbors_1),
    .io_neighbors_2(Cell_50_io_neighbors_2),
    .io_neighbors_3(Cell_50_io_neighbors_3),
    .io_neighbors_4(Cell_50_io_neighbors_4),
    .io_neighbors_5(Cell_50_io_neighbors_5),
    .io_neighbors_6(Cell_50_io_neighbors_6),
    .io_neighbors_7(Cell_50_io_neighbors_7),
    .io_out(Cell_50_io_out),
    .io_running(Cell_50_io_running),
    .io_writeEnable(Cell_50_io_writeEnable),
    .io_writeValue(Cell_50_io_writeValue)
  );
  Cell Cell_51 ( // @[Life.scala 59:52]
    .clock(Cell_51_clock),
    .reset(Cell_51_reset),
    .io_neighbors_0(Cell_51_io_neighbors_0),
    .io_neighbors_1(Cell_51_io_neighbors_1),
    .io_neighbors_2(Cell_51_io_neighbors_2),
    .io_neighbors_3(Cell_51_io_neighbors_3),
    .io_neighbors_4(Cell_51_io_neighbors_4),
    .io_neighbors_5(Cell_51_io_neighbors_5),
    .io_neighbors_6(Cell_51_io_neighbors_6),
    .io_neighbors_7(Cell_51_io_neighbors_7),
    .io_out(Cell_51_io_out),
    .io_running(Cell_51_io_running),
    .io_writeEnable(Cell_51_io_writeEnable),
    .io_writeValue(Cell_51_io_writeValue)
  );
  Cell Cell_52 ( // @[Life.scala 59:52]
    .clock(Cell_52_clock),
    .reset(Cell_52_reset),
    .io_neighbors_0(Cell_52_io_neighbors_0),
    .io_neighbors_1(Cell_52_io_neighbors_1),
    .io_neighbors_2(Cell_52_io_neighbors_2),
    .io_neighbors_3(Cell_52_io_neighbors_3),
    .io_neighbors_4(Cell_52_io_neighbors_4),
    .io_neighbors_5(Cell_52_io_neighbors_5),
    .io_neighbors_6(Cell_52_io_neighbors_6),
    .io_neighbors_7(Cell_52_io_neighbors_7),
    .io_out(Cell_52_io_out),
    .io_running(Cell_52_io_running),
    .io_writeEnable(Cell_52_io_writeEnable),
    .io_writeValue(Cell_52_io_writeValue)
  );
  Cell Cell_53 ( // @[Life.scala 59:52]
    .clock(Cell_53_clock),
    .reset(Cell_53_reset),
    .io_neighbors_0(Cell_53_io_neighbors_0),
    .io_neighbors_1(Cell_53_io_neighbors_1),
    .io_neighbors_2(Cell_53_io_neighbors_2),
    .io_neighbors_3(Cell_53_io_neighbors_3),
    .io_neighbors_4(Cell_53_io_neighbors_4),
    .io_neighbors_5(Cell_53_io_neighbors_5),
    .io_neighbors_6(Cell_53_io_neighbors_6),
    .io_neighbors_7(Cell_53_io_neighbors_7),
    .io_out(Cell_53_io_out),
    .io_running(Cell_53_io_running),
    .io_writeEnable(Cell_53_io_writeEnable),
    .io_writeValue(Cell_53_io_writeValue)
  );
  Cell Cell_54 ( // @[Life.scala 59:52]
    .clock(Cell_54_clock),
    .reset(Cell_54_reset),
    .io_neighbors_0(Cell_54_io_neighbors_0),
    .io_neighbors_1(Cell_54_io_neighbors_1),
    .io_neighbors_2(Cell_54_io_neighbors_2),
    .io_neighbors_3(Cell_54_io_neighbors_3),
    .io_neighbors_4(Cell_54_io_neighbors_4),
    .io_neighbors_5(Cell_54_io_neighbors_5),
    .io_neighbors_6(Cell_54_io_neighbors_6),
    .io_neighbors_7(Cell_54_io_neighbors_7),
    .io_out(Cell_54_io_out),
    .io_running(Cell_54_io_running),
    .io_writeEnable(Cell_54_io_writeEnable),
    .io_writeValue(Cell_54_io_writeValue)
  );
  Cell Cell_55 ( // @[Life.scala 59:52]
    .clock(Cell_55_clock),
    .reset(Cell_55_reset),
    .io_neighbors_0(Cell_55_io_neighbors_0),
    .io_neighbors_1(Cell_55_io_neighbors_1),
    .io_neighbors_2(Cell_55_io_neighbors_2),
    .io_neighbors_3(Cell_55_io_neighbors_3),
    .io_neighbors_4(Cell_55_io_neighbors_4),
    .io_neighbors_5(Cell_55_io_neighbors_5),
    .io_neighbors_6(Cell_55_io_neighbors_6),
    .io_neighbors_7(Cell_55_io_neighbors_7),
    .io_out(Cell_55_io_out),
    .io_running(Cell_55_io_running),
    .io_writeEnable(Cell_55_io_writeEnable),
    .io_writeValue(Cell_55_io_writeValue)
  );
  Cell Cell_56 ( // @[Life.scala 59:52]
    .clock(Cell_56_clock),
    .reset(Cell_56_reset),
    .io_neighbors_0(Cell_56_io_neighbors_0),
    .io_neighbors_1(Cell_56_io_neighbors_1),
    .io_neighbors_2(Cell_56_io_neighbors_2),
    .io_neighbors_3(Cell_56_io_neighbors_3),
    .io_neighbors_4(Cell_56_io_neighbors_4),
    .io_neighbors_5(Cell_56_io_neighbors_5),
    .io_neighbors_6(Cell_56_io_neighbors_6),
    .io_neighbors_7(Cell_56_io_neighbors_7),
    .io_out(Cell_56_io_out),
    .io_running(Cell_56_io_running),
    .io_writeEnable(Cell_56_io_writeEnable),
    .io_writeValue(Cell_56_io_writeValue)
  );
  Cell Cell_57 ( // @[Life.scala 59:52]
    .clock(Cell_57_clock),
    .reset(Cell_57_reset),
    .io_neighbors_0(Cell_57_io_neighbors_0),
    .io_neighbors_1(Cell_57_io_neighbors_1),
    .io_neighbors_2(Cell_57_io_neighbors_2),
    .io_neighbors_3(Cell_57_io_neighbors_3),
    .io_neighbors_4(Cell_57_io_neighbors_4),
    .io_neighbors_5(Cell_57_io_neighbors_5),
    .io_neighbors_6(Cell_57_io_neighbors_6),
    .io_neighbors_7(Cell_57_io_neighbors_7),
    .io_out(Cell_57_io_out),
    .io_running(Cell_57_io_running),
    .io_writeEnable(Cell_57_io_writeEnable),
    .io_writeValue(Cell_57_io_writeValue)
  );
  Cell Cell_58 ( // @[Life.scala 59:52]
    .clock(Cell_58_clock),
    .reset(Cell_58_reset),
    .io_neighbors_0(Cell_58_io_neighbors_0),
    .io_neighbors_1(Cell_58_io_neighbors_1),
    .io_neighbors_2(Cell_58_io_neighbors_2),
    .io_neighbors_3(Cell_58_io_neighbors_3),
    .io_neighbors_4(Cell_58_io_neighbors_4),
    .io_neighbors_5(Cell_58_io_neighbors_5),
    .io_neighbors_6(Cell_58_io_neighbors_6),
    .io_neighbors_7(Cell_58_io_neighbors_7),
    .io_out(Cell_58_io_out),
    .io_running(Cell_58_io_running),
    .io_writeEnable(Cell_58_io_writeEnable),
    .io_writeValue(Cell_58_io_writeValue)
  );
  Cell Cell_59 ( // @[Life.scala 59:52]
    .clock(Cell_59_clock),
    .reset(Cell_59_reset),
    .io_neighbors_0(Cell_59_io_neighbors_0),
    .io_neighbors_1(Cell_59_io_neighbors_1),
    .io_neighbors_2(Cell_59_io_neighbors_2),
    .io_neighbors_3(Cell_59_io_neighbors_3),
    .io_neighbors_4(Cell_59_io_neighbors_4),
    .io_neighbors_5(Cell_59_io_neighbors_5),
    .io_neighbors_6(Cell_59_io_neighbors_6),
    .io_neighbors_7(Cell_59_io_neighbors_7),
    .io_out(Cell_59_io_out),
    .io_running(Cell_59_io_running),
    .io_writeEnable(Cell_59_io_writeEnable),
    .io_writeValue(Cell_59_io_writeValue)
  );
  Cell Cell_60 ( // @[Life.scala 59:52]
    .clock(Cell_60_clock),
    .reset(Cell_60_reset),
    .io_neighbors_0(Cell_60_io_neighbors_0),
    .io_neighbors_1(Cell_60_io_neighbors_1),
    .io_neighbors_2(Cell_60_io_neighbors_2),
    .io_neighbors_3(Cell_60_io_neighbors_3),
    .io_neighbors_4(Cell_60_io_neighbors_4),
    .io_neighbors_5(Cell_60_io_neighbors_5),
    .io_neighbors_6(Cell_60_io_neighbors_6),
    .io_neighbors_7(Cell_60_io_neighbors_7),
    .io_out(Cell_60_io_out),
    .io_running(Cell_60_io_running),
    .io_writeEnable(Cell_60_io_writeEnable),
    .io_writeValue(Cell_60_io_writeValue)
  );
  Cell Cell_61 ( // @[Life.scala 59:52]
    .clock(Cell_61_clock),
    .reset(Cell_61_reset),
    .io_neighbors_0(Cell_61_io_neighbors_0),
    .io_neighbors_1(Cell_61_io_neighbors_1),
    .io_neighbors_2(Cell_61_io_neighbors_2),
    .io_neighbors_3(Cell_61_io_neighbors_3),
    .io_neighbors_4(Cell_61_io_neighbors_4),
    .io_neighbors_5(Cell_61_io_neighbors_5),
    .io_neighbors_6(Cell_61_io_neighbors_6),
    .io_neighbors_7(Cell_61_io_neighbors_7),
    .io_out(Cell_61_io_out),
    .io_running(Cell_61_io_running),
    .io_writeEnable(Cell_61_io_writeEnable),
    .io_writeValue(Cell_61_io_writeValue)
  );
  Cell Cell_62 ( // @[Life.scala 59:52]
    .clock(Cell_62_clock),
    .reset(Cell_62_reset),
    .io_neighbors_0(Cell_62_io_neighbors_0),
    .io_neighbors_1(Cell_62_io_neighbors_1),
    .io_neighbors_2(Cell_62_io_neighbors_2),
    .io_neighbors_3(Cell_62_io_neighbors_3),
    .io_neighbors_4(Cell_62_io_neighbors_4),
    .io_neighbors_5(Cell_62_io_neighbors_5),
    .io_neighbors_6(Cell_62_io_neighbors_6),
    .io_neighbors_7(Cell_62_io_neighbors_7),
    .io_out(Cell_62_io_out),
    .io_running(Cell_62_io_running),
    .io_writeEnable(Cell_62_io_writeEnable),
    .io_writeValue(Cell_62_io_writeValue)
  );
  Cell Cell_63 ( // @[Life.scala 59:52]
    .clock(Cell_63_clock),
    .reset(Cell_63_reset),
    .io_neighbors_0(Cell_63_io_neighbors_0),
    .io_neighbors_1(Cell_63_io_neighbors_1),
    .io_neighbors_2(Cell_63_io_neighbors_2),
    .io_neighbors_3(Cell_63_io_neighbors_3),
    .io_neighbors_4(Cell_63_io_neighbors_4),
    .io_neighbors_5(Cell_63_io_neighbors_5),
    .io_neighbors_6(Cell_63_io_neighbors_6),
    .io_neighbors_7(Cell_63_io_neighbors_7),
    .io_out(Cell_63_io_out),
    .io_running(Cell_63_io_running),
    .io_writeEnable(Cell_63_io_writeEnable),
    .io_writeValue(Cell_63_io_writeValue)
  );
  Cell Cell_64 ( // @[Life.scala 59:52]
    .clock(Cell_64_clock),
    .reset(Cell_64_reset),
    .io_neighbors_0(Cell_64_io_neighbors_0),
    .io_neighbors_1(Cell_64_io_neighbors_1),
    .io_neighbors_2(Cell_64_io_neighbors_2),
    .io_neighbors_3(Cell_64_io_neighbors_3),
    .io_neighbors_4(Cell_64_io_neighbors_4),
    .io_neighbors_5(Cell_64_io_neighbors_5),
    .io_neighbors_6(Cell_64_io_neighbors_6),
    .io_neighbors_7(Cell_64_io_neighbors_7),
    .io_out(Cell_64_io_out),
    .io_running(Cell_64_io_running),
    .io_writeEnable(Cell_64_io_writeEnable),
    .io_writeValue(Cell_64_io_writeValue)
  );
  Cell Cell_65 ( // @[Life.scala 59:52]
    .clock(Cell_65_clock),
    .reset(Cell_65_reset),
    .io_neighbors_0(Cell_65_io_neighbors_0),
    .io_neighbors_1(Cell_65_io_neighbors_1),
    .io_neighbors_2(Cell_65_io_neighbors_2),
    .io_neighbors_3(Cell_65_io_neighbors_3),
    .io_neighbors_4(Cell_65_io_neighbors_4),
    .io_neighbors_5(Cell_65_io_neighbors_5),
    .io_neighbors_6(Cell_65_io_neighbors_6),
    .io_neighbors_7(Cell_65_io_neighbors_7),
    .io_out(Cell_65_io_out),
    .io_running(Cell_65_io_running),
    .io_writeEnable(Cell_65_io_writeEnable),
    .io_writeValue(Cell_65_io_writeValue)
  );
  Cell Cell_66 ( // @[Life.scala 59:52]
    .clock(Cell_66_clock),
    .reset(Cell_66_reset),
    .io_neighbors_0(Cell_66_io_neighbors_0),
    .io_neighbors_1(Cell_66_io_neighbors_1),
    .io_neighbors_2(Cell_66_io_neighbors_2),
    .io_neighbors_3(Cell_66_io_neighbors_3),
    .io_neighbors_4(Cell_66_io_neighbors_4),
    .io_neighbors_5(Cell_66_io_neighbors_5),
    .io_neighbors_6(Cell_66_io_neighbors_6),
    .io_neighbors_7(Cell_66_io_neighbors_7),
    .io_out(Cell_66_io_out),
    .io_running(Cell_66_io_running),
    .io_writeEnable(Cell_66_io_writeEnable),
    .io_writeValue(Cell_66_io_writeValue)
  );
  Cell Cell_67 ( // @[Life.scala 59:52]
    .clock(Cell_67_clock),
    .reset(Cell_67_reset),
    .io_neighbors_0(Cell_67_io_neighbors_0),
    .io_neighbors_1(Cell_67_io_neighbors_1),
    .io_neighbors_2(Cell_67_io_neighbors_2),
    .io_neighbors_3(Cell_67_io_neighbors_3),
    .io_neighbors_4(Cell_67_io_neighbors_4),
    .io_neighbors_5(Cell_67_io_neighbors_5),
    .io_neighbors_6(Cell_67_io_neighbors_6),
    .io_neighbors_7(Cell_67_io_neighbors_7),
    .io_out(Cell_67_io_out),
    .io_running(Cell_67_io_running),
    .io_writeEnable(Cell_67_io_writeEnable),
    .io_writeValue(Cell_67_io_writeValue)
  );
  Cell Cell_68 ( // @[Life.scala 59:52]
    .clock(Cell_68_clock),
    .reset(Cell_68_reset),
    .io_neighbors_0(Cell_68_io_neighbors_0),
    .io_neighbors_1(Cell_68_io_neighbors_1),
    .io_neighbors_2(Cell_68_io_neighbors_2),
    .io_neighbors_3(Cell_68_io_neighbors_3),
    .io_neighbors_4(Cell_68_io_neighbors_4),
    .io_neighbors_5(Cell_68_io_neighbors_5),
    .io_neighbors_6(Cell_68_io_neighbors_6),
    .io_neighbors_7(Cell_68_io_neighbors_7),
    .io_out(Cell_68_io_out),
    .io_running(Cell_68_io_running),
    .io_writeEnable(Cell_68_io_writeEnable),
    .io_writeValue(Cell_68_io_writeValue)
  );
  Cell Cell_69 ( // @[Life.scala 59:52]
    .clock(Cell_69_clock),
    .reset(Cell_69_reset),
    .io_neighbors_0(Cell_69_io_neighbors_0),
    .io_neighbors_1(Cell_69_io_neighbors_1),
    .io_neighbors_2(Cell_69_io_neighbors_2),
    .io_neighbors_3(Cell_69_io_neighbors_3),
    .io_neighbors_4(Cell_69_io_neighbors_4),
    .io_neighbors_5(Cell_69_io_neighbors_5),
    .io_neighbors_6(Cell_69_io_neighbors_6),
    .io_neighbors_7(Cell_69_io_neighbors_7),
    .io_out(Cell_69_io_out),
    .io_running(Cell_69_io_running),
    .io_writeEnable(Cell_69_io_writeEnable),
    .io_writeValue(Cell_69_io_writeValue)
  );
  Cell Cell_70 ( // @[Life.scala 59:52]
    .clock(Cell_70_clock),
    .reset(Cell_70_reset),
    .io_neighbors_0(Cell_70_io_neighbors_0),
    .io_neighbors_1(Cell_70_io_neighbors_1),
    .io_neighbors_2(Cell_70_io_neighbors_2),
    .io_neighbors_3(Cell_70_io_neighbors_3),
    .io_neighbors_4(Cell_70_io_neighbors_4),
    .io_neighbors_5(Cell_70_io_neighbors_5),
    .io_neighbors_6(Cell_70_io_neighbors_6),
    .io_neighbors_7(Cell_70_io_neighbors_7),
    .io_out(Cell_70_io_out),
    .io_running(Cell_70_io_running),
    .io_writeEnable(Cell_70_io_writeEnable),
    .io_writeValue(Cell_70_io_writeValue)
  );
  Cell Cell_71 ( // @[Life.scala 59:52]
    .clock(Cell_71_clock),
    .reset(Cell_71_reset),
    .io_neighbors_0(Cell_71_io_neighbors_0),
    .io_neighbors_1(Cell_71_io_neighbors_1),
    .io_neighbors_2(Cell_71_io_neighbors_2),
    .io_neighbors_3(Cell_71_io_neighbors_3),
    .io_neighbors_4(Cell_71_io_neighbors_4),
    .io_neighbors_5(Cell_71_io_neighbors_5),
    .io_neighbors_6(Cell_71_io_neighbors_6),
    .io_neighbors_7(Cell_71_io_neighbors_7),
    .io_out(Cell_71_io_out),
    .io_running(Cell_71_io_running),
    .io_writeEnable(Cell_71_io_writeEnable),
    .io_writeValue(Cell_71_io_writeValue)
  );
  Cell Cell_72 ( // @[Life.scala 59:52]
    .clock(Cell_72_clock),
    .reset(Cell_72_reset),
    .io_neighbors_0(Cell_72_io_neighbors_0),
    .io_neighbors_1(Cell_72_io_neighbors_1),
    .io_neighbors_2(Cell_72_io_neighbors_2),
    .io_neighbors_3(Cell_72_io_neighbors_3),
    .io_neighbors_4(Cell_72_io_neighbors_4),
    .io_neighbors_5(Cell_72_io_neighbors_5),
    .io_neighbors_6(Cell_72_io_neighbors_6),
    .io_neighbors_7(Cell_72_io_neighbors_7),
    .io_out(Cell_72_io_out),
    .io_running(Cell_72_io_running),
    .io_writeEnable(Cell_72_io_writeEnable),
    .io_writeValue(Cell_72_io_writeValue)
  );
  Cell Cell_73 ( // @[Life.scala 59:52]
    .clock(Cell_73_clock),
    .reset(Cell_73_reset),
    .io_neighbors_0(Cell_73_io_neighbors_0),
    .io_neighbors_1(Cell_73_io_neighbors_1),
    .io_neighbors_2(Cell_73_io_neighbors_2),
    .io_neighbors_3(Cell_73_io_neighbors_3),
    .io_neighbors_4(Cell_73_io_neighbors_4),
    .io_neighbors_5(Cell_73_io_neighbors_5),
    .io_neighbors_6(Cell_73_io_neighbors_6),
    .io_neighbors_7(Cell_73_io_neighbors_7),
    .io_out(Cell_73_io_out),
    .io_running(Cell_73_io_running),
    .io_writeEnable(Cell_73_io_writeEnable),
    .io_writeValue(Cell_73_io_writeValue)
  );
  Cell Cell_74 ( // @[Life.scala 59:52]
    .clock(Cell_74_clock),
    .reset(Cell_74_reset),
    .io_neighbors_0(Cell_74_io_neighbors_0),
    .io_neighbors_1(Cell_74_io_neighbors_1),
    .io_neighbors_2(Cell_74_io_neighbors_2),
    .io_neighbors_3(Cell_74_io_neighbors_3),
    .io_neighbors_4(Cell_74_io_neighbors_4),
    .io_neighbors_5(Cell_74_io_neighbors_5),
    .io_neighbors_6(Cell_74_io_neighbors_6),
    .io_neighbors_7(Cell_74_io_neighbors_7),
    .io_out(Cell_74_io_out),
    .io_running(Cell_74_io_running),
    .io_writeEnable(Cell_74_io_writeEnable),
    .io_writeValue(Cell_74_io_writeValue)
  );
  Cell Cell_75 ( // @[Life.scala 59:52]
    .clock(Cell_75_clock),
    .reset(Cell_75_reset),
    .io_neighbors_0(Cell_75_io_neighbors_0),
    .io_neighbors_1(Cell_75_io_neighbors_1),
    .io_neighbors_2(Cell_75_io_neighbors_2),
    .io_neighbors_3(Cell_75_io_neighbors_3),
    .io_neighbors_4(Cell_75_io_neighbors_4),
    .io_neighbors_5(Cell_75_io_neighbors_5),
    .io_neighbors_6(Cell_75_io_neighbors_6),
    .io_neighbors_7(Cell_75_io_neighbors_7),
    .io_out(Cell_75_io_out),
    .io_running(Cell_75_io_running),
    .io_writeEnable(Cell_75_io_writeEnable),
    .io_writeValue(Cell_75_io_writeValue)
  );
  Cell Cell_76 ( // @[Life.scala 59:52]
    .clock(Cell_76_clock),
    .reset(Cell_76_reset),
    .io_neighbors_0(Cell_76_io_neighbors_0),
    .io_neighbors_1(Cell_76_io_neighbors_1),
    .io_neighbors_2(Cell_76_io_neighbors_2),
    .io_neighbors_3(Cell_76_io_neighbors_3),
    .io_neighbors_4(Cell_76_io_neighbors_4),
    .io_neighbors_5(Cell_76_io_neighbors_5),
    .io_neighbors_6(Cell_76_io_neighbors_6),
    .io_neighbors_7(Cell_76_io_neighbors_7),
    .io_out(Cell_76_io_out),
    .io_running(Cell_76_io_running),
    .io_writeEnable(Cell_76_io_writeEnable),
    .io_writeValue(Cell_76_io_writeValue)
  );
  Cell Cell_77 ( // @[Life.scala 59:52]
    .clock(Cell_77_clock),
    .reset(Cell_77_reset),
    .io_neighbors_0(Cell_77_io_neighbors_0),
    .io_neighbors_1(Cell_77_io_neighbors_1),
    .io_neighbors_2(Cell_77_io_neighbors_2),
    .io_neighbors_3(Cell_77_io_neighbors_3),
    .io_neighbors_4(Cell_77_io_neighbors_4),
    .io_neighbors_5(Cell_77_io_neighbors_5),
    .io_neighbors_6(Cell_77_io_neighbors_6),
    .io_neighbors_7(Cell_77_io_neighbors_7),
    .io_out(Cell_77_io_out),
    .io_running(Cell_77_io_running),
    .io_writeEnable(Cell_77_io_writeEnable),
    .io_writeValue(Cell_77_io_writeValue)
  );
  Cell Cell_78 ( // @[Life.scala 59:52]
    .clock(Cell_78_clock),
    .reset(Cell_78_reset),
    .io_neighbors_0(Cell_78_io_neighbors_0),
    .io_neighbors_1(Cell_78_io_neighbors_1),
    .io_neighbors_2(Cell_78_io_neighbors_2),
    .io_neighbors_3(Cell_78_io_neighbors_3),
    .io_neighbors_4(Cell_78_io_neighbors_4),
    .io_neighbors_5(Cell_78_io_neighbors_5),
    .io_neighbors_6(Cell_78_io_neighbors_6),
    .io_neighbors_7(Cell_78_io_neighbors_7),
    .io_out(Cell_78_io_out),
    .io_running(Cell_78_io_running),
    .io_writeEnable(Cell_78_io_writeEnable),
    .io_writeValue(Cell_78_io_writeValue)
  );
  Cell Cell_79 ( // @[Life.scala 59:52]
    .clock(Cell_79_clock),
    .reset(Cell_79_reset),
    .io_neighbors_0(Cell_79_io_neighbors_0),
    .io_neighbors_1(Cell_79_io_neighbors_1),
    .io_neighbors_2(Cell_79_io_neighbors_2),
    .io_neighbors_3(Cell_79_io_neighbors_3),
    .io_neighbors_4(Cell_79_io_neighbors_4),
    .io_neighbors_5(Cell_79_io_neighbors_5),
    .io_neighbors_6(Cell_79_io_neighbors_6),
    .io_neighbors_7(Cell_79_io_neighbors_7),
    .io_out(Cell_79_io_out),
    .io_running(Cell_79_io_running),
    .io_writeEnable(Cell_79_io_writeEnable),
    .io_writeValue(Cell_79_io_writeValue)
  );
  Cell Cell_80 ( // @[Life.scala 59:52]
    .clock(Cell_80_clock),
    .reset(Cell_80_reset),
    .io_neighbors_0(Cell_80_io_neighbors_0),
    .io_neighbors_1(Cell_80_io_neighbors_1),
    .io_neighbors_2(Cell_80_io_neighbors_2),
    .io_neighbors_3(Cell_80_io_neighbors_3),
    .io_neighbors_4(Cell_80_io_neighbors_4),
    .io_neighbors_5(Cell_80_io_neighbors_5),
    .io_neighbors_6(Cell_80_io_neighbors_6),
    .io_neighbors_7(Cell_80_io_neighbors_7),
    .io_out(Cell_80_io_out),
    .io_running(Cell_80_io_running),
    .io_writeEnable(Cell_80_io_writeEnable),
    .io_writeValue(Cell_80_io_writeValue)
  );
  Cell Cell_81 ( // @[Life.scala 59:52]
    .clock(Cell_81_clock),
    .reset(Cell_81_reset),
    .io_neighbors_0(Cell_81_io_neighbors_0),
    .io_neighbors_1(Cell_81_io_neighbors_1),
    .io_neighbors_2(Cell_81_io_neighbors_2),
    .io_neighbors_3(Cell_81_io_neighbors_3),
    .io_neighbors_4(Cell_81_io_neighbors_4),
    .io_neighbors_5(Cell_81_io_neighbors_5),
    .io_neighbors_6(Cell_81_io_neighbors_6),
    .io_neighbors_7(Cell_81_io_neighbors_7),
    .io_out(Cell_81_io_out),
    .io_running(Cell_81_io_running),
    .io_writeEnable(Cell_81_io_writeEnable),
    .io_writeValue(Cell_81_io_writeValue)
  );
  Cell Cell_82 ( // @[Life.scala 59:52]
    .clock(Cell_82_clock),
    .reset(Cell_82_reset),
    .io_neighbors_0(Cell_82_io_neighbors_0),
    .io_neighbors_1(Cell_82_io_neighbors_1),
    .io_neighbors_2(Cell_82_io_neighbors_2),
    .io_neighbors_3(Cell_82_io_neighbors_3),
    .io_neighbors_4(Cell_82_io_neighbors_4),
    .io_neighbors_5(Cell_82_io_neighbors_5),
    .io_neighbors_6(Cell_82_io_neighbors_6),
    .io_neighbors_7(Cell_82_io_neighbors_7),
    .io_out(Cell_82_io_out),
    .io_running(Cell_82_io_running),
    .io_writeEnable(Cell_82_io_writeEnable),
    .io_writeValue(Cell_82_io_writeValue)
  );
  Cell Cell_83 ( // @[Life.scala 59:52]
    .clock(Cell_83_clock),
    .reset(Cell_83_reset),
    .io_neighbors_0(Cell_83_io_neighbors_0),
    .io_neighbors_1(Cell_83_io_neighbors_1),
    .io_neighbors_2(Cell_83_io_neighbors_2),
    .io_neighbors_3(Cell_83_io_neighbors_3),
    .io_neighbors_4(Cell_83_io_neighbors_4),
    .io_neighbors_5(Cell_83_io_neighbors_5),
    .io_neighbors_6(Cell_83_io_neighbors_6),
    .io_neighbors_7(Cell_83_io_neighbors_7),
    .io_out(Cell_83_io_out),
    .io_running(Cell_83_io_running),
    .io_writeEnable(Cell_83_io_writeEnable),
    .io_writeValue(Cell_83_io_writeValue)
  );
  Cell Cell_84 ( // @[Life.scala 59:52]
    .clock(Cell_84_clock),
    .reset(Cell_84_reset),
    .io_neighbors_0(Cell_84_io_neighbors_0),
    .io_neighbors_1(Cell_84_io_neighbors_1),
    .io_neighbors_2(Cell_84_io_neighbors_2),
    .io_neighbors_3(Cell_84_io_neighbors_3),
    .io_neighbors_4(Cell_84_io_neighbors_4),
    .io_neighbors_5(Cell_84_io_neighbors_5),
    .io_neighbors_6(Cell_84_io_neighbors_6),
    .io_neighbors_7(Cell_84_io_neighbors_7),
    .io_out(Cell_84_io_out),
    .io_running(Cell_84_io_running),
    .io_writeEnable(Cell_84_io_writeEnable),
    .io_writeValue(Cell_84_io_writeValue)
  );
  Cell Cell_85 ( // @[Life.scala 59:52]
    .clock(Cell_85_clock),
    .reset(Cell_85_reset),
    .io_neighbors_0(Cell_85_io_neighbors_0),
    .io_neighbors_1(Cell_85_io_neighbors_1),
    .io_neighbors_2(Cell_85_io_neighbors_2),
    .io_neighbors_3(Cell_85_io_neighbors_3),
    .io_neighbors_4(Cell_85_io_neighbors_4),
    .io_neighbors_5(Cell_85_io_neighbors_5),
    .io_neighbors_6(Cell_85_io_neighbors_6),
    .io_neighbors_7(Cell_85_io_neighbors_7),
    .io_out(Cell_85_io_out),
    .io_running(Cell_85_io_running),
    .io_writeEnable(Cell_85_io_writeEnable),
    .io_writeValue(Cell_85_io_writeValue)
  );
  Cell Cell_86 ( // @[Life.scala 59:52]
    .clock(Cell_86_clock),
    .reset(Cell_86_reset),
    .io_neighbors_0(Cell_86_io_neighbors_0),
    .io_neighbors_1(Cell_86_io_neighbors_1),
    .io_neighbors_2(Cell_86_io_neighbors_2),
    .io_neighbors_3(Cell_86_io_neighbors_3),
    .io_neighbors_4(Cell_86_io_neighbors_4),
    .io_neighbors_5(Cell_86_io_neighbors_5),
    .io_neighbors_6(Cell_86_io_neighbors_6),
    .io_neighbors_7(Cell_86_io_neighbors_7),
    .io_out(Cell_86_io_out),
    .io_running(Cell_86_io_running),
    .io_writeEnable(Cell_86_io_writeEnable),
    .io_writeValue(Cell_86_io_writeValue)
  );
  Cell Cell_87 ( // @[Life.scala 59:52]
    .clock(Cell_87_clock),
    .reset(Cell_87_reset),
    .io_neighbors_0(Cell_87_io_neighbors_0),
    .io_neighbors_1(Cell_87_io_neighbors_1),
    .io_neighbors_2(Cell_87_io_neighbors_2),
    .io_neighbors_3(Cell_87_io_neighbors_3),
    .io_neighbors_4(Cell_87_io_neighbors_4),
    .io_neighbors_5(Cell_87_io_neighbors_5),
    .io_neighbors_6(Cell_87_io_neighbors_6),
    .io_neighbors_7(Cell_87_io_neighbors_7),
    .io_out(Cell_87_io_out),
    .io_running(Cell_87_io_running),
    .io_writeEnable(Cell_87_io_writeEnable),
    .io_writeValue(Cell_87_io_writeValue)
  );
  Cell Cell_88 ( // @[Life.scala 59:52]
    .clock(Cell_88_clock),
    .reset(Cell_88_reset),
    .io_neighbors_0(Cell_88_io_neighbors_0),
    .io_neighbors_1(Cell_88_io_neighbors_1),
    .io_neighbors_2(Cell_88_io_neighbors_2),
    .io_neighbors_3(Cell_88_io_neighbors_3),
    .io_neighbors_4(Cell_88_io_neighbors_4),
    .io_neighbors_5(Cell_88_io_neighbors_5),
    .io_neighbors_6(Cell_88_io_neighbors_6),
    .io_neighbors_7(Cell_88_io_neighbors_7),
    .io_out(Cell_88_io_out),
    .io_running(Cell_88_io_running),
    .io_writeEnable(Cell_88_io_writeEnable),
    .io_writeValue(Cell_88_io_writeValue)
  );
  Cell Cell_89 ( // @[Life.scala 59:52]
    .clock(Cell_89_clock),
    .reset(Cell_89_reset),
    .io_neighbors_0(Cell_89_io_neighbors_0),
    .io_neighbors_1(Cell_89_io_neighbors_1),
    .io_neighbors_2(Cell_89_io_neighbors_2),
    .io_neighbors_3(Cell_89_io_neighbors_3),
    .io_neighbors_4(Cell_89_io_neighbors_4),
    .io_neighbors_5(Cell_89_io_neighbors_5),
    .io_neighbors_6(Cell_89_io_neighbors_6),
    .io_neighbors_7(Cell_89_io_neighbors_7),
    .io_out(Cell_89_io_out),
    .io_running(Cell_89_io_running),
    .io_writeEnable(Cell_89_io_writeEnable),
    .io_writeValue(Cell_89_io_writeValue)
  );
  Cell Cell_90 ( // @[Life.scala 59:52]
    .clock(Cell_90_clock),
    .reset(Cell_90_reset),
    .io_neighbors_0(Cell_90_io_neighbors_0),
    .io_neighbors_1(Cell_90_io_neighbors_1),
    .io_neighbors_2(Cell_90_io_neighbors_2),
    .io_neighbors_3(Cell_90_io_neighbors_3),
    .io_neighbors_4(Cell_90_io_neighbors_4),
    .io_neighbors_5(Cell_90_io_neighbors_5),
    .io_neighbors_6(Cell_90_io_neighbors_6),
    .io_neighbors_7(Cell_90_io_neighbors_7),
    .io_out(Cell_90_io_out),
    .io_running(Cell_90_io_running),
    .io_writeEnable(Cell_90_io_writeEnable),
    .io_writeValue(Cell_90_io_writeValue)
  );
  Cell Cell_91 ( // @[Life.scala 59:52]
    .clock(Cell_91_clock),
    .reset(Cell_91_reset),
    .io_neighbors_0(Cell_91_io_neighbors_0),
    .io_neighbors_1(Cell_91_io_neighbors_1),
    .io_neighbors_2(Cell_91_io_neighbors_2),
    .io_neighbors_3(Cell_91_io_neighbors_3),
    .io_neighbors_4(Cell_91_io_neighbors_4),
    .io_neighbors_5(Cell_91_io_neighbors_5),
    .io_neighbors_6(Cell_91_io_neighbors_6),
    .io_neighbors_7(Cell_91_io_neighbors_7),
    .io_out(Cell_91_io_out),
    .io_running(Cell_91_io_running),
    .io_writeEnable(Cell_91_io_writeEnable),
    .io_writeValue(Cell_91_io_writeValue)
  );
  Cell Cell_92 ( // @[Life.scala 59:52]
    .clock(Cell_92_clock),
    .reset(Cell_92_reset),
    .io_neighbors_0(Cell_92_io_neighbors_0),
    .io_neighbors_1(Cell_92_io_neighbors_1),
    .io_neighbors_2(Cell_92_io_neighbors_2),
    .io_neighbors_3(Cell_92_io_neighbors_3),
    .io_neighbors_4(Cell_92_io_neighbors_4),
    .io_neighbors_5(Cell_92_io_neighbors_5),
    .io_neighbors_6(Cell_92_io_neighbors_6),
    .io_neighbors_7(Cell_92_io_neighbors_7),
    .io_out(Cell_92_io_out),
    .io_running(Cell_92_io_running),
    .io_writeEnable(Cell_92_io_writeEnable),
    .io_writeValue(Cell_92_io_writeValue)
  );
  Cell Cell_93 ( // @[Life.scala 59:52]
    .clock(Cell_93_clock),
    .reset(Cell_93_reset),
    .io_neighbors_0(Cell_93_io_neighbors_0),
    .io_neighbors_1(Cell_93_io_neighbors_1),
    .io_neighbors_2(Cell_93_io_neighbors_2),
    .io_neighbors_3(Cell_93_io_neighbors_3),
    .io_neighbors_4(Cell_93_io_neighbors_4),
    .io_neighbors_5(Cell_93_io_neighbors_5),
    .io_neighbors_6(Cell_93_io_neighbors_6),
    .io_neighbors_7(Cell_93_io_neighbors_7),
    .io_out(Cell_93_io_out),
    .io_running(Cell_93_io_running),
    .io_writeEnable(Cell_93_io_writeEnable),
    .io_writeValue(Cell_93_io_writeValue)
  );
  Cell Cell_94 ( // @[Life.scala 59:52]
    .clock(Cell_94_clock),
    .reset(Cell_94_reset),
    .io_neighbors_0(Cell_94_io_neighbors_0),
    .io_neighbors_1(Cell_94_io_neighbors_1),
    .io_neighbors_2(Cell_94_io_neighbors_2),
    .io_neighbors_3(Cell_94_io_neighbors_3),
    .io_neighbors_4(Cell_94_io_neighbors_4),
    .io_neighbors_5(Cell_94_io_neighbors_5),
    .io_neighbors_6(Cell_94_io_neighbors_6),
    .io_neighbors_7(Cell_94_io_neighbors_7),
    .io_out(Cell_94_io_out),
    .io_running(Cell_94_io_running),
    .io_writeEnable(Cell_94_io_writeEnable),
    .io_writeValue(Cell_94_io_writeValue)
  );
  Cell Cell_95 ( // @[Life.scala 59:52]
    .clock(Cell_95_clock),
    .reset(Cell_95_reset),
    .io_neighbors_0(Cell_95_io_neighbors_0),
    .io_neighbors_1(Cell_95_io_neighbors_1),
    .io_neighbors_2(Cell_95_io_neighbors_2),
    .io_neighbors_3(Cell_95_io_neighbors_3),
    .io_neighbors_4(Cell_95_io_neighbors_4),
    .io_neighbors_5(Cell_95_io_neighbors_5),
    .io_neighbors_6(Cell_95_io_neighbors_6),
    .io_neighbors_7(Cell_95_io_neighbors_7),
    .io_out(Cell_95_io_out),
    .io_running(Cell_95_io_running),
    .io_writeEnable(Cell_95_io_writeEnable),
    .io_writeValue(Cell_95_io_writeValue)
  );
  Cell Cell_96 ( // @[Life.scala 59:52]
    .clock(Cell_96_clock),
    .reset(Cell_96_reset),
    .io_neighbors_0(Cell_96_io_neighbors_0),
    .io_neighbors_1(Cell_96_io_neighbors_1),
    .io_neighbors_2(Cell_96_io_neighbors_2),
    .io_neighbors_3(Cell_96_io_neighbors_3),
    .io_neighbors_4(Cell_96_io_neighbors_4),
    .io_neighbors_5(Cell_96_io_neighbors_5),
    .io_neighbors_6(Cell_96_io_neighbors_6),
    .io_neighbors_7(Cell_96_io_neighbors_7),
    .io_out(Cell_96_io_out),
    .io_running(Cell_96_io_running),
    .io_writeEnable(Cell_96_io_writeEnable),
    .io_writeValue(Cell_96_io_writeValue)
  );
  Cell Cell_97 ( // @[Life.scala 59:52]
    .clock(Cell_97_clock),
    .reset(Cell_97_reset),
    .io_neighbors_0(Cell_97_io_neighbors_0),
    .io_neighbors_1(Cell_97_io_neighbors_1),
    .io_neighbors_2(Cell_97_io_neighbors_2),
    .io_neighbors_3(Cell_97_io_neighbors_3),
    .io_neighbors_4(Cell_97_io_neighbors_4),
    .io_neighbors_5(Cell_97_io_neighbors_5),
    .io_neighbors_6(Cell_97_io_neighbors_6),
    .io_neighbors_7(Cell_97_io_neighbors_7),
    .io_out(Cell_97_io_out),
    .io_running(Cell_97_io_running),
    .io_writeEnable(Cell_97_io_writeEnable),
    .io_writeValue(Cell_97_io_writeValue)
  );
  Cell Cell_98 ( // @[Life.scala 59:52]
    .clock(Cell_98_clock),
    .reset(Cell_98_reset),
    .io_neighbors_0(Cell_98_io_neighbors_0),
    .io_neighbors_1(Cell_98_io_neighbors_1),
    .io_neighbors_2(Cell_98_io_neighbors_2),
    .io_neighbors_3(Cell_98_io_neighbors_3),
    .io_neighbors_4(Cell_98_io_neighbors_4),
    .io_neighbors_5(Cell_98_io_neighbors_5),
    .io_neighbors_6(Cell_98_io_neighbors_6),
    .io_neighbors_7(Cell_98_io_neighbors_7),
    .io_out(Cell_98_io_out),
    .io_running(Cell_98_io_running),
    .io_writeEnable(Cell_98_io_writeEnable),
    .io_writeValue(Cell_98_io_writeValue)
  );
  Cell Cell_99 ( // @[Life.scala 59:52]
    .clock(Cell_99_clock),
    .reset(Cell_99_reset),
    .io_neighbors_0(Cell_99_io_neighbors_0),
    .io_neighbors_1(Cell_99_io_neighbors_1),
    .io_neighbors_2(Cell_99_io_neighbors_2),
    .io_neighbors_3(Cell_99_io_neighbors_3),
    .io_neighbors_4(Cell_99_io_neighbors_4),
    .io_neighbors_5(Cell_99_io_neighbors_5),
    .io_neighbors_6(Cell_99_io_neighbors_6),
    .io_neighbors_7(Cell_99_io_neighbors_7),
    .io_out(Cell_99_io_out),
    .io_running(Cell_99_io_running),
    .io_writeEnable(Cell_99_io_writeEnable),
    .io_writeValue(Cell_99_io_writeValue)
  );
  Cell Cell_100 ( // @[Life.scala 59:52]
    .clock(Cell_100_clock),
    .reset(Cell_100_reset),
    .io_neighbors_0(Cell_100_io_neighbors_0),
    .io_neighbors_1(Cell_100_io_neighbors_1),
    .io_neighbors_2(Cell_100_io_neighbors_2),
    .io_neighbors_3(Cell_100_io_neighbors_3),
    .io_neighbors_4(Cell_100_io_neighbors_4),
    .io_neighbors_5(Cell_100_io_neighbors_5),
    .io_neighbors_6(Cell_100_io_neighbors_6),
    .io_neighbors_7(Cell_100_io_neighbors_7),
    .io_out(Cell_100_io_out),
    .io_running(Cell_100_io_running),
    .io_writeEnable(Cell_100_io_writeEnable),
    .io_writeValue(Cell_100_io_writeValue)
  );
  Cell Cell_101 ( // @[Life.scala 59:52]
    .clock(Cell_101_clock),
    .reset(Cell_101_reset),
    .io_neighbors_0(Cell_101_io_neighbors_0),
    .io_neighbors_1(Cell_101_io_neighbors_1),
    .io_neighbors_2(Cell_101_io_neighbors_2),
    .io_neighbors_3(Cell_101_io_neighbors_3),
    .io_neighbors_4(Cell_101_io_neighbors_4),
    .io_neighbors_5(Cell_101_io_neighbors_5),
    .io_neighbors_6(Cell_101_io_neighbors_6),
    .io_neighbors_7(Cell_101_io_neighbors_7),
    .io_out(Cell_101_io_out),
    .io_running(Cell_101_io_running),
    .io_writeEnable(Cell_101_io_writeEnable),
    .io_writeValue(Cell_101_io_writeValue)
  );
  Cell Cell_102 ( // @[Life.scala 59:52]
    .clock(Cell_102_clock),
    .reset(Cell_102_reset),
    .io_neighbors_0(Cell_102_io_neighbors_0),
    .io_neighbors_1(Cell_102_io_neighbors_1),
    .io_neighbors_2(Cell_102_io_neighbors_2),
    .io_neighbors_3(Cell_102_io_neighbors_3),
    .io_neighbors_4(Cell_102_io_neighbors_4),
    .io_neighbors_5(Cell_102_io_neighbors_5),
    .io_neighbors_6(Cell_102_io_neighbors_6),
    .io_neighbors_7(Cell_102_io_neighbors_7),
    .io_out(Cell_102_io_out),
    .io_running(Cell_102_io_running),
    .io_writeEnable(Cell_102_io_writeEnable),
    .io_writeValue(Cell_102_io_writeValue)
  );
  Cell Cell_103 ( // @[Life.scala 59:52]
    .clock(Cell_103_clock),
    .reset(Cell_103_reset),
    .io_neighbors_0(Cell_103_io_neighbors_0),
    .io_neighbors_1(Cell_103_io_neighbors_1),
    .io_neighbors_2(Cell_103_io_neighbors_2),
    .io_neighbors_3(Cell_103_io_neighbors_3),
    .io_neighbors_4(Cell_103_io_neighbors_4),
    .io_neighbors_5(Cell_103_io_neighbors_5),
    .io_neighbors_6(Cell_103_io_neighbors_6),
    .io_neighbors_7(Cell_103_io_neighbors_7),
    .io_out(Cell_103_io_out),
    .io_running(Cell_103_io_running),
    .io_writeEnable(Cell_103_io_writeEnable),
    .io_writeValue(Cell_103_io_writeValue)
  );
  Cell Cell_104 ( // @[Life.scala 59:52]
    .clock(Cell_104_clock),
    .reset(Cell_104_reset),
    .io_neighbors_0(Cell_104_io_neighbors_0),
    .io_neighbors_1(Cell_104_io_neighbors_1),
    .io_neighbors_2(Cell_104_io_neighbors_2),
    .io_neighbors_3(Cell_104_io_neighbors_3),
    .io_neighbors_4(Cell_104_io_neighbors_4),
    .io_neighbors_5(Cell_104_io_neighbors_5),
    .io_neighbors_6(Cell_104_io_neighbors_6),
    .io_neighbors_7(Cell_104_io_neighbors_7),
    .io_out(Cell_104_io_out),
    .io_running(Cell_104_io_running),
    .io_writeEnable(Cell_104_io_writeEnable),
    .io_writeValue(Cell_104_io_writeValue)
  );
  Cell Cell_105 ( // @[Life.scala 59:52]
    .clock(Cell_105_clock),
    .reset(Cell_105_reset),
    .io_neighbors_0(Cell_105_io_neighbors_0),
    .io_neighbors_1(Cell_105_io_neighbors_1),
    .io_neighbors_2(Cell_105_io_neighbors_2),
    .io_neighbors_3(Cell_105_io_neighbors_3),
    .io_neighbors_4(Cell_105_io_neighbors_4),
    .io_neighbors_5(Cell_105_io_neighbors_5),
    .io_neighbors_6(Cell_105_io_neighbors_6),
    .io_neighbors_7(Cell_105_io_neighbors_7),
    .io_out(Cell_105_io_out),
    .io_running(Cell_105_io_running),
    .io_writeEnable(Cell_105_io_writeEnable),
    .io_writeValue(Cell_105_io_writeValue)
  );
  Cell Cell_106 ( // @[Life.scala 59:52]
    .clock(Cell_106_clock),
    .reset(Cell_106_reset),
    .io_neighbors_0(Cell_106_io_neighbors_0),
    .io_neighbors_1(Cell_106_io_neighbors_1),
    .io_neighbors_2(Cell_106_io_neighbors_2),
    .io_neighbors_3(Cell_106_io_neighbors_3),
    .io_neighbors_4(Cell_106_io_neighbors_4),
    .io_neighbors_5(Cell_106_io_neighbors_5),
    .io_neighbors_6(Cell_106_io_neighbors_6),
    .io_neighbors_7(Cell_106_io_neighbors_7),
    .io_out(Cell_106_io_out),
    .io_running(Cell_106_io_running),
    .io_writeEnable(Cell_106_io_writeEnable),
    .io_writeValue(Cell_106_io_writeValue)
  );
  Cell Cell_107 ( // @[Life.scala 59:52]
    .clock(Cell_107_clock),
    .reset(Cell_107_reset),
    .io_neighbors_0(Cell_107_io_neighbors_0),
    .io_neighbors_1(Cell_107_io_neighbors_1),
    .io_neighbors_2(Cell_107_io_neighbors_2),
    .io_neighbors_3(Cell_107_io_neighbors_3),
    .io_neighbors_4(Cell_107_io_neighbors_4),
    .io_neighbors_5(Cell_107_io_neighbors_5),
    .io_neighbors_6(Cell_107_io_neighbors_6),
    .io_neighbors_7(Cell_107_io_neighbors_7),
    .io_out(Cell_107_io_out),
    .io_running(Cell_107_io_running),
    .io_writeEnable(Cell_107_io_writeEnable),
    .io_writeValue(Cell_107_io_writeValue)
  );
  Cell Cell_108 ( // @[Life.scala 59:52]
    .clock(Cell_108_clock),
    .reset(Cell_108_reset),
    .io_neighbors_0(Cell_108_io_neighbors_0),
    .io_neighbors_1(Cell_108_io_neighbors_1),
    .io_neighbors_2(Cell_108_io_neighbors_2),
    .io_neighbors_3(Cell_108_io_neighbors_3),
    .io_neighbors_4(Cell_108_io_neighbors_4),
    .io_neighbors_5(Cell_108_io_neighbors_5),
    .io_neighbors_6(Cell_108_io_neighbors_6),
    .io_neighbors_7(Cell_108_io_neighbors_7),
    .io_out(Cell_108_io_out),
    .io_running(Cell_108_io_running),
    .io_writeEnable(Cell_108_io_writeEnable),
    .io_writeValue(Cell_108_io_writeValue)
  );
  Cell Cell_109 ( // @[Life.scala 59:52]
    .clock(Cell_109_clock),
    .reset(Cell_109_reset),
    .io_neighbors_0(Cell_109_io_neighbors_0),
    .io_neighbors_1(Cell_109_io_neighbors_1),
    .io_neighbors_2(Cell_109_io_neighbors_2),
    .io_neighbors_3(Cell_109_io_neighbors_3),
    .io_neighbors_4(Cell_109_io_neighbors_4),
    .io_neighbors_5(Cell_109_io_neighbors_5),
    .io_neighbors_6(Cell_109_io_neighbors_6),
    .io_neighbors_7(Cell_109_io_neighbors_7),
    .io_out(Cell_109_io_out),
    .io_running(Cell_109_io_running),
    .io_writeEnable(Cell_109_io_writeEnable),
    .io_writeValue(Cell_109_io_writeValue)
  );
  Cell Cell_110 ( // @[Life.scala 59:52]
    .clock(Cell_110_clock),
    .reset(Cell_110_reset),
    .io_neighbors_0(Cell_110_io_neighbors_0),
    .io_neighbors_1(Cell_110_io_neighbors_1),
    .io_neighbors_2(Cell_110_io_neighbors_2),
    .io_neighbors_3(Cell_110_io_neighbors_3),
    .io_neighbors_4(Cell_110_io_neighbors_4),
    .io_neighbors_5(Cell_110_io_neighbors_5),
    .io_neighbors_6(Cell_110_io_neighbors_6),
    .io_neighbors_7(Cell_110_io_neighbors_7),
    .io_out(Cell_110_io_out),
    .io_running(Cell_110_io_running),
    .io_writeEnable(Cell_110_io_writeEnable),
    .io_writeValue(Cell_110_io_writeValue)
  );
  Cell Cell_111 ( // @[Life.scala 59:52]
    .clock(Cell_111_clock),
    .reset(Cell_111_reset),
    .io_neighbors_0(Cell_111_io_neighbors_0),
    .io_neighbors_1(Cell_111_io_neighbors_1),
    .io_neighbors_2(Cell_111_io_neighbors_2),
    .io_neighbors_3(Cell_111_io_neighbors_3),
    .io_neighbors_4(Cell_111_io_neighbors_4),
    .io_neighbors_5(Cell_111_io_neighbors_5),
    .io_neighbors_6(Cell_111_io_neighbors_6),
    .io_neighbors_7(Cell_111_io_neighbors_7),
    .io_out(Cell_111_io_out),
    .io_running(Cell_111_io_running),
    .io_writeEnable(Cell_111_io_writeEnable),
    .io_writeValue(Cell_111_io_writeValue)
  );
  Cell Cell_112 ( // @[Life.scala 59:52]
    .clock(Cell_112_clock),
    .reset(Cell_112_reset),
    .io_neighbors_0(Cell_112_io_neighbors_0),
    .io_neighbors_1(Cell_112_io_neighbors_1),
    .io_neighbors_2(Cell_112_io_neighbors_2),
    .io_neighbors_3(Cell_112_io_neighbors_3),
    .io_neighbors_4(Cell_112_io_neighbors_4),
    .io_neighbors_5(Cell_112_io_neighbors_5),
    .io_neighbors_6(Cell_112_io_neighbors_6),
    .io_neighbors_7(Cell_112_io_neighbors_7),
    .io_out(Cell_112_io_out),
    .io_running(Cell_112_io_running),
    .io_writeEnable(Cell_112_io_writeEnable),
    .io_writeValue(Cell_112_io_writeValue)
  );
  Cell Cell_113 ( // @[Life.scala 59:52]
    .clock(Cell_113_clock),
    .reset(Cell_113_reset),
    .io_neighbors_0(Cell_113_io_neighbors_0),
    .io_neighbors_1(Cell_113_io_neighbors_1),
    .io_neighbors_2(Cell_113_io_neighbors_2),
    .io_neighbors_3(Cell_113_io_neighbors_3),
    .io_neighbors_4(Cell_113_io_neighbors_4),
    .io_neighbors_5(Cell_113_io_neighbors_5),
    .io_neighbors_6(Cell_113_io_neighbors_6),
    .io_neighbors_7(Cell_113_io_neighbors_7),
    .io_out(Cell_113_io_out),
    .io_running(Cell_113_io_running),
    .io_writeEnable(Cell_113_io_writeEnable),
    .io_writeValue(Cell_113_io_writeValue)
  );
  Cell Cell_114 ( // @[Life.scala 59:52]
    .clock(Cell_114_clock),
    .reset(Cell_114_reset),
    .io_neighbors_0(Cell_114_io_neighbors_0),
    .io_neighbors_1(Cell_114_io_neighbors_1),
    .io_neighbors_2(Cell_114_io_neighbors_2),
    .io_neighbors_3(Cell_114_io_neighbors_3),
    .io_neighbors_4(Cell_114_io_neighbors_4),
    .io_neighbors_5(Cell_114_io_neighbors_5),
    .io_neighbors_6(Cell_114_io_neighbors_6),
    .io_neighbors_7(Cell_114_io_neighbors_7),
    .io_out(Cell_114_io_out),
    .io_running(Cell_114_io_running),
    .io_writeEnable(Cell_114_io_writeEnable),
    .io_writeValue(Cell_114_io_writeValue)
  );
  Cell Cell_115 ( // @[Life.scala 59:52]
    .clock(Cell_115_clock),
    .reset(Cell_115_reset),
    .io_neighbors_0(Cell_115_io_neighbors_0),
    .io_neighbors_1(Cell_115_io_neighbors_1),
    .io_neighbors_2(Cell_115_io_neighbors_2),
    .io_neighbors_3(Cell_115_io_neighbors_3),
    .io_neighbors_4(Cell_115_io_neighbors_4),
    .io_neighbors_5(Cell_115_io_neighbors_5),
    .io_neighbors_6(Cell_115_io_neighbors_6),
    .io_neighbors_7(Cell_115_io_neighbors_7),
    .io_out(Cell_115_io_out),
    .io_running(Cell_115_io_running),
    .io_writeEnable(Cell_115_io_writeEnable),
    .io_writeValue(Cell_115_io_writeValue)
  );
  Cell Cell_116 ( // @[Life.scala 59:52]
    .clock(Cell_116_clock),
    .reset(Cell_116_reset),
    .io_neighbors_0(Cell_116_io_neighbors_0),
    .io_neighbors_1(Cell_116_io_neighbors_1),
    .io_neighbors_2(Cell_116_io_neighbors_2),
    .io_neighbors_3(Cell_116_io_neighbors_3),
    .io_neighbors_4(Cell_116_io_neighbors_4),
    .io_neighbors_5(Cell_116_io_neighbors_5),
    .io_neighbors_6(Cell_116_io_neighbors_6),
    .io_neighbors_7(Cell_116_io_neighbors_7),
    .io_out(Cell_116_io_out),
    .io_running(Cell_116_io_running),
    .io_writeEnable(Cell_116_io_writeEnable),
    .io_writeValue(Cell_116_io_writeValue)
  );
  Cell Cell_117 ( // @[Life.scala 59:52]
    .clock(Cell_117_clock),
    .reset(Cell_117_reset),
    .io_neighbors_0(Cell_117_io_neighbors_0),
    .io_neighbors_1(Cell_117_io_neighbors_1),
    .io_neighbors_2(Cell_117_io_neighbors_2),
    .io_neighbors_3(Cell_117_io_neighbors_3),
    .io_neighbors_4(Cell_117_io_neighbors_4),
    .io_neighbors_5(Cell_117_io_neighbors_5),
    .io_neighbors_6(Cell_117_io_neighbors_6),
    .io_neighbors_7(Cell_117_io_neighbors_7),
    .io_out(Cell_117_io_out),
    .io_running(Cell_117_io_running),
    .io_writeEnable(Cell_117_io_writeEnable),
    .io_writeValue(Cell_117_io_writeValue)
  );
  Cell Cell_118 ( // @[Life.scala 59:52]
    .clock(Cell_118_clock),
    .reset(Cell_118_reset),
    .io_neighbors_0(Cell_118_io_neighbors_0),
    .io_neighbors_1(Cell_118_io_neighbors_1),
    .io_neighbors_2(Cell_118_io_neighbors_2),
    .io_neighbors_3(Cell_118_io_neighbors_3),
    .io_neighbors_4(Cell_118_io_neighbors_4),
    .io_neighbors_5(Cell_118_io_neighbors_5),
    .io_neighbors_6(Cell_118_io_neighbors_6),
    .io_neighbors_7(Cell_118_io_neighbors_7),
    .io_out(Cell_118_io_out),
    .io_running(Cell_118_io_running),
    .io_writeEnable(Cell_118_io_writeEnable),
    .io_writeValue(Cell_118_io_writeValue)
  );
  Cell Cell_119 ( // @[Life.scala 59:52]
    .clock(Cell_119_clock),
    .reset(Cell_119_reset),
    .io_neighbors_0(Cell_119_io_neighbors_0),
    .io_neighbors_1(Cell_119_io_neighbors_1),
    .io_neighbors_2(Cell_119_io_neighbors_2),
    .io_neighbors_3(Cell_119_io_neighbors_3),
    .io_neighbors_4(Cell_119_io_neighbors_4),
    .io_neighbors_5(Cell_119_io_neighbors_5),
    .io_neighbors_6(Cell_119_io_neighbors_6),
    .io_neighbors_7(Cell_119_io_neighbors_7),
    .io_out(Cell_119_io_out),
    .io_running(Cell_119_io_running),
    .io_writeEnable(Cell_119_io_writeEnable),
    .io_writeValue(Cell_119_io_writeValue)
  );
  Cell Cell_120 ( // @[Life.scala 59:52]
    .clock(Cell_120_clock),
    .reset(Cell_120_reset),
    .io_neighbors_0(Cell_120_io_neighbors_0),
    .io_neighbors_1(Cell_120_io_neighbors_1),
    .io_neighbors_2(Cell_120_io_neighbors_2),
    .io_neighbors_3(Cell_120_io_neighbors_3),
    .io_neighbors_4(Cell_120_io_neighbors_4),
    .io_neighbors_5(Cell_120_io_neighbors_5),
    .io_neighbors_6(Cell_120_io_neighbors_6),
    .io_neighbors_7(Cell_120_io_neighbors_7),
    .io_out(Cell_120_io_out),
    .io_running(Cell_120_io_running),
    .io_writeEnable(Cell_120_io_writeEnable),
    .io_writeValue(Cell_120_io_writeValue)
  );
  Cell Cell_121 ( // @[Life.scala 59:52]
    .clock(Cell_121_clock),
    .reset(Cell_121_reset),
    .io_neighbors_0(Cell_121_io_neighbors_0),
    .io_neighbors_1(Cell_121_io_neighbors_1),
    .io_neighbors_2(Cell_121_io_neighbors_2),
    .io_neighbors_3(Cell_121_io_neighbors_3),
    .io_neighbors_4(Cell_121_io_neighbors_4),
    .io_neighbors_5(Cell_121_io_neighbors_5),
    .io_neighbors_6(Cell_121_io_neighbors_6),
    .io_neighbors_7(Cell_121_io_neighbors_7),
    .io_out(Cell_121_io_out),
    .io_running(Cell_121_io_running),
    .io_writeEnable(Cell_121_io_writeEnable),
    .io_writeValue(Cell_121_io_writeValue)
  );
  Cell Cell_122 ( // @[Life.scala 59:52]
    .clock(Cell_122_clock),
    .reset(Cell_122_reset),
    .io_neighbors_0(Cell_122_io_neighbors_0),
    .io_neighbors_1(Cell_122_io_neighbors_1),
    .io_neighbors_2(Cell_122_io_neighbors_2),
    .io_neighbors_3(Cell_122_io_neighbors_3),
    .io_neighbors_4(Cell_122_io_neighbors_4),
    .io_neighbors_5(Cell_122_io_neighbors_5),
    .io_neighbors_6(Cell_122_io_neighbors_6),
    .io_neighbors_7(Cell_122_io_neighbors_7),
    .io_out(Cell_122_io_out),
    .io_running(Cell_122_io_running),
    .io_writeEnable(Cell_122_io_writeEnable),
    .io_writeValue(Cell_122_io_writeValue)
  );
  Cell Cell_123 ( // @[Life.scala 59:52]
    .clock(Cell_123_clock),
    .reset(Cell_123_reset),
    .io_neighbors_0(Cell_123_io_neighbors_0),
    .io_neighbors_1(Cell_123_io_neighbors_1),
    .io_neighbors_2(Cell_123_io_neighbors_2),
    .io_neighbors_3(Cell_123_io_neighbors_3),
    .io_neighbors_4(Cell_123_io_neighbors_4),
    .io_neighbors_5(Cell_123_io_neighbors_5),
    .io_neighbors_6(Cell_123_io_neighbors_6),
    .io_neighbors_7(Cell_123_io_neighbors_7),
    .io_out(Cell_123_io_out),
    .io_running(Cell_123_io_running),
    .io_writeEnable(Cell_123_io_writeEnable),
    .io_writeValue(Cell_123_io_writeValue)
  );
  Cell Cell_124 ( // @[Life.scala 59:52]
    .clock(Cell_124_clock),
    .reset(Cell_124_reset),
    .io_neighbors_0(Cell_124_io_neighbors_0),
    .io_neighbors_1(Cell_124_io_neighbors_1),
    .io_neighbors_2(Cell_124_io_neighbors_2),
    .io_neighbors_3(Cell_124_io_neighbors_3),
    .io_neighbors_4(Cell_124_io_neighbors_4),
    .io_neighbors_5(Cell_124_io_neighbors_5),
    .io_neighbors_6(Cell_124_io_neighbors_6),
    .io_neighbors_7(Cell_124_io_neighbors_7),
    .io_out(Cell_124_io_out),
    .io_running(Cell_124_io_running),
    .io_writeEnable(Cell_124_io_writeEnable),
    .io_writeValue(Cell_124_io_writeValue)
  );
  Cell Cell_125 ( // @[Life.scala 59:52]
    .clock(Cell_125_clock),
    .reset(Cell_125_reset),
    .io_neighbors_0(Cell_125_io_neighbors_0),
    .io_neighbors_1(Cell_125_io_neighbors_1),
    .io_neighbors_2(Cell_125_io_neighbors_2),
    .io_neighbors_3(Cell_125_io_neighbors_3),
    .io_neighbors_4(Cell_125_io_neighbors_4),
    .io_neighbors_5(Cell_125_io_neighbors_5),
    .io_neighbors_6(Cell_125_io_neighbors_6),
    .io_neighbors_7(Cell_125_io_neighbors_7),
    .io_out(Cell_125_io_out),
    .io_running(Cell_125_io_running),
    .io_writeEnable(Cell_125_io_writeEnable),
    .io_writeValue(Cell_125_io_writeValue)
  );
  Cell Cell_126 ( // @[Life.scala 59:52]
    .clock(Cell_126_clock),
    .reset(Cell_126_reset),
    .io_neighbors_0(Cell_126_io_neighbors_0),
    .io_neighbors_1(Cell_126_io_neighbors_1),
    .io_neighbors_2(Cell_126_io_neighbors_2),
    .io_neighbors_3(Cell_126_io_neighbors_3),
    .io_neighbors_4(Cell_126_io_neighbors_4),
    .io_neighbors_5(Cell_126_io_neighbors_5),
    .io_neighbors_6(Cell_126_io_neighbors_6),
    .io_neighbors_7(Cell_126_io_neighbors_7),
    .io_out(Cell_126_io_out),
    .io_running(Cell_126_io_running),
    .io_writeEnable(Cell_126_io_writeEnable),
    .io_writeValue(Cell_126_io_writeValue)
  );
  Cell Cell_127 ( // @[Life.scala 59:52]
    .clock(Cell_127_clock),
    .reset(Cell_127_reset),
    .io_neighbors_0(Cell_127_io_neighbors_0),
    .io_neighbors_1(Cell_127_io_neighbors_1),
    .io_neighbors_2(Cell_127_io_neighbors_2),
    .io_neighbors_3(Cell_127_io_neighbors_3),
    .io_neighbors_4(Cell_127_io_neighbors_4),
    .io_neighbors_5(Cell_127_io_neighbors_5),
    .io_neighbors_6(Cell_127_io_neighbors_6),
    .io_neighbors_7(Cell_127_io_neighbors_7),
    .io_out(Cell_127_io_out),
    .io_running(Cell_127_io_running),
    .io_writeEnable(Cell_127_io_writeEnable),
    .io_writeValue(Cell_127_io_writeValue)
  );
  Cell Cell_128 ( // @[Life.scala 59:52]
    .clock(Cell_128_clock),
    .reset(Cell_128_reset),
    .io_neighbors_0(Cell_128_io_neighbors_0),
    .io_neighbors_1(Cell_128_io_neighbors_1),
    .io_neighbors_2(Cell_128_io_neighbors_2),
    .io_neighbors_3(Cell_128_io_neighbors_3),
    .io_neighbors_4(Cell_128_io_neighbors_4),
    .io_neighbors_5(Cell_128_io_neighbors_5),
    .io_neighbors_6(Cell_128_io_neighbors_6),
    .io_neighbors_7(Cell_128_io_neighbors_7),
    .io_out(Cell_128_io_out),
    .io_running(Cell_128_io_running),
    .io_writeEnable(Cell_128_io_writeEnable),
    .io_writeValue(Cell_128_io_writeValue)
  );
  Cell Cell_129 ( // @[Life.scala 59:52]
    .clock(Cell_129_clock),
    .reset(Cell_129_reset),
    .io_neighbors_0(Cell_129_io_neighbors_0),
    .io_neighbors_1(Cell_129_io_neighbors_1),
    .io_neighbors_2(Cell_129_io_neighbors_2),
    .io_neighbors_3(Cell_129_io_neighbors_3),
    .io_neighbors_4(Cell_129_io_neighbors_4),
    .io_neighbors_5(Cell_129_io_neighbors_5),
    .io_neighbors_6(Cell_129_io_neighbors_6),
    .io_neighbors_7(Cell_129_io_neighbors_7),
    .io_out(Cell_129_io_out),
    .io_running(Cell_129_io_running),
    .io_writeEnable(Cell_129_io_writeEnable),
    .io_writeValue(Cell_129_io_writeValue)
  );
  Cell Cell_130 ( // @[Life.scala 59:52]
    .clock(Cell_130_clock),
    .reset(Cell_130_reset),
    .io_neighbors_0(Cell_130_io_neighbors_0),
    .io_neighbors_1(Cell_130_io_neighbors_1),
    .io_neighbors_2(Cell_130_io_neighbors_2),
    .io_neighbors_3(Cell_130_io_neighbors_3),
    .io_neighbors_4(Cell_130_io_neighbors_4),
    .io_neighbors_5(Cell_130_io_neighbors_5),
    .io_neighbors_6(Cell_130_io_neighbors_6),
    .io_neighbors_7(Cell_130_io_neighbors_7),
    .io_out(Cell_130_io_out),
    .io_running(Cell_130_io_running),
    .io_writeEnable(Cell_130_io_writeEnable),
    .io_writeValue(Cell_130_io_writeValue)
  );
  Cell Cell_131 ( // @[Life.scala 59:52]
    .clock(Cell_131_clock),
    .reset(Cell_131_reset),
    .io_neighbors_0(Cell_131_io_neighbors_0),
    .io_neighbors_1(Cell_131_io_neighbors_1),
    .io_neighbors_2(Cell_131_io_neighbors_2),
    .io_neighbors_3(Cell_131_io_neighbors_3),
    .io_neighbors_4(Cell_131_io_neighbors_4),
    .io_neighbors_5(Cell_131_io_neighbors_5),
    .io_neighbors_6(Cell_131_io_neighbors_6),
    .io_neighbors_7(Cell_131_io_neighbors_7),
    .io_out(Cell_131_io_out),
    .io_running(Cell_131_io_running),
    .io_writeEnable(Cell_131_io_writeEnable),
    .io_writeValue(Cell_131_io_writeValue)
  );
  Cell Cell_132 ( // @[Life.scala 59:52]
    .clock(Cell_132_clock),
    .reset(Cell_132_reset),
    .io_neighbors_0(Cell_132_io_neighbors_0),
    .io_neighbors_1(Cell_132_io_neighbors_1),
    .io_neighbors_2(Cell_132_io_neighbors_2),
    .io_neighbors_3(Cell_132_io_neighbors_3),
    .io_neighbors_4(Cell_132_io_neighbors_4),
    .io_neighbors_5(Cell_132_io_neighbors_5),
    .io_neighbors_6(Cell_132_io_neighbors_6),
    .io_neighbors_7(Cell_132_io_neighbors_7),
    .io_out(Cell_132_io_out),
    .io_running(Cell_132_io_running),
    .io_writeEnable(Cell_132_io_writeEnable),
    .io_writeValue(Cell_132_io_writeValue)
  );
  Cell Cell_133 ( // @[Life.scala 59:52]
    .clock(Cell_133_clock),
    .reset(Cell_133_reset),
    .io_neighbors_0(Cell_133_io_neighbors_0),
    .io_neighbors_1(Cell_133_io_neighbors_1),
    .io_neighbors_2(Cell_133_io_neighbors_2),
    .io_neighbors_3(Cell_133_io_neighbors_3),
    .io_neighbors_4(Cell_133_io_neighbors_4),
    .io_neighbors_5(Cell_133_io_neighbors_5),
    .io_neighbors_6(Cell_133_io_neighbors_6),
    .io_neighbors_7(Cell_133_io_neighbors_7),
    .io_out(Cell_133_io_out),
    .io_running(Cell_133_io_running),
    .io_writeEnable(Cell_133_io_writeEnable),
    .io_writeValue(Cell_133_io_writeValue)
  );
  Cell Cell_134 ( // @[Life.scala 59:52]
    .clock(Cell_134_clock),
    .reset(Cell_134_reset),
    .io_neighbors_0(Cell_134_io_neighbors_0),
    .io_neighbors_1(Cell_134_io_neighbors_1),
    .io_neighbors_2(Cell_134_io_neighbors_2),
    .io_neighbors_3(Cell_134_io_neighbors_3),
    .io_neighbors_4(Cell_134_io_neighbors_4),
    .io_neighbors_5(Cell_134_io_neighbors_5),
    .io_neighbors_6(Cell_134_io_neighbors_6),
    .io_neighbors_7(Cell_134_io_neighbors_7),
    .io_out(Cell_134_io_out),
    .io_running(Cell_134_io_running),
    .io_writeEnable(Cell_134_io_writeEnable),
    .io_writeValue(Cell_134_io_writeValue)
  );
  Cell Cell_135 ( // @[Life.scala 59:52]
    .clock(Cell_135_clock),
    .reset(Cell_135_reset),
    .io_neighbors_0(Cell_135_io_neighbors_0),
    .io_neighbors_1(Cell_135_io_neighbors_1),
    .io_neighbors_2(Cell_135_io_neighbors_2),
    .io_neighbors_3(Cell_135_io_neighbors_3),
    .io_neighbors_4(Cell_135_io_neighbors_4),
    .io_neighbors_5(Cell_135_io_neighbors_5),
    .io_neighbors_6(Cell_135_io_neighbors_6),
    .io_neighbors_7(Cell_135_io_neighbors_7),
    .io_out(Cell_135_io_out),
    .io_running(Cell_135_io_running),
    .io_writeEnable(Cell_135_io_writeEnable),
    .io_writeValue(Cell_135_io_writeValue)
  );
  Cell Cell_136 ( // @[Life.scala 59:52]
    .clock(Cell_136_clock),
    .reset(Cell_136_reset),
    .io_neighbors_0(Cell_136_io_neighbors_0),
    .io_neighbors_1(Cell_136_io_neighbors_1),
    .io_neighbors_2(Cell_136_io_neighbors_2),
    .io_neighbors_3(Cell_136_io_neighbors_3),
    .io_neighbors_4(Cell_136_io_neighbors_4),
    .io_neighbors_5(Cell_136_io_neighbors_5),
    .io_neighbors_6(Cell_136_io_neighbors_6),
    .io_neighbors_7(Cell_136_io_neighbors_7),
    .io_out(Cell_136_io_out),
    .io_running(Cell_136_io_running),
    .io_writeEnable(Cell_136_io_writeEnable),
    .io_writeValue(Cell_136_io_writeValue)
  );
  Cell Cell_137 ( // @[Life.scala 59:52]
    .clock(Cell_137_clock),
    .reset(Cell_137_reset),
    .io_neighbors_0(Cell_137_io_neighbors_0),
    .io_neighbors_1(Cell_137_io_neighbors_1),
    .io_neighbors_2(Cell_137_io_neighbors_2),
    .io_neighbors_3(Cell_137_io_neighbors_3),
    .io_neighbors_4(Cell_137_io_neighbors_4),
    .io_neighbors_5(Cell_137_io_neighbors_5),
    .io_neighbors_6(Cell_137_io_neighbors_6),
    .io_neighbors_7(Cell_137_io_neighbors_7),
    .io_out(Cell_137_io_out),
    .io_running(Cell_137_io_running),
    .io_writeEnable(Cell_137_io_writeEnable),
    .io_writeValue(Cell_137_io_writeValue)
  );
  Cell Cell_138 ( // @[Life.scala 59:52]
    .clock(Cell_138_clock),
    .reset(Cell_138_reset),
    .io_neighbors_0(Cell_138_io_neighbors_0),
    .io_neighbors_1(Cell_138_io_neighbors_1),
    .io_neighbors_2(Cell_138_io_neighbors_2),
    .io_neighbors_3(Cell_138_io_neighbors_3),
    .io_neighbors_4(Cell_138_io_neighbors_4),
    .io_neighbors_5(Cell_138_io_neighbors_5),
    .io_neighbors_6(Cell_138_io_neighbors_6),
    .io_neighbors_7(Cell_138_io_neighbors_7),
    .io_out(Cell_138_io_out),
    .io_running(Cell_138_io_running),
    .io_writeEnable(Cell_138_io_writeEnable),
    .io_writeValue(Cell_138_io_writeValue)
  );
  Cell Cell_139 ( // @[Life.scala 59:52]
    .clock(Cell_139_clock),
    .reset(Cell_139_reset),
    .io_neighbors_0(Cell_139_io_neighbors_0),
    .io_neighbors_1(Cell_139_io_neighbors_1),
    .io_neighbors_2(Cell_139_io_neighbors_2),
    .io_neighbors_3(Cell_139_io_neighbors_3),
    .io_neighbors_4(Cell_139_io_neighbors_4),
    .io_neighbors_5(Cell_139_io_neighbors_5),
    .io_neighbors_6(Cell_139_io_neighbors_6),
    .io_neighbors_7(Cell_139_io_neighbors_7),
    .io_out(Cell_139_io_out),
    .io_running(Cell_139_io_running),
    .io_writeEnable(Cell_139_io_writeEnable),
    .io_writeValue(Cell_139_io_writeValue)
  );
  Cell Cell_140 ( // @[Life.scala 59:52]
    .clock(Cell_140_clock),
    .reset(Cell_140_reset),
    .io_neighbors_0(Cell_140_io_neighbors_0),
    .io_neighbors_1(Cell_140_io_neighbors_1),
    .io_neighbors_2(Cell_140_io_neighbors_2),
    .io_neighbors_3(Cell_140_io_neighbors_3),
    .io_neighbors_4(Cell_140_io_neighbors_4),
    .io_neighbors_5(Cell_140_io_neighbors_5),
    .io_neighbors_6(Cell_140_io_neighbors_6),
    .io_neighbors_7(Cell_140_io_neighbors_7),
    .io_out(Cell_140_io_out),
    .io_running(Cell_140_io_running),
    .io_writeEnable(Cell_140_io_writeEnable),
    .io_writeValue(Cell_140_io_writeValue)
  );
  Cell Cell_141 ( // @[Life.scala 59:52]
    .clock(Cell_141_clock),
    .reset(Cell_141_reset),
    .io_neighbors_0(Cell_141_io_neighbors_0),
    .io_neighbors_1(Cell_141_io_neighbors_1),
    .io_neighbors_2(Cell_141_io_neighbors_2),
    .io_neighbors_3(Cell_141_io_neighbors_3),
    .io_neighbors_4(Cell_141_io_neighbors_4),
    .io_neighbors_5(Cell_141_io_neighbors_5),
    .io_neighbors_6(Cell_141_io_neighbors_6),
    .io_neighbors_7(Cell_141_io_neighbors_7),
    .io_out(Cell_141_io_out),
    .io_running(Cell_141_io_running),
    .io_writeEnable(Cell_141_io_writeEnable),
    .io_writeValue(Cell_141_io_writeValue)
  );
  Cell Cell_142 ( // @[Life.scala 59:52]
    .clock(Cell_142_clock),
    .reset(Cell_142_reset),
    .io_neighbors_0(Cell_142_io_neighbors_0),
    .io_neighbors_1(Cell_142_io_neighbors_1),
    .io_neighbors_2(Cell_142_io_neighbors_2),
    .io_neighbors_3(Cell_142_io_neighbors_3),
    .io_neighbors_4(Cell_142_io_neighbors_4),
    .io_neighbors_5(Cell_142_io_neighbors_5),
    .io_neighbors_6(Cell_142_io_neighbors_6),
    .io_neighbors_7(Cell_142_io_neighbors_7),
    .io_out(Cell_142_io_out),
    .io_running(Cell_142_io_running),
    .io_writeEnable(Cell_142_io_writeEnable),
    .io_writeValue(Cell_142_io_writeValue)
  );
  Cell Cell_143 ( // @[Life.scala 59:52]
    .clock(Cell_143_clock),
    .reset(Cell_143_reset),
    .io_neighbors_0(Cell_143_io_neighbors_0),
    .io_neighbors_1(Cell_143_io_neighbors_1),
    .io_neighbors_2(Cell_143_io_neighbors_2),
    .io_neighbors_3(Cell_143_io_neighbors_3),
    .io_neighbors_4(Cell_143_io_neighbors_4),
    .io_neighbors_5(Cell_143_io_neighbors_5),
    .io_neighbors_6(Cell_143_io_neighbors_6),
    .io_neighbors_7(Cell_143_io_neighbors_7),
    .io_out(Cell_143_io_out),
    .io_running(Cell_143_io_running),
    .io_writeEnable(Cell_143_io_writeEnable),
    .io_writeValue(Cell_143_io_writeValue)
  );
  assign io_state_0_0 = Cell_io_out; // @[Life.scala 65:24]
  assign io_state_0_1 = Cell_1_io_out; // @[Life.scala 65:24]
  assign io_state_0_2 = Cell_2_io_out; // @[Life.scala 65:24]
  assign io_state_0_3 = Cell_3_io_out; // @[Life.scala 65:24]
  assign io_state_0_4 = Cell_4_io_out; // @[Life.scala 65:24]
  assign io_state_0_5 = Cell_5_io_out; // @[Life.scala 65:24]
  assign io_state_0_6 = Cell_6_io_out; // @[Life.scala 65:24]
  assign io_state_0_7 = Cell_7_io_out; // @[Life.scala 65:24]
  assign io_state_0_8 = Cell_8_io_out; // @[Life.scala 65:24]
  assign io_state_0_9 = Cell_9_io_out; // @[Life.scala 65:24]
  assign io_state_0_10 = Cell_10_io_out; // @[Life.scala 65:24]
  assign io_state_0_11 = Cell_11_io_out; // @[Life.scala 65:24]
  assign io_state_1_0 = Cell_12_io_out; // @[Life.scala 65:24]
  assign io_state_1_1 = Cell_13_io_out; // @[Life.scala 65:24]
  assign io_state_1_2 = Cell_14_io_out; // @[Life.scala 65:24]
  assign io_state_1_3 = Cell_15_io_out; // @[Life.scala 65:24]
  assign io_state_1_4 = Cell_16_io_out; // @[Life.scala 65:24]
  assign io_state_1_5 = Cell_17_io_out; // @[Life.scala 65:24]
  assign io_state_1_6 = Cell_18_io_out; // @[Life.scala 65:24]
  assign io_state_1_7 = Cell_19_io_out; // @[Life.scala 65:24]
  assign io_state_1_8 = Cell_20_io_out; // @[Life.scala 65:24]
  assign io_state_1_9 = Cell_21_io_out; // @[Life.scala 65:24]
  assign io_state_1_10 = Cell_22_io_out; // @[Life.scala 65:24]
  assign io_state_1_11 = Cell_23_io_out; // @[Life.scala 65:24]
  assign io_state_2_0 = Cell_24_io_out; // @[Life.scala 65:24]
  assign io_state_2_1 = Cell_25_io_out; // @[Life.scala 65:24]
  assign io_state_2_2 = Cell_26_io_out; // @[Life.scala 65:24]
  assign io_state_2_3 = Cell_27_io_out; // @[Life.scala 65:24]
  assign io_state_2_4 = Cell_28_io_out; // @[Life.scala 65:24]
  assign io_state_2_5 = Cell_29_io_out; // @[Life.scala 65:24]
  assign io_state_2_6 = Cell_30_io_out; // @[Life.scala 65:24]
  assign io_state_2_7 = Cell_31_io_out; // @[Life.scala 65:24]
  assign io_state_2_8 = Cell_32_io_out; // @[Life.scala 65:24]
  assign io_state_2_9 = Cell_33_io_out; // @[Life.scala 65:24]
  assign io_state_2_10 = Cell_34_io_out; // @[Life.scala 65:24]
  assign io_state_2_11 = Cell_35_io_out; // @[Life.scala 65:24]
  assign io_state_3_0 = Cell_36_io_out; // @[Life.scala 65:24]
  assign io_state_3_1 = Cell_37_io_out; // @[Life.scala 65:24]
  assign io_state_3_2 = Cell_38_io_out; // @[Life.scala 65:24]
  assign io_state_3_3 = Cell_39_io_out; // @[Life.scala 65:24]
  assign io_state_3_4 = Cell_40_io_out; // @[Life.scala 65:24]
  assign io_state_3_5 = Cell_41_io_out; // @[Life.scala 65:24]
  assign io_state_3_6 = Cell_42_io_out; // @[Life.scala 65:24]
  assign io_state_3_7 = Cell_43_io_out; // @[Life.scala 65:24]
  assign io_state_3_8 = Cell_44_io_out; // @[Life.scala 65:24]
  assign io_state_3_9 = Cell_45_io_out; // @[Life.scala 65:24]
  assign io_state_3_10 = Cell_46_io_out; // @[Life.scala 65:24]
  assign io_state_3_11 = Cell_47_io_out; // @[Life.scala 65:24]
  assign io_state_4_0 = Cell_48_io_out; // @[Life.scala 65:24]
  assign io_state_4_1 = Cell_49_io_out; // @[Life.scala 65:24]
  assign io_state_4_2 = Cell_50_io_out; // @[Life.scala 65:24]
  assign io_state_4_3 = Cell_51_io_out; // @[Life.scala 65:24]
  assign io_state_4_4 = Cell_52_io_out; // @[Life.scala 65:24]
  assign io_state_4_5 = Cell_53_io_out; // @[Life.scala 65:24]
  assign io_state_4_6 = Cell_54_io_out; // @[Life.scala 65:24]
  assign io_state_4_7 = Cell_55_io_out; // @[Life.scala 65:24]
  assign io_state_4_8 = Cell_56_io_out; // @[Life.scala 65:24]
  assign io_state_4_9 = Cell_57_io_out; // @[Life.scala 65:24]
  assign io_state_4_10 = Cell_58_io_out; // @[Life.scala 65:24]
  assign io_state_4_11 = Cell_59_io_out; // @[Life.scala 65:24]
  assign io_state_5_0 = Cell_60_io_out; // @[Life.scala 65:24]
  assign io_state_5_1 = Cell_61_io_out; // @[Life.scala 65:24]
  assign io_state_5_2 = Cell_62_io_out; // @[Life.scala 65:24]
  assign io_state_5_3 = Cell_63_io_out; // @[Life.scala 65:24]
  assign io_state_5_4 = Cell_64_io_out; // @[Life.scala 65:24]
  assign io_state_5_5 = Cell_65_io_out; // @[Life.scala 65:24]
  assign io_state_5_6 = Cell_66_io_out; // @[Life.scala 65:24]
  assign io_state_5_7 = Cell_67_io_out; // @[Life.scala 65:24]
  assign io_state_5_8 = Cell_68_io_out; // @[Life.scala 65:24]
  assign io_state_5_9 = Cell_69_io_out; // @[Life.scala 65:24]
  assign io_state_5_10 = Cell_70_io_out; // @[Life.scala 65:24]
  assign io_state_5_11 = Cell_71_io_out; // @[Life.scala 65:24]
  assign io_state_6_0 = Cell_72_io_out; // @[Life.scala 65:24]
  assign io_state_6_1 = Cell_73_io_out; // @[Life.scala 65:24]
  assign io_state_6_2 = Cell_74_io_out; // @[Life.scala 65:24]
  assign io_state_6_3 = Cell_75_io_out; // @[Life.scala 65:24]
  assign io_state_6_4 = Cell_76_io_out; // @[Life.scala 65:24]
  assign io_state_6_5 = Cell_77_io_out; // @[Life.scala 65:24]
  assign io_state_6_6 = Cell_78_io_out; // @[Life.scala 65:24]
  assign io_state_6_7 = Cell_79_io_out; // @[Life.scala 65:24]
  assign io_state_6_8 = Cell_80_io_out; // @[Life.scala 65:24]
  assign io_state_6_9 = Cell_81_io_out; // @[Life.scala 65:24]
  assign io_state_6_10 = Cell_82_io_out; // @[Life.scala 65:24]
  assign io_state_6_11 = Cell_83_io_out; // @[Life.scala 65:24]
  assign io_state_7_0 = Cell_84_io_out; // @[Life.scala 65:24]
  assign io_state_7_1 = Cell_85_io_out; // @[Life.scala 65:24]
  assign io_state_7_2 = Cell_86_io_out; // @[Life.scala 65:24]
  assign io_state_7_3 = Cell_87_io_out; // @[Life.scala 65:24]
  assign io_state_7_4 = Cell_88_io_out; // @[Life.scala 65:24]
  assign io_state_7_5 = Cell_89_io_out; // @[Life.scala 65:24]
  assign io_state_7_6 = Cell_90_io_out; // @[Life.scala 65:24]
  assign io_state_7_7 = Cell_91_io_out; // @[Life.scala 65:24]
  assign io_state_7_8 = Cell_92_io_out; // @[Life.scala 65:24]
  assign io_state_7_9 = Cell_93_io_out; // @[Life.scala 65:24]
  assign io_state_7_10 = Cell_94_io_out; // @[Life.scala 65:24]
  assign io_state_7_11 = Cell_95_io_out; // @[Life.scala 65:24]
  assign io_state_8_0 = Cell_96_io_out; // @[Life.scala 65:24]
  assign io_state_8_1 = Cell_97_io_out; // @[Life.scala 65:24]
  assign io_state_8_2 = Cell_98_io_out; // @[Life.scala 65:24]
  assign io_state_8_3 = Cell_99_io_out; // @[Life.scala 65:24]
  assign io_state_8_4 = Cell_100_io_out; // @[Life.scala 65:24]
  assign io_state_8_5 = Cell_101_io_out; // @[Life.scala 65:24]
  assign io_state_8_6 = Cell_102_io_out; // @[Life.scala 65:24]
  assign io_state_8_7 = Cell_103_io_out; // @[Life.scala 65:24]
  assign io_state_8_8 = Cell_104_io_out; // @[Life.scala 65:24]
  assign io_state_8_9 = Cell_105_io_out; // @[Life.scala 65:24]
  assign io_state_8_10 = Cell_106_io_out; // @[Life.scala 65:24]
  assign io_state_8_11 = Cell_107_io_out; // @[Life.scala 65:24]
  assign io_state_9_0 = Cell_108_io_out; // @[Life.scala 65:24]
  assign io_state_9_1 = Cell_109_io_out; // @[Life.scala 65:24]
  assign io_state_9_2 = Cell_110_io_out; // @[Life.scala 65:24]
  assign io_state_9_3 = Cell_111_io_out; // @[Life.scala 65:24]
  assign io_state_9_4 = Cell_112_io_out; // @[Life.scala 65:24]
  assign io_state_9_5 = Cell_113_io_out; // @[Life.scala 65:24]
  assign io_state_9_6 = Cell_114_io_out; // @[Life.scala 65:24]
  assign io_state_9_7 = Cell_115_io_out; // @[Life.scala 65:24]
  assign io_state_9_8 = Cell_116_io_out; // @[Life.scala 65:24]
  assign io_state_9_9 = Cell_117_io_out; // @[Life.scala 65:24]
  assign io_state_9_10 = Cell_118_io_out; // @[Life.scala 65:24]
  assign io_state_9_11 = Cell_119_io_out; // @[Life.scala 65:24]
  assign io_state_10_0 = Cell_120_io_out; // @[Life.scala 65:24]
  assign io_state_10_1 = Cell_121_io_out; // @[Life.scala 65:24]
  assign io_state_10_2 = Cell_122_io_out; // @[Life.scala 65:24]
  assign io_state_10_3 = Cell_123_io_out; // @[Life.scala 65:24]
  assign io_state_10_4 = Cell_124_io_out; // @[Life.scala 65:24]
  assign io_state_10_5 = Cell_125_io_out; // @[Life.scala 65:24]
  assign io_state_10_6 = Cell_126_io_out; // @[Life.scala 65:24]
  assign io_state_10_7 = Cell_127_io_out; // @[Life.scala 65:24]
  assign io_state_10_8 = Cell_128_io_out; // @[Life.scala 65:24]
  assign io_state_10_9 = Cell_129_io_out; // @[Life.scala 65:24]
  assign io_state_10_10 = Cell_130_io_out; // @[Life.scala 65:24]
  assign io_state_10_11 = Cell_131_io_out; // @[Life.scala 65:24]
  assign io_state_11_0 = Cell_132_io_out; // @[Life.scala 65:24]
  assign io_state_11_1 = Cell_133_io_out; // @[Life.scala 65:24]
  assign io_state_11_2 = Cell_134_io_out; // @[Life.scala 65:24]
  assign io_state_11_3 = Cell_135_io_out; // @[Life.scala 65:24]
  assign io_state_11_4 = Cell_136_io_out; // @[Life.scala 65:24]
  assign io_state_11_5 = Cell_137_io_out; // @[Life.scala 65:24]
  assign io_state_11_6 = Cell_138_io_out; // @[Life.scala 65:24]
  assign io_state_11_7 = Cell_139_io_out; // @[Life.scala 65:24]
  assign io_state_11_8 = Cell_140_io_out; // @[Life.scala 65:24]
  assign io_state_11_9 = Cell_141_io_out; // @[Life.scala 65:24]
  assign io_state_11_10 = Cell_142_io_out; // @[Life.scala 65:24]
  assign io_state_11_11 = Cell_143_io_out; // @[Life.scala 65:24]
  assign Cell_clock = clock;
  assign Cell_reset = reset;
  assign Cell_io_neighbors_0 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_1 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_2 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_3 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_4 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_5 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_6 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_io_neighbors_7 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_1_clock = clock;
  assign Cell_1_reset = reset;
  assign Cell_1_io_neighbors_0 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_1 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_2 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_3 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_4 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_5 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_6 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_neighbors_7 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_1_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_1_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_1_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_2_clock = clock;
  assign Cell_2_reset = reset;
  assign Cell_2_io_neighbors_0 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_1 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_2 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_3 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_4 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_5 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_6 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_neighbors_7 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_2_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_2_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_2_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_3_clock = clock;
  assign Cell_3_reset = reset;
  assign Cell_3_io_neighbors_0 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_1 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_2 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_3 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_4 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_5 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_6 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_neighbors_7 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_3_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_3_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_3_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_4_clock = clock;
  assign Cell_4_reset = reset;
  assign Cell_4_io_neighbors_0 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_1 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_2 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_3 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_4 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_5 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_6 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_neighbors_7 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_4_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_4_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_4_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_5_clock = clock;
  assign Cell_5_reset = reset;
  assign Cell_5_io_neighbors_0 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_1 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_2 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_3 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_4 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_5 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_6 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_neighbors_7 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_5_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_5_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_5_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_6_clock = clock;
  assign Cell_6_reset = reset;
  assign Cell_6_io_neighbors_0 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_1 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_2 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_3 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_4 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_5 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_6 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_neighbors_7 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_6_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_6_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_6_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_7_clock = clock;
  assign Cell_7_reset = reset;
  assign Cell_7_io_neighbors_0 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_1 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_2 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_3 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_4 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_5 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_6 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_neighbors_7 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_7_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_7_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_7_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_8_clock = clock;
  assign Cell_8_reset = reset;
  assign Cell_8_io_neighbors_0 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_1 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_2 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_3 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_4 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_5 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_6 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_neighbors_7 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_8_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_8_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_8_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_9_clock = clock;
  assign Cell_9_reset = reset;
  assign Cell_9_io_neighbors_0 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_1 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_2 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_3 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_4 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_5 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_6 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_neighbors_7 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_9_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_9_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_9_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_10_clock = clock;
  assign Cell_10_reset = reset;
  assign Cell_10_io_neighbors_0 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_1 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_2 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_3 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_4 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_5 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_6 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_neighbors_7 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_10_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_10_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_10_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_11_clock = clock;
  assign Cell_11_reset = reset;
  assign Cell_11_io_neighbors_0 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_1 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_2 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_3 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_4 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_5 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_6 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_neighbors_7 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_11_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_11_io_writeEnable = io_writeRowAddress == 4'h0 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_11_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_12_clock = clock;
  assign Cell_12_reset = reset;
  assign Cell_12_io_neighbors_0 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_1 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_2 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_3 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_4 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_5 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_6 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_neighbors_7 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_12_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_12_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_12_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_13_clock = clock;
  assign Cell_13_reset = reset;
  assign Cell_13_io_neighbors_0 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_1 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_2 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_3 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_4 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_5 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_6 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_neighbors_7 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_13_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_13_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_13_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_14_clock = clock;
  assign Cell_14_reset = reset;
  assign Cell_14_io_neighbors_0 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_1 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_2 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_3 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_4 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_5 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_6 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_neighbors_7 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_14_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_14_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_14_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_15_clock = clock;
  assign Cell_15_reset = reset;
  assign Cell_15_io_neighbors_0 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_1 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_2 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_3 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_4 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_5 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_6 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_neighbors_7 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_15_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_15_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_15_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_16_clock = clock;
  assign Cell_16_reset = reset;
  assign Cell_16_io_neighbors_0 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_1 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_2 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_3 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_4 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_5 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_6 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_neighbors_7 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_16_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_16_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_16_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_17_clock = clock;
  assign Cell_17_reset = reset;
  assign Cell_17_io_neighbors_0 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_1 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_2 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_3 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_4 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_5 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_6 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_neighbors_7 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_17_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_17_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_17_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_18_clock = clock;
  assign Cell_18_reset = reset;
  assign Cell_18_io_neighbors_0 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_1 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_2 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_3 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_4 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_5 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_6 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_neighbors_7 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_18_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_18_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_18_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_19_clock = clock;
  assign Cell_19_reset = reset;
  assign Cell_19_io_neighbors_0 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_1 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_2 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_3 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_4 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_5 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_6 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_neighbors_7 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_19_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_19_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_19_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_20_clock = clock;
  assign Cell_20_reset = reset;
  assign Cell_20_io_neighbors_0 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_1 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_2 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_3 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_4 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_5 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_6 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_neighbors_7 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_20_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_20_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_20_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_21_clock = clock;
  assign Cell_21_reset = reset;
  assign Cell_21_io_neighbors_0 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_1 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_2 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_3 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_4 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_5 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_6 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_neighbors_7 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_21_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_21_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_21_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_22_clock = clock;
  assign Cell_22_reset = reset;
  assign Cell_22_io_neighbors_0 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_1 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_2 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_3 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_4 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_5 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_6 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_neighbors_7 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_22_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_22_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_22_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_23_clock = clock;
  assign Cell_23_reset = reset;
  assign Cell_23_io_neighbors_0 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_1 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_2 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_3 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_4 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_5 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_6 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_neighbors_7 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_23_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_23_io_writeEnable = io_writeRowAddress == 4'h1 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_23_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_24_clock = clock;
  assign Cell_24_reset = reset;
  assign Cell_24_io_neighbors_0 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_1 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_2 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_3 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_4 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_5 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_6 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_neighbors_7 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_24_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_24_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_24_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_25_clock = clock;
  assign Cell_25_reset = reset;
  assign Cell_25_io_neighbors_0 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_1 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_2 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_3 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_4 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_5 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_6 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_neighbors_7 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_25_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_25_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_25_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_26_clock = clock;
  assign Cell_26_reset = reset;
  assign Cell_26_io_neighbors_0 = Cell_13_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_1 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_2 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_3 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_4 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_5 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_6 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_neighbors_7 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_26_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_26_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_26_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_27_clock = clock;
  assign Cell_27_reset = reset;
  assign Cell_27_io_neighbors_0 = Cell_14_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_1 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_2 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_3 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_4 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_5 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_6 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_neighbors_7 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_27_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_27_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_27_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_28_clock = clock;
  assign Cell_28_reset = reset;
  assign Cell_28_io_neighbors_0 = Cell_15_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_1 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_2 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_3 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_4 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_5 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_6 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_neighbors_7 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_28_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_28_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_28_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_29_clock = clock;
  assign Cell_29_reset = reset;
  assign Cell_29_io_neighbors_0 = Cell_16_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_1 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_2 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_3 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_4 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_5 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_6 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_neighbors_7 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_29_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_29_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_29_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_30_clock = clock;
  assign Cell_30_reset = reset;
  assign Cell_30_io_neighbors_0 = Cell_17_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_1 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_2 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_3 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_4 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_5 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_6 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_neighbors_7 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_30_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_30_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_30_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_31_clock = clock;
  assign Cell_31_reset = reset;
  assign Cell_31_io_neighbors_0 = Cell_18_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_1 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_2 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_3 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_4 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_5 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_6 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_neighbors_7 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_31_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_31_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_31_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_32_clock = clock;
  assign Cell_32_reset = reset;
  assign Cell_32_io_neighbors_0 = Cell_19_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_1 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_2 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_3 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_4 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_5 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_6 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_neighbors_7 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_32_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_32_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_32_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_33_clock = clock;
  assign Cell_33_reset = reset;
  assign Cell_33_io_neighbors_0 = Cell_20_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_1 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_2 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_3 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_4 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_5 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_6 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_neighbors_7 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_33_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_33_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_33_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_34_clock = clock;
  assign Cell_34_reset = reset;
  assign Cell_34_io_neighbors_0 = Cell_21_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_1 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_2 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_3 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_4 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_5 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_6 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_neighbors_7 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_34_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_34_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_34_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_35_clock = clock;
  assign Cell_35_reset = reset;
  assign Cell_35_io_neighbors_0 = Cell_22_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_1 = Cell_23_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_2 = Cell_12_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_3 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_4 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_5 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_6 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_neighbors_7 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_35_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_35_io_writeEnable = io_writeRowAddress == 4'h2 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_35_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_36_clock = clock;
  assign Cell_36_reset = reset;
  assign Cell_36_io_neighbors_0 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_1 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_2 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_3 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_4 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_5 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_6 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_neighbors_7 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_36_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_36_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_36_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_37_clock = clock;
  assign Cell_37_reset = reset;
  assign Cell_37_io_neighbors_0 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_1 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_2 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_3 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_4 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_5 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_6 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_neighbors_7 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_37_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_37_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_37_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_38_clock = clock;
  assign Cell_38_reset = reset;
  assign Cell_38_io_neighbors_0 = Cell_25_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_1 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_2 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_3 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_4 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_5 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_6 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_neighbors_7 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_38_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_38_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_38_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_39_clock = clock;
  assign Cell_39_reset = reset;
  assign Cell_39_io_neighbors_0 = Cell_26_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_1 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_2 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_3 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_4 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_5 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_6 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_neighbors_7 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_39_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_39_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_39_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_40_clock = clock;
  assign Cell_40_reset = reset;
  assign Cell_40_io_neighbors_0 = Cell_27_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_1 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_2 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_3 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_4 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_5 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_6 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_neighbors_7 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_40_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_40_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_40_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_41_clock = clock;
  assign Cell_41_reset = reset;
  assign Cell_41_io_neighbors_0 = Cell_28_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_1 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_2 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_3 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_4 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_5 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_6 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_neighbors_7 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_41_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_41_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_41_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_42_clock = clock;
  assign Cell_42_reset = reset;
  assign Cell_42_io_neighbors_0 = Cell_29_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_1 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_2 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_3 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_4 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_5 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_6 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_neighbors_7 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_42_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_42_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_42_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_43_clock = clock;
  assign Cell_43_reset = reset;
  assign Cell_43_io_neighbors_0 = Cell_30_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_1 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_2 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_3 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_4 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_5 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_6 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_neighbors_7 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_43_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_43_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_43_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_44_clock = clock;
  assign Cell_44_reset = reset;
  assign Cell_44_io_neighbors_0 = Cell_31_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_1 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_2 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_3 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_4 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_5 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_6 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_neighbors_7 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_44_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_44_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_44_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_45_clock = clock;
  assign Cell_45_reset = reset;
  assign Cell_45_io_neighbors_0 = Cell_32_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_1 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_2 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_3 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_4 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_5 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_6 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_neighbors_7 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_45_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_45_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_45_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_46_clock = clock;
  assign Cell_46_reset = reset;
  assign Cell_46_io_neighbors_0 = Cell_33_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_1 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_2 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_3 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_4 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_5 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_6 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_neighbors_7 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_46_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_46_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_46_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_47_clock = clock;
  assign Cell_47_reset = reset;
  assign Cell_47_io_neighbors_0 = Cell_34_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_1 = Cell_35_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_2 = Cell_24_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_3 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_4 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_5 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_6 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_neighbors_7 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_47_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_47_io_writeEnable = io_writeRowAddress == 4'h3 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_47_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_48_clock = clock;
  assign Cell_48_reset = reset;
  assign Cell_48_io_neighbors_0 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_1 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_2 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_3 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_4 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_5 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_6 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_neighbors_7 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_48_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_48_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_48_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_49_clock = clock;
  assign Cell_49_reset = reset;
  assign Cell_49_io_neighbors_0 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_1 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_2 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_3 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_4 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_5 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_6 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_neighbors_7 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_49_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_49_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_49_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_50_clock = clock;
  assign Cell_50_reset = reset;
  assign Cell_50_io_neighbors_0 = Cell_37_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_1 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_2 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_3 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_4 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_5 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_6 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_neighbors_7 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_50_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_50_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_50_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_51_clock = clock;
  assign Cell_51_reset = reset;
  assign Cell_51_io_neighbors_0 = Cell_38_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_1 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_2 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_3 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_4 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_5 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_6 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_neighbors_7 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_51_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_51_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_51_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_52_clock = clock;
  assign Cell_52_reset = reset;
  assign Cell_52_io_neighbors_0 = Cell_39_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_1 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_2 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_3 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_4 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_5 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_6 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_neighbors_7 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_52_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_52_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_52_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_53_clock = clock;
  assign Cell_53_reset = reset;
  assign Cell_53_io_neighbors_0 = Cell_40_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_1 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_2 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_3 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_4 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_5 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_6 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_neighbors_7 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_53_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_53_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_53_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_54_clock = clock;
  assign Cell_54_reset = reset;
  assign Cell_54_io_neighbors_0 = Cell_41_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_1 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_2 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_3 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_4 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_5 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_6 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_neighbors_7 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_54_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_54_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_54_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_55_clock = clock;
  assign Cell_55_reset = reset;
  assign Cell_55_io_neighbors_0 = Cell_42_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_1 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_2 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_3 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_4 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_5 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_6 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_neighbors_7 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_55_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_55_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_55_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_56_clock = clock;
  assign Cell_56_reset = reset;
  assign Cell_56_io_neighbors_0 = Cell_43_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_1 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_2 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_3 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_4 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_5 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_6 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_neighbors_7 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_56_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_56_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_56_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_57_clock = clock;
  assign Cell_57_reset = reset;
  assign Cell_57_io_neighbors_0 = Cell_44_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_1 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_2 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_3 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_4 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_5 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_6 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_neighbors_7 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_57_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_57_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_57_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_58_clock = clock;
  assign Cell_58_reset = reset;
  assign Cell_58_io_neighbors_0 = Cell_45_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_1 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_2 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_3 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_4 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_5 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_6 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_neighbors_7 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_58_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_58_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_58_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_59_clock = clock;
  assign Cell_59_reset = reset;
  assign Cell_59_io_neighbors_0 = Cell_46_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_1 = Cell_47_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_2 = Cell_36_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_3 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_4 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_5 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_6 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_neighbors_7 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_59_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_59_io_writeEnable = io_writeRowAddress == 4'h4 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_59_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_60_clock = clock;
  assign Cell_60_reset = reset;
  assign Cell_60_io_neighbors_0 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_1 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_2 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_3 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_4 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_5 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_6 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_neighbors_7 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_60_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_60_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_60_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_61_clock = clock;
  assign Cell_61_reset = reset;
  assign Cell_61_io_neighbors_0 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_1 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_2 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_3 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_4 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_5 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_6 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_neighbors_7 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_61_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_61_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_61_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_62_clock = clock;
  assign Cell_62_reset = reset;
  assign Cell_62_io_neighbors_0 = Cell_49_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_1 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_2 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_3 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_4 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_5 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_6 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_neighbors_7 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_62_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_62_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_62_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_63_clock = clock;
  assign Cell_63_reset = reset;
  assign Cell_63_io_neighbors_0 = Cell_50_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_1 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_2 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_3 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_4 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_5 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_6 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_neighbors_7 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_63_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_63_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_63_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_64_clock = clock;
  assign Cell_64_reset = reset;
  assign Cell_64_io_neighbors_0 = Cell_51_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_1 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_2 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_3 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_4 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_5 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_6 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_neighbors_7 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_64_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_64_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_64_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_65_clock = clock;
  assign Cell_65_reset = reset;
  assign Cell_65_io_neighbors_0 = Cell_52_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_1 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_2 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_3 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_4 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_5 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_6 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_neighbors_7 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_65_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_65_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_65_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_66_clock = clock;
  assign Cell_66_reset = reset;
  assign Cell_66_io_neighbors_0 = Cell_53_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_1 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_2 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_3 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_4 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_5 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_6 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_neighbors_7 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_66_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_66_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_66_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_67_clock = clock;
  assign Cell_67_reset = reset;
  assign Cell_67_io_neighbors_0 = Cell_54_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_1 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_2 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_3 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_4 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_5 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_6 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_neighbors_7 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_67_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_67_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_67_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_68_clock = clock;
  assign Cell_68_reset = reset;
  assign Cell_68_io_neighbors_0 = Cell_55_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_1 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_2 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_3 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_4 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_5 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_6 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_neighbors_7 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_68_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_68_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_68_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_69_clock = clock;
  assign Cell_69_reset = reset;
  assign Cell_69_io_neighbors_0 = Cell_56_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_1 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_2 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_3 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_4 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_5 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_6 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_neighbors_7 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_69_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_69_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_69_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_70_clock = clock;
  assign Cell_70_reset = reset;
  assign Cell_70_io_neighbors_0 = Cell_57_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_1 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_2 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_3 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_4 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_5 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_6 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_neighbors_7 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_70_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_70_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_70_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_71_clock = clock;
  assign Cell_71_reset = reset;
  assign Cell_71_io_neighbors_0 = Cell_58_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_1 = Cell_59_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_2 = Cell_48_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_3 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_4 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_5 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_6 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_neighbors_7 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_71_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_71_io_writeEnable = io_writeRowAddress == 4'h5 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_71_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_72_clock = clock;
  assign Cell_72_reset = reset;
  assign Cell_72_io_neighbors_0 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_1 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_2 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_3 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_4 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_5 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_6 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_neighbors_7 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_72_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_72_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_72_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_73_clock = clock;
  assign Cell_73_reset = reset;
  assign Cell_73_io_neighbors_0 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_1 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_2 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_3 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_4 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_5 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_6 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_neighbors_7 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_73_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_73_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_73_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_74_clock = clock;
  assign Cell_74_reset = reset;
  assign Cell_74_io_neighbors_0 = Cell_61_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_1 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_2 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_3 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_4 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_5 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_6 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_neighbors_7 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_74_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_74_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_74_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_75_clock = clock;
  assign Cell_75_reset = reset;
  assign Cell_75_io_neighbors_0 = Cell_62_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_1 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_2 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_3 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_4 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_5 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_6 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_neighbors_7 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_75_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_75_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_75_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_76_clock = clock;
  assign Cell_76_reset = reset;
  assign Cell_76_io_neighbors_0 = Cell_63_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_1 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_2 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_3 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_4 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_5 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_6 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_neighbors_7 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_76_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_76_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_76_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_77_clock = clock;
  assign Cell_77_reset = reset;
  assign Cell_77_io_neighbors_0 = Cell_64_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_1 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_2 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_3 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_4 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_5 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_6 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_neighbors_7 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_77_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_77_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_77_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_78_clock = clock;
  assign Cell_78_reset = reset;
  assign Cell_78_io_neighbors_0 = Cell_65_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_1 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_2 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_3 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_4 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_5 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_6 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_neighbors_7 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_78_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_78_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_78_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_79_clock = clock;
  assign Cell_79_reset = reset;
  assign Cell_79_io_neighbors_0 = Cell_66_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_1 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_2 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_3 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_4 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_5 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_6 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_neighbors_7 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_79_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_79_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_79_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_80_clock = clock;
  assign Cell_80_reset = reset;
  assign Cell_80_io_neighbors_0 = Cell_67_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_1 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_2 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_3 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_4 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_5 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_6 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_neighbors_7 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_80_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_80_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_80_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_81_clock = clock;
  assign Cell_81_reset = reset;
  assign Cell_81_io_neighbors_0 = Cell_68_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_1 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_2 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_3 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_4 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_5 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_6 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_neighbors_7 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_81_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_81_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_81_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_82_clock = clock;
  assign Cell_82_reset = reset;
  assign Cell_82_io_neighbors_0 = Cell_69_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_1 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_2 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_3 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_4 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_5 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_6 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_neighbors_7 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_82_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_82_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_82_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_83_clock = clock;
  assign Cell_83_reset = reset;
  assign Cell_83_io_neighbors_0 = Cell_70_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_1 = Cell_71_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_2 = Cell_60_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_3 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_4 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_5 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_6 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_neighbors_7 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_83_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_83_io_writeEnable = io_writeRowAddress == 4'h6 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_83_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_84_clock = clock;
  assign Cell_84_reset = reset;
  assign Cell_84_io_neighbors_0 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_1 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_2 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_3 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_4 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_5 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_6 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_neighbors_7 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_84_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_84_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_84_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_85_clock = clock;
  assign Cell_85_reset = reset;
  assign Cell_85_io_neighbors_0 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_1 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_2 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_3 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_4 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_5 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_6 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_neighbors_7 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_85_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_85_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_85_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_86_clock = clock;
  assign Cell_86_reset = reset;
  assign Cell_86_io_neighbors_0 = Cell_73_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_1 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_2 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_3 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_4 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_5 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_6 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_neighbors_7 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_86_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_86_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_86_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_87_clock = clock;
  assign Cell_87_reset = reset;
  assign Cell_87_io_neighbors_0 = Cell_74_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_1 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_2 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_3 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_4 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_5 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_6 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_neighbors_7 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_87_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_87_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_87_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_88_clock = clock;
  assign Cell_88_reset = reset;
  assign Cell_88_io_neighbors_0 = Cell_75_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_1 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_2 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_3 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_4 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_5 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_6 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_neighbors_7 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_88_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_88_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_88_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_89_clock = clock;
  assign Cell_89_reset = reset;
  assign Cell_89_io_neighbors_0 = Cell_76_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_1 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_2 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_3 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_4 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_5 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_6 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_neighbors_7 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_89_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_89_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_89_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_90_clock = clock;
  assign Cell_90_reset = reset;
  assign Cell_90_io_neighbors_0 = Cell_77_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_1 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_2 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_3 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_4 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_5 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_6 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_neighbors_7 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_90_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_90_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_90_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_91_clock = clock;
  assign Cell_91_reset = reset;
  assign Cell_91_io_neighbors_0 = Cell_78_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_1 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_2 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_3 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_4 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_5 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_6 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_neighbors_7 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_91_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_91_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_91_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_92_clock = clock;
  assign Cell_92_reset = reset;
  assign Cell_92_io_neighbors_0 = Cell_79_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_1 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_2 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_3 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_4 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_5 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_6 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_neighbors_7 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_92_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_92_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_92_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_93_clock = clock;
  assign Cell_93_reset = reset;
  assign Cell_93_io_neighbors_0 = Cell_80_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_1 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_2 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_3 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_4 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_5 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_6 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_neighbors_7 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_93_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_93_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_93_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_94_clock = clock;
  assign Cell_94_reset = reset;
  assign Cell_94_io_neighbors_0 = Cell_81_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_1 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_2 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_3 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_4 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_5 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_6 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_neighbors_7 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_94_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_94_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_94_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_95_clock = clock;
  assign Cell_95_reset = reset;
  assign Cell_95_io_neighbors_0 = Cell_82_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_1 = Cell_83_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_2 = Cell_72_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_3 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_4 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_5 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_6 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_neighbors_7 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_95_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_95_io_writeEnable = io_writeRowAddress == 4'h7 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_95_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_96_clock = clock;
  assign Cell_96_reset = reset;
  assign Cell_96_io_neighbors_0 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_1 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_2 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_3 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_4 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_5 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_6 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_neighbors_7 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_96_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_96_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_96_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_97_clock = clock;
  assign Cell_97_reset = reset;
  assign Cell_97_io_neighbors_0 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_1 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_2 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_3 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_4 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_5 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_6 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_neighbors_7 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_97_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_97_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_97_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_98_clock = clock;
  assign Cell_98_reset = reset;
  assign Cell_98_io_neighbors_0 = Cell_85_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_1 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_2 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_3 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_4 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_5 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_6 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_neighbors_7 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_98_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_98_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_98_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_99_clock = clock;
  assign Cell_99_reset = reset;
  assign Cell_99_io_neighbors_0 = Cell_86_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_1 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_2 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_3 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_4 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_5 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_6 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_neighbors_7 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_99_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_99_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_99_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_100_clock = clock;
  assign Cell_100_reset = reset;
  assign Cell_100_io_neighbors_0 = Cell_87_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_1 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_2 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_3 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_4 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_5 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_6 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_neighbors_7 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_100_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_100_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_100_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_101_clock = clock;
  assign Cell_101_reset = reset;
  assign Cell_101_io_neighbors_0 = Cell_88_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_1 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_2 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_3 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_4 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_5 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_6 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_neighbors_7 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_101_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_101_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_101_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_102_clock = clock;
  assign Cell_102_reset = reset;
  assign Cell_102_io_neighbors_0 = Cell_89_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_1 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_2 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_3 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_4 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_5 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_6 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_neighbors_7 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_102_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_102_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_102_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_103_clock = clock;
  assign Cell_103_reset = reset;
  assign Cell_103_io_neighbors_0 = Cell_90_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_1 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_2 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_3 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_4 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_5 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_6 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_neighbors_7 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_103_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_103_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_103_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_104_clock = clock;
  assign Cell_104_reset = reset;
  assign Cell_104_io_neighbors_0 = Cell_91_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_1 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_2 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_3 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_4 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_5 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_6 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_neighbors_7 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_104_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_104_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_104_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_105_clock = clock;
  assign Cell_105_reset = reset;
  assign Cell_105_io_neighbors_0 = Cell_92_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_1 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_2 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_3 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_4 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_5 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_6 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_neighbors_7 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_105_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_105_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_105_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_106_clock = clock;
  assign Cell_106_reset = reset;
  assign Cell_106_io_neighbors_0 = Cell_93_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_1 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_2 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_3 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_4 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_5 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_6 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_neighbors_7 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_106_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_106_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_106_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_107_clock = clock;
  assign Cell_107_reset = reset;
  assign Cell_107_io_neighbors_0 = Cell_94_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_1 = Cell_95_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_2 = Cell_84_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_3 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_4 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_5 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_6 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_neighbors_7 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_107_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_107_io_writeEnable = io_writeRowAddress == 4'h8 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_107_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_108_clock = clock;
  assign Cell_108_reset = reset;
  assign Cell_108_io_neighbors_0 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_1 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_2 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_3 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_4 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_5 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_6 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_neighbors_7 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_108_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_108_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_108_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_109_clock = clock;
  assign Cell_109_reset = reset;
  assign Cell_109_io_neighbors_0 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_1 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_2 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_3 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_4 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_5 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_6 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_neighbors_7 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_109_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_109_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_109_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_110_clock = clock;
  assign Cell_110_reset = reset;
  assign Cell_110_io_neighbors_0 = Cell_97_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_1 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_2 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_3 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_4 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_5 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_6 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_neighbors_7 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_110_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_110_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_110_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_111_clock = clock;
  assign Cell_111_reset = reset;
  assign Cell_111_io_neighbors_0 = Cell_98_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_1 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_2 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_3 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_4 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_5 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_6 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_neighbors_7 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_111_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_111_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_111_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_112_clock = clock;
  assign Cell_112_reset = reset;
  assign Cell_112_io_neighbors_0 = Cell_99_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_1 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_2 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_3 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_4 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_5 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_6 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_neighbors_7 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_112_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_112_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_112_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_113_clock = clock;
  assign Cell_113_reset = reset;
  assign Cell_113_io_neighbors_0 = Cell_100_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_1 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_2 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_3 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_4 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_5 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_6 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_neighbors_7 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_113_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_113_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_113_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_114_clock = clock;
  assign Cell_114_reset = reset;
  assign Cell_114_io_neighbors_0 = Cell_101_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_1 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_2 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_3 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_4 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_5 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_6 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_neighbors_7 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_114_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_114_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_114_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_115_clock = clock;
  assign Cell_115_reset = reset;
  assign Cell_115_io_neighbors_0 = Cell_102_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_1 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_2 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_3 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_4 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_5 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_6 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_neighbors_7 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_115_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_115_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_115_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_116_clock = clock;
  assign Cell_116_reset = reset;
  assign Cell_116_io_neighbors_0 = Cell_103_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_1 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_2 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_3 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_4 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_5 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_6 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_neighbors_7 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_116_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_116_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_116_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_117_clock = clock;
  assign Cell_117_reset = reset;
  assign Cell_117_io_neighbors_0 = Cell_104_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_1 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_2 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_3 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_4 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_5 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_6 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_neighbors_7 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_117_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_117_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_117_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_118_clock = clock;
  assign Cell_118_reset = reset;
  assign Cell_118_io_neighbors_0 = Cell_105_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_1 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_2 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_3 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_4 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_5 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_6 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_neighbors_7 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_118_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_118_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_118_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_119_clock = clock;
  assign Cell_119_reset = reset;
  assign Cell_119_io_neighbors_0 = Cell_106_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_1 = Cell_107_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_2 = Cell_96_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_3 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_4 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_5 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_6 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_neighbors_7 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_119_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_119_io_writeEnable = io_writeRowAddress == 4'h9 & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_119_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_120_clock = clock;
  assign Cell_120_reset = reset;
  assign Cell_120_io_neighbors_0 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_1 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_2 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_3 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_4 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_5 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_6 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_neighbors_7 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_120_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_120_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_120_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_121_clock = clock;
  assign Cell_121_reset = reset;
  assign Cell_121_io_neighbors_0 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_1 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_2 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_3 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_4 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_5 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_6 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_neighbors_7 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_121_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_121_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_121_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_122_clock = clock;
  assign Cell_122_reset = reset;
  assign Cell_122_io_neighbors_0 = Cell_109_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_1 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_2 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_3 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_4 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_5 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_6 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_neighbors_7 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_122_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_122_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_122_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_123_clock = clock;
  assign Cell_123_reset = reset;
  assign Cell_123_io_neighbors_0 = Cell_110_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_1 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_2 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_3 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_4 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_5 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_6 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_neighbors_7 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_123_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_123_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_123_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_124_clock = clock;
  assign Cell_124_reset = reset;
  assign Cell_124_io_neighbors_0 = Cell_111_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_1 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_2 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_3 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_4 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_5 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_6 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_neighbors_7 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_124_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_124_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_124_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_125_clock = clock;
  assign Cell_125_reset = reset;
  assign Cell_125_io_neighbors_0 = Cell_112_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_1 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_2 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_3 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_4 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_5 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_6 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_neighbors_7 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_125_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_125_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_125_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_126_clock = clock;
  assign Cell_126_reset = reset;
  assign Cell_126_io_neighbors_0 = Cell_113_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_1 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_2 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_3 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_4 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_5 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_6 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_neighbors_7 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_126_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_126_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_126_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_127_clock = clock;
  assign Cell_127_reset = reset;
  assign Cell_127_io_neighbors_0 = Cell_114_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_1 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_2 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_3 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_4 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_5 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_6 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_neighbors_7 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_127_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_127_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_127_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_128_clock = clock;
  assign Cell_128_reset = reset;
  assign Cell_128_io_neighbors_0 = Cell_115_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_1 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_2 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_3 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_4 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_5 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_6 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_neighbors_7 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_128_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_128_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_128_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_129_clock = clock;
  assign Cell_129_reset = reset;
  assign Cell_129_io_neighbors_0 = Cell_116_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_1 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_2 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_3 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_4 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_5 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_6 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_neighbors_7 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_129_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_129_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_129_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_130_clock = clock;
  assign Cell_130_reset = reset;
  assign Cell_130_io_neighbors_0 = Cell_117_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_1 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_2 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_3 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_4 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_5 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_6 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_neighbors_7 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_130_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_130_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_130_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_131_clock = clock;
  assign Cell_131_reset = reset;
  assign Cell_131_io_neighbors_0 = Cell_118_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_1 = Cell_119_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_2 = Cell_108_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_3 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_4 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_5 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_6 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_neighbors_7 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_131_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_131_io_writeEnable = io_writeRowAddress == 4'ha & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_131_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_132_clock = clock;
  assign Cell_132_reset = reset;
  assign Cell_132_io_neighbors_0 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_1 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_2 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_3 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_4 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_5 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_6 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_neighbors_7 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_132_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_132_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h0; // @[Life.scala 68:68]
  assign Cell_132_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_133_clock = clock;
  assign Cell_133_reset = reset;
  assign Cell_133_io_neighbors_0 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_1 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_2 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_3 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_4 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_5 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_6 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_neighbors_7 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_133_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_133_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h1; // @[Life.scala 68:68]
  assign Cell_133_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_134_clock = clock;
  assign Cell_134_reset = reset;
  assign Cell_134_io_neighbors_0 = Cell_121_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_1 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_2 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_3 = Cell_133_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_4 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_5 = Cell_1_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_6 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_neighbors_7 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_134_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_134_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h2; // @[Life.scala 68:68]
  assign Cell_134_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_135_clock = clock;
  assign Cell_135_reset = reset;
  assign Cell_135_io_neighbors_0 = Cell_122_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_1 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_2 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_3 = Cell_134_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_4 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_5 = Cell_2_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_6 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_neighbors_7 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_135_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_135_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h3; // @[Life.scala 68:68]
  assign Cell_135_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_136_clock = clock;
  assign Cell_136_reset = reset;
  assign Cell_136_io_neighbors_0 = Cell_123_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_1 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_2 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_3 = Cell_135_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_4 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_5 = Cell_3_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_6 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_neighbors_7 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_136_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_136_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h4; // @[Life.scala 68:68]
  assign Cell_136_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_137_clock = clock;
  assign Cell_137_reset = reset;
  assign Cell_137_io_neighbors_0 = Cell_124_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_1 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_2 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_3 = Cell_136_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_4 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_5 = Cell_4_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_6 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_neighbors_7 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_137_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_137_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h5; // @[Life.scala 68:68]
  assign Cell_137_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_138_clock = clock;
  assign Cell_138_reset = reset;
  assign Cell_138_io_neighbors_0 = Cell_125_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_1 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_2 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_3 = Cell_137_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_4 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_5 = Cell_5_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_6 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_neighbors_7 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_138_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_138_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h6; // @[Life.scala 68:68]
  assign Cell_138_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_139_clock = clock;
  assign Cell_139_reset = reset;
  assign Cell_139_io_neighbors_0 = Cell_126_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_1 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_2 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_3 = Cell_138_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_4 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_5 = Cell_6_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_6 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_neighbors_7 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_139_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_139_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h7; // @[Life.scala 68:68]
  assign Cell_139_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_140_clock = clock;
  assign Cell_140_reset = reset;
  assign Cell_140_io_neighbors_0 = Cell_127_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_1 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_2 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_3 = Cell_139_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_4 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_5 = Cell_7_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_6 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_neighbors_7 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_140_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_140_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h8; // @[Life.scala 68:68]
  assign Cell_140_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_141_clock = clock;
  assign Cell_141_reset = reset;
  assign Cell_141_io_neighbors_0 = Cell_128_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_1 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_2 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_3 = Cell_140_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_4 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_5 = Cell_8_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_6 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_neighbors_7 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_141_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_141_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'h9; // @[Life.scala 68:68]
  assign Cell_141_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_142_clock = clock;
  assign Cell_142_reset = reset;
  assign Cell_142_io_neighbors_0 = Cell_129_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_1 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_2 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_3 = Cell_141_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_4 = Cell_143_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_5 = Cell_9_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_6 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_neighbors_7 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_142_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_142_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'ha; // @[Life.scala 68:68]
  assign Cell_142_io_writeValue = io_writeValue; // @[Life.scala 67:35]
  assign Cell_143_clock = clock;
  assign Cell_143_reset = reset;
  assign Cell_143_io_neighbors_0 = Cell_130_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_1 = Cell_131_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_2 = Cell_120_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_3 = Cell_142_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_4 = Cell_132_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_5 = Cell_10_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_6 = Cell_11_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_neighbors_7 = Cell_io_out; // @[Life.scala 89:46]
  assign Cell_143_io_running = io_running; // @[Life.scala 66:32]
  assign Cell_143_io_writeEnable = io_writeRowAddress == 4'hb & io_writeColAddress == 4'hb; // @[Life.scala 68:68]
  assign Cell_143_io_writeValue = io_writeValue; // @[Life.scala 67:35]
endmodule
