module RVCExpander_2(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire [6:0] _T_4 = |io_in[12:5] ? 7'h13 : 7'h1f; // @[RVC.scala 54:20]
  wire [4:0] _T_14 = {2'h1,io_in[4:2]}; // @[Cat.scala 29:58]
  wire [29:0] _T_18 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_4}; // @[Cat.scala 29:58]
  wire [7:0] _T_28 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [4:0] _T_30 = {2'h1,io_in[9:7]}; // @[Cat.scala 29:58]
  wire [27:0] _T_36 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [6:0] _T_50 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [27:0] _T_78 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [26:0] _T_109 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58]
  wire [27:0] _T_136 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _T_167 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _T_194 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [6:0] _T_205 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_207 = {_T_205,io_in[6:2]}; // @[Cat.scala 29:58]
  wire [31:0] _T_213 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_221 = |io_in[11:7]; // @[RVC.scala 78:24]
  wire [6:0] _T_222 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[RVC.scala 78:20]
  wire [31:0] _T_233 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],_T_222}; // @[Cat.scala 29:58]
  wire [31:0] _T_249 = {_T_205,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_260 = |_T_207; // @[RVC.scala 91:29]
  wire [6:0] _T_261 = |_T_207 ? 7'h37 : 7'h3f; // @[RVC.scala 91:20]
  wire [14:0] _T_264 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_267 = {_T_264,io_in[6:2],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_271 = {_T_267[31:12],io_in[11:7],_T_261}; // @[Cat.scala 29:58]
  wire [6:0] _T_289 = _T_260 ? 7'h13 : 7'h1f; // @[RVC.scala 87:20]
  wire [2:0] _T_292 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_307 = {_T_292,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_289}; // @[Cat.scala 29:58]
  wire [31:0] _T_314_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? _T_307 : _T_271; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rd = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rs2 = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? _T_14 : _T_14; // @[RVC.scala 93:10]
  wire [4:0] _T_314_rs3 = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 93:10]
  wire [25:0] _T_325 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_0 = {{5'd0}, _T_325}; // @[RVC.scala 100:23]
  wire [30:0] _T_337 = _GEN_0 | 31'h40000000; // @[RVC.scala 100:23]
  wire [31:0] _T_350 = {_T_205,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [2:0] _T_353 = {io_in[12],io_in[6:5]}; // @[Cat.scala 29:58]
  wire [2:0] _T_355 = _T_353 == 3'h1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  wire [2:0] _T_357 = _T_353 == 3'h2 ? 3'h6 : _T_355; // @[package.scala 32:76]
  wire [2:0] _T_359 = _T_353 == 3'h3 ? 3'h7 : _T_357; // @[package.scala 32:76]
  wire [2:0] _T_361 = _T_353 == 3'h4 ? 3'h0 : _T_359; // @[package.scala 32:76]
  wire [2:0] _T_363 = _T_353 == 3'h5 ? 3'h0 : _T_361; // @[package.scala 32:76]
  wire [2:0] _T_365 = _T_353 == 3'h6 ? 3'h2 : _T_363; // @[package.scala 32:76]
  wire [2:0] _T_367 = _T_353 == 3'h7 ? 3'h3 : _T_365; // @[package.scala 32:76]
  wire [30:0] _T_370 = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[RVC.scala 104:22]
  wire [6:0] _T_372 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 105:22]
  wire [24:0] _T_382 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_T_367,2'h1,io_in[9:7],_T_372}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_1 = {{6'd0}, _T_382}; // @[RVC.scala 106:43]
  wire [30:0] _T_383 = _GEN_1 | _T_370; // @[RVC.scala 106:43]
  wire [30:0] _T_386 = io_in[11:10] == 2'h1 ? _T_337 : {{5'd0}, _T_325}; // @[package.scala 32:76]
  wire [31:0] _T_388 = io_in[11:10] == 2'h2 ? _T_350 : {{1'd0}, _T_386}; // @[package.scala 32:76]
  wire [31:0] _T_390 = io_in[11:10] == 2'h3 ? {{1'd0}, _T_383} : _T_388; // @[package.scala 32:76]
  wire [9:0] _T_401 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire [20:0] _T_416 = {_T_401,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_479 = {_T_416[20],_T_416[10:1],_T_416[11],_T_416[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] _T_488 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _T_497 = {_T_488,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_546 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58]
  wire [31:0] _T_613 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58]
  wire [6:0] _T_620 = _T_221 ? 7'h3 : 7'h1f; // @[RVC.scala 114:23]
  wire [25:0] _T_629 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _T_645 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [27:0] _T_660 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_620}; // @[Cat.scala 29:58]
  wire [28:0] _T_675 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],_T_620}; // @[Cat.scala 29:58]
  wire [24:0] _T_685 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_696 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_707 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [24:0] _T_709 = {_T_707[24:7],7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _T_712 = _T_221 ? _T_707 : _T_709; // @[RVC.scala 135:33]
  wire  _T_718 = |io_in[6:2]; // @[RVC.scala 136:27]
  wire [31:0] _T_689_bits = {{7'd0}, _T_685}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_716_bits = {{7'd0}, _T_712}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_719_bits = |io_in[6:2] ? _T_689_bits : _T_716_bits; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rd = |io_in[6:2] ? io_in[11:7] : 5'h0; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs1 = |io_in[6:2] ? 5'h0 : io_in[11:7]; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs2 = |io_in[6:2] ? io_in[6:2] : io_in[6:2]; // @[RVC.scala 136:22]
  wire [4:0] _T_719_rs3 = |io_in[6:2] ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 136:22]
  wire [24:0] _T_725 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _T_727 = {_T_707[24:7],7'h73}; // @[Cat.scala 29:58]
  wire [24:0] _T_728 = _T_727 | 25'h100000; // @[RVC.scala 138:46]
  wire [24:0] _T_731 = _T_221 ? _T_725 : _T_728; // @[RVC.scala 139:33]
  wire [31:0] _T_701_bits = {{7'd0}, _T_696}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_735_bits = {{7'd0}, _T_731}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_738_bits = _T_718 ? _T_701_bits : _T_735_bits; // @[RVC.scala 140:25]
  wire [4:0] _T_738_rd = _T_718 ? io_in[11:7] : 5'h1; // @[RVC.scala 140:25]
  wire [4:0] _T_738_rs1 = _T_718 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 140:25]
  wire [31:0] _T_740_bits = io_in[12] ? _T_738_bits : _T_719_bits; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rd = io_in[12] ? _T_738_rd : _T_719_rd; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs1 = io_in[12] ? _T_738_rs1 : _T_719_rs1; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs2 = io_in[12] ? _T_719_rs2 : _T_719_rs2; // @[RVC.scala 141:10]
  wire [4:0] _T_740_rs3 = io_in[12] ? _T_719_rs3 : _T_719_rs3; // @[RVC.scala 141:10]
  wire [8:0] _T_744 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [28:0] _T_756 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [7:0] _T_764 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_776 = {_T_764[7:5],io_in[6:2],5'h2,3'h2,_T_764[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [28:0] _T_796 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [4:0] _T_843 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 29:58]
  wire [31:0] _T_44_bits = {{4'd0}, _T_36}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_24_bits = {{2'd0}, _T_18}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_845_bits = _T_843 == 5'h1 ? _T_44_bits : _T_24_bits; // @[package.scala 32:76]
  wire [4:0] _T_845_rd = _T_843 == 5'h1 ? _T_14 : _T_14; // @[package.scala 32:76]
  wire [4:0] _T_845_rs1 = _T_843 == 5'h1 ? _T_30 : 5'h2; // @[package.scala 32:76]
  wire [4:0] _T_845_rs3 = _T_843 == 5'h1 ? io_in[31:27] : io_in[31:27]; // @[package.scala 32:76]
  wire [31:0] _T_66_bits = {{5'd0}, _T_58}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_847_bits = _T_843 == 5'h2 ? _T_66_bits : _T_845_bits; // @[package.scala 32:76]
  wire [4:0] _T_847_rd = _T_843 == 5'h2 ? _T_14 : _T_845_rd; // @[package.scala 32:76]
  wire [4:0] _T_847_rs1 = _T_843 == 5'h2 ? _T_30 : _T_845_rs1; // @[package.scala 32:76]
  wire [4:0] _T_847_rs3 = _T_843 == 5'h2 ? io_in[31:27] : _T_845_rs3; // @[package.scala 32:76]
  wire [31:0] _T_86_bits = {{4'd0}, _T_78}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_849_bits = _T_843 == 5'h3 ? _T_86_bits : _T_847_bits; // @[package.scala 32:76]
  wire [4:0] _T_849_rd = _T_843 == 5'h3 ? _T_14 : _T_847_rd; // @[package.scala 32:76]
  wire [4:0] _T_849_rs1 = _T_843 == 5'h3 ? _T_30 : _T_847_rs1; // @[package.scala 32:76]
  wire [4:0] _T_849_rs3 = _T_843 == 5'h3 ? io_in[31:27] : _T_847_rs3; // @[package.scala 32:76]
  wire [31:0] _T_117_bits = {{5'd0}, _T_109}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_851_bits = _T_843 == 5'h4 ? _T_117_bits : _T_849_bits; // @[package.scala 32:76]
  wire [4:0] _T_851_rd = _T_843 == 5'h4 ? _T_14 : _T_849_rd; // @[package.scala 32:76]
  wire [4:0] _T_851_rs1 = _T_843 == 5'h4 ? _T_30 : _T_849_rs1; // @[package.scala 32:76]
  wire [4:0] _T_851_rs3 = _T_843 == 5'h4 ? io_in[31:27] : _T_849_rs3; // @[package.scala 32:76]
  wire [31:0] _T_144_bits = {{4'd0}, _T_136}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_853_bits = _T_843 == 5'h5 ? _T_144_bits : _T_851_bits; // @[package.scala 32:76]
  wire [4:0] _T_853_rd = _T_843 == 5'h5 ? _T_14 : _T_851_rd; // @[package.scala 32:76]
  wire [4:0] _T_853_rs1 = _T_843 == 5'h5 ? _T_30 : _T_851_rs1; // @[package.scala 32:76]
  wire [4:0] _T_853_rs3 = _T_843 == 5'h5 ? io_in[31:27] : _T_851_rs3; // @[package.scala 32:76]
  wire [31:0] _T_175_bits = {{5'd0}, _T_167}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_855_bits = _T_843 == 5'h6 ? _T_175_bits : _T_853_bits; // @[package.scala 32:76]
  wire [4:0] _T_855_rd = _T_843 == 5'h6 ? _T_14 : _T_853_rd; // @[package.scala 32:76]
  wire [4:0] _T_855_rs1 = _T_843 == 5'h6 ? _T_30 : _T_853_rs1; // @[package.scala 32:76]
  wire [4:0] _T_855_rs3 = _T_843 == 5'h6 ? io_in[31:27] : _T_853_rs3; // @[package.scala 32:76]
  wire [31:0] _T_202_bits = {{4'd0}, _T_194}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_857_bits = _T_843 == 5'h7 ? _T_202_bits : _T_855_bits; // @[package.scala 32:76]
  wire [4:0] _T_857_rd = _T_843 == 5'h7 ? _T_14 : _T_855_rd; // @[package.scala 32:76]
  wire [4:0] _T_857_rs1 = _T_843 == 5'h7 ? _T_30 : _T_855_rs1; // @[package.scala 32:76]
  wire [4:0] _T_857_rs3 = _T_843 == 5'h7 ? io_in[31:27] : _T_855_rs3; // @[package.scala 32:76]
  wire [31:0] _T_859_bits = _T_843 == 5'h8 ? _T_213 : _T_857_bits; // @[package.scala 32:76]
  wire [4:0] _T_859_rd = _T_843 == 5'h8 ? io_in[11:7] : _T_857_rd; // @[package.scala 32:76]
  wire [4:0] _T_859_rs1 = _T_843 == 5'h8 ? io_in[11:7] : _T_857_rs1; // @[package.scala 32:76]
  wire [4:0] _T_859_rs2 = _T_843 == 5'h8 ? _T_14 : _T_857_rd; // @[package.scala 32:76]
  wire [4:0] _T_859_rs3 = _T_843 == 5'h8 ? io_in[31:27] : _T_857_rs3; // @[package.scala 32:76]
  wire [31:0] _T_861_bits = _T_843 == 5'h9 ? _T_233 : _T_859_bits; // @[package.scala 32:76]
  wire [4:0] _T_861_rd = _T_843 == 5'h9 ? io_in[11:7] : _T_859_rd; // @[package.scala 32:76]
  wire [4:0] _T_861_rs1 = _T_843 == 5'h9 ? io_in[11:7] : _T_859_rs1; // @[package.scala 32:76]
  wire [4:0] _T_861_rs2 = _T_843 == 5'h9 ? _T_14 : _T_859_rs2; // @[package.scala 32:76]
  wire [4:0] _T_861_rs3 = _T_843 == 5'h9 ? io_in[31:27] : _T_859_rs3; // @[package.scala 32:76]
  wire [31:0] _T_863_bits = _T_843 == 5'ha ? _T_249 : _T_861_bits; // @[package.scala 32:76]
  wire [4:0] _T_863_rd = _T_843 == 5'ha ? io_in[11:7] : _T_861_rd; // @[package.scala 32:76]
  wire [4:0] _T_863_rs1 = _T_843 == 5'ha ? 5'h0 : _T_861_rs1; // @[package.scala 32:76]
  wire [4:0] _T_863_rs2 = _T_843 == 5'ha ? _T_14 : _T_861_rs2; // @[package.scala 32:76]
  wire [4:0] _T_863_rs3 = _T_843 == 5'ha ? io_in[31:27] : _T_861_rs3; // @[package.scala 32:76]
  wire [31:0] _T_865_bits = _T_843 == 5'hb ? _T_314_bits : _T_863_bits; // @[package.scala 32:76]
  wire [4:0] _T_865_rd = _T_843 == 5'hb ? _T_314_rd : _T_863_rd; // @[package.scala 32:76]
  wire [4:0] _T_865_rs1 = _T_843 == 5'hb ? _T_314_rd : _T_863_rs1; // @[package.scala 32:76]
  wire [4:0] _T_865_rs2 = _T_843 == 5'hb ? _T_314_rs2 : _T_863_rs2; // @[package.scala 32:76]
  wire [4:0] _T_865_rs3 = _T_843 == 5'hb ? _T_314_rs3 : _T_863_rs3; // @[package.scala 32:76]
  wire [31:0] _T_867_bits = _T_843 == 5'hc ? _T_390 : _T_865_bits; // @[package.scala 32:76]
  wire [4:0] _T_867_rd = _T_843 == 5'hc ? _T_30 : _T_865_rd; // @[package.scala 32:76]
  wire [4:0] _T_867_rs1 = _T_843 == 5'hc ? _T_30 : _T_865_rs1; // @[package.scala 32:76]
  wire [4:0] _T_867_rs2 = _T_843 == 5'hc ? _T_14 : _T_865_rs2; // @[package.scala 32:76]
  wire [4:0] _T_867_rs3 = _T_843 == 5'hc ? io_in[31:27] : _T_865_rs3; // @[package.scala 32:76]
  wire [31:0] _T_869_bits = _T_843 == 5'hd ? _T_479 : _T_867_bits; // @[package.scala 32:76]
  wire [4:0] _T_869_rd = _T_843 == 5'hd ? 5'h0 : _T_867_rd; // @[package.scala 32:76]
  wire [4:0] _T_869_rs1 = _T_843 == 5'hd ? _T_30 : _T_867_rs1; // @[package.scala 32:76]
  wire [4:0] _T_869_rs2 = _T_843 == 5'hd ? _T_14 : _T_867_rs2; // @[package.scala 32:76]
  wire [4:0] _T_869_rs3 = _T_843 == 5'hd ? io_in[31:27] : _T_867_rs3; // @[package.scala 32:76]
  wire [31:0] _T_871_bits = _T_843 == 5'he ? _T_546 : _T_869_bits; // @[package.scala 32:76]
  wire [4:0] _T_871_rd = _T_843 == 5'he ? _T_30 : _T_869_rd; // @[package.scala 32:76]
  wire [4:0] _T_871_rs1 = _T_843 == 5'he ? _T_30 : _T_869_rs1; // @[package.scala 32:76]
  wire [4:0] _T_871_rs2 = _T_843 == 5'he ? 5'h0 : _T_869_rs2; // @[package.scala 32:76]
  wire [4:0] _T_871_rs3 = _T_843 == 5'he ? io_in[31:27] : _T_869_rs3; // @[package.scala 32:76]
  wire [31:0] _T_873_bits = _T_843 == 5'hf ? _T_613 : _T_871_bits; // @[package.scala 32:76]
  wire [4:0] _T_873_rd = _T_843 == 5'hf ? 5'h0 : _T_871_rd; // @[package.scala 32:76]
  wire [4:0] _T_873_rs1 = _T_843 == 5'hf ? _T_30 : _T_871_rs1; // @[package.scala 32:76]
  wire [4:0] _T_873_rs2 = _T_843 == 5'hf ? 5'h0 : _T_871_rs2; // @[package.scala 32:76]
  wire [4:0] _T_873_rs3 = _T_843 == 5'hf ? io_in[31:27] : _T_871_rs3; // @[package.scala 32:76]
  wire [31:0] _T_634_bits = {{6'd0}, _T_629}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_875_bits = _T_843 == 5'h10 ? _T_634_bits : _T_873_bits; // @[package.scala 32:76]
  wire [4:0] _T_875_rd = _T_843 == 5'h10 ? io_in[11:7] : _T_873_rd; // @[package.scala 32:76]
  wire [4:0] _T_875_rs1 = _T_843 == 5'h10 ? io_in[11:7] : _T_873_rs1; // @[package.scala 32:76]
  wire [4:0] _T_875_rs2 = _T_843 == 5'h10 ? io_in[6:2] : _T_873_rs2; // @[package.scala 32:76]
  wire [4:0] _T_875_rs3 = _T_843 == 5'h10 ? io_in[31:27] : _T_873_rs3; // @[package.scala 32:76]
  wire [31:0] _T_649_bits = {{3'd0}, _T_645}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_877_bits = _T_843 == 5'h11 ? _T_649_bits : _T_875_bits; // @[package.scala 32:76]
  wire [4:0] _T_877_rd = _T_843 == 5'h11 ? io_in[11:7] : _T_875_rd; // @[package.scala 32:76]
  wire [4:0] _T_877_rs1 = _T_843 == 5'h11 ? 5'h2 : _T_875_rs1; // @[package.scala 32:76]
  wire [4:0] _T_877_rs2 = _T_843 == 5'h11 ? io_in[6:2] : _T_875_rs2; // @[package.scala 32:76]
  wire [4:0] _T_877_rs3 = _T_843 == 5'h11 ? io_in[31:27] : _T_875_rs3; // @[package.scala 32:76]
  wire [31:0] _T_664_bits = {{4'd0}, _T_660}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_879_bits = _T_843 == 5'h12 ? _T_664_bits : _T_877_bits; // @[package.scala 32:76]
  wire [4:0] _T_879_rd = _T_843 == 5'h12 ? io_in[11:7] : _T_877_rd; // @[package.scala 32:76]
  wire [4:0] _T_879_rs1 = _T_843 == 5'h12 ? 5'h2 : _T_877_rs1; // @[package.scala 32:76]
  wire [4:0] _T_879_rs2 = _T_843 == 5'h12 ? io_in[6:2] : _T_877_rs2; // @[package.scala 32:76]
  wire [4:0] _T_879_rs3 = _T_843 == 5'h12 ? io_in[31:27] : _T_877_rs3; // @[package.scala 32:76]
  wire [31:0] _T_679_bits = {{3'd0}, _T_675}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_881_bits = _T_843 == 5'h13 ? _T_679_bits : _T_879_bits; // @[package.scala 32:76]
  wire [4:0] _T_881_rd = _T_843 == 5'h13 ? io_in[11:7] : _T_879_rd; // @[package.scala 32:76]
  wire [4:0] _T_881_rs1 = _T_843 == 5'h13 ? 5'h2 : _T_879_rs1; // @[package.scala 32:76]
  wire [4:0] _T_881_rs2 = _T_843 == 5'h13 ? io_in[6:2] : _T_879_rs2; // @[package.scala 32:76]
  wire [4:0] _T_881_rs3 = _T_843 == 5'h13 ? io_in[31:27] : _T_879_rs3; // @[package.scala 32:76]
  wire [31:0] _T_883_bits = _T_843 == 5'h14 ? _T_740_bits : _T_881_bits; // @[package.scala 32:76]
  wire [4:0] _T_883_rd = _T_843 == 5'h14 ? _T_740_rd : _T_881_rd; // @[package.scala 32:76]
  wire [4:0] _T_883_rs1 = _T_843 == 5'h14 ? _T_740_rs1 : _T_881_rs1; // @[package.scala 32:76]
  wire [4:0] _T_883_rs2 = _T_843 == 5'h14 ? _T_740_rs2 : _T_881_rs2; // @[package.scala 32:76]
  wire [4:0] _T_883_rs3 = _T_843 == 5'h14 ? _T_740_rs3 : _T_881_rs3; // @[package.scala 32:76]
  wire [31:0] _T_760_bits = {{3'd0}, _T_756}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_885_bits = _T_843 == 5'h15 ? _T_760_bits : _T_883_bits; // @[package.scala 32:76]
  wire [4:0] _T_885_rd = _T_843 == 5'h15 ? io_in[11:7] : _T_883_rd; // @[package.scala 32:76]
  wire [4:0] _T_885_rs1 = _T_843 == 5'h15 ? 5'h2 : _T_883_rs1; // @[package.scala 32:76]
  wire [4:0] _T_885_rs2 = _T_843 == 5'h15 ? io_in[6:2] : _T_883_rs2; // @[package.scala 32:76]
  wire [4:0] _T_885_rs3 = _T_843 == 5'h15 ? io_in[31:27] : _T_883_rs3; // @[package.scala 32:76]
  wire [31:0] _T_780_bits = {{4'd0}, _T_776}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_887_bits = _T_843 == 5'h16 ? _T_780_bits : _T_885_bits; // @[package.scala 32:76]
  wire [4:0] _T_887_rd = _T_843 == 5'h16 ? io_in[11:7] : _T_885_rd; // @[package.scala 32:76]
  wire [4:0] _T_887_rs1 = _T_843 == 5'h16 ? 5'h2 : _T_885_rs1; // @[package.scala 32:76]
  wire [4:0] _T_887_rs2 = _T_843 == 5'h16 ? io_in[6:2] : _T_885_rs2; // @[package.scala 32:76]
  wire [4:0] _T_887_rs3 = _T_843 == 5'h16 ? io_in[31:27] : _T_885_rs3; // @[package.scala 32:76]
  wire [31:0] _T_800_bits = {{3'd0}, _T_796}; // @[RVC.scala 22:19 23:14]
  wire [31:0] _T_889_bits = _T_843 == 5'h17 ? _T_800_bits : _T_887_bits; // @[package.scala 32:76]
  wire [4:0] _T_889_rd = _T_843 == 5'h17 ? io_in[11:7] : _T_887_rd; // @[package.scala 32:76]
  wire [4:0] _T_889_rs1 = _T_843 == 5'h17 ? 5'h2 : _T_887_rs1; // @[package.scala 32:76]
  wire [4:0] _T_889_rs2 = _T_843 == 5'h17 ? io_in[6:2] : _T_887_rs2; // @[package.scala 32:76]
  wire [4:0] _T_889_rs3 = _T_843 == 5'h17 ? io_in[31:27] : _T_887_rs3; // @[package.scala 32:76]
  wire [31:0] _T_891_bits = _T_843 == 5'h18 ? io_in : _T_889_bits; // @[package.scala 32:76]
  wire [4:0] _T_891_rd = _T_843 == 5'h18 ? io_in[11:7] : _T_889_rd; // @[package.scala 32:76]
  wire [4:0] _T_891_rs1 = _T_843 == 5'h18 ? io_in[19:15] : _T_889_rs1; // @[package.scala 32:76]
  wire [4:0] _T_891_rs2 = _T_843 == 5'h18 ? io_in[24:20] : _T_889_rs2; // @[package.scala 32:76]
  wire [4:0] _T_891_rs3 = _T_843 == 5'h18 ? io_in[31:27] : _T_889_rs3; // @[package.scala 32:76]
  wire [31:0] _T_893_bits = _T_843 == 5'h19 ? io_in : _T_891_bits; // @[package.scala 32:76]
  wire [4:0] _T_893_rd = _T_843 == 5'h19 ? io_in[11:7] : _T_891_rd; // @[package.scala 32:76]
  wire [4:0] _T_893_rs1 = _T_843 == 5'h19 ? io_in[19:15] : _T_891_rs1; // @[package.scala 32:76]
  wire [4:0] _T_893_rs2 = _T_843 == 5'h19 ? io_in[24:20] : _T_891_rs2; // @[package.scala 32:76]
  wire [4:0] _T_893_rs3 = _T_843 == 5'h19 ? io_in[31:27] : _T_891_rs3; // @[package.scala 32:76]
  wire [31:0] _T_895_bits = _T_843 == 5'h1a ? io_in : _T_893_bits; // @[package.scala 32:76]
  wire [4:0] _T_895_rd = _T_843 == 5'h1a ? io_in[11:7] : _T_893_rd; // @[package.scala 32:76]
  wire [4:0] _T_895_rs1 = _T_843 == 5'h1a ? io_in[19:15] : _T_893_rs1; // @[package.scala 32:76]
  wire [4:0] _T_895_rs2 = _T_843 == 5'h1a ? io_in[24:20] : _T_893_rs2; // @[package.scala 32:76]
  wire [4:0] _T_895_rs3 = _T_843 == 5'h1a ? io_in[31:27] : _T_893_rs3; // @[package.scala 32:76]
  wire [31:0] _T_897_bits = _T_843 == 5'h1b ? io_in : _T_895_bits; // @[package.scala 32:76]
  wire [4:0] _T_897_rd = _T_843 == 5'h1b ? io_in[11:7] : _T_895_rd; // @[package.scala 32:76]
  wire [4:0] _T_897_rs1 = _T_843 == 5'h1b ? io_in[19:15] : _T_895_rs1; // @[package.scala 32:76]
  wire [4:0] _T_897_rs2 = _T_843 == 5'h1b ? io_in[24:20] : _T_895_rs2; // @[package.scala 32:76]
  wire [4:0] _T_897_rs3 = _T_843 == 5'h1b ? io_in[31:27] : _T_895_rs3; // @[package.scala 32:76]
  wire [31:0] _T_899_bits = _T_843 == 5'h1c ? io_in : _T_897_bits; // @[package.scala 32:76]
  wire [4:0] _T_899_rd = _T_843 == 5'h1c ? io_in[11:7] : _T_897_rd; // @[package.scala 32:76]
  wire [4:0] _T_899_rs1 = _T_843 == 5'h1c ? io_in[19:15] : _T_897_rs1; // @[package.scala 32:76]
  wire [4:0] _T_899_rs2 = _T_843 == 5'h1c ? io_in[24:20] : _T_897_rs2; // @[package.scala 32:76]
  wire [4:0] _T_899_rs3 = _T_843 == 5'h1c ? io_in[31:27] : _T_897_rs3; // @[package.scala 32:76]
  wire [31:0] _T_901_bits = _T_843 == 5'h1d ? io_in : _T_899_bits; // @[package.scala 32:76]
  wire [4:0] _T_901_rd = _T_843 == 5'h1d ? io_in[11:7] : _T_899_rd; // @[package.scala 32:76]
  wire [4:0] _T_901_rs1 = _T_843 == 5'h1d ? io_in[19:15] : _T_899_rs1; // @[package.scala 32:76]
  wire [4:0] _T_901_rs2 = _T_843 == 5'h1d ? io_in[24:20] : _T_899_rs2; // @[package.scala 32:76]
  wire [4:0] _T_901_rs3 = _T_843 == 5'h1d ? io_in[31:27] : _T_899_rs3; // @[package.scala 32:76]
  wire [31:0] _T_903_bits = _T_843 == 5'h1e ? io_in : _T_901_bits; // @[package.scala 32:76]
  wire [4:0] _T_903_rd = _T_843 == 5'h1e ? io_in[11:7] : _T_901_rd; // @[package.scala 32:76]
  wire [4:0] _T_903_rs1 = _T_843 == 5'h1e ? io_in[19:15] : _T_901_rs1; // @[package.scala 32:76]
  wire [4:0] _T_903_rs2 = _T_843 == 5'h1e ? io_in[24:20] : _T_901_rs2; // @[package.scala 32:76]
  wire [4:0] _T_903_rs3 = _T_843 == 5'h1e ? io_in[31:27] : _T_901_rs3; // @[package.scala 32:76]
  assign io_out_bits = _T_843 == 5'h1f ? io_in : _T_903_bits; // @[package.scala 32:76]
  assign io_out_rd = _T_843 == 5'h1f ? io_in[11:7] : _T_903_rd; // @[package.scala 32:76]
  assign io_out_rs1 = _T_843 == 5'h1f ? io_in[19:15] : _T_903_rs1; // @[package.scala 32:76]
  assign io_out_rs2 = _T_843 == 5'h1f ? io_in[24:20] : _T_903_rs2; // @[package.scala 32:76]
  assign io_out_rs3 = _T_843 == 5'h1f ? io_in[31:27] : _T_903_rs3; // @[package.scala 32:76]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 164:26]
endmodule
