
module trivial_and (input [1:0] a, input [1:0] b, output [1:0] g);

assign g = a & b;

endmodule

