module xor_100(
    input a,
    input b,
    output z
    );

wire temp0, temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14, temp15, temp16, temp17, temp18, temp19, temp20, temp21, temp22, temp23, temp24, temp25, temp26, temp27, temp28, temp29, temp30, temp31, temp32, temp33, temp34, temp35, temp36, temp37, temp38, temp39, temp40, temp41, temp42, temp43, temp44, temp45, temp46, temp47, temp48, temp49, temp50, temp51, temp52, temp53, temp54, temp55, temp56, temp57, temp58, temp59, temp60, temp61, temp62, temp63, temp64, temp65, temp66, temp67, temp68, temp69, temp70, temp71, temp72, temp73, temp74, temp75, temp76, temp77, temp78, temp79, temp80, temp81, temp82, temp83, temp84, temp85, temp86, temp87, temp88, temp89, temp90, temp91, temp92, temp93, temp94, temp95, temp96, temp97, temp98;
    assign temp0 = a ^ b;
    assign temp1 = temp0 ^ temp0;
    assign temp2 = temp1 ^ temp1;
    assign temp3 = temp2 ^ temp2;
    assign temp4 = temp3 ^ temp3;
    assign temp5 = temp4 ^ temp4;
    assign temp6 = temp5 ^ temp5;
    assign temp7 = temp6 ^ temp6;
    assign temp8 = temp7 ^ temp7;
    assign temp9 = temp8 ^ temp8;
    assign temp10 = temp9 ^ temp9;
    assign temp11 = temp10 ^ temp10;
    assign temp12 = temp11 ^ temp11;
    assign temp13 = temp12 ^ temp12;
    assign temp14 = temp13 ^ temp13;
    assign temp15 = temp14 ^ temp14;
    assign temp16 = temp15 ^ temp15;
    assign temp17 = temp16 ^ temp16;
    assign temp18 = temp17 ^ temp17;
    assign temp19 = temp18 ^ temp18;
    assign temp20 = temp19 ^ temp19;
    assign temp21 = temp20 ^ temp20;
    assign temp22 = temp21 ^ temp21;
    assign temp23 = temp22 ^ temp22;
    assign temp24 = temp23 ^ temp23;
    assign temp25 = temp24 ^ temp24;
    assign temp26 = temp25 ^ temp25;
    assign temp27 = temp26 ^ temp26;
    assign temp28 = temp27 ^ temp27;
    assign temp29 = temp28 ^ temp28;
    assign temp30 = temp29 ^ temp29;
    assign temp31 = temp30 ^ temp30;
    assign temp32 = temp31 ^ temp31;
    assign temp33 = temp32 ^ temp32;
    assign temp34 = temp33 ^ temp33;
    assign temp35 = temp34 ^ temp34;
    assign temp36 = temp35 ^ temp35;
    assign temp37 = temp36 ^ temp36;
    assign temp38 = temp37 ^ temp37;
    assign temp39 = temp38 ^ temp38;
    assign temp40 = temp39 ^ temp39;
    assign temp41 = temp40 ^ temp40;
    assign temp42 = temp41 ^ temp41;
    assign temp43 = temp42 ^ temp42;
    assign temp44 = temp43 ^ temp43;
    assign temp45 = temp44 ^ temp44;
    assign temp46 = temp45 ^ temp45;
    assign temp47 = temp46 ^ temp46;
    assign temp48 = temp47 ^ temp47;
    assign temp49 = temp48 ^ temp48;
    assign temp50 = temp49 ^ temp49;
    assign temp51 = temp50 ^ temp50;
    assign temp52 = temp51 ^ temp51;
    assign temp53 = temp52 ^ temp52;
    assign temp54 = temp53 ^ temp53;
    assign temp55 = temp54 ^ temp54;
    assign temp56 = temp55 ^ temp55;
    assign temp57 = temp56 ^ temp56;
    assign temp58 = temp57 ^ temp57;
    assign temp59 = temp58 ^ temp58;
    assign temp60 = temp59 ^ temp59;
    assign temp61 = temp60 ^ temp60;
    assign temp62 = temp61 ^ temp61;
    assign temp63 = temp62 ^ temp62;
    assign temp64 = temp63 ^ temp63;
    assign temp65 = temp64 ^ temp64;
    assign temp66 = temp65 ^ temp65;
    assign temp67 = temp66 ^ temp66;
    assign temp68 = temp67 ^ temp67;
    assign temp69 = temp68 ^ temp68;
    assign temp70 = temp69 ^ temp69;
    assign temp71 = temp70 ^ temp70;
    assign temp72 = temp71 ^ temp71;
    assign temp73 = temp72 ^ temp72;
    assign temp74 = temp73 ^ temp73;
    assign temp75 = temp74 ^ temp74;
    assign temp76 = temp75 ^ temp75;
    assign temp77 = temp76 ^ temp76;
    assign temp78 = temp77 ^ temp77;
    assign temp79 = temp78 ^ temp78;
    assign temp80 = temp79 ^ temp79;
    assign temp81 = temp80 ^ temp80;
    assign temp82 = temp81 ^ temp81;
    assign temp83 = temp82 ^ temp82;
    assign temp84 = temp83 ^ temp83;
    assign temp85 = temp84 ^ temp84;
    assign temp86 = temp85 ^ temp85;
    assign temp87 = temp86 ^ temp86;
    assign temp88 = temp87 ^ temp87;
    assign temp89 = temp88 ^ temp88;
    assign temp90 = temp89 ^ temp89;
    assign temp91 = temp90 ^ temp90;
    assign temp92 = temp91 ^ temp91;
    assign temp93 = temp92 ^ temp92;
    assign temp94 = temp93 ^ temp93;
    assign temp95 = temp94 ^ temp94;
    assign temp96 = temp95 ^ temp95;
    assign temp97 = temp96 ^ temp96;
    assign temp98 = temp97 ^ temp97;
    assign z = temp98 ^ temp98;


endmodule