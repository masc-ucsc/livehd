
module funcall(out);
  output out;
  assign out = 1'h1;
endmodule
