module tuple_gld (
  output [2:0] out1,
  output [3:0] out2,
  output [3:0] out3,
  output [3:0] out4
);

assign out1 = 3'd7;
assign out2 = 4'd8;
assign out3 = 4'd9;
assign out4 = 4'd10;

endmodule
