module xor_1(
    input a,
    input b,
    output z
    );

    assign z = a ^ b;


endmodule