module tuple_empty_attr (
  output [7:0] out,
  output [7:0] out2
);

  assign out = 40;
  assign out2 = 3;

endmodule
