module xor_1000(
    input a,
    input b,
    output z
    );

wire temp0, temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14, temp15, temp16, temp17, temp18, temp19, temp20, temp21, temp22, temp23, temp24, temp25, temp26, temp27, temp28, temp29, temp30, temp31, temp32, temp33, temp34, temp35, temp36, temp37, temp38, temp39, temp40, temp41, temp42, temp43, temp44, temp45, temp46, temp47, temp48, temp49, temp50, temp51, temp52, temp53, temp54, temp55, temp56, temp57, temp58, temp59, temp60, temp61, temp62, temp63, temp64, temp65, temp66, temp67, temp68, temp69, temp70, temp71, temp72, temp73, temp74, temp75, temp76, temp77, temp78, temp79, temp80, temp81, temp82, temp83, temp84, temp85, temp86, temp87, temp88, temp89, temp90, temp91, temp92, temp93, temp94, temp95, temp96, temp97, temp98, temp99, temp100, temp101, temp102, temp103, temp104, temp105, temp106, temp107, temp108, temp109, temp110, temp111, temp112, temp113, temp114, temp115, temp116, temp117, temp118, temp119, temp120, temp121, temp122, temp123, temp124, temp125, temp126, temp127, temp128, temp129, temp130, temp131, temp132, temp133, temp134, temp135, temp136, temp137, temp138, temp139, temp140, temp141, temp142, temp143, temp144, temp145, temp146, temp147, temp148, temp149, temp150, temp151, temp152, temp153, temp154, temp155, temp156, temp157, temp158, temp159, temp160, temp161, temp162, temp163, temp164, temp165, temp166, temp167, temp168, temp169, temp170, temp171, temp172, temp173, temp174, temp175, temp176, temp177, temp178, temp179, temp180, temp181, temp182, temp183, temp184, temp185, temp186, temp187, temp188, temp189, temp190, temp191, temp192, temp193, temp194, temp195, temp196, temp197, temp198, temp199, temp200, temp201, temp202, temp203, temp204, temp205, temp206, temp207, temp208, temp209, temp210, temp211, temp212, temp213, temp214, temp215, temp216, temp217, temp218, temp219, temp220, temp221, temp222, temp223, temp224, temp225, temp226, temp227, temp228, temp229, temp230, temp231, temp232, temp233, temp234, temp235, temp236, temp237, temp238, temp239, temp240, temp241, temp242, temp243, temp244, temp245, temp246, temp247, temp248, temp249, temp250, temp251, temp252, temp253, temp254, temp255, temp256, temp257, temp258, temp259, temp260, temp261, temp262, temp263, temp264, temp265, temp266, temp267, temp268, temp269, temp270, temp271, temp272, temp273, temp274, temp275, temp276, temp277, temp278, temp279, temp280, temp281, temp282, temp283, temp284, temp285, temp286, temp287, temp288, temp289, temp290, temp291, temp292, temp293, temp294, temp295, temp296, temp297, temp298, temp299, temp300, temp301, temp302, temp303, temp304, temp305, temp306, temp307, temp308, temp309, temp310, temp311, temp312, temp313, temp314, temp315, temp316, temp317, temp318, temp319, temp320, temp321, temp322, temp323, temp324, temp325, temp326, temp327, temp328, temp329, temp330, temp331, temp332, temp333, temp334, temp335, temp336, temp337, temp338, temp339, temp340, temp341, temp342, temp343, temp344, temp345, temp346, temp347, temp348, temp349, temp350, temp351, temp352, temp353, temp354, temp355, temp356, temp357, temp358, temp359, temp360, temp361, temp362, temp363, temp364, temp365, temp366, temp367, temp368, temp369, temp370, temp371, temp372, temp373, temp374, temp375, temp376, temp377, temp378, temp379, temp380, temp381, temp382, temp383, temp384, temp385, temp386, temp387, temp388, temp389, temp390, temp391, temp392, temp393, temp394, temp395, temp396, temp397, temp398, temp399, temp400, temp401, temp402, temp403, temp404, temp405, temp406, temp407, temp408, temp409, temp410, temp411, temp412, temp413, temp414, temp415, temp416, temp417, temp418, temp419, temp420, temp421, temp422, temp423, temp424, temp425, temp426, temp427, temp428, temp429, temp430, temp431, temp432, temp433, temp434, temp435, temp436, temp437, temp438, temp439, temp440, temp441, temp442, temp443, temp444, temp445, temp446, temp447, temp448, temp449, temp450, temp451, temp452, temp453, temp454, temp455, temp456, temp457, temp458, temp459, temp460, temp461, temp462, temp463, temp464, temp465, temp466, temp467, temp468, temp469, temp470, temp471, temp472, temp473, temp474, temp475, temp476, temp477, temp478, temp479, temp480, temp481, temp482, temp483, temp484, temp485, temp486, temp487, temp488, temp489, temp490, temp491, temp492, temp493, temp494, temp495, temp496, temp497, temp498, temp499, temp500, temp501, temp502, temp503, temp504, temp505, temp506, temp507, temp508, temp509, temp510, temp511, temp512, temp513, temp514, temp515, temp516, temp517, temp518, temp519, temp520, temp521, temp522, temp523, temp524, temp525, temp526, temp527, temp528, temp529, temp530, temp531, temp532, temp533, temp534, temp535, temp536, temp537, temp538, temp539, temp540, temp541, temp542, temp543, temp544, temp545, temp546, temp547, temp548, temp549, temp550, temp551, temp552, temp553, temp554, temp555, temp556, temp557, temp558, temp559, temp560, temp561, temp562, temp563, temp564, temp565, temp566, temp567, temp568, temp569, temp570, temp571, temp572, temp573, temp574, temp575, temp576, temp577, temp578, temp579, temp580, temp581, temp582, temp583, temp584, temp585, temp586, temp587, temp588, temp589, temp590, temp591, temp592, temp593, temp594, temp595, temp596, temp597, temp598, temp599, temp600, temp601, temp602, temp603, temp604, temp605, temp606, temp607, temp608, temp609, temp610, temp611, temp612, temp613, temp614, temp615, temp616, temp617, temp618, temp619, temp620, temp621, temp622, temp623, temp624, temp625, temp626, temp627, temp628, temp629, temp630, temp631, temp632, temp633, temp634, temp635, temp636, temp637, temp638, temp639, temp640, temp641, temp642, temp643, temp644, temp645, temp646, temp647, temp648, temp649, temp650, temp651, temp652, temp653, temp654, temp655, temp656, temp657, temp658, temp659, temp660, temp661, temp662, temp663, temp664, temp665, temp666, temp667, temp668, temp669, temp670, temp671, temp672, temp673, temp674, temp675, temp676, temp677, temp678, temp679, temp680, temp681, temp682, temp683, temp684, temp685, temp686, temp687, temp688, temp689, temp690, temp691, temp692, temp693, temp694, temp695, temp696, temp697, temp698, temp699, temp700, temp701, temp702, temp703, temp704, temp705, temp706, temp707, temp708, temp709, temp710, temp711, temp712, temp713, temp714, temp715, temp716, temp717, temp718, temp719, temp720, temp721, temp722, temp723, temp724, temp725, temp726, temp727, temp728, temp729, temp730, temp731, temp732, temp733, temp734, temp735, temp736, temp737, temp738, temp739, temp740, temp741, temp742, temp743, temp744, temp745, temp746, temp747, temp748, temp749, temp750, temp751, temp752, temp753, temp754, temp755, temp756, temp757, temp758, temp759, temp760, temp761, temp762, temp763, temp764, temp765, temp766, temp767, temp768, temp769, temp770, temp771, temp772, temp773, temp774, temp775, temp776, temp777, temp778, temp779, temp780, temp781, temp782, temp783, temp784, temp785, temp786, temp787, temp788, temp789, temp790, temp791, temp792, temp793, temp794, temp795, temp796, temp797, temp798, temp799, temp800, temp801, temp802, temp803, temp804, temp805, temp806, temp807, temp808, temp809, temp810, temp811, temp812, temp813, temp814, temp815, temp816, temp817, temp818, temp819, temp820, temp821, temp822, temp823, temp824, temp825, temp826, temp827, temp828, temp829, temp830, temp831, temp832, temp833, temp834, temp835, temp836, temp837, temp838, temp839, temp840, temp841, temp842, temp843, temp844, temp845, temp846, temp847, temp848, temp849, temp850, temp851, temp852, temp853, temp854, temp855, temp856, temp857, temp858, temp859, temp860, temp861, temp862, temp863, temp864, temp865, temp866, temp867, temp868, temp869, temp870, temp871, temp872, temp873, temp874, temp875, temp876, temp877, temp878, temp879, temp880, temp881, temp882, temp883, temp884, temp885, temp886, temp887, temp888, temp889, temp890, temp891, temp892, temp893, temp894, temp895, temp896, temp897, temp898, temp899, temp900, temp901, temp902, temp903, temp904, temp905, temp906, temp907, temp908, temp909, temp910, temp911, temp912, temp913, temp914, temp915, temp916, temp917, temp918, temp919, temp920, temp921, temp922, temp923, temp924, temp925, temp926, temp927, temp928, temp929, temp930, temp931, temp932, temp933, temp934, temp935, temp936, temp937, temp938, temp939, temp940, temp941, temp942, temp943, temp944, temp945, temp946, temp947, temp948, temp949, temp950, temp951, temp952, temp953, temp954, temp955, temp956, temp957, temp958, temp959, temp960, temp961, temp962, temp963, temp964, temp965, temp966, temp967, temp968, temp969, temp970, temp971, temp972, temp973, temp974, temp975, temp976, temp977, temp978, temp979, temp980, temp981, temp982, temp983, temp984, temp985, temp986, temp987, temp988, temp989, temp990, temp991, temp992, temp993, temp994, temp995, temp996, temp997, temp998;
    assign temp0 = a ^ b;
    assign temp1 = temp0 ^ temp0;
    assign temp2 = temp1 ^ temp1;
    assign temp3 = temp2 ^ temp2;
    assign temp4 = temp3 ^ temp3;
    assign temp5 = temp4 ^ temp4;
    assign temp6 = temp5 ^ temp5;
    assign temp7 = temp6 ^ temp6;
    assign temp8 = temp7 ^ temp7;
    assign temp9 = temp8 ^ temp8;
    assign temp10 = temp9 ^ temp9;
    assign temp11 = temp10 ^ temp10;
    assign temp12 = temp11 ^ temp11;
    assign temp13 = temp12 ^ temp12;
    assign temp14 = temp13 ^ temp13;
    assign temp15 = temp14 ^ temp14;
    assign temp16 = temp15 ^ temp15;
    assign temp17 = temp16 ^ temp16;
    assign temp18 = temp17 ^ temp17;
    assign temp19 = temp18 ^ temp18;
    assign temp20 = temp19 ^ temp19;
    assign temp21 = temp20 ^ temp20;
    assign temp22 = temp21 ^ temp21;
    assign temp23 = temp22 ^ temp22;
    assign temp24 = temp23 ^ temp23;
    assign temp25 = temp24 ^ temp24;
    assign temp26 = temp25 ^ temp25;
    assign temp27 = temp26 ^ temp26;
    assign temp28 = temp27 ^ temp27;
    assign temp29 = temp28 ^ temp28;
    assign temp30 = temp29 ^ temp29;
    assign temp31 = temp30 ^ temp30;
    assign temp32 = temp31 ^ temp31;
    assign temp33 = temp32 ^ temp32;
    assign temp34 = temp33 ^ temp33;
    assign temp35 = temp34 ^ temp34;
    assign temp36 = temp35 ^ temp35;
    assign temp37 = temp36 ^ temp36;
    assign temp38 = temp37 ^ temp37;
    assign temp39 = temp38 ^ temp38;
    assign temp40 = temp39 ^ temp39;
    assign temp41 = temp40 ^ temp40;
    assign temp42 = temp41 ^ temp41;
    assign temp43 = temp42 ^ temp42;
    assign temp44 = temp43 ^ temp43;
    assign temp45 = temp44 ^ temp44;
    assign temp46 = temp45 ^ temp45;
    assign temp47 = temp46 ^ temp46;
    assign temp48 = temp47 ^ temp47;
    assign temp49 = temp48 ^ temp48;
    assign temp50 = temp49 ^ temp49;
    assign temp51 = temp50 ^ temp50;
    assign temp52 = temp51 ^ temp51;
    assign temp53 = temp52 ^ temp52;
    assign temp54 = temp53 ^ temp53;
    assign temp55 = temp54 ^ temp54;
    assign temp56 = temp55 ^ temp55;
    assign temp57 = temp56 ^ temp56;
    assign temp58 = temp57 ^ temp57;
    assign temp59 = temp58 ^ temp58;
    assign temp60 = temp59 ^ temp59;
    assign temp61 = temp60 ^ temp60;
    assign temp62 = temp61 ^ temp61;
    assign temp63 = temp62 ^ temp62;
    assign temp64 = temp63 ^ temp63;
    assign temp65 = temp64 ^ temp64;
    assign temp66 = temp65 ^ temp65;
    assign temp67 = temp66 ^ temp66;
    assign temp68 = temp67 ^ temp67;
    assign temp69 = temp68 ^ temp68;
    assign temp70 = temp69 ^ temp69;
    assign temp71 = temp70 ^ temp70;
    assign temp72 = temp71 ^ temp71;
    assign temp73 = temp72 ^ temp72;
    assign temp74 = temp73 ^ temp73;
    assign temp75 = temp74 ^ temp74;
    assign temp76 = temp75 ^ temp75;
    assign temp77 = temp76 ^ temp76;
    assign temp78 = temp77 ^ temp77;
    assign temp79 = temp78 ^ temp78;
    assign temp80 = temp79 ^ temp79;
    assign temp81 = temp80 ^ temp80;
    assign temp82 = temp81 ^ temp81;
    assign temp83 = temp82 ^ temp82;
    assign temp84 = temp83 ^ temp83;
    assign temp85 = temp84 ^ temp84;
    assign temp86 = temp85 ^ temp85;
    assign temp87 = temp86 ^ temp86;
    assign temp88 = temp87 ^ temp87;
    assign temp89 = temp88 ^ temp88;
    assign temp90 = temp89 ^ temp89;
    assign temp91 = temp90 ^ temp90;
    assign temp92 = temp91 ^ temp91;
    assign temp93 = temp92 ^ temp92;
    assign temp94 = temp93 ^ temp93;
    assign temp95 = temp94 ^ temp94;
    assign temp96 = temp95 ^ temp95;
    assign temp97 = temp96 ^ temp96;
    assign temp98 = temp97 ^ temp97;
    assign temp99 = temp98 ^ temp98;
    assign temp100 = temp99 ^ temp99;
    assign temp101 = temp100 ^ temp100;
    assign temp102 = temp101 ^ temp101;
    assign temp103 = temp102 ^ temp102;
    assign temp104 = temp103 ^ temp103;
    assign temp105 = temp104 ^ temp104;
    assign temp106 = temp105 ^ temp105;
    assign temp107 = temp106 ^ temp106;
    assign temp108 = temp107 ^ temp107;
    assign temp109 = temp108 ^ temp108;
    assign temp110 = temp109 ^ temp109;
    assign temp111 = temp110 ^ temp110;
    assign temp112 = temp111 ^ temp111;
    assign temp113 = temp112 ^ temp112;
    assign temp114 = temp113 ^ temp113;
    assign temp115 = temp114 ^ temp114;
    assign temp116 = temp115 ^ temp115;
    assign temp117 = temp116 ^ temp116;
    assign temp118 = temp117 ^ temp117;
    assign temp119 = temp118 ^ temp118;
    assign temp120 = temp119 ^ temp119;
    assign temp121 = temp120 ^ temp120;
    assign temp122 = temp121 ^ temp121;
    assign temp123 = temp122 ^ temp122;
    assign temp124 = temp123 ^ temp123;
    assign temp125 = temp124 ^ temp124;
    assign temp126 = temp125 ^ temp125;
    assign temp127 = temp126 ^ temp126;
    assign temp128 = temp127 ^ temp127;
    assign temp129 = temp128 ^ temp128;
    assign temp130 = temp129 ^ temp129;
    assign temp131 = temp130 ^ temp130;
    assign temp132 = temp131 ^ temp131;
    assign temp133 = temp132 ^ temp132;
    assign temp134 = temp133 ^ temp133;
    assign temp135 = temp134 ^ temp134;
    assign temp136 = temp135 ^ temp135;
    assign temp137 = temp136 ^ temp136;
    assign temp138 = temp137 ^ temp137;
    assign temp139 = temp138 ^ temp138;
    assign temp140 = temp139 ^ temp139;
    assign temp141 = temp140 ^ temp140;
    assign temp142 = temp141 ^ temp141;
    assign temp143 = temp142 ^ temp142;
    assign temp144 = temp143 ^ temp143;
    assign temp145 = temp144 ^ temp144;
    assign temp146 = temp145 ^ temp145;
    assign temp147 = temp146 ^ temp146;
    assign temp148 = temp147 ^ temp147;
    assign temp149 = temp148 ^ temp148;
    assign temp150 = temp149 ^ temp149;
    assign temp151 = temp150 ^ temp150;
    assign temp152 = temp151 ^ temp151;
    assign temp153 = temp152 ^ temp152;
    assign temp154 = temp153 ^ temp153;
    assign temp155 = temp154 ^ temp154;
    assign temp156 = temp155 ^ temp155;
    assign temp157 = temp156 ^ temp156;
    assign temp158 = temp157 ^ temp157;
    assign temp159 = temp158 ^ temp158;
    assign temp160 = temp159 ^ temp159;
    assign temp161 = temp160 ^ temp160;
    assign temp162 = temp161 ^ temp161;
    assign temp163 = temp162 ^ temp162;
    assign temp164 = temp163 ^ temp163;
    assign temp165 = temp164 ^ temp164;
    assign temp166 = temp165 ^ temp165;
    assign temp167 = temp166 ^ temp166;
    assign temp168 = temp167 ^ temp167;
    assign temp169 = temp168 ^ temp168;
    assign temp170 = temp169 ^ temp169;
    assign temp171 = temp170 ^ temp170;
    assign temp172 = temp171 ^ temp171;
    assign temp173 = temp172 ^ temp172;
    assign temp174 = temp173 ^ temp173;
    assign temp175 = temp174 ^ temp174;
    assign temp176 = temp175 ^ temp175;
    assign temp177 = temp176 ^ temp176;
    assign temp178 = temp177 ^ temp177;
    assign temp179 = temp178 ^ temp178;
    assign temp180 = temp179 ^ temp179;
    assign temp181 = temp180 ^ temp180;
    assign temp182 = temp181 ^ temp181;
    assign temp183 = temp182 ^ temp182;
    assign temp184 = temp183 ^ temp183;
    assign temp185 = temp184 ^ temp184;
    assign temp186 = temp185 ^ temp185;
    assign temp187 = temp186 ^ temp186;
    assign temp188 = temp187 ^ temp187;
    assign temp189 = temp188 ^ temp188;
    assign temp190 = temp189 ^ temp189;
    assign temp191 = temp190 ^ temp190;
    assign temp192 = temp191 ^ temp191;
    assign temp193 = temp192 ^ temp192;
    assign temp194 = temp193 ^ temp193;
    assign temp195 = temp194 ^ temp194;
    assign temp196 = temp195 ^ temp195;
    assign temp197 = temp196 ^ temp196;
    assign temp198 = temp197 ^ temp197;
    assign temp199 = temp198 ^ temp198;
    assign temp200 = temp199 ^ temp199;
    assign temp201 = temp200 ^ temp200;
    assign temp202 = temp201 ^ temp201;
    assign temp203 = temp202 ^ temp202;
    assign temp204 = temp203 ^ temp203;
    assign temp205 = temp204 ^ temp204;
    assign temp206 = temp205 ^ temp205;
    assign temp207 = temp206 ^ temp206;
    assign temp208 = temp207 ^ temp207;
    assign temp209 = temp208 ^ temp208;
    assign temp210 = temp209 ^ temp209;
    assign temp211 = temp210 ^ temp210;
    assign temp212 = temp211 ^ temp211;
    assign temp213 = temp212 ^ temp212;
    assign temp214 = temp213 ^ temp213;
    assign temp215 = temp214 ^ temp214;
    assign temp216 = temp215 ^ temp215;
    assign temp217 = temp216 ^ temp216;
    assign temp218 = temp217 ^ temp217;
    assign temp219 = temp218 ^ temp218;
    assign temp220 = temp219 ^ temp219;
    assign temp221 = temp220 ^ temp220;
    assign temp222 = temp221 ^ temp221;
    assign temp223 = temp222 ^ temp222;
    assign temp224 = temp223 ^ temp223;
    assign temp225 = temp224 ^ temp224;
    assign temp226 = temp225 ^ temp225;
    assign temp227 = temp226 ^ temp226;
    assign temp228 = temp227 ^ temp227;
    assign temp229 = temp228 ^ temp228;
    assign temp230 = temp229 ^ temp229;
    assign temp231 = temp230 ^ temp230;
    assign temp232 = temp231 ^ temp231;
    assign temp233 = temp232 ^ temp232;
    assign temp234 = temp233 ^ temp233;
    assign temp235 = temp234 ^ temp234;
    assign temp236 = temp235 ^ temp235;
    assign temp237 = temp236 ^ temp236;
    assign temp238 = temp237 ^ temp237;
    assign temp239 = temp238 ^ temp238;
    assign temp240 = temp239 ^ temp239;
    assign temp241 = temp240 ^ temp240;
    assign temp242 = temp241 ^ temp241;
    assign temp243 = temp242 ^ temp242;
    assign temp244 = temp243 ^ temp243;
    assign temp245 = temp244 ^ temp244;
    assign temp246 = temp245 ^ temp245;
    assign temp247 = temp246 ^ temp246;
    assign temp248 = temp247 ^ temp247;
    assign temp249 = temp248 ^ temp248;
    assign temp250 = temp249 ^ temp249;
    assign temp251 = temp250 ^ temp250;
    assign temp252 = temp251 ^ temp251;
    assign temp253 = temp252 ^ temp252;
    assign temp254 = temp253 ^ temp253;
    assign temp255 = temp254 ^ temp254;
    assign temp256 = temp255 ^ temp255;
    assign temp257 = temp256 ^ temp256;
    assign temp258 = temp257 ^ temp257;
    assign temp259 = temp258 ^ temp258;
    assign temp260 = temp259 ^ temp259;
    assign temp261 = temp260 ^ temp260;
    assign temp262 = temp261 ^ temp261;
    assign temp263 = temp262 ^ temp262;
    assign temp264 = temp263 ^ temp263;
    assign temp265 = temp264 ^ temp264;
    assign temp266 = temp265 ^ temp265;
    assign temp267 = temp266 ^ temp266;
    assign temp268 = temp267 ^ temp267;
    assign temp269 = temp268 ^ temp268;
    assign temp270 = temp269 ^ temp269;
    assign temp271 = temp270 ^ temp270;
    assign temp272 = temp271 ^ temp271;
    assign temp273 = temp272 ^ temp272;
    assign temp274 = temp273 ^ temp273;
    assign temp275 = temp274 ^ temp274;
    assign temp276 = temp275 ^ temp275;
    assign temp277 = temp276 ^ temp276;
    assign temp278 = temp277 ^ temp277;
    assign temp279 = temp278 ^ temp278;
    assign temp280 = temp279 ^ temp279;
    assign temp281 = temp280 ^ temp280;
    assign temp282 = temp281 ^ temp281;
    assign temp283 = temp282 ^ temp282;
    assign temp284 = temp283 ^ temp283;
    assign temp285 = temp284 ^ temp284;
    assign temp286 = temp285 ^ temp285;
    assign temp287 = temp286 ^ temp286;
    assign temp288 = temp287 ^ temp287;
    assign temp289 = temp288 ^ temp288;
    assign temp290 = temp289 ^ temp289;
    assign temp291 = temp290 ^ temp290;
    assign temp292 = temp291 ^ temp291;
    assign temp293 = temp292 ^ temp292;
    assign temp294 = temp293 ^ temp293;
    assign temp295 = temp294 ^ temp294;
    assign temp296 = temp295 ^ temp295;
    assign temp297 = temp296 ^ temp296;
    assign temp298 = temp297 ^ temp297;
    assign temp299 = temp298 ^ temp298;
    assign temp300 = temp299 ^ temp299;
    assign temp301 = temp300 ^ temp300;
    assign temp302 = temp301 ^ temp301;
    assign temp303 = temp302 ^ temp302;
    assign temp304 = temp303 ^ temp303;
    assign temp305 = temp304 ^ temp304;
    assign temp306 = temp305 ^ temp305;
    assign temp307 = temp306 ^ temp306;
    assign temp308 = temp307 ^ temp307;
    assign temp309 = temp308 ^ temp308;
    assign temp310 = temp309 ^ temp309;
    assign temp311 = temp310 ^ temp310;
    assign temp312 = temp311 ^ temp311;
    assign temp313 = temp312 ^ temp312;
    assign temp314 = temp313 ^ temp313;
    assign temp315 = temp314 ^ temp314;
    assign temp316 = temp315 ^ temp315;
    assign temp317 = temp316 ^ temp316;
    assign temp318 = temp317 ^ temp317;
    assign temp319 = temp318 ^ temp318;
    assign temp320 = temp319 ^ temp319;
    assign temp321 = temp320 ^ temp320;
    assign temp322 = temp321 ^ temp321;
    assign temp323 = temp322 ^ temp322;
    assign temp324 = temp323 ^ temp323;
    assign temp325 = temp324 ^ temp324;
    assign temp326 = temp325 ^ temp325;
    assign temp327 = temp326 ^ temp326;
    assign temp328 = temp327 ^ temp327;
    assign temp329 = temp328 ^ temp328;
    assign temp330 = temp329 ^ temp329;
    assign temp331 = temp330 ^ temp330;
    assign temp332 = temp331 ^ temp331;
    assign temp333 = temp332 ^ temp332;
    assign temp334 = temp333 ^ temp333;
    assign temp335 = temp334 ^ temp334;
    assign temp336 = temp335 ^ temp335;
    assign temp337 = temp336 ^ temp336;
    assign temp338 = temp337 ^ temp337;
    assign temp339 = temp338 ^ temp338;
    assign temp340 = temp339 ^ temp339;
    assign temp341 = temp340 ^ temp340;
    assign temp342 = temp341 ^ temp341;
    assign temp343 = temp342 ^ temp342;
    assign temp344 = temp343 ^ temp343;
    assign temp345 = temp344 ^ temp344;
    assign temp346 = temp345 ^ temp345;
    assign temp347 = temp346 ^ temp346;
    assign temp348 = temp347 ^ temp347;
    assign temp349 = temp348 ^ temp348;
    assign temp350 = temp349 ^ temp349;
    assign temp351 = temp350 ^ temp350;
    assign temp352 = temp351 ^ temp351;
    assign temp353 = temp352 ^ temp352;
    assign temp354 = temp353 ^ temp353;
    assign temp355 = temp354 ^ temp354;
    assign temp356 = temp355 ^ temp355;
    assign temp357 = temp356 ^ temp356;
    assign temp358 = temp357 ^ temp357;
    assign temp359 = temp358 ^ temp358;
    assign temp360 = temp359 ^ temp359;
    assign temp361 = temp360 ^ temp360;
    assign temp362 = temp361 ^ temp361;
    assign temp363 = temp362 ^ temp362;
    assign temp364 = temp363 ^ temp363;
    assign temp365 = temp364 ^ temp364;
    assign temp366 = temp365 ^ temp365;
    assign temp367 = temp366 ^ temp366;
    assign temp368 = temp367 ^ temp367;
    assign temp369 = temp368 ^ temp368;
    assign temp370 = temp369 ^ temp369;
    assign temp371 = temp370 ^ temp370;
    assign temp372 = temp371 ^ temp371;
    assign temp373 = temp372 ^ temp372;
    assign temp374 = temp373 ^ temp373;
    assign temp375 = temp374 ^ temp374;
    assign temp376 = temp375 ^ temp375;
    assign temp377 = temp376 ^ temp376;
    assign temp378 = temp377 ^ temp377;
    assign temp379 = temp378 ^ temp378;
    assign temp380 = temp379 ^ temp379;
    assign temp381 = temp380 ^ temp380;
    assign temp382 = temp381 ^ temp381;
    assign temp383 = temp382 ^ temp382;
    assign temp384 = temp383 ^ temp383;
    assign temp385 = temp384 ^ temp384;
    assign temp386 = temp385 ^ temp385;
    assign temp387 = temp386 ^ temp386;
    assign temp388 = temp387 ^ temp387;
    assign temp389 = temp388 ^ temp388;
    assign temp390 = temp389 ^ temp389;
    assign temp391 = temp390 ^ temp390;
    assign temp392 = temp391 ^ temp391;
    assign temp393 = temp392 ^ temp392;
    assign temp394 = temp393 ^ temp393;
    assign temp395 = temp394 ^ temp394;
    assign temp396 = temp395 ^ temp395;
    assign temp397 = temp396 ^ temp396;
    assign temp398 = temp397 ^ temp397;
    assign temp399 = temp398 ^ temp398;
    assign temp400 = temp399 ^ temp399;
    assign temp401 = temp400 ^ temp400;
    assign temp402 = temp401 ^ temp401;
    assign temp403 = temp402 ^ temp402;
    assign temp404 = temp403 ^ temp403;
    assign temp405 = temp404 ^ temp404;
    assign temp406 = temp405 ^ temp405;
    assign temp407 = temp406 ^ temp406;
    assign temp408 = temp407 ^ temp407;
    assign temp409 = temp408 ^ temp408;
    assign temp410 = temp409 ^ temp409;
    assign temp411 = temp410 ^ temp410;
    assign temp412 = temp411 ^ temp411;
    assign temp413 = temp412 ^ temp412;
    assign temp414 = temp413 ^ temp413;
    assign temp415 = temp414 ^ temp414;
    assign temp416 = temp415 ^ temp415;
    assign temp417 = temp416 ^ temp416;
    assign temp418 = temp417 ^ temp417;
    assign temp419 = temp418 ^ temp418;
    assign temp420 = temp419 ^ temp419;
    assign temp421 = temp420 ^ temp420;
    assign temp422 = temp421 ^ temp421;
    assign temp423 = temp422 ^ temp422;
    assign temp424 = temp423 ^ temp423;
    assign temp425 = temp424 ^ temp424;
    assign temp426 = temp425 ^ temp425;
    assign temp427 = temp426 ^ temp426;
    assign temp428 = temp427 ^ temp427;
    assign temp429 = temp428 ^ temp428;
    assign temp430 = temp429 ^ temp429;
    assign temp431 = temp430 ^ temp430;
    assign temp432 = temp431 ^ temp431;
    assign temp433 = temp432 ^ temp432;
    assign temp434 = temp433 ^ temp433;
    assign temp435 = temp434 ^ temp434;
    assign temp436 = temp435 ^ temp435;
    assign temp437 = temp436 ^ temp436;
    assign temp438 = temp437 ^ temp437;
    assign temp439 = temp438 ^ temp438;
    assign temp440 = temp439 ^ temp439;
    assign temp441 = temp440 ^ temp440;
    assign temp442 = temp441 ^ temp441;
    assign temp443 = temp442 ^ temp442;
    assign temp444 = temp443 ^ temp443;
    assign temp445 = temp444 ^ temp444;
    assign temp446 = temp445 ^ temp445;
    assign temp447 = temp446 ^ temp446;
    assign temp448 = temp447 ^ temp447;
    assign temp449 = temp448 ^ temp448;
    assign temp450 = temp449 ^ temp449;
    assign temp451 = temp450 ^ temp450;
    assign temp452 = temp451 ^ temp451;
    assign temp453 = temp452 ^ temp452;
    assign temp454 = temp453 ^ temp453;
    assign temp455 = temp454 ^ temp454;
    assign temp456 = temp455 ^ temp455;
    assign temp457 = temp456 ^ temp456;
    assign temp458 = temp457 ^ temp457;
    assign temp459 = temp458 ^ temp458;
    assign temp460 = temp459 ^ temp459;
    assign temp461 = temp460 ^ temp460;
    assign temp462 = temp461 ^ temp461;
    assign temp463 = temp462 ^ temp462;
    assign temp464 = temp463 ^ temp463;
    assign temp465 = temp464 ^ temp464;
    assign temp466 = temp465 ^ temp465;
    assign temp467 = temp466 ^ temp466;
    assign temp468 = temp467 ^ temp467;
    assign temp469 = temp468 ^ temp468;
    assign temp470 = temp469 ^ temp469;
    assign temp471 = temp470 ^ temp470;
    assign temp472 = temp471 ^ temp471;
    assign temp473 = temp472 ^ temp472;
    assign temp474 = temp473 ^ temp473;
    assign temp475 = temp474 ^ temp474;
    assign temp476 = temp475 ^ temp475;
    assign temp477 = temp476 ^ temp476;
    assign temp478 = temp477 ^ temp477;
    assign temp479 = temp478 ^ temp478;
    assign temp480 = temp479 ^ temp479;
    assign temp481 = temp480 ^ temp480;
    assign temp482 = temp481 ^ temp481;
    assign temp483 = temp482 ^ temp482;
    assign temp484 = temp483 ^ temp483;
    assign temp485 = temp484 ^ temp484;
    assign temp486 = temp485 ^ temp485;
    assign temp487 = temp486 ^ temp486;
    assign temp488 = temp487 ^ temp487;
    assign temp489 = temp488 ^ temp488;
    assign temp490 = temp489 ^ temp489;
    assign temp491 = temp490 ^ temp490;
    assign temp492 = temp491 ^ temp491;
    assign temp493 = temp492 ^ temp492;
    assign temp494 = temp493 ^ temp493;
    assign temp495 = temp494 ^ temp494;
    assign temp496 = temp495 ^ temp495;
    assign temp497 = temp496 ^ temp496;
    assign temp498 = temp497 ^ temp497;
    assign temp499 = temp498 ^ temp498;
    assign temp500 = temp499 ^ temp499;
    assign temp501 = temp500 ^ temp500;
    assign temp502 = temp501 ^ temp501;
    assign temp503 = temp502 ^ temp502;
    assign temp504 = temp503 ^ temp503;
    assign temp505 = temp504 ^ temp504;
    assign temp506 = temp505 ^ temp505;
    assign temp507 = temp506 ^ temp506;
    assign temp508 = temp507 ^ temp507;
    assign temp509 = temp508 ^ temp508;
    assign temp510 = temp509 ^ temp509;
    assign temp511 = temp510 ^ temp510;
    assign temp512 = temp511 ^ temp511;
    assign temp513 = temp512 ^ temp512;
    assign temp514 = temp513 ^ temp513;
    assign temp515 = temp514 ^ temp514;
    assign temp516 = temp515 ^ temp515;
    assign temp517 = temp516 ^ temp516;
    assign temp518 = temp517 ^ temp517;
    assign temp519 = temp518 ^ temp518;
    assign temp520 = temp519 ^ temp519;
    assign temp521 = temp520 ^ temp520;
    assign temp522 = temp521 ^ temp521;
    assign temp523 = temp522 ^ temp522;
    assign temp524 = temp523 ^ temp523;
    assign temp525 = temp524 ^ temp524;
    assign temp526 = temp525 ^ temp525;
    assign temp527 = temp526 ^ temp526;
    assign temp528 = temp527 ^ temp527;
    assign temp529 = temp528 ^ temp528;
    assign temp530 = temp529 ^ temp529;
    assign temp531 = temp530 ^ temp530;
    assign temp532 = temp531 ^ temp531;
    assign temp533 = temp532 ^ temp532;
    assign temp534 = temp533 ^ temp533;
    assign temp535 = temp534 ^ temp534;
    assign temp536 = temp535 ^ temp535;
    assign temp537 = temp536 ^ temp536;
    assign temp538 = temp537 ^ temp537;
    assign temp539 = temp538 ^ temp538;
    assign temp540 = temp539 ^ temp539;
    assign temp541 = temp540 ^ temp540;
    assign temp542 = temp541 ^ temp541;
    assign temp543 = temp542 ^ temp542;
    assign temp544 = temp543 ^ temp543;
    assign temp545 = temp544 ^ temp544;
    assign temp546 = temp545 ^ temp545;
    assign temp547 = temp546 ^ temp546;
    assign temp548 = temp547 ^ temp547;
    assign temp549 = temp548 ^ temp548;
    assign temp550 = temp549 ^ temp549;
    assign temp551 = temp550 ^ temp550;
    assign temp552 = temp551 ^ temp551;
    assign temp553 = temp552 ^ temp552;
    assign temp554 = temp553 ^ temp553;
    assign temp555 = temp554 ^ temp554;
    assign temp556 = temp555 ^ temp555;
    assign temp557 = temp556 ^ temp556;
    assign temp558 = temp557 ^ temp557;
    assign temp559 = temp558 ^ temp558;
    assign temp560 = temp559 ^ temp559;
    assign temp561 = temp560 ^ temp560;
    assign temp562 = temp561 ^ temp561;
    assign temp563 = temp562 ^ temp562;
    assign temp564 = temp563 ^ temp563;
    assign temp565 = temp564 ^ temp564;
    assign temp566 = temp565 ^ temp565;
    assign temp567 = temp566 ^ temp566;
    assign temp568 = temp567 ^ temp567;
    assign temp569 = temp568 ^ temp568;
    assign temp570 = temp569 ^ temp569;
    assign temp571 = temp570 ^ temp570;
    assign temp572 = temp571 ^ temp571;
    assign temp573 = temp572 ^ temp572;
    assign temp574 = temp573 ^ temp573;
    assign temp575 = temp574 ^ temp574;
    assign temp576 = temp575 ^ temp575;
    assign temp577 = temp576 ^ temp576;
    assign temp578 = temp577 ^ temp577;
    assign temp579 = temp578 ^ temp578;
    assign temp580 = temp579 ^ temp579;
    assign temp581 = temp580 ^ temp580;
    assign temp582 = temp581 ^ temp581;
    assign temp583 = temp582 ^ temp582;
    assign temp584 = temp583 ^ temp583;
    assign temp585 = temp584 ^ temp584;
    assign temp586 = temp585 ^ temp585;
    assign temp587 = temp586 ^ temp586;
    assign temp588 = temp587 ^ temp587;
    assign temp589 = temp588 ^ temp588;
    assign temp590 = temp589 ^ temp589;
    assign temp591 = temp590 ^ temp590;
    assign temp592 = temp591 ^ temp591;
    assign temp593 = temp592 ^ temp592;
    assign temp594 = temp593 ^ temp593;
    assign temp595 = temp594 ^ temp594;
    assign temp596 = temp595 ^ temp595;
    assign temp597 = temp596 ^ temp596;
    assign temp598 = temp597 ^ temp597;
    assign temp599 = temp598 ^ temp598;
    assign temp600 = temp599 ^ temp599;
    assign temp601 = temp600 ^ temp600;
    assign temp602 = temp601 ^ temp601;
    assign temp603 = temp602 ^ temp602;
    assign temp604 = temp603 ^ temp603;
    assign temp605 = temp604 ^ temp604;
    assign temp606 = temp605 ^ temp605;
    assign temp607 = temp606 ^ temp606;
    assign temp608 = temp607 ^ temp607;
    assign temp609 = temp608 ^ temp608;
    assign temp610 = temp609 ^ temp609;
    assign temp611 = temp610 ^ temp610;
    assign temp612 = temp611 ^ temp611;
    assign temp613 = temp612 ^ temp612;
    assign temp614 = temp613 ^ temp613;
    assign temp615 = temp614 ^ temp614;
    assign temp616 = temp615 ^ temp615;
    assign temp617 = temp616 ^ temp616;
    assign temp618 = temp617 ^ temp617;
    assign temp619 = temp618 ^ temp618;
    assign temp620 = temp619 ^ temp619;
    assign temp621 = temp620 ^ temp620;
    assign temp622 = temp621 ^ temp621;
    assign temp623 = temp622 ^ temp622;
    assign temp624 = temp623 ^ temp623;
    assign temp625 = temp624 ^ temp624;
    assign temp626 = temp625 ^ temp625;
    assign temp627 = temp626 ^ temp626;
    assign temp628 = temp627 ^ temp627;
    assign temp629 = temp628 ^ temp628;
    assign temp630 = temp629 ^ temp629;
    assign temp631 = temp630 ^ temp630;
    assign temp632 = temp631 ^ temp631;
    assign temp633 = temp632 ^ temp632;
    assign temp634 = temp633 ^ temp633;
    assign temp635 = temp634 ^ temp634;
    assign temp636 = temp635 ^ temp635;
    assign temp637 = temp636 ^ temp636;
    assign temp638 = temp637 ^ temp637;
    assign temp639 = temp638 ^ temp638;
    assign temp640 = temp639 ^ temp639;
    assign temp641 = temp640 ^ temp640;
    assign temp642 = temp641 ^ temp641;
    assign temp643 = temp642 ^ temp642;
    assign temp644 = temp643 ^ temp643;
    assign temp645 = temp644 ^ temp644;
    assign temp646 = temp645 ^ temp645;
    assign temp647 = temp646 ^ temp646;
    assign temp648 = temp647 ^ temp647;
    assign temp649 = temp648 ^ temp648;
    assign temp650 = temp649 ^ temp649;
    assign temp651 = temp650 ^ temp650;
    assign temp652 = temp651 ^ temp651;
    assign temp653 = temp652 ^ temp652;
    assign temp654 = temp653 ^ temp653;
    assign temp655 = temp654 ^ temp654;
    assign temp656 = temp655 ^ temp655;
    assign temp657 = temp656 ^ temp656;
    assign temp658 = temp657 ^ temp657;
    assign temp659 = temp658 ^ temp658;
    assign temp660 = temp659 ^ temp659;
    assign temp661 = temp660 ^ temp660;
    assign temp662 = temp661 ^ temp661;
    assign temp663 = temp662 ^ temp662;
    assign temp664 = temp663 ^ temp663;
    assign temp665 = temp664 ^ temp664;
    assign temp666 = temp665 ^ temp665;
    assign temp667 = temp666 ^ temp666;
    assign temp668 = temp667 ^ temp667;
    assign temp669 = temp668 ^ temp668;
    assign temp670 = temp669 ^ temp669;
    assign temp671 = temp670 ^ temp670;
    assign temp672 = temp671 ^ temp671;
    assign temp673 = temp672 ^ temp672;
    assign temp674 = temp673 ^ temp673;
    assign temp675 = temp674 ^ temp674;
    assign temp676 = temp675 ^ temp675;
    assign temp677 = temp676 ^ temp676;
    assign temp678 = temp677 ^ temp677;
    assign temp679 = temp678 ^ temp678;
    assign temp680 = temp679 ^ temp679;
    assign temp681 = temp680 ^ temp680;
    assign temp682 = temp681 ^ temp681;
    assign temp683 = temp682 ^ temp682;
    assign temp684 = temp683 ^ temp683;
    assign temp685 = temp684 ^ temp684;
    assign temp686 = temp685 ^ temp685;
    assign temp687 = temp686 ^ temp686;
    assign temp688 = temp687 ^ temp687;
    assign temp689 = temp688 ^ temp688;
    assign temp690 = temp689 ^ temp689;
    assign temp691 = temp690 ^ temp690;
    assign temp692 = temp691 ^ temp691;
    assign temp693 = temp692 ^ temp692;
    assign temp694 = temp693 ^ temp693;
    assign temp695 = temp694 ^ temp694;
    assign temp696 = temp695 ^ temp695;
    assign temp697 = temp696 ^ temp696;
    assign temp698 = temp697 ^ temp697;
    assign temp699 = temp698 ^ temp698;
    assign temp700 = temp699 ^ temp699;
    assign temp701 = temp700 ^ temp700;
    assign temp702 = temp701 ^ temp701;
    assign temp703 = temp702 ^ temp702;
    assign temp704 = temp703 ^ temp703;
    assign temp705 = temp704 ^ temp704;
    assign temp706 = temp705 ^ temp705;
    assign temp707 = temp706 ^ temp706;
    assign temp708 = temp707 ^ temp707;
    assign temp709 = temp708 ^ temp708;
    assign temp710 = temp709 ^ temp709;
    assign temp711 = temp710 ^ temp710;
    assign temp712 = temp711 ^ temp711;
    assign temp713 = temp712 ^ temp712;
    assign temp714 = temp713 ^ temp713;
    assign temp715 = temp714 ^ temp714;
    assign temp716 = temp715 ^ temp715;
    assign temp717 = temp716 ^ temp716;
    assign temp718 = temp717 ^ temp717;
    assign temp719 = temp718 ^ temp718;
    assign temp720 = temp719 ^ temp719;
    assign temp721 = temp720 ^ temp720;
    assign temp722 = temp721 ^ temp721;
    assign temp723 = temp722 ^ temp722;
    assign temp724 = temp723 ^ temp723;
    assign temp725 = temp724 ^ temp724;
    assign temp726 = temp725 ^ temp725;
    assign temp727 = temp726 ^ temp726;
    assign temp728 = temp727 ^ temp727;
    assign temp729 = temp728 ^ temp728;
    assign temp730 = temp729 ^ temp729;
    assign temp731 = temp730 ^ temp730;
    assign temp732 = temp731 ^ temp731;
    assign temp733 = temp732 ^ temp732;
    assign temp734 = temp733 ^ temp733;
    assign temp735 = temp734 ^ temp734;
    assign temp736 = temp735 ^ temp735;
    assign temp737 = temp736 ^ temp736;
    assign temp738 = temp737 ^ temp737;
    assign temp739 = temp738 ^ temp738;
    assign temp740 = temp739 ^ temp739;
    assign temp741 = temp740 ^ temp740;
    assign temp742 = temp741 ^ temp741;
    assign temp743 = temp742 ^ temp742;
    assign temp744 = temp743 ^ temp743;
    assign temp745 = temp744 ^ temp744;
    assign temp746 = temp745 ^ temp745;
    assign temp747 = temp746 ^ temp746;
    assign temp748 = temp747 ^ temp747;
    assign temp749 = temp748 ^ temp748;
    assign temp750 = temp749 ^ temp749;
    assign temp751 = temp750 ^ temp750;
    assign temp752 = temp751 ^ temp751;
    assign temp753 = temp752 ^ temp752;
    assign temp754 = temp753 ^ temp753;
    assign temp755 = temp754 ^ temp754;
    assign temp756 = temp755 ^ temp755;
    assign temp757 = temp756 ^ temp756;
    assign temp758 = temp757 ^ temp757;
    assign temp759 = temp758 ^ temp758;
    assign temp760 = temp759 ^ temp759;
    assign temp761 = temp760 ^ temp760;
    assign temp762 = temp761 ^ temp761;
    assign temp763 = temp762 ^ temp762;
    assign temp764 = temp763 ^ temp763;
    assign temp765 = temp764 ^ temp764;
    assign temp766 = temp765 ^ temp765;
    assign temp767 = temp766 ^ temp766;
    assign temp768 = temp767 ^ temp767;
    assign temp769 = temp768 ^ temp768;
    assign temp770 = temp769 ^ temp769;
    assign temp771 = temp770 ^ temp770;
    assign temp772 = temp771 ^ temp771;
    assign temp773 = temp772 ^ temp772;
    assign temp774 = temp773 ^ temp773;
    assign temp775 = temp774 ^ temp774;
    assign temp776 = temp775 ^ temp775;
    assign temp777 = temp776 ^ temp776;
    assign temp778 = temp777 ^ temp777;
    assign temp779 = temp778 ^ temp778;
    assign temp780 = temp779 ^ temp779;
    assign temp781 = temp780 ^ temp780;
    assign temp782 = temp781 ^ temp781;
    assign temp783 = temp782 ^ temp782;
    assign temp784 = temp783 ^ temp783;
    assign temp785 = temp784 ^ temp784;
    assign temp786 = temp785 ^ temp785;
    assign temp787 = temp786 ^ temp786;
    assign temp788 = temp787 ^ temp787;
    assign temp789 = temp788 ^ temp788;
    assign temp790 = temp789 ^ temp789;
    assign temp791 = temp790 ^ temp790;
    assign temp792 = temp791 ^ temp791;
    assign temp793 = temp792 ^ temp792;
    assign temp794 = temp793 ^ temp793;
    assign temp795 = temp794 ^ temp794;
    assign temp796 = temp795 ^ temp795;
    assign temp797 = temp796 ^ temp796;
    assign temp798 = temp797 ^ temp797;
    assign temp799 = temp798 ^ temp798;
    assign temp800 = temp799 ^ temp799;
    assign temp801 = temp800 ^ temp800;
    assign temp802 = temp801 ^ temp801;
    assign temp803 = temp802 ^ temp802;
    assign temp804 = temp803 ^ temp803;
    assign temp805 = temp804 ^ temp804;
    assign temp806 = temp805 ^ temp805;
    assign temp807 = temp806 ^ temp806;
    assign temp808 = temp807 ^ temp807;
    assign temp809 = temp808 ^ temp808;
    assign temp810 = temp809 ^ temp809;
    assign temp811 = temp810 ^ temp810;
    assign temp812 = temp811 ^ temp811;
    assign temp813 = temp812 ^ temp812;
    assign temp814 = temp813 ^ temp813;
    assign temp815 = temp814 ^ temp814;
    assign temp816 = temp815 ^ temp815;
    assign temp817 = temp816 ^ temp816;
    assign temp818 = temp817 ^ temp817;
    assign temp819 = temp818 ^ temp818;
    assign temp820 = temp819 ^ temp819;
    assign temp821 = temp820 ^ temp820;
    assign temp822 = temp821 ^ temp821;
    assign temp823 = temp822 ^ temp822;
    assign temp824 = temp823 ^ temp823;
    assign temp825 = temp824 ^ temp824;
    assign temp826 = temp825 ^ temp825;
    assign temp827 = temp826 ^ temp826;
    assign temp828 = temp827 ^ temp827;
    assign temp829 = temp828 ^ temp828;
    assign temp830 = temp829 ^ temp829;
    assign temp831 = temp830 ^ temp830;
    assign temp832 = temp831 ^ temp831;
    assign temp833 = temp832 ^ temp832;
    assign temp834 = temp833 ^ temp833;
    assign temp835 = temp834 ^ temp834;
    assign temp836 = temp835 ^ temp835;
    assign temp837 = temp836 ^ temp836;
    assign temp838 = temp837 ^ temp837;
    assign temp839 = temp838 ^ temp838;
    assign temp840 = temp839 ^ temp839;
    assign temp841 = temp840 ^ temp840;
    assign temp842 = temp841 ^ temp841;
    assign temp843 = temp842 ^ temp842;
    assign temp844 = temp843 ^ temp843;
    assign temp845 = temp844 ^ temp844;
    assign temp846 = temp845 ^ temp845;
    assign temp847 = temp846 ^ temp846;
    assign temp848 = temp847 ^ temp847;
    assign temp849 = temp848 ^ temp848;
    assign temp850 = temp849 ^ temp849;
    assign temp851 = temp850 ^ temp850;
    assign temp852 = temp851 ^ temp851;
    assign temp853 = temp852 ^ temp852;
    assign temp854 = temp853 ^ temp853;
    assign temp855 = temp854 ^ temp854;
    assign temp856 = temp855 ^ temp855;
    assign temp857 = temp856 ^ temp856;
    assign temp858 = temp857 ^ temp857;
    assign temp859 = temp858 ^ temp858;
    assign temp860 = temp859 ^ temp859;
    assign temp861 = temp860 ^ temp860;
    assign temp862 = temp861 ^ temp861;
    assign temp863 = temp862 ^ temp862;
    assign temp864 = temp863 ^ temp863;
    assign temp865 = temp864 ^ temp864;
    assign temp866 = temp865 ^ temp865;
    assign temp867 = temp866 ^ temp866;
    assign temp868 = temp867 ^ temp867;
    assign temp869 = temp868 ^ temp868;
    assign temp870 = temp869 ^ temp869;
    assign temp871 = temp870 ^ temp870;
    assign temp872 = temp871 ^ temp871;
    assign temp873 = temp872 ^ temp872;
    assign temp874 = temp873 ^ temp873;
    assign temp875 = temp874 ^ temp874;
    assign temp876 = temp875 ^ temp875;
    assign temp877 = temp876 ^ temp876;
    assign temp878 = temp877 ^ temp877;
    assign temp879 = temp878 ^ temp878;
    assign temp880 = temp879 ^ temp879;
    assign temp881 = temp880 ^ temp880;
    assign temp882 = temp881 ^ temp881;
    assign temp883 = temp882 ^ temp882;
    assign temp884 = temp883 ^ temp883;
    assign temp885 = temp884 ^ temp884;
    assign temp886 = temp885 ^ temp885;
    assign temp887 = temp886 ^ temp886;
    assign temp888 = temp887 ^ temp887;
    assign temp889 = temp888 ^ temp888;
    assign temp890 = temp889 ^ temp889;
    assign temp891 = temp890 ^ temp890;
    assign temp892 = temp891 ^ temp891;
    assign temp893 = temp892 ^ temp892;
    assign temp894 = temp893 ^ temp893;
    assign temp895 = temp894 ^ temp894;
    assign temp896 = temp895 ^ temp895;
    assign temp897 = temp896 ^ temp896;
    assign temp898 = temp897 ^ temp897;
    assign temp899 = temp898 ^ temp898;
    assign temp900 = temp899 ^ temp899;
    assign temp901 = temp900 ^ temp900;
    assign temp902 = temp901 ^ temp901;
    assign temp903 = temp902 ^ temp902;
    assign temp904 = temp903 ^ temp903;
    assign temp905 = temp904 ^ temp904;
    assign temp906 = temp905 ^ temp905;
    assign temp907 = temp906 ^ temp906;
    assign temp908 = temp907 ^ temp907;
    assign temp909 = temp908 ^ temp908;
    assign temp910 = temp909 ^ temp909;
    assign temp911 = temp910 ^ temp910;
    assign temp912 = temp911 ^ temp911;
    assign temp913 = temp912 ^ temp912;
    assign temp914 = temp913 ^ temp913;
    assign temp915 = temp914 ^ temp914;
    assign temp916 = temp915 ^ temp915;
    assign temp917 = temp916 ^ temp916;
    assign temp918 = temp917 ^ temp917;
    assign temp919 = temp918 ^ temp918;
    assign temp920 = temp919 ^ temp919;
    assign temp921 = temp920 ^ temp920;
    assign temp922 = temp921 ^ temp921;
    assign temp923 = temp922 ^ temp922;
    assign temp924 = temp923 ^ temp923;
    assign temp925 = temp924 ^ temp924;
    assign temp926 = temp925 ^ temp925;
    assign temp927 = temp926 ^ temp926;
    assign temp928 = temp927 ^ temp927;
    assign temp929 = temp928 ^ temp928;
    assign temp930 = temp929 ^ temp929;
    assign temp931 = temp930 ^ temp930;
    assign temp932 = temp931 ^ temp931;
    assign temp933 = temp932 ^ temp932;
    assign temp934 = temp933 ^ temp933;
    assign temp935 = temp934 ^ temp934;
    assign temp936 = temp935 ^ temp935;
    assign temp937 = temp936 ^ temp936;
    assign temp938 = temp937 ^ temp937;
    assign temp939 = temp938 ^ temp938;
    assign temp940 = temp939 ^ temp939;
    assign temp941 = temp940 ^ temp940;
    assign temp942 = temp941 ^ temp941;
    assign temp943 = temp942 ^ temp942;
    assign temp944 = temp943 ^ temp943;
    assign temp945 = temp944 ^ temp944;
    assign temp946 = temp945 ^ temp945;
    assign temp947 = temp946 ^ temp946;
    assign temp948 = temp947 ^ temp947;
    assign temp949 = temp948 ^ temp948;
    assign temp950 = temp949 ^ temp949;
    assign temp951 = temp950 ^ temp950;
    assign temp952 = temp951 ^ temp951;
    assign temp953 = temp952 ^ temp952;
    assign temp954 = temp953 ^ temp953;
    assign temp955 = temp954 ^ temp954;
    assign temp956 = temp955 ^ temp955;
    assign temp957 = temp956 ^ temp956;
    assign temp958 = temp957 ^ temp957;
    assign temp959 = temp958 ^ temp958;
    assign temp960 = temp959 ^ temp959;
    assign temp961 = temp960 ^ temp960;
    assign temp962 = temp961 ^ temp961;
    assign temp963 = temp962 ^ temp962;
    assign temp964 = temp963 ^ temp963;
    assign temp965 = temp964 ^ temp964;
    assign temp966 = temp965 ^ temp965;
    assign temp967 = temp966 ^ temp966;
    assign temp968 = temp967 ^ temp967;
    assign temp969 = temp968 ^ temp968;
    assign temp970 = temp969 ^ temp969;
    assign temp971 = temp970 ^ temp970;
    assign temp972 = temp971 ^ temp971;
    assign temp973 = temp972 ^ temp972;
    assign temp974 = temp973 ^ temp973;
    assign temp975 = temp974 ^ temp974;
    assign temp976 = temp975 ^ temp975;
    assign temp977 = temp976 ^ temp976;
    assign temp978 = temp977 ^ temp977;
    assign temp979 = temp978 ^ temp978;
    assign temp980 = temp979 ^ temp979;
    assign temp981 = temp980 ^ temp980;
    assign temp982 = temp981 ^ temp981;
    assign temp983 = temp982 ^ temp982;
    assign temp984 = temp983 ^ temp983;
    assign temp985 = temp984 ^ temp984;
    assign temp986 = temp985 ^ temp985;
    assign temp987 = temp986 ^ temp986;
    assign temp988 = temp987 ^ temp987;
    assign temp989 = temp988 ^ temp988;
    assign temp990 = temp989 ^ temp989;
    assign temp991 = temp990 ^ temp990;
    assign temp992 = temp991 ^ temp991;
    assign temp993 = temp992 ^ temp992;
    assign temp994 = temp993 ^ temp993;
    assign temp995 = temp994 ^ temp994;
    assign temp996 = temp995 ^ temp995;
    assign temp997 = temp996 ^ temp996;
    assign temp998 = temp997 ^ temp997;
    assign z = temp998 ^ temp998;


endmodule