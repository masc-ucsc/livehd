
module punch.gld(output logic [3:0] total);

  assign total = 9;

endmodule
