

module blackbox(input a, input b, output c);

  potato potato1(.a(a), .b(b), .c(c));

endmodule

